module housekeeping (debug_in,
    debug_mode,
    debug_oeb,
    debug_out,
    pad_flash_clk,
    pad_flash_clk_oeb,
    pad_flash_csb,
    pad_flash_csb_oeb,
    pad_flash_io0_di,
    pad_flash_io0_do,
    pad_flash_io0_ieb,
    pad_flash_io0_oeb,
    pad_flash_io1_di,
    pad_flash_io1_do,
    pad_flash_io1_ieb,
    pad_flash_io1_oeb,
    pll_bypass,
    pll_dco_ena,
    pll_ena,
    porb,
    qspi_enabled,
    reset,
    ser_rx,
    ser_tx,
    serial_clock,
    serial_data_1,
    serial_data_2,
    serial_load,
    serial_resetn,
    spi_csb,
    spi_enabled,
    spi_sck,
    spi_sdi,
    spi_sdo,
    spi_sdoenb,
    spimemio_flash_clk,
    spimemio_flash_csb,
    spimemio_flash_io0_di,
    spimemio_flash_io0_do,
    spimemio_flash_io0_oeb,
    spimemio_flash_io1_di,
    spimemio_flash_io1_do,
    spimemio_flash_io1_oeb,
    spimemio_flash_io2_di,
    spimemio_flash_io2_do,
    spimemio_flash_io2_oeb,
    spimemio_flash_io3_di,
    spimemio_flash_io3_do,
    spimemio_flash_io3_oeb,
    sram_ro_clk,
    sram_ro_csb,
    trap,
    uart_enabled,
    user_clock,
    usr1_vcc_pwrgood,
    usr1_vdd_pwrgood,
    usr2_vcc_pwrgood,
    usr2_vdd_pwrgood,
    wb_ack_o,
    wb_clk_i,
    wb_cyc_i,
    wb_rstn_i,
    wb_stb_i,
    wb_we_i,
    irq,
    mask_rev_in,
    mgmt_gpio_in,
    mgmt_gpio_oeb,
    mgmt_gpio_out,
    pll90_sel,
    pll_div,
    pll_sel,
    pll_trim,
    pwr_ctrl_out,
    sram_ro_addr,
    sram_ro_data,
    wb_adr_i,
    wb_dat_i,
    wb_dat_o,
    wb_sel_i);
 output debug_in;
 input debug_mode;
 input debug_oeb;
 input debug_out;
 output pad_flash_clk;
 output pad_flash_clk_oeb;
 output pad_flash_csb;
 output pad_flash_csb_oeb;
 input pad_flash_io0_di;
 output pad_flash_io0_do;
 output pad_flash_io0_ieb;
 output pad_flash_io0_oeb;
 input pad_flash_io1_di;
 output pad_flash_io1_do;
 output pad_flash_io1_ieb;
 output pad_flash_io1_oeb;
 output pll_bypass;
 output pll_dco_ena;
 output pll_ena;
 input porb;
 input qspi_enabled;
 output reset;
 output ser_rx;
 input ser_tx;
 output serial_clock;
 output serial_data_1;
 output serial_data_2;
 output serial_load;
 output serial_resetn;
 input spi_csb;
 input spi_enabled;
 input spi_sck;
 output spi_sdi;
 input spi_sdo;
 input spi_sdoenb;
 input spimemio_flash_clk;
 input spimemio_flash_csb;
 output spimemio_flash_io0_di;
 input spimemio_flash_io0_do;
 input spimemio_flash_io0_oeb;
 output spimemio_flash_io1_di;
 input spimemio_flash_io1_do;
 input spimemio_flash_io1_oeb;
 output spimemio_flash_io2_di;
 input spimemio_flash_io2_do;
 input spimemio_flash_io2_oeb;
 output spimemio_flash_io3_di;
 input spimemio_flash_io3_do;
 input spimemio_flash_io3_oeb;
 output sram_ro_clk;
 output sram_ro_csb;
 input trap;
 input uart_enabled;
 input user_clock;
 input usr1_vcc_pwrgood;
 input usr1_vdd_pwrgood;
 input usr2_vcc_pwrgood;
 input usr2_vdd_pwrgood;
 output wb_ack_o;
 input wb_clk_i;
 input wb_cyc_i;
 input wb_rstn_i;
 input wb_stb_i;
 input wb_we_i;
 output [2:0] irq;
 input [31:0] mask_rev_in;
 input [37:0] mgmt_gpio_in;
 output [37:0] mgmt_gpio_oeb;
 output [37:0] mgmt_gpio_out;
 output [2:0] pll90_sel;
 output [4:0] pll_div;
 output [2:0] pll_sel;
 output [25:0] pll_trim;
 output [3:0] pwr_ctrl_out;
 output [7:0] sram_ro_addr;
 input [31:0] sram_ro_data;
 input [31:0] wb_adr_i;
 input [31:0] wb_dat_i;
 output [31:0] wb_dat_o;
 input [3:0] wb_sel_i;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire clknet_0_wb_clk_i;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire _1610_;
 wire _1611_;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire _1618_;
 wire _1619_;
 wire _1620_;
 wire _1621_;
 wire _1622_;
 wire _1623_;
 wire _1624_;
 wire _1625_;
 wire _1626_;
 wire _1627_;
 wire _1628_;
 wire _1629_;
 wire _1630_;
 wire _1631_;
 wire _1632_;
 wire _1633_;
 wire _1634_;
 wire _1635_;
 wire _1636_;
 wire _1637_;
 wire _1638_;
 wire _1639_;
 wire _1640_;
 wire _1641_;
 wire _1642_;
 wire _1643_;
 wire _1644_;
 wire _1645_;
 wire _1646_;
 wire _1647_;
 wire _1648_;
 wire _1649_;
 wire _1650_;
 wire _1651_;
 wire _1652_;
 wire _1653_;
 wire _1654_;
 wire _1655_;
 wire _1656_;
 wire _1657_;
 wire _1658_;
 wire _1659_;
 wire _1660_;
 wire _1661_;
 wire _1662_;
 wire _1663_;
 wire _1664_;
 wire _1665_;
 wire _1666_;
 wire _1667_;
 wire _1668_;
 wire _1669_;
 wire _1670_;
 wire _1671_;
 wire _1672_;
 wire _1673_;
 wire _1674_;
 wire _1675_;
 wire _1676_;
 wire _1677_;
 wire _1678_;
 wire _1679_;
 wire _1680_;
 wire _1681_;
 wire _1682_;
 wire _1683_;
 wire _1684_;
 wire _1685_;
 wire _1686_;
 wire _1687_;
 wire _1688_;
 wire _1689_;
 wire _1690_;
 wire _1691_;
 wire _1692_;
 wire _1693_;
 wire _1694_;
 wire _1695_;
 wire _1696_;
 wire _1697_;
 wire _1698_;
 wire _1699_;
 wire _1700_;
 wire _1701_;
 wire _1702_;
 wire _1703_;
 wire _1704_;
 wire _1705_;
 wire _1706_;
 wire _1707_;
 wire _1708_;
 wire _1709_;
 wire _1710_;
 wire _1711_;
 wire _1712_;
 wire _1713_;
 wire _1714_;
 wire _1715_;
 wire _1716_;
 wire _1717_;
 wire _1718_;
 wire _1719_;
 wire _1720_;
 wire _1721_;
 wire _1722_;
 wire _1723_;
 wire _1724_;
 wire _1725_;
 wire _1726_;
 wire _1727_;
 wire _1728_;
 wire _1729_;
 wire _1730_;
 wire _1731_;
 wire _1732_;
 wire _1733_;
 wire _1734_;
 wire _1735_;
 wire _1736_;
 wire _1737_;
 wire _1738_;
 wire _1739_;
 wire _1740_;
 wire _1741_;
 wire _1742_;
 wire _1743_;
 wire _1744_;
 wire _1745_;
 wire _1746_;
 wire _1747_;
 wire _1748_;
 wire _1749_;
 wire _1750_;
 wire _1751_;
 wire _1752_;
 wire _1753_;
 wire _1754_;
 wire _1755_;
 wire _1756_;
 wire _1757_;
 wire _1758_;
 wire _1759_;
 wire _1760_;
 wire _1761_;
 wire _1762_;
 wire _1763_;
 wire _1764_;
 wire _1765_;
 wire _1766_;
 wire _1767_;
 wire _1768_;
 wire _1769_;
 wire _1770_;
 wire _1771_;
 wire _1772_;
 wire _1773_;
 wire _1774_;
 wire _1775_;
 wire _1776_;
 wire _1777_;
 wire _1778_;
 wire _1779_;
 wire _1780_;
 wire _1781_;
 wire _1782_;
 wire _1783_;
 wire _1784_;
 wire _1785_;
 wire _1786_;
 wire _1787_;
 wire _1788_;
 wire _1789_;
 wire _1790_;
 wire _1791_;
 wire _1792_;
 wire _1793_;
 wire _1794_;
 wire _1795_;
 wire _1796_;
 wire _1797_;
 wire _1798_;
 wire _1799_;
 wire _1800_;
 wire _1801_;
 wire _1802_;
 wire _1803_;
 wire _1804_;
 wire _1805_;
 wire _1806_;
 wire _1807_;
 wire _1808_;
 wire _1809_;
 wire _1810_;
 wire _1811_;
 wire _1812_;
 wire _1813_;
 wire _1814_;
 wire _1815_;
 wire _1816_;
 wire _1817_;
 wire _1818_;
 wire _1819_;
 wire _1820_;
 wire _1821_;
 wire _1822_;
 wire _1823_;
 wire _1824_;
 wire _1825_;
 wire _1826_;
 wire _1827_;
 wire _1828_;
 wire _1829_;
 wire _1830_;
 wire _1831_;
 wire _1832_;
 wire _1833_;
 wire _1834_;
 wire _1835_;
 wire _1836_;
 wire _1837_;
 wire _1838_;
 wire _1839_;
 wire _1840_;
 wire _1841_;
 wire _1842_;
 wire _1843_;
 wire _1844_;
 wire _1845_;
 wire _1846_;
 wire _1847_;
 wire _1848_;
 wire _1849_;
 wire _1850_;
 wire _1851_;
 wire _1852_;
 wire _1853_;
 wire _1854_;
 wire _1855_;
 wire _1856_;
 wire _1857_;
 wire _1858_;
 wire _1859_;
 wire _1860_;
 wire _1861_;
 wire _1862_;
 wire _1863_;
 wire _1864_;
 wire _1865_;
 wire _1866_;
 wire _1867_;
 wire _1868_;
 wire _1869_;
 wire _1870_;
 wire _1871_;
 wire _1872_;
 wire _1873_;
 wire _1874_;
 wire _1875_;
 wire _1876_;
 wire _1877_;
 wire _1878_;
 wire _1879_;
 wire _1880_;
 wire _1881_;
 wire _1882_;
 wire _1883_;
 wire _1884_;
 wire _1885_;
 wire _1886_;
 wire _1887_;
 wire _1888_;
 wire _1889_;
 wire _1890_;
 wire _1891_;
 wire _1892_;
 wire _1893_;
 wire _1894_;
 wire _1895_;
 wire _1896_;
 wire _1897_;
 wire _1898_;
 wire _1899_;
 wire _1900_;
 wire _1901_;
 wire _1902_;
 wire _1903_;
 wire _1904_;
 wire _1905_;
 wire _1906_;
 wire _1907_;
 wire _1908_;
 wire _1909_;
 wire _1910_;
 wire _1911_;
 wire _1912_;
 wire _1913_;
 wire _1914_;
 wire _1915_;
 wire _1916_;
 wire _1917_;
 wire _1918_;
 wire _1919_;
 wire _1920_;
 wire _1921_;
 wire _1922_;
 wire _1923_;
 wire _1924_;
 wire _1925_;
 wire _1926_;
 wire _1927_;
 wire _1928_;
 wire _1929_;
 wire _1930_;
 wire _1931_;
 wire _1932_;
 wire _1933_;
 wire _1934_;
 wire _1935_;
 wire _1936_;
 wire _1937_;
 wire _1938_;
 wire _1939_;
 wire _1940_;
 wire _1941_;
 wire _1942_;
 wire _1943_;
 wire _1944_;
 wire _1945_;
 wire _1946_;
 wire _1947_;
 wire _1948_;
 wire _1949_;
 wire _1950_;
 wire _1951_;
 wire _1952_;
 wire _1953_;
 wire _1954_;
 wire _1955_;
 wire _1956_;
 wire _1957_;
 wire _1958_;
 wire _1959_;
 wire _1960_;
 wire _1961_;
 wire _1962_;
 wire _1963_;
 wire _1964_;
 wire _1965_;
 wire _1966_;
 wire _1967_;
 wire _1968_;
 wire _1969_;
 wire _1970_;
 wire _1971_;
 wire _1972_;
 wire _1973_;
 wire _1974_;
 wire _1975_;
 wire _1976_;
 wire _1977_;
 wire _1978_;
 wire _1979_;
 wire _1980_;
 wire _1981_;
 wire _1982_;
 wire _1983_;
 wire _1984_;
 wire _1985_;
 wire _1986_;
 wire _1987_;
 wire _1988_;
 wire _1989_;
 wire _1990_;
 wire _1991_;
 wire _1992_;
 wire _1993_;
 wire _1994_;
 wire _1995_;
 wire _1996_;
 wire _1997_;
 wire _1998_;
 wire _1999_;
 wire _2000_;
 wire _2001_;
 wire _2002_;
 wire _2003_;
 wire _2004_;
 wire _2005_;
 wire _2006_;
 wire _2007_;
 wire _2008_;
 wire _2009_;
 wire _2010_;
 wire _2011_;
 wire _2012_;
 wire _2013_;
 wire _2014_;
 wire _2015_;
 wire _2016_;
 wire _2017_;
 wire _2018_;
 wire _2019_;
 wire _2020_;
 wire _2021_;
 wire _2022_;
 wire _2023_;
 wire _2024_;
 wire _2025_;
 wire _2026_;
 wire _2027_;
 wire _2028_;
 wire _2029_;
 wire _2030_;
 wire _2031_;
 wire _2032_;
 wire _2033_;
 wire _2034_;
 wire _2035_;
 wire _2036_;
 wire _2037_;
 wire _2038_;
 wire _2039_;
 wire _2040_;
 wire _2041_;
 wire _2042_;
 wire _2043_;
 wire _2044_;
 wire _2045_;
 wire _2046_;
 wire _2047_;
 wire _2048_;
 wire _2049_;
 wire _2050_;
 wire _2051_;
 wire _2052_;
 wire _2053_;
 wire _2054_;
 wire _2055_;
 wire _2056_;
 wire _2057_;
 wire _2058_;
 wire _2059_;
 wire _2060_;
 wire _2061_;
 wire _2062_;
 wire _2063_;
 wire _2064_;
 wire _2065_;
 wire _2066_;
 wire _2067_;
 wire _2068_;
 wire _2069_;
 wire _2070_;
 wire _2071_;
 wire _2072_;
 wire _2073_;
 wire _2074_;
 wire _2075_;
 wire _2076_;
 wire _2077_;
 wire _2078_;
 wire _2079_;
 wire _2080_;
 wire _2081_;
 wire _2082_;
 wire _2083_;
 wire _2084_;
 wire _2085_;
 wire _2086_;
 wire _2087_;
 wire _2088_;
 wire _2089_;
 wire _2090_;
 wire _2091_;
 wire _2092_;
 wire _2093_;
 wire _2094_;
 wire _2095_;
 wire _2096_;
 wire _2097_;
 wire _2098_;
 wire _2099_;
 wire _2100_;
 wire _2101_;
 wire _2102_;
 wire _2103_;
 wire _2104_;
 wire _2105_;
 wire _2106_;
 wire _2107_;
 wire _2108_;
 wire _2109_;
 wire _2110_;
 wire _2111_;
 wire _2112_;
 wire _2113_;
 wire _2114_;
 wire _2115_;
 wire _2116_;
 wire _2117_;
 wire _2118_;
 wire _2119_;
 wire _2120_;
 wire _2121_;
 wire _2122_;
 wire _2123_;
 wire _2124_;
 wire _2125_;
 wire _2126_;
 wire _2127_;
 wire _2128_;
 wire _2129_;
 wire _2130_;
 wire _2131_;
 wire _2132_;
 wire _2133_;
 wire _2134_;
 wire _2135_;
 wire _2136_;
 wire _2137_;
 wire _2138_;
 wire _2139_;
 wire _2140_;
 wire _2141_;
 wire _2142_;
 wire _2143_;
 wire _2144_;
 wire _2145_;
 wire _2146_;
 wire _2147_;
 wire _2148_;
 wire _2149_;
 wire _2150_;
 wire _2151_;
 wire _2152_;
 wire _2153_;
 wire _2154_;
 wire _2155_;
 wire _2156_;
 wire _2157_;
 wire _2158_;
 wire _2159_;
 wire _2160_;
 wire _2161_;
 wire _2162_;
 wire _2163_;
 wire _2164_;
 wire _2165_;
 wire _2166_;
 wire _2167_;
 wire _2168_;
 wire _2169_;
 wire _2170_;
 wire _2171_;
 wire _2172_;
 wire _2173_;
 wire _2174_;
 wire _2175_;
 wire _2176_;
 wire _2177_;
 wire _2178_;
 wire _2179_;
 wire _2180_;
 wire _2181_;
 wire _2182_;
 wire _2183_;
 wire _2184_;
 wire _2185_;
 wire _2186_;
 wire _2187_;
 wire _2188_;
 wire _2189_;
 wire _2190_;
 wire _2191_;
 wire _2192_;
 wire _2193_;
 wire _2194_;
 wire _2195_;
 wire _2196_;
 wire _2197_;
 wire _2198_;
 wire _2199_;
 wire _2200_;
 wire _2201_;
 wire _2202_;
 wire _2203_;
 wire _2204_;
 wire _2205_;
 wire _2206_;
 wire _2207_;
 wire _2208_;
 wire _2209_;
 wire _2210_;
 wire _2211_;
 wire _2212_;
 wire _2213_;
 wire _2214_;
 wire _2215_;
 wire _2216_;
 wire _2217_;
 wire _2218_;
 wire _2219_;
 wire _2220_;
 wire _2221_;
 wire _2222_;
 wire _2223_;
 wire _2224_;
 wire _2225_;
 wire _2226_;
 wire _2227_;
 wire _2228_;
 wire _2229_;
 wire _2230_;
 wire _2231_;
 wire _2232_;
 wire _2233_;
 wire _2234_;
 wire _2235_;
 wire _2236_;
 wire _2237_;
 wire _2238_;
 wire _2239_;
 wire _2240_;
 wire _2241_;
 wire _2242_;
 wire _2243_;
 wire _2244_;
 wire _2245_;
 wire _2246_;
 wire _2247_;
 wire _2248_;
 wire _2249_;
 wire _2250_;
 wire _2251_;
 wire _2252_;
 wire _2253_;
 wire _2254_;
 wire _2255_;
 wire _2256_;
 wire _2257_;
 wire _2258_;
 wire _2259_;
 wire _2260_;
 wire _2261_;
 wire _2262_;
 wire _2263_;
 wire _2264_;
 wire _2265_;
 wire _2266_;
 wire _2267_;
 wire _2268_;
 wire _2269_;
 wire _2270_;
 wire _2271_;
 wire _2272_;
 wire _2273_;
 wire _2274_;
 wire _2275_;
 wire _2276_;
 wire _2277_;
 wire _2278_;
 wire _2279_;
 wire _2280_;
 wire _2281_;
 wire _2282_;
 wire _2283_;
 wire _2284_;
 wire _2285_;
 wire _2286_;
 wire _2287_;
 wire _2288_;
 wire _2289_;
 wire _2290_;
 wire _2291_;
 wire _2292_;
 wire _2293_;
 wire _2294_;
 wire _2295_;
 wire _2296_;
 wire _2297_;
 wire _2298_;
 wire _2299_;
 wire _2300_;
 wire _2301_;
 wire _2302_;
 wire _2303_;
 wire _2304_;
 wire _2305_;
 wire _2306_;
 wire _2307_;
 wire _2308_;
 wire _2309_;
 wire _2310_;
 wire _2311_;
 wire _2312_;
 wire _2313_;
 wire _2314_;
 wire _2315_;
 wire _2316_;
 wire _2317_;
 wire _2318_;
 wire _2319_;
 wire _2320_;
 wire _2321_;
 wire _2322_;
 wire _2323_;
 wire _2324_;
 wire _2325_;
 wire _2326_;
 wire _2327_;
 wire _2328_;
 wire _2329_;
 wire _2330_;
 wire _2331_;
 wire _2332_;
 wire _2333_;
 wire _2334_;
 wire _2335_;
 wire _2336_;
 wire _2337_;
 wire _2338_;
 wire _2339_;
 wire _2340_;
 wire _2341_;
 wire _2342_;
 wire _2343_;
 wire _2344_;
 wire _2345_;
 wire _2346_;
 wire _2347_;
 wire _2348_;
 wire _2349_;
 wire _2350_;
 wire _2351_;
 wire _2352_;
 wire _2353_;
 wire _2354_;
 wire _2355_;
 wire _2356_;
 wire _2357_;
 wire _2358_;
 wire _2359_;
 wire _2360_;
 wire _2361_;
 wire _2362_;
 wire _2363_;
 wire _2364_;
 wire _2365_;
 wire _2366_;
 wire _2367_;
 wire _2368_;
 wire _2369_;
 wire _2370_;
 wire _2371_;
 wire _2372_;
 wire _2373_;
 wire _2374_;
 wire _2375_;
 wire _2376_;
 wire _2377_;
 wire _2378_;
 wire _2379_;
 wire _2380_;
 wire _2381_;
 wire _2382_;
 wire _2383_;
 wire _2384_;
 wire _2385_;
 wire _2386_;
 wire _2387_;
 wire _2388_;
 wire _2389_;
 wire _2390_;
 wire _2391_;
 wire _2392_;
 wire _2393_;
 wire _2394_;
 wire _2395_;
 wire _2396_;
 wire _2397_;
 wire _2398_;
 wire _2399_;
 wire _2400_;
 wire _2401_;
 wire _2402_;
 wire _2403_;
 wire _2404_;
 wire _2405_;
 wire _2406_;
 wire _2407_;
 wire _2408_;
 wire _2409_;
 wire _2410_;
 wire _2411_;
 wire _2412_;
 wire _2413_;
 wire _2414_;
 wire _2415_;
 wire _2416_;
 wire _2417_;
 wire _2418_;
 wire _2419_;
 wire _2420_;
 wire _2421_;
 wire _2422_;
 wire _2423_;
 wire _2424_;
 wire _2425_;
 wire _2426_;
 wire _2427_;
 wire _2428_;
 wire _2429_;
 wire _2430_;
 wire _2431_;
 wire _2432_;
 wire _2433_;
 wire _2434_;
 wire _2435_;
 wire _2436_;
 wire _2437_;
 wire _2438_;
 wire _2439_;
 wire _2440_;
 wire _2441_;
 wire _2442_;
 wire _2443_;
 wire _2444_;
 wire _2445_;
 wire _2446_;
 wire _2447_;
 wire _2448_;
 wire _2449_;
 wire _2450_;
 wire _2451_;
 wire _2452_;
 wire _2453_;
 wire _2454_;
 wire _2455_;
 wire _2456_;
 wire _2457_;
 wire _2458_;
 wire _2459_;
 wire _2460_;
 wire _2461_;
 wire _2462_;
 wire _2463_;
 wire _2464_;
 wire _2465_;
 wire _2466_;
 wire _2467_;
 wire _2468_;
 wire _2469_;
 wire _2470_;
 wire _2471_;
 wire _2472_;
 wire _2473_;
 wire _2474_;
 wire _2475_;
 wire _2476_;
 wire _2477_;
 wire _2478_;
 wire _2479_;
 wire _2480_;
 wire _2481_;
 wire _2482_;
 wire _2483_;
 wire _2484_;
 wire _2485_;
 wire _2486_;
 wire _2487_;
 wire _2488_;
 wire _2489_;
 wire _2490_;
 wire _2491_;
 wire _2492_;
 wire _2493_;
 wire _2494_;
 wire _2495_;
 wire _2496_;
 wire _2497_;
 wire _2498_;
 wire _2499_;
 wire _2500_;
 wire _2501_;
 wire _2502_;
 wire _2503_;
 wire _2504_;
 wire _2505_;
 wire _2506_;
 wire _2507_;
 wire _2508_;
 wire _2509_;
 wire _2510_;
 wire _2511_;
 wire _2512_;
 wire _2513_;
 wire _2514_;
 wire _2515_;
 wire _2516_;
 wire _2517_;
 wire _2518_;
 wire _2519_;
 wire _2520_;
 wire _2521_;
 wire _2522_;
 wire _2523_;
 wire _2524_;
 wire _2525_;
 wire _2526_;
 wire _2527_;
 wire _2528_;
 wire _2529_;
 wire _2530_;
 wire _2531_;
 wire _2532_;
 wire _2533_;
 wire _2534_;
 wire _2535_;
 wire _2536_;
 wire _2537_;
 wire _2538_;
 wire _2539_;
 wire _2540_;
 wire _2541_;
 wire _2542_;
 wire _2543_;
 wire _2544_;
 wire _2545_;
 wire _2546_;
 wire _2547_;
 wire _2548_;
 wire _2549_;
 wire _2550_;
 wire _2551_;
 wire _2552_;
 wire _2553_;
 wire _2554_;
 wire _2555_;
 wire _2556_;
 wire _2557_;
 wire _2558_;
 wire _2559_;
 wire _2560_;
 wire _2561_;
 wire _2562_;
 wire _2563_;
 wire _2564_;
 wire _2565_;
 wire _2566_;
 wire _2567_;
 wire _2568_;
 wire _2569_;
 wire _2570_;
 wire _2571_;
 wire _2572_;
 wire _2573_;
 wire _2574_;
 wire _2575_;
 wire _2576_;
 wire _2577_;
 wire _2578_;
 wire _2579_;
 wire _2580_;
 wire _2581_;
 wire _2582_;
 wire _2583_;
 wire _2584_;
 wire _2585_;
 wire _2586_;
 wire _2587_;
 wire _2588_;
 wire _2589_;
 wire _2590_;
 wire _2591_;
 wire _2592_;
 wire _2593_;
 wire _2594_;
 wire _2595_;
 wire _2596_;
 wire _2597_;
 wire _2598_;
 wire _2599_;
 wire _2600_;
 wire _2601_;
 wire _2602_;
 wire _2603_;
 wire _2604_;
 wire _2605_;
 wire _2606_;
 wire _2607_;
 wire _2608_;
 wire _2609_;
 wire _2610_;
 wire _2611_;
 wire _2612_;
 wire _2613_;
 wire _2614_;
 wire _2615_;
 wire _2616_;
 wire _2617_;
 wire _2618_;
 wire _2619_;
 wire _2620_;
 wire _2621_;
 wire _2622_;
 wire _2623_;
 wire _2624_;
 wire _2625_;
 wire _2626_;
 wire _2627_;
 wire _2628_;
 wire _2629_;
 wire _2630_;
 wire _2631_;
 wire _2632_;
 wire _2633_;
 wire _2634_;
 wire _2635_;
 wire _2636_;
 wire _2637_;
 wire _2638_;
 wire _2639_;
 wire _2640_;
 wire _2641_;
 wire _2642_;
 wire _2643_;
 wire _2644_;
 wire _2645_;
 wire _2646_;
 wire _2647_;
 wire _2648_;
 wire _2649_;
 wire _2650_;
 wire _2651_;
 wire _2652_;
 wire _2653_;
 wire _2654_;
 wire _2655_;
 wire _2656_;
 wire _2657_;
 wire _2658_;
 wire _2659_;
 wire _2660_;
 wire _2661_;
 wire _2662_;
 wire _2663_;
 wire _2664_;
 wire _2665_;
 wire _2666_;
 wire _2667_;
 wire _2668_;
 wire _2669_;
 wire _2670_;
 wire _2671_;
 wire _2672_;
 wire _2673_;
 wire _2674_;
 wire _2675_;
 wire _2676_;
 wire _2677_;
 wire _2678_;
 wire _2679_;
 wire _2680_;
 wire _2681_;
 wire _2682_;
 wire _2683_;
 wire _2684_;
 wire _2685_;
 wire _2686_;
 wire _2687_;
 wire _2688_;
 wire _2689_;
 wire _2690_;
 wire _2691_;
 wire _2692_;
 wire _2693_;
 wire _2694_;
 wire _2695_;
 wire _2696_;
 wire _2697_;
 wire _2698_;
 wire _2699_;
 wire _2700_;
 wire _2701_;
 wire _2702_;
 wire _2703_;
 wire _2704_;
 wire _2705_;
 wire _2706_;
 wire _2707_;
 wire _2708_;
 wire _2709_;
 wire _2710_;
 wire _2711_;
 wire _2712_;
 wire _2713_;
 wire _2714_;
 wire _2715_;
 wire _2716_;
 wire _2717_;
 wire _2718_;
 wire _2719_;
 wire _2720_;
 wire _2721_;
 wire _2722_;
 wire _2723_;
 wire _2724_;
 wire _2725_;
 wire _2726_;
 wire _2727_;
 wire _2728_;
 wire _2729_;
 wire _2730_;
 wire _2731_;
 wire _2732_;
 wire _2733_;
 wire _2734_;
 wire _2735_;
 wire _2736_;
 wire _2737_;
 wire _2738_;
 wire _2739_;
 wire _2740_;
 wire _2741_;
 wire _2742_;
 wire _2743_;
 wire _2744_;
 wire _2745_;
 wire _2746_;
 wire _2747_;
 wire _2748_;
 wire _2749_;
 wire _2750_;
 wire _2751_;
 wire _2752_;
 wire _2753_;
 wire _2754_;
 wire _2755_;
 wire _2756_;
 wire _2757_;
 wire _2758_;
 wire _2759_;
 wire _2760_;
 wire _2761_;
 wire _2762_;
 wire _2763_;
 wire _2764_;
 wire _2765_;
 wire _2766_;
 wire _2767_;
 wire _2768_;
 wire _2769_;
 wire _2770_;
 wire _2771_;
 wire _2772_;
 wire _2773_;
 wire _2774_;
 wire _2775_;
 wire _2776_;
 wire _2777_;
 wire _2778_;
 wire _2779_;
 wire _2780_;
 wire _2781_;
 wire _2782_;
 wire _2783_;
 wire _2784_;
 wire _2785_;
 wire _2786_;
 wire _2787_;
 wire _2788_;
 wire _2789_;
 wire _2790_;
 wire _2791_;
 wire _2792_;
 wire _2793_;
 wire _2794_;
 wire _2795_;
 wire _2796_;
 wire _2797_;
 wire _2798_;
 wire _2799_;
 wire _2800_;
 wire _2801_;
 wire _2802_;
 wire _2803_;
 wire _2804_;
 wire _2805_;
 wire _2806_;
 wire _2807_;
 wire _2808_;
 wire _2809_;
 wire _2810_;
 wire _2811_;
 wire _2812_;
 wire _2813_;
 wire _2814_;
 wire _2815_;
 wire _2816_;
 wire _2817_;
 wire _2818_;
 wire _2819_;
 wire _2820_;
 wire _2821_;
 wire _2822_;
 wire _2823_;
 wire _2824_;
 wire _2825_;
 wire _2826_;
 wire _2827_;
 wire _2828_;
 wire _2829_;
 wire _2830_;
 wire _2831_;
 wire _2832_;
 wire _2833_;
 wire _2834_;
 wire _2835_;
 wire _2836_;
 wire _2837_;
 wire _2838_;
 wire _2839_;
 wire _2840_;
 wire _2841_;
 wire _2842_;
 wire _2843_;
 wire _2844_;
 wire _2845_;
 wire _2846_;
 wire _2847_;
 wire _2848_;
 wire _2849_;
 wire _2850_;
 wire _2851_;
 wire _2852_;
 wire _2853_;
 wire _2854_;
 wire _2855_;
 wire _2856_;
 wire _2857_;
 wire _2858_;
 wire _2859_;
 wire _2860_;
 wire _2861_;
 wire _2862_;
 wire _2863_;
 wire _2864_;
 wire _2865_;
 wire _2866_;
 wire _2867_;
 wire _2868_;
 wire _2869_;
 wire _2870_;
 wire _2871_;
 wire _2872_;
 wire _2873_;
 wire _2874_;
 wire _2875_;
 wire _2876_;
 wire _2877_;
 wire _2878_;
 wire _2879_;
 wire _2880_;
 wire _2881_;
 wire _2882_;
 wire _2883_;
 wire _2884_;
 wire _2885_;
 wire _2886_;
 wire _2887_;
 wire _2888_;
 wire _2889_;
 wire _2890_;
 wire _2891_;
 wire _2892_;
 wire _2893_;
 wire _2894_;
 wire _2895_;
 wire _2896_;
 wire _2897_;
 wire _2898_;
 wire _2899_;
 wire _2900_;
 wire _2901_;
 wire _2902_;
 wire _2903_;
 wire _2904_;
 wire _2905_;
 wire _2906_;
 wire _2907_;
 wire _2908_;
 wire _2909_;
 wire _2910_;
 wire _2911_;
 wire _2912_;
 wire _2913_;
 wire _2914_;
 wire _2915_;
 wire _2916_;
 wire _2917_;
 wire _2918_;
 wire _2919_;
 wire _2920_;
 wire _2921_;
 wire _2922_;
 wire _2923_;
 wire _2924_;
 wire _2925_;
 wire _2926_;
 wire _2927_;
 wire _2928_;
 wire _2929_;
 wire _2930_;
 wire _2931_;
 wire _2932_;
 wire _2933_;
 wire _2934_;
 wire _2935_;
 wire _2936_;
 wire _2937_;
 wire _2938_;
 wire _2939_;
 wire _2940_;
 wire _2941_;
 wire _2942_;
 wire _2943_;
 wire _2944_;
 wire _2945_;
 wire _2946_;
 wire _2947_;
 wire _2948_;
 wire _2949_;
 wire _2950_;
 wire _2951_;
 wire _2952_;
 wire _2953_;
 wire _2954_;
 wire _2955_;
 wire _2956_;
 wire _2957_;
 wire _2958_;
 wire _2959_;
 wire _2960_;
 wire _2961_;
 wire _2962_;
 wire _2963_;
 wire _2964_;
 wire _2965_;
 wire _2966_;
 wire _2967_;
 wire _2968_;
 wire _2969_;
 wire _2970_;
 wire _2971_;
 wire _2972_;
 wire _2973_;
 wire _2974_;
 wire _2975_;
 wire _2976_;
 wire _2977_;
 wire _2978_;
 wire _2979_;
 wire _2980_;
 wire _2981_;
 wire _2982_;
 wire _2983_;
 wire _2984_;
 wire _2985_;
 wire _2986_;
 wire _2987_;
 wire _2988_;
 wire _2989_;
 wire _2990_;
 wire _2991_;
 wire _2992_;
 wire _2993_;
 wire _2994_;
 wire _2995_;
 wire _2996_;
 wire _2997_;
 wire _2998_;
 wire _2999_;
 wire _3000_;
 wire _3001_;
 wire _3002_;
 wire _3003_;
 wire _3004_;
 wire _3005_;
 wire _3006_;
 wire _3007_;
 wire _3008_;
 wire _3009_;
 wire _3010_;
 wire _3011_;
 wire _3012_;
 wire _3013_;
 wire _3014_;
 wire _3015_;
 wire _3016_;
 wire _3017_;
 wire _3018_;
 wire _3019_;
 wire _3020_;
 wire _3021_;
 wire _3022_;
 wire _3023_;
 wire _3024_;
 wire _3025_;
 wire _3026_;
 wire _3027_;
 wire _3028_;
 wire _3029_;
 wire _3030_;
 wire _3031_;
 wire _3032_;
 wire _3033_;
 wire _3034_;
 wire _3035_;
 wire _3036_;
 wire _3037_;
 wire _3038_;
 wire _3039_;
 wire _3040_;
 wire _3041_;
 wire _3042_;
 wire _3043_;
 wire _3044_;
 wire _3045_;
 wire _3046_;
 wire _3047_;
 wire _3048_;
 wire _3049_;
 wire _3050_;
 wire _3051_;
 wire _3052_;
 wire _3053_;
 wire _3054_;
 wire _3055_;
 wire _3056_;
 wire _3057_;
 wire _3058_;
 wire _3059_;
 wire _3060_;
 wire _3061_;
 wire _3062_;
 wire _3063_;
 wire _3064_;
 wire _3065_;
 wire _3066_;
 wire _3067_;
 wire _3068_;
 wire _3069_;
 wire _3070_;
 wire _3071_;
 wire _3072_;
 wire _3073_;
 wire _3074_;
 wire _3075_;
 wire _3076_;
 wire _3077_;
 wire _3078_;
 wire _3079_;
 wire _3080_;
 wire _3081_;
 wire _3082_;
 wire _3083_;
 wire _3084_;
 wire _3085_;
 wire _3086_;
 wire _3087_;
 wire _3088_;
 wire _3089_;
 wire _3090_;
 wire _3091_;
 wire _3092_;
 wire _3093_;
 wire _3094_;
 wire _3095_;
 wire _3096_;
 wire _3097_;
 wire _3098_;
 wire _3099_;
 wire _3100_;
 wire _3101_;
 wire _3102_;
 wire _3103_;
 wire _3104_;
 wire _3105_;
 wire _3106_;
 wire _3107_;
 wire _3108_;
 wire _3109_;
 wire _3110_;
 wire _3111_;
 wire _3112_;
 wire _3113_;
 wire _3114_;
 wire _3115_;
 wire _3116_;
 wire _3117_;
 wire _3118_;
 wire _3119_;
 wire _3120_;
 wire _3121_;
 wire _3122_;
 wire _3123_;
 wire _3124_;
 wire _3125_;
 wire _3126_;
 wire _3127_;
 wire _3128_;
 wire _3129_;
 wire _3130_;
 wire _3131_;
 wire _3132_;
 wire _3133_;
 wire _3134_;
 wire _3135_;
 wire _3136_;
 wire _3137_;
 wire _3138_;
 wire _3139_;
 wire _3140_;
 wire _3141_;
 wire _3142_;
 wire _3143_;
 wire _3144_;
 wire _3145_;
 wire _3146_;
 wire _3147_;
 wire _3148_;
 wire _3149_;
 wire _3150_;
 wire _3151_;
 wire _3152_;
 wire _3153_;
 wire _3154_;
 wire _3155_;
 wire _3156_;
 wire _3157_;
 wire _3158_;
 wire _3159_;
 wire _3160_;
 wire _3161_;
 wire _3162_;
 wire _3163_;
 wire _3164_;
 wire _3165_;
 wire _3166_;
 wire _3167_;
 wire _3168_;
 wire _3169_;
 wire _3170_;
 wire _3171_;
 wire _3172_;
 wire _3173_;
 wire _3174_;
 wire _3175_;
 wire _3176_;
 wire _3177_;
 wire _3178_;
 wire _3179_;
 wire _3180_;
 wire _3181_;
 wire _3182_;
 wire _3183_;
 wire _3184_;
 wire _3185_;
 wire _3186_;
 wire _3187_;
 wire _3188_;
 wire _3189_;
 wire _3190_;
 wire _3191_;
 wire _3192_;
 wire _3193_;
 wire _3194_;
 wire _3195_;
 wire _3196_;
 wire _3197_;
 wire _3198_;
 wire _3199_;
 wire _3200_;
 wire _3201_;
 wire _3202_;
 wire _3203_;
 wire _3204_;
 wire _3205_;
 wire _3206_;
 wire _3207_;
 wire _3208_;
 wire _3209_;
 wire _3210_;
 wire _3211_;
 wire _3212_;
 wire _3213_;
 wire _3214_;
 wire _3215_;
 wire _3216_;
 wire _3217_;
 wire _3218_;
 wire _3219_;
 wire _3220_;
 wire _3221_;
 wire _3222_;
 wire _3223_;
 wire _3224_;
 wire _3225_;
 wire _3226_;
 wire _3227_;
 wire _3228_;
 wire _3229_;
 wire _3230_;
 wire _3231_;
 wire _3232_;
 wire _3233_;
 wire _3234_;
 wire _3235_;
 wire _3236_;
 wire _3237_;
 wire _3238_;
 wire _3239_;
 wire _3240_;
 wire _3241_;
 wire _3242_;
 wire _3243_;
 wire _3244_;
 wire _3245_;
 wire _3246_;
 wire _3247_;
 wire _3248_;
 wire _3249_;
 wire _3250_;
 wire _3251_;
 wire _3252_;
 wire _3253_;
 wire _3254_;
 wire _3255_;
 wire _3256_;
 wire _3257_;
 wire _3258_;
 wire _3259_;
 wire _3260_;
 wire _3261_;
 wire _3262_;
 wire _3263_;
 wire _3264_;
 wire _3265_;
 wire _3266_;
 wire _3267_;
 wire _3268_;
 wire _3269_;
 wire _3270_;
 wire _3271_;
 wire _3272_;
 wire _3273_;
 wire _3274_;
 wire _3275_;
 wire _3276_;
 wire _3277_;
 wire _3278_;
 wire _3279_;
 wire _3280_;
 wire _3281_;
 wire _3282_;
 wire _3283_;
 wire _3284_;
 wire _3285_;
 wire _3286_;
 wire _3287_;
 wire _3288_;
 wire _3289_;
 wire _3290_;
 wire _3291_;
 wire _3292_;
 wire _3293_;
 wire _3294_;
 wire _3295_;
 wire _3296_;
 wire _3297_;
 wire _3298_;
 wire _3299_;
 wire _3300_;
 wire _3301_;
 wire _3302_;
 wire _3303_;
 wire _3304_;
 wire _3305_;
 wire _3306_;
 wire _3307_;
 wire _3308_;
 wire _3309_;
 wire _3310_;
 wire _3311_;
 wire _3312_;
 wire _3313_;
 wire _3314_;
 wire _3315_;
 wire _3316_;
 wire _3317_;
 wire _3318_;
 wire _3319_;
 wire _3320_;
 wire _3321_;
 wire _3322_;
 wire _3323_;
 wire _3324_;
 wire _3325_;
 wire _3326_;
 wire _3327_;
 wire _3328_;
 wire _3329_;
 wire _3330_;
 wire _3331_;
 wire _3332_;
 wire _3333_;
 wire _3334_;
 wire _3335_;
 wire _3336_;
 wire _3337_;
 wire _3338_;
 wire _3339_;
 wire _3340_;
 wire _3341_;
 wire _3342_;
 wire _3343_;
 wire _3344_;
 wire _3345_;
 wire _3346_;
 wire _3347_;
 wire _3348_;
 wire _3349_;
 wire _3350_;
 wire _3351_;
 wire _3352_;
 wire _3353_;
 wire _3354_;
 wire _3355_;
 wire _3356_;
 wire _3357_;
 wire _3358_;
 wire _3359_;
 wire _3360_;
 wire _3361_;
 wire _3362_;
 wire _3363_;
 wire _3364_;
 wire _3365_;
 wire _3366_;
 wire _3367_;
 wire _3368_;
 wire _3369_;
 wire _3370_;
 wire _3371_;
 wire _3372_;
 wire _3373_;
 wire _3374_;
 wire _3375_;
 wire _3376_;
 wire _3377_;
 wire _3378_;
 wire _3379_;
 wire _3380_;
 wire _3381_;
 wire _3382_;
 wire _3383_;
 wire _3384_;
 wire _3385_;
 wire _3386_;
 wire _3387_;
 wire _3388_;
 wire _3389_;
 wire _3390_;
 wire _3391_;
 wire _3392_;
 wire _3393_;
 wire _3394_;
 wire _3395_;
 wire _3396_;
 wire _3397_;
 wire _3398_;
 wire _3399_;
 wire _3400_;
 wire _3401_;
 wire _3402_;
 wire _3403_;
 wire _3404_;
 wire _3405_;
 wire _3406_;
 wire _3407_;
 wire _3408_;
 wire _3409_;
 wire _3410_;
 wire _3411_;
 wire _3412_;
 wire _3413_;
 wire _3414_;
 wire _3415_;
 wire _3416_;
 wire _3417_;
 wire _3418_;
 wire _3419_;
 wire _3420_;
 wire _3421_;
 wire _3422_;
 wire _3423_;
 wire _3424_;
 wire _3425_;
 wire _3426_;
 wire _3427_;
 wire _3428_;
 wire _3429_;
 wire _3430_;
 wire _3431_;
 wire _3432_;
 wire _3433_;
 wire _3434_;
 wire _3435_;
 wire _3436_;
 wire _3437_;
 wire _3438_;
 wire _3439_;
 wire _3440_;
 wire _3441_;
 wire _3442_;
 wire _3443_;
 wire _3444_;
 wire _3445_;
 wire _3446_;
 wire _3447_;
 wire _3448_;
 wire _3449_;
 wire _3450_;
 wire _3451_;
 wire _3452_;
 wire _3453_;
 wire _3454_;
 wire _3455_;
 wire _3456_;
 wire _3457_;
 wire _3458_;
 wire _3459_;
 wire _3460_;
 wire _3461_;
 wire _3462_;
 wire _3463_;
 wire _3464_;
 wire _3465_;
 wire _3466_;
 wire _3467_;
 wire _3468_;
 wire _3469_;
 wire _3470_;
 wire _3471_;
 wire _3472_;
 wire _3473_;
 wire _3474_;
 wire _3475_;
 wire _3476_;
 wire _3477_;
 wire _3478_;
 wire _3479_;
 wire _3480_;
 wire _3481_;
 wire _3482_;
 wire _3483_;
 wire _3484_;
 wire _3485_;
 wire _3486_;
 wire _3487_;
 wire _3488_;
 wire _3489_;
 wire _3490_;
 wire _3491_;
 wire _3492_;
 wire _3493_;
 wire _3494_;
 wire _3495_;
 wire _3496_;
 wire _3497_;
 wire _3498_;
 wire _3499_;
 wire _3500_;
 wire _3501_;
 wire _3502_;
 wire _3503_;
 wire _3504_;
 wire _3505_;
 wire _3506_;
 wire _3507_;
 wire _3508_;
 wire _3509_;
 wire _3510_;
 wire _3511_;
 wire _3512_;
 wire _3513_;
 wire _3514_;
 wire _3515_;
 wire _3516_;
 wire _3517_;
 wire _3518_;
 wire _3519_;
 wire _3520_;
 wire _3521_;
 wire _3522_;
 wire _3523_;
 wire _3524_;
 wire _3525_;
 wire _3526_;
 wire _3527_;
 wire _3528_;
 wire _3529_;
 wire _3530_;
 wire _3531_;
 wire _3532_;
 wire _3533_;
 wire _3534_;
 wire _3535_;
 wire _3536_;
 wire _3537_;
 wire _3538_;
 wire _3539_;
 wire _3540_;
 wire _3541_;
 wire _3542_;
 wire _3543_;
 wire _3544_;
 wire _3545_;
 wire _3546_;
 wire _3547_;
 wire _3548_;
 wire _3549_;
 wire _3550_;
 wire _3551_;
 wire _3552_;
 wire _3553_;
 wire _3554_;
 wire _3555_;
 wire _3556_;
 wire _3557_;
 wire _3558_;
 wire _3559_;
 wire _3560_;
 wire _3561_;
 wire _3562_;
 wire _3563_;
 wire _3564_;
 wire _3565_;
 wire _3566_;
 wire _3567_;
 wire _3568_;
 wire _3569_;
 wire _3570_;
 wire _3571_;
 wire _3572_;
 wire _3573_;
 wire _3574_;
 wire _3575_;
 wire _3576_;
 wire _3577_;
 wire _3578_;
 wire _3579_;
 wire _3580_;
 wire _3581_;
 wire _3582_;
 wire _3583_;
 wire _3584_;
 wire _3585_;
 wire _3586_;
 wire _3587_;
 wire _3588_;
 wire _3589_;
 wire _3590_;
 wire _3591_;
 wire _3592_;
 wire _3593_;
 wire _3594_;
 wire _3595_;
 wire _3596_;
 wire _3597_;
 wire _3598_;
 wire _3599_;
 wire _3600_;
 wire _3601_;
 wire _3602_;
 wire _3603_;
 wire _3604_;
 wire _3605_;
 wire _3606_;
 wire _3607_;
 wire _3608_;
 wire _3609_;
 wire _3610_;
 wire _3611_;
 wire _3612_;
 wire _3613_;
 wire _3614_;
 wire _3615_;
 wire _3616_;
 wire _3617_;
 wire _3618_;
 wire _3619_;
 wire _3620_;
 wire _3621_;
 wire _3622_;
 wire _3623_;
 wire _3624_;
 wire _3625_;
 wire _3626_;
 wire _3627_;
 wire _3628_;
 wire _3629_;
 wire _3630_;
 wire _3631_;
 wire _3632_;
 wire _3633_;
 wire _3634_;
 wire _3635_;
 wire _3636_;
 wire _3637_;
 wire _3638_;
 wire _3639_;
 wire _3640_;
 wire _3641_;
 wire _3642_;
 wire _3643_;
 wire _3644_;
 wire _3645_;
 wire _3646_;
 wire _3647_;
 wire _3648_;
 wire _3649_;
 wire _3650_;
 wire _3651_;
 wire _3652_;
 wire _3653_;
 wire _3654_;
 wire _3655_;
 wire _3656_;
 wire _3657_;
 wire _3658_;
 wire _3659_;
 wire _3660_;
 wire _3661_;
 wire _3662_;
 wire _3663_;
 wire _3664_;
 wire _3665_;
 wire _3666_;
 wire _3667_;
 wire _3668_;
 wire _3669_;
 wire _3670_;
 wire _3671_;
 wire _3672_;
 wire _3673_;
 wire _3674_;
 wire _3675_;
 wire _3676_;
 wire _3677_;
 wire _3678_;
 wire _3679_;
 wire _3680_;
 wire _3681_;
 wire _3682_;
 wire _3683_;
 wire _3684_;
 wire _3685_;
 wire _3686_;
 wire _3687_;
 wire _3688_;
 wire _3689_;
 wire _3690_;
 wire _3691_;
 wire _3692_;
 wire _3693_;
 wire _3694_;
 wire _3695_;
 wire _3696_;
 wire _3697_;
 wire _3698_;
 wire _3699_;
 wire _3700_;
 wire _3701_;
 wire _3702_;
 wire _3703_;
 wire _3704_;
 wire _3705_;
 wire _3706_;
 wire _3707_;
 wire _3708_;
 wire _3709_;
 wire _3710_;
 wire _3711_;
 wire _3712_;
 wire _3713_;
 wire _3714_;
 wire _3715_;
 wire _3716_;
 wire _3717_;
 wire _3718_;
 wire _3719_;
 wire _3720_;
 wire _3721_;
 wire _3722_;
 wire _3723_;
 wire _3724_;
 wire _3725_;
 wire _3726_;
 wire _3727_;
 wire _3728_;
 wire _3729_;
 wire _3730_;
 wire _3731_;
 wire _3732_;
 wire _3733_;
 wire _3734_;
 wire _3735_;
 wire _3736_;
 wire _3737_;
 wire _3738_;
 wire _3739_;
 wire _3740_;
 wire _3741_;
 wire _3742_;
 wire _3743_;
 wire _3744_;
 wire _3745_;
 wire _3746_;
 wire _3747_;
 wire _3748_;
 wire _3749_;
 wire _3750_;
 wire _3751_;
 wire _3752_;
 wire _3753_;
 wire _3754_;
 wire _3755_;
 wire _3756_;
 wire _3757_;
 wire _3758_;
 wire _3759_;
 wire _3760_;
 wire _3761_;
 wire _3762_;
 wire _3763_;
 wire _3764_;
 wire _3765_;
 wire _3766_;
 wire _3767_;
 wire _3768_;
 wire _3769_;
 wire _3770_;
 wire _3771_;
 wire _3772_;
 wire _3773_;
 wire _3774_;
 wire _3775_;
 wire _3776_;
 wire _3777_;
 wire _3778_;
 wire _3779_;
 wire _3780_;
 wire _3781_;
 wire _3782_;
 wire _3783_;
 wire _3784_;
 wire _3785_;
 wire _3786_;
 wire _3787_;
 wire _3788_;
 wire _3789_;
 wire _3790_;
 wire _3791_;
 wire _3792_;
 wire _3793_;
 wire _3794_;
 wire _3795_;
 wire _3796_;
 wire _3797_;
 wire _3798_;
 wire _3799_;
 wire _3800_;
 wire _3801_;
 wire _3802_;
 wire _3803_;
 wire _3804_;
 wire _3805_;
 wire _3806_;
 wire _3807_;
 wire _3808_;
 wire _3809_;
 wire _3810_;
 wire _3811_;
 wire _3812_;
 wire _3813_;
 wire _3814_;
 wire _3815_;
 wire _3816_;
 wire _3817_;
 wire _3818_;
 wire _3819_;
 wire _3820_;
 wire _3821_;
 wire _3822_;
 wire _3823_;
 wire _3824_;
 wire _3825_;
 wire _3826_;
 wire _3827_;
 wire _3828_;
 wire _3829_;
 wire _3830_;
 wire _3831_;
 wire _3832_;
 wire _3833_;
 wire _3834_;
 wire _3835_;
 wire _3836_;
 wire _3837_;
 wire _3838_;
 wire _3839_;
 wire _3840_;
 wire _3841_;
 wire _3842_;
 wire _3843_;
 wire _3844_;
 wire _3845_;
 wire _3846_;
 wire _3847_;
 wire _3848_;
 wire _3849_;
 wire _3850_;
 wire _3851_;
 wire _3852_;
 wire _3853_;
 wire _3854_;
 wire _3855_;
 wire _3856_;
 wire _3857_;
 wire _3858_;
 wire _3859_;
 wire _3860_;
 wire _3861_;
 wire _3862_;
 wire _3863_;
 wire _3864_;
 wire _3865_;
 wire _3866_;
 wire _3867_;
 wire _3868_;
 wire _3869_;
 wire _3870_;
 wire _3871_;
 wire _3872_;
 wire _3873_;
 wire _3874_;
 wire _3875_;
 wire _3876_;
 wire _3877_;
 wire _3878_;
 wire _3879_;
 wire _3880_;
 wire _3881_;
 wire _3882_;
 wire _3883_;
 wire _3884_;
 wire _3885_;
 wire _3886_;
 wire _3887_;
 wire _3888_;
 wire _3889_;
 wire _3890_;
 wire _3891_;
 wire _3892_;
 wire _3893_;
 wire _3894_;
 wire _3895_;
 wire _3896_;
 wire _3897_;
 wire _3898_;
 wire _3899_;
 wire _3900_;
 wire _3901_;
 wire _3902_;
 wire _3903_;
 wire _3904_;
 wire _3905_;
 wire _3906_;
 wire _3907_;
 wire _3908_;
 wire _3909_;
 wire _3910_;
 wire _3911_;
 wire _3912_;
 wire _3913_;
 wire _3914_;
 wire _3915_;
 wire _3916_;
 wire _3917_;
 wire _3918_;
 wire _3919_;
 wire _3920_;
 wire _3921_;
 wire _3922_;
 wire _3923_;
 wire _3924_;
 wire _3925_;
 wire _3926_;
 wire _3927_;
 wire _3928_;
 wire _3929_;
 wire _3930_;
 wire _3931_;
 wire _3932_;
 wire _3933_;
 wire _3934_;
 wire _3935_;
 wire _3936_;
 wire _3937_;
 wire _3938_;
 wire _3939_;
 wire _3940_;
 wire _3941_;
 wire _3942_;
 wire _3943_;
 wire _3944_;
 wire _3945_;
 wire _3946_;
 wire _3947_;
 wire _3948_;
 wire _3949_;
 wire _3950_;
 wire _3951_;
 wire _3952_;
 wire _3953_;
 wire _3954_;
 wire _3955_;
 wire _3956_;
 wire _3957_;
 wire _3958_;
 wire _3959_;
 wire _3960_;
 wire _3961_;
 wire _3962_;
 wire _3963_;
 wire _3964_;
 wire _3965_;
 wire _3966_;
 wire _3967_;
 wire _3968_;
 wire _3969_;
 wire _3970_;
 wire _3971_;
 wire _3972_;
 wire _3973_;
 wire _3974_;
 wire _3975_;
 wire _3976_;
 wire _3977_;
 wire _3978_;
 wire _3979_;
 wire _3980_;
 wire _3981_;
 wire _3982_;
 wire _3983_;
 wire _3984_;
 wire _3985_;
 wire _3986_;
 wire _3987_;
 wire _3988_;
 wire _3989_;
 wire _3990_;
 wire _3991_;
 wire _3992_;
 wire _3993_;
 wire _3994_;
 wire _3995_;
 wire _3996_;
 wire _3997_;
 wire _3998_;
 wire _3999_;
 wire _4000_;
 wire _4001_;
 wire _4002_;
 wire _4003_;
 wire _4004_;
 wire _4005_;
 wire _4006_;
 wire _4007_;
 wire _4008_;
 wire _4009_;
 wire _4010_;
 wire _4011_;
 wire _4012_;
 wire _4013_;
 wire _4014_;
 wire _4015_;
 wire _4016_;
 wire _4017_;
 wire _4018_;
 wire _4019_;
 wire _4020_;
 wire _4021_;
 wire _4022_;
 wire _4023_;
 wire _4024_;
 wire _4025_;
 wire _4026_;
 wire _4027_;
 wire _4028_;
 wire _4029_;
 wire _4030_;
 wire _4031_;
 wire _4032_;
 wire _4033_;
 wire _4034_;
 wire _4035_;
 wire _4036_;
 wire _4037_;
 wire _4038_;
 wire _4039_;
 wire _4040_;
 wire _4041_;
 wire _4042_;
 wire _4043_;
 wire _4044_;
 wire _4045_;
 wire _4046_;
 wire _4047_;
 wire _4048_;
 wire _4049_;
 wire _4050_;
 wire _4051_;
 wire _4052_;
 wire _4053_;
 wire _4054_;
 wire _4055_;
 wire _4056_;
 wire _4057_;
 wire _4058_;
 wire _4059_;
 wire _4060_;
 wire _4061_;
 wire _4062_;
 wire _4063_;
 wire _4064_;
 wire _4065_;
 wire _4066_;
 wire _4067_;
 wire _4068_;
 wire _4069_;
 wire _4070_;
 wire _4071_;
 wire _4072_;
 wire _4073_;
 wire _4074_;
 wire _4075_;
 wire _4076_;
 wire _4077_;
 wire _4078_;
 wire _4079_;
 wire _4080_;
 wire _4081_;
 wire _4082_;
 wire _4083_;
 wire _4084_;
 wire _4085_;
 wire _4086_;
 wire _4087_;
 wire _4088_;
 wire _4089_;
 wire _4090_;
 wire _4091_;
 wire _4092_;
 wire _4093_;
 wire _4094_;
 wire _4095_;
 wire _4096_;
 wire _4097_;
 wire _4098_;
 wire _4099_;
 wire _4100_;
 wire _4101_;
 wire _4102_;
 wire _4103_;
 wire _4104_;
 wire _4105_;
 wire _4106_;
 wire _4107_;
 wire _4108_;
 wire _4109_;
 wire _4110_;
 wire _4111_;
 wire _4112_;
 wire _4113_;
 wire _4114_;
 wire _4115_;
 wire _4116_;
 wire _4117_;
 wire _4118_;
 wire _4119_;
 wire _4120_;
 wire _4121_;
 wire _4122_;
 wire _4123_;
 wire _4124_;
 wire _4125_;
 wire _4126_;
 wire _4127_;
 wire _4128_;
 wire _4129_;
 wire _4130_;
 wire _4131_;
 wire _4132_;
 wire _4133_;
 wire _4134_;
 wire _4135_;
 wire _4136_;
 wire _4137_;
 wire _4138_;
 wire _4139_;
 wire _4140_;
 wire _4141_;
 wire _4142_;
 wire _4143_;
 wire _4144_;
 wire _4145_;
 wire _4146_;
 wire _4147_;
 wire _4148_;
 wire _4149_;
 wire _4150_;
 wire _4151_;
 wire _4152_;
 wire _4153_;
 wire _4154_;
 wire _4155_;
 wire _4156_;
 wire _4157_;
 wire _4158_;
 wire _4159_;
 wire _4160_;
 wire _4161_;
 wire _4162_;
 wire _4163_;
 wire _4164_;
 wire _4165_;
 wire _4166_;
 wire _4167_;
 wire _4168_;
 wire _4169_;
 wire _4170_;
 wire _4171_;
 wire _4172_;
 wire _4173_;
 wire _4174_;
 wire _4175_;
 wire _4176_;
 wire _4177_;
 wire _4178_;
 wire _4179_;
 wire _4180_;
 wire _4181_;
 wire _4182_;
 wire _4183_;
 wire _4184_;
 wire _4185_;
 wire _4186_;
 wire _4187_;
 wire _4188_;
 wire _4189_;
 wire _4190_;
 wire _4191_;
 wire _4192_;
 wire _4193_;
 wire _4194_;
 wire _4195_;
 wire _4196_;
 wire _4197_;
 wire _4198_;
 wire _4199_;
 wire _4200_;
 wire _4201_;
 wire _4202_;
 wire _4203_;
 wire _4204_;
 wire _4205_;
 wire _4206_;
 wire _4207_;
 wire _4208_;
 wire _4209_;
 wire _4210_;
 wire _4211_;
 wire _4212_;
 wire _4213_;
 wire _4214_;
 wire _4215_;
 wire _4216_;
 wire _4217_;
 wire _4218_;
 wire _4219_;
 wire _4220_;
 wire _4221_;
 wire _4222_;
 wire _4223_;
 wire _4224_;
 wire _4225_;
 wire _4226_;
 wire _4227_;
 wire _4228_;
 wire _4229_;
 wire _4230_;
 wire _4231_;
 wire _4232_;
 wire _4233_;
 wire _4234_;
 wire _4235_;
 wire _4236_;
 wire _4237_;
 wire _4238_;
 wire _4239_;
 wire _4240_;
 wire _4241_;
 wire _4242_;
 wire _4243_;
 wire _4244_;
 wire _4245_;
 wire _4246_;
 wire _4247_;
 wire _4248_;
 wire _4249_;
 wire _4250_;
 wire _4251_;
 wire _4252_;
 wire _4253_;
 wire _4254_;
 wire _4255_;
 wire _4256_;
 wire _4257_;
 wire _4258_;
 wire _4259_;
 wire _4260_;
 wire _4261_;
 wire _4262_;
 wire _4263_;
 wire _4264_;
 wire _4265_;
 wire _4266_;
 wire _4267_;
 wire _4268_;
 wire _4269_;
 wire _4270_;
 wire _4271_;
 wire _4272_;
 wire _4273_;
 wire _4274_;
 wire _4275_;
 wire _4276_;
 wire _4277_;
 wire _4278_;
 wire _4279_;
 wire _4280_;
 wire _4281_;
 wire _4282_;
 wire _4283_;
 wire _4284_;
 wire _4285_;
 wire _4286_;
 wire _4287_;
 wire _4288_;
 wire _4289_;
 wire _4290_;
 wire _4291_;
 wire _4292_;
 wire _4293_;
 wire _4294_;
 wire _4295_;
 wire _4296_;
 wire _4297_;
 wire _4298_;
 wire _4299_;
 wire _4300_;
 wire _4301_;
 wire _4302_;
 wire _4303_;
 wire _4304_;
 wire _4305_;
 wire _4306_;
 wire _4307_;
 wire _4308_;
 wire _4309_;
 wire _4310_;
 wire _4311_;
 wire _4312_;
 wire _4313_;
 wire _4314_;
 wire _4315_;
 wire _4316_;
 wire _4317_;
 wire _4318_;
 wire _4319_;
 wire _4320_;
 wire _4321_;
 wire _4322_;
 wire _4323_;
 wire _4324_;
 wire _4325_;
 wire _4326_;
 wire _4327_;
 wire _4328_;
 wire _4329_;
 wire _4330_;
 wire _4331_;
 wire _4332_;
 wire _4333_;
 wire _4334_;
 wire _4335_;
 wire _4336_;
 wire _4337_;
 wire _4338_;
 wire _4339_;
 wire _4340_;
 wire _4341_;
 wire _4342_;
 wire _4343_;
 wire _4344_;
 wire _4345_;
 wire _4346_;
 wire _4347_;
 wire net505;
 wire clk1_output_dest;
 wire clk2_output_dest;
 wire csclk;
 wire \gpio_configure[0][0] ;
 wire \gpio_configure[0][10] ;
 wire \gpio_configure[0][11] ;
 wire \gpio_configure[0][12] ;
 wire \gpio_configure[0][1] ;
 wire \gpio_configure[0][2] ;
 wire \gpio_configure[0][3] ;
 wire \gpio_configure[0][4] ;
 wire \gpio_configure[0][5] ;
 wire \gpio_configure[0][6] ;
 wire \gpio_configure[0][7] ;
 wire \gpio_configure[0][8] ;
 wire \gpio_configure[0][9] ;
 wire \gpio_configure[10][0] ;
 wire \gpio_configure[10][10] ;
 wire \gpio_configure[10][11] ;
 wire \gpio_configure[10][12] ;
 wire \gpio_configure[10][1] ;
 wire \gpio_configure[10][2] ;
 wire \gpio_configure[10][3] ;
 wire \gpio_configure[10][4] ;
 wire \gpio_configure[10][5] ;
 wire \gpio_configure[10][6] ;
 wire \gpio_configure[10][7] ;
 wire \gpio_configure[10][8] ;
 wire \gpio_configure[10][9] ;
 wire \gpio_configure[11][0] ;
 wire \gpio_configure[11][10] ;
 wire \gpio_configure[11][11] ;
 wire \gpio_configure[11][12] ;
 wire \gpio_configure[11][1] ;
 wire \gpio_configure[11][2] ;
 wire \gpio_configure[11][3] ;
 wire \gpio_configure[11][4] ;
 wire \gpio_configure[11][5] ;
 wire \gpio_configure[11][6] ;
 wire \gpio_configure[11][7] ;
 wire \gpio_configure[11][8] ;
 wire \gpio_configure[11][9] ;
 wire \gpio_configure[12][0] ;
 wire \gpio_configure[12][10] ;
 wire \gpio_configure[12][11] ;
 wire \gpio_configure[12][12] ;
 wire \gpio_configure[12][1] ;
 wire \gpio_configure[12][2] ;
 wire \gpio_configure[12][3] ;
 wire \gpio_configure[12][4] ;
 wire \gpio_configure[12][5] ;
 wire \gpio_configure[12][6] ;
 wire \gpio_configure[12][7] ;
 wire \gpio_configure[12][8] ;
 wire \gpio_configure[12][9] ;
 wire \gpio_configure[13][0] ;
 wire \gpio_configure[13][10] ;
 wire \gpio_configure[13][11] ;
 wire \gpio_configure[13][12] ;
 wire \gpio_configure[13][1] ;
 wire \gpio_configure[13][2] ;
 wire \gpio_configure[13][3] ;
 wire \gpio_configure[13][4] ;
 wire \gpio_configure[13][5] ;
 wire \gpio_configure[13][6] ;
 wire \gpio_configure[13][7] ;
 wire \gpio_configure[13][8] ;
 wire \gpio_configure[13][9] ;
 wire \gpio_configure[14][0] ;
 wire \gpio_configure[14][10] ;
 wire \gpio_configure[14][11] ;
 wire \gpio_configure[14][12] ;
 wire \gpio_configure[14][1] ;
 wire \gpio_configure[14][2] ;
 wire \gpio_configure[14][3] ;
 wire \gpio_configure[14][4] ;
 wire \gpio_configure[14][5] ;
 wire \gpio_configure[14][6] ;
 wire \gpio_configure[14][7] ;
 wire \gpio_configure[14][8] ;
 wire \gpio_configure[14][9] ;
 wire \gpio_configure[15][0] ;
 wire \gpio_configure[15][10] ;
 wire \gpio_configure[15][11] ;
 wire \gpio_configure[15][12] ;
 wire \gpio_configure[15][1] ;
 wire \gpio_configure[15][2] ;
 wire \gpio_configure[15][3] ;
 wire \gpio_configure[15][4] ;
 wire \gpio_configure[15][5] ;
 wire \gpio_configure[15][6] ;
 wire \gpio_configure[15][7] ;
 wire \gpio_configure[15][8] ;
 wire \gpio_configure[15][9] ;
 wire \gpio_configure[16][0] ;
 wire \gpio_configure[16][10] ;
 wire \gpio_configure[16][11] ;
 wire \gpio_configure[16][12] ;
 wire \gpio_configure[16][1] ;
 wire \gpio_configure[16][2] ;
 wire \gpio_configure[16][3] ;
 wire \gpio_configure[16][4] ;
 wire \gpio_configure[16][5] ;
 wire \gpio_configure[16][6] ;
 wire \gpio_configure[16][7] ;
 wire \gpio_configure[16][8] ;
 wire \gpio_configure[16][9] ;
 wire \gpio_configure[17][0] ;
 wire \gpio_configure[17][10] ;
 wire \gpio_configure[17][11] ;
 wire \gpio_configure[17][12] ;
 wire \gpio_configure[17][1] ;
 wire \gpio_configure[17][2] ;
 wire \gpio_configure[17][3] ;
 wire \gpio_configure[17][4] ;
 wire \gpio_configure[17][5] ;
 wire \gpio_configure[17][6] ;
 wire \gpio_configure[17][7] ;
 wire \gpio_configure[17][8] ;
 wire \gpio_configure[17][9] ;
 wire \gpio_configure[18][0] ;
 wire \gpio_configure[18][10] ;
 wire \gpio_configure[18][11] ;
 wire \gpio_configure[18][12] ;
 wire \gpio_configure[18][1] ;
 wire \gpio_configure[18][2] ;
 wire \gpio_configure[18][3] ;
 wire \gpio_configure[18][4] ;
 wire \gpio_configure[18][5] ;
 wire \gpio_configure[18][6] ;
 wire \gpio_configure[18][7] ;
 wire \gpio_configure[18][8] ;
 wire \gpio_configure[18][9] ;
 wire \gpio_configure[19][0] ;
 wire \gpio_configure[19][10] ;
 wire \gpio_configure[19][11] ;
 wire \gpio_configure[19][12] ;
 wire \gpio_configure[19][1] ;
 wire \gpio_configure[19][2] ;
 wire \gpio_configure[19][3] ;
 wire \gpio_configure[19][4] ;
 wire \gpio_configure[19][5] ;
 wire \gpio_configure[19][6] ;
 wire \gpio_configure[19][7] ;
 wire \gpio_configure[19][8] ;
 wire \gpio_configure[19][9] ;
 wire \gpio_configure[1][0] ;
 wire \gpio_configure[1][10] ;
 wire \gpio_configure[1][11] ;
 wire \gpio_configure[1][12] ;
 wire \gpio_configure[1][1] ;
 wire \gpio_configure[1][2] ;
 wire \gpio_configure[1][3] ;
 wire \gpio_configure[1][4] ;
 wire \gpio_configure[1][5] ;
 wire \gpio_configure[1][6] ;
 wire \gpio_configure[1][7] ;
 wire \gpio_configure[1][8] ;
 wire \gpio_configure[1][9] ;
 wire \gpio_configure[20][0] ;
 wire \gpio_configure[20][10] ;
 wire \gpio_configure[20][11] ;
 wire \gpio_configure[20][12] ;
 wire \gpio_configure[20][1] ;
 wire \gpio_configure[20][2] ;
 wire \gpio_configure[20][3] ;
 wire \gpio_configure[20][4] ;
 wire \gpio_configure[20][5] ;
 wire \gpio_configure[20][6] ;
 wire \gpio_configure[20][7] ;
 wire \gpio_configure[20][8] ;
 wire \gpio_configure[20][9] ;
 wire \gpio_configure[21][0] ;
 wire \gpio_configure[21][10] ;
 wire \gpio_configure[21][11] ;
 wire \gpio_configure[21][12] ;
 wire \gpio_configure[21][1] ;
 wire \gpio_configure[21][2] ;
 wire \gpio_configure[21][3] ;
 wire \gpio_configure[21][4] ;
 wire \gpio_configure[21][5] ;
 wire \gpio_configure[21][6] ;
 wire \gpio_configure[21][7] ;
 wire \gpio_configure[21][8] ;
 wire \gpio_configure[21][9] ;
 wire \gpio_configure[22][0] ;
 wire \gpio_configure[22][10] ;
 wire \gpio_configure[22][11] ;
 wire \gpio_configure[22][12] ;
 wire \gpio_configure[22][1] ;
 wire \gpio_configure[22][2] ;
 wire \gpio_configure[22][3] ;
 wire \gpio_configure[22][4] ;
 wire \gpio_configure[22][5] ;
 wire \gpio_configure[22][6] ;
 wire \gpio_configure[22][7] ;
 wire \gpio_configure[22][8] ;
 wire \gpio_configure[22][9] ;
 wire \gpio_configure[23][0] ;
 wire \gpio_configure[23][10] ;
 wire \gpio_configure[23][11] ;
 wire \gpio_configure[23][12] ;
 wire \gpio_configure[23][1] ;
 wire \gpio_configure[23][2] ;
 wire \gpio_configure[23][3] ;
 wire \gpio_configure[23][4] ;
 wire \gpio_configure[23][5] ;
 wire \gpio_configure[23][6] ;
 wire \gpio_configure[23][7] ;
 wire \gpio_configure[23][8] ;
 wire \gpio_configure[23][9] ;
 wire \gpio_configure[24][0] ;
 wire \gpio_configure[24][10] ;
 wire \gpio_configure[24][11] ;
 wire \gpio_configure[24][12] ;
 wire \gpio_configure[24][1] ;
 wire \gpio_configure[24][2] ;
 wire \gpio_configure[24][3] ;
 wire \gpio_configure[24][4] ;
 wire \gpio_configure[24][5] ;
 wire \gpio_configure[24][6] ;
 wire \gpio_configure[24][7] ;
 wire \gpio_configure[24][8] ;
 wire \gpio_configure[24][9] ;
 wire \gpio_configure[25][0] ;
 wire \gpio_configure[25][10] ;
 wire \gpio_configure[25][11] ;
 wire \gpio_configure[25][12] ;
 wire \gpio_configure[25][1] ;
 wire \gpio_configure[25][2] ;
 wire \gpio_configure[25][3] ;
 wire \gpio_configure[25][4] ;
 wire \gpio_configure[25][5] ;
 wire \gpio_configure[25][6] ;
 wire \gpio_configure[25][7] ;
 wire \gpio_configure[25][8] ;
 wire \gpio_configure[25][9] ;
 wire \gpio_configure[26][0] ;
 wire \gpio_configure[26][10] ;
 wire \gpio_configure[26][11] ;
 wire \gpio_configure[26][12] ;
 wire \gpio_configure[26][1] ;
 wire \gpio_configure[26][2] ;
 wire \gpio_configure[26][3] ;
 wire \gpio_configure[26][4] ;
 wire \gpio_configure[26][5] ;
 wire \gpio_configure[26][6] ;
 wire \gpio_configure[26][7] ;
 wire \gpio_configure[26][8] ;
 wire \gpio_configure[26][9] ;
 wire \gpio_configure[27][0] ;
 wire \gpio_configure[27][10] ;
 wire \gpio_configure[27][11] ;
 wire \gpio_configure[27][12] ;
 wire \gpio_configure[27][1] ;
 wire \gpio_configure[27][2] ;
 wire \gpio_configure[27][3] ;
 wire \gpio_configure[27][4] ;
 wire \gpio_configure[27][5] ;
 wire \gpio_configure[27][6] ;
 wire \gpio_configure[27][7] ;
 wire \gpio_configure[27][8] ;
 wire \gpio_configure[27][9] ;
 wire \gpio_configure[28][0] ;
 wire \gpio_configure[28][10] ;
 wire \gpio_configure[28][11] ;
 wire \gpio_configure[28][12] ;
 wire \gpio_configure[28][1] ;
 wire \gpio_configure[28][2] ;
 wire \gpio_configure[28][3] ;
 wire \gpio_configure[28][4] ;
 wire \gpio_configure[28][5] ;
 wire \gpio_configure[28][6] ;
 wire \gpio_configure[28][7] ;
 wire \gpio_configure[28][8] ;
 wire \gpio_configure[28][9] ;
 wire \gpio_configure[29][0] ;
 wire \gpio_configure[29][10] ;
 wire \gpio_configure[29][11] ;
 wire \gpio_configure[29][12] ;
 wire \gpio_configure[29][1] ;
 wire \gpio_configure[29][2] ;
 wire \gpio_configure[29][3] ;
 wire \gpio_configure[29][4] ;
 wire \gpio_configure[29][5] ;
 wire \gpio_configure[29][6] ;
 wire \gpio_configure[29][7] ;
 wire \gpio_configure[29][8] ;
 wire \gpio_configure[29][9] ;
 wire \gpio_configure[2][0] ;
 wire \gpio_configure[2][10] ;
 wire \gpio_configure[2][11] ;
 wire \gpio_configure[2][12] ;
 wire \gpio_configure[2][1] ;
 wire \gpio_configure[2][2] ;
 wire \gpio_configure[2][3] ;
 wire \gpio_configure[2][4] ;
 wire \gpio_configure[2][5] ;
 wire \gpio_configure[2][6] ;
 wire \gpio_configure[2][7] ;
 wire \gpio_configure[2][8] ;
 wire \gpio_configure[2][9] ;
 wire \gpio_configure[30][0] ;
 wire \gpio_configure[30][10] ;
 wire \gpio_configure[30][11] ;
 wire \gpio_configure[30][12] ;
 wire \gpio_configure[30][1] ;
 wire \gpio_configure[30][2] ;
 wire \gpio_configure[30][3] ;
 wire \gpio_configure[30][4] ;
 wire \gpio_configure[30][5] ;
 wire \gpio_configure[30][6] ;
 wire \gpio_configure[30][7] ;
 wire \gpio_configure[30][8] ;
 wire \gpio_configure[30][9] ;
 wire \gpio_configure[31][0] ;
 wire \gpio_configure[31][10] ;
 wire \gpio_configure[31][11] ;
 wire \gpio_configure[31][12] ;
 wire \gpio_configure[31][1] ;
 wire \gpio_configure[31][2] ;
 wire \gpio_configure[31][3] ;
 wire \gpio_configure[31][4] ;
 wire \gpio_configure[31][5] ;
 wire \gpio_configure[31][6] ;
 wire \gpio_configure[31][7] ;
 wire \gpio_configure[31][8] ;
 wire \gpio_configure[31][9] ;
 wire \gpio_configure[32][0] ;
 wire \gpio_configure[32][10] ;
 wire \gpio_configure[32][11] ;
 wire \gpio_configure[32][12] ;
 wire \gpio_configure[32][1] ;
 wire \gpio_configure[32][2] ;
 wire \gpio_configure[32][3] ;
 wire \gpio_configure[32][4] ;
 wire \gpio_configure[32][5] ;
 wire \gpio_configure[32][6] ;
 wire \gpio_configure[32][7] ;
 wire \gpio_configure[32][8] ;
 wire \gpio_configure[32][9] ;
 wire \gpio_configure[33][0] ;
 wire \gpio_configure[33][10] ;
 wire \gpio_configure[33][11] ;
 wire \gpio_configure[33][12] ;
 wire \gpio_configure[33][1] ;
 wire \gpio_configure[33][2] ;
 wire \gpio_configure[33][3] ;
 wire \gpio_configure[33][4] ;
 wire \gpio_configure[33][5] ;
 wire \gpio_configure[33][6] ;
 wire \gpio_configure[33][7] ;
 wire \gpio_configure[33][8] ;
 wire \gpio_configure[33][9] ;
 wire \gpio_configure[34][0] ;
 wire \gpio_configure[34][10] ;
 wire \gpio_configure[34][11] ;
 wire \gpio_configure[34][12] ;
 wire \gpio_configure[34][1] ;
 wire \gpio_configure[34][2] ;
 wire \gpio_configure[34][3] ;
 wire \gpio_configure[34][4] ;
 wire \gpio_configure[34][5] ;
 wire \gpio_configure[34][6] ;
 wire \gpio_configure[34][7] ;
 wire \gpio_configure[34][8] ;
 wire \gpio_configure[34][9] ;
 wire \gpio_configure[35][0] ;
 wire \gpio_configure[35][10] ;
 wire \gpio_configure[35][11] ;
 wire \gpio_configure[35][12] ;
 wire \gpio_configure[35][1] ;
 wire \gpio_configure[35][2] ;
 wire \gpio_configure[35][3] ;
 wire \gpio_configure[35][4] ;
 wire \gpio_configure[35][5] ;
 wire \gpio_configure[35][6] ;
 wire \gpio_configure[35][7] ;
 wire \gpio_configure[35][8] ;
 wire \gpio_configure[35][9] ;
 wire \gpio_configure[36][0] ;
 wire \gpio_configure[36][10] ;
 wire \gpio_configure[36][11] ;
 wire \gpio_configure[36][12] ;
 wire \gpio_configure[36][1] ;
 wire \gpio_configure[36][2] ;
 wire \gpio_configure[36][3] ;
 wire \gpio_configure[36][4] ;
 wire \gpio_configure[36][5] ;
 wire \gpio_configure[36][6] ;
 wire \gpio_configure[36][7] ;
 wire \gpio_configure[36][8] ;
 wire \gpio_configure[36][9] ;
 wire \gpio_configure[37][0] ;
 wire \gpio_configure[37][10] ;
 wire \gpio_configure[37][11] ;
 wire \gpio_configure[37][12] ;
 wire \gpio_configure[37][1] ;
 wire \gpio_configure[37][2] ;
 wire \gpio_configure[37][3] ;
 wire \gpio_configure[37][4] ;
 wire \gpio_configure[37][5] ;
 wire \gpio_configure[37][6] ;
 wire \gpio_configure[37][7] ;
 wire \gpio_configure[37][8] ;
 wire \gpio_configure[37][9] ;
 wire \gpio_configure[3][0] ;
 wire \gpio_configure[3][10] ;
 wire \gpio_configure[3][11] ;
 wire \gpio_configure[3][12] ;
 wire \gpio_configure[3][1] ;
 wire \gpio_configure[3][2] ;
 wire \gpio_configure[3][3] ;
 wire \gpio_configure[3][4] ;
 wire \gpio_configure[3][5] ;
 wire \gpio_configure[3][6] ;
 wire \gpio_configure[3][7] ;
 wire \gpio_configure[3][8] ;
 wire \gpio_configure[3][9] ;
 wire \gpio_configure[4][0] ;
 wire \gpio_configure[4][10] ;
 wire \gpio_configure[4][11] ;
 wire \gpio_configure[4][12] ;
 wire \gpio_configure[4][1] ;
 wire \gpio_configure[4][2] ;
 wire \gpio_configure[4][3] ;
 wire \gpio_configure[4][4] ;
 wire \gpio_configure[4][5] ;
 wire \gpio_configure[4][6] ;
 wire \gpio_configure[4][7] ;
 wire \gpio_configure[4][8] ;
 wire \gpio_configure[4][9] ;
 wire \gpio_configure[5][0] ;
 wire \gpio_configure[5][10] ;
 wire \gpio_configure[5][11] ;
 wire \gpio_configure[5][12] ;
 wire \gpio_configure[5][1] ;
 wire \gpio_configure[5][2] ;
 wire \gpio_configure[5][3] ;
 wire \gpio_configure[5][4] ;
 wire \gpio_configure[5][5] ;
 wire \gpio_configure[5][6] ;
 wire \gpio_configure[5][7] ;
 wire \gpio_configure[5][8] ;
 wire \gpio_configure[5][9] ;
 wire \gpio_configure[6][0] ;
 wire \gpio_configure[6][10] ;
 wire \gpio_configure[6][11] ;
 wire \gpio_configure[6][12] ;
 wire \gpio_configure[6][1] ;
 wire \gpio_configure[6][2] ;
 wire \gpio_configure[6][3] ;
 wire \gpio_configure[6][4] ;
 wire \gpio_configure[6][5] ;
 wire \gpio_configure[6][6] ;
 wire \gpio_configure[6][7] ;
 wire \gpio_configure[6][8] ;
 wire \gpio_configure[6][9] ;
 wire \gpio_configure[7][0] ;
 wire \gpio_configure[7][10] ;
 wire \gpio_configure[7][11] ;
 wire \gpio_configure[7][12] ;
 wire \gpio_configure[7][1] ;
 wire \gpio_configure[7][2] ;
 wire \gpio_configure[7][3] ;
 wire \gpio_configure[7][4] ;
 wire \gpio_configure[7][5] ;
 wire \gpio_configure[7][6] ;
 wire \gpio_configure[7][7] ;
 wire \gpio_configure[7][8] ;
 wire \gpio_configure[7][9] ;
 wire \gpio_configure[8][0] ;
 wire \gpio_configure[8][10] ;
 wire \gpio_configure[8][11] ;
 wire \gpio_configure[8][12] ;
 wire \gpio_configure[8][1] ;
 wire \gpio_configure[8][2] ;
 wire \gpio_configure[8][3] ;
 wire \gpio_configure[8][4] ;
 wire \gpio_configure[8][5] ;
 wire \gpio_configure[8][6] ;
 wire \gpio_configure[8][7] ;
 wire \gpio_configure[8][8] ;
 wire \gpio_configure[8][9] ;
 wire \gpio_configure[9][0] ;
 wire \gpio_configure[9][10] ;
 wire \gpio_configure[9][11] ;
 wire \gpio_configure[9][12] ;
 wire \gpio_configure[9][1] ;
 wire \gpio_configure[9][2] ;
 wire \gpio_configure[9][3] ;
 wire \gpio_configure[9][4] ;
 wire \gpio_configure[9][5] ;
 wire \gpio_configure[9][6] ;
 wire \gpio_configure[9][7] ;
 wire \gpio_configure[9][8] ;
 wire \gpio_configure[9][9] ;
 wire \hkspi.SDO ;
 wire \hkspi.addr[0] ;
 wire \hkspi.addr[1] ;
 wire \hkspi.addr[2] ;
 wire \hkspi.addr[3] ;
 wire \hkspi.addr[4] ;
 wire \hkspi.addr[5] ;
 wire \hkspi.addr[6] ;
 wire \hkspi.addr[7] ;
 wire \hkspi.count[0] ;
 wire \hkspi.count[1] ;
 wire \hkspi.count[2] ;
 wire \hkspi.fixed[0] ;
 wire \hkspi.fixed[1] ;
 wire \hkspi.fixed[2] ;
 wire \hkspi.ldata[0] ;
 wire \hkspi.ldata[1] ;
 wire \hkspi.ldata[2] ;
 wire \hkspi.ldata[3] ;
 wire \hkspi.ldata[4] ;
 wire \hkspi.ldata[5] ;
 wire \hkspi.ldata[6] ;
 wire \hkspi.odata[1] ;
 wire \hkspi.odata[2] ;
 wire \hkspi.odata[3] ;
 wire \hkspi.odata[4] ;
 wire \hkspi.odata[5] ;
 wire \hkspi.odata[6] ;
 wire \hkspi.odata[7] ;
 wire \hkspi.pass_thru_mgmt ;
 wire \hkspi.pass_thru_mgmt_delay ;
 wire \hkspi.pass_thru_user ;
 wire \hkspi.pass_thru_user_delay ;
 wire \hkspi.pre_pass_thru_mgmt ;
 wire \hkspi.pre_pass_thru_user ;
 wire \hkspi.rdstb ;
 wire \hkspi.readmode ;
 wire \hkspi.sdoenb ;
 wire \hkspi.state[0] ;
 wire \hkspi.state[1] ;
 wire \hkspi.state[2] ;
 wire \hkspi.state[3] ;
 wire \hkspi.state[4] ;
 wire \hkspi.writemode ;
 wire \hkspi.wrstb ;
 wire hkspi_disable;
 wire irq_1_inputsrc;
 wire irq_2_inputsrc;
 wire \mgmt_gpio_data[0] ;
 wire \mgmt_gpio_data[10] ;
 wire \mgmt_gpio_data[11] ;
 wire \mgmt_gpio_data[12] ;
 wire \mgmt_gpio_data[13] ;
 wire \mgmt_gpio_data[14] ;
 wire \mgmt_gpio_data[15] ;
 wire \mgmt_gpio_data[16] ;
 wire \mgmt_gpio_data[17] ;
 wire \mgmt_gpio_data[18] ;
 wire \mgmt_gpio_data[19] ;
 wire \mgmt_gpio_data[1] ;
 wire \mgmt_gpio_data[20] ;
 wire \mgmt_gpio_data[21] ;
 wire \mgmt_gpio_data[22] ;
 wire \mgmt_gpio_data[23] ;
 wire \mgmt_gpio_data[24] ;
 wire \mgmt_gpio_data[25] ;
 wire \mgmt_gpio_data[26] ;
 wire \mgmt_gpio_data[27] ;
 wire \mgmt_gpio_data[28] ;
 wire \mgmt_gpio_data[29] ;
 wire \mgmt_gpio_data[2] ;
 wire \mgmt_gpio_data[30] ;
 wire \mgmt_gpio_data[31] ;
 wire \mgmt_gpio_data[32] ;
 wire \mgmt_gpio_data[33] ;
 wire \mgmt_gpio_data[34] ;
 wire \mgmt_gpio_data[35] ;
 wire \mgmt_gpio_data[36] ;
 wire \mgmt_gpio_data[37] ;
 wire \mgmt_gpio_data[3] ;
 wire \mgmt_gpio_data[4] ;
 wire \mgmt_gpio_data[5] ;
 wire \mgmt_gpio_data[6] ;
 wire \mgmt_gpio_data[7] ;
 wire \mgmt_gpio_data[8] ;
 wire \mgmt_gpio_data[9] ;
 wire \mgmt_gpio_data_buf[0] ;
 wire \mgmt_gpio_data_buf[10] ;
 wire \mgmt_gpio_data_buf[11] ;
 wire \mgmt_gpio_data_buf[12] ;
 wire \mgmt_gpio_data_buf[13] ;
 wire \mgmt_gpio_data_buf[14] ;
 wire \mgmt_gpio_data_buf[15] ;
 wire \mgmt_gpio_data_buf[16] ;
 wire \mgmt_gpio_data_buf[17] ;
 wire \mgmt_gpio_data_buf[18] ;
 wire \mgmt_gpio_data_buf[19] ;
 wire \mgmt_gpio_data_buf[1] ;
 wire \mgmt_gpio_data_buf[20] ;
 wire \mgmt_gpio_data_buf[21] ;
 wire \mgmt_gpio_data_buf[22] ;
 wire \mgmt_gpio_data_buf[23] ;
 wire \mgmt_gpio_data_buf[2] ;
 wire \mgmt_gpio_data_buf[3] ;
 wire \mgmt_gpio_data_buf[4] ;
 wire \mgmt_gpio_data_buf[5] ;
 wire \mgmt_gpio_data_buf[6] ;
 wire \mgmt_gpio_data_buf[7] ;
 wire \mgmt_gpio_data_buf[8] ;
 wire \mgmt_gpio_data_buf[9] ;
 wire \mgmt_gpio_out_pre[10] ;
 wire \mgmt_gpio_out_pre[13] ;
 wire \mgmt_gpio_out_pre[14] ;
 wire \mgmt_gpio_out_pre[15] ;
 wire \mgmt_gpio_out_pre[32] ;
 wire \mgmt_gpio_out_pre[33] ;
 wire \mgmt_gpio_out_pre[6] ;
 wire \mgmt_gpio_out_pre[8] ;
 wire \mgmt_gpio_out_pre[9] ;
 wire \pad_count_1[0] ;
 wire \pad_count_1[1] ;
 wire \pad_count_1[2] ;
 wire \pad_count_1[3] ;
 wire \pad_count_1[4] ;
 wire \pad_count_2[0] ;
 wire \pad_count_2[1] ;
 wire \pad_count_2[2] ;
 wire \pad_count_2[3] ;
 wire \pad_count_2[4] ;
 wire \pad_count_2[5] ;
 wire reset_reg;
 wire serial_bb_clock;
 wire serial_bb_data_1;
 wire serial_bb_data_2;
 wire serial_bb_enable;
 wire serial_bb_load;
 wire serial_bb_resetn;
 wire serial_busy;
 wire serial_clock_pre;
 wire \serial_data_staging_1[0] ;
 wire \serial_data_staging_1[10] ;
 wire \serial_data_staging_1[11] ;
 wire \serial_data_staging_1[12] ;
 wire \serial_data_staging_1[1] ;
 wire \serial_data_staging_1[2] ;
 wire \serial_data_staging_1[3] ;
 wire \serial_data_staging_1[4] ;
 wire \serial_data_staging_1[5] ;
 wire \serial_data_staging_1[6] ;
 wire \serial_data_staging_1[7] ;
 wire \serial_data_staging_1[8] ;
 wire \serial_data_staging_1[9] ;
 wire \serial_data_staging_2[0] ;
 wire \serial_data_staging_2[10] ;
 wire \serial_data_staging_2[11] ;
 wire \serial_data_staging_2[12] ;
 wire \serial_data_staging_2[1] ;
 wire \serial_data_staging_2[2] ;
 wire \serial_data_staging_2[3] ;
 wire \serial_data_staging_2[4] ;
 wire \serial_data_staging_2[5] ;
 wire \serial_data_staging_2[6] ;
 wire \serial_data_staging_2[7] ;
 wire \serial_data_staging_2[8] ;
 wire \serial_data_staging_2[9] ;
 wire serial_load_pre;
 wire serial_resetn_pre;
 wire serial_xfer;
 wire trap_output_dest;
 wire \wbbd_addr[0] ;
 wire \wbbd_addr[1] ;
 wire \wbbd_addr[2] ;
 wire \wbbd_addr[3] ;
 wire \wbbd_addr[4] ;
 wire \wbbd_addr[5] ;
 wire \wbbd_addr[6] ;
 wire wbbd_busy;
 wire \wbbd_data[0] ;
 wire \wbbd_data[1] ;
 wire \wbbd_data[2] ;
 wire \wbbd_data[3] ;
 wire \wbbd_data[4] ;
 wire \wbbd_data[5] ;
 wire \wbbd_data[6] ;
 wire \wbbd_data[7] ;
 wire wbbd_sck;
 wire \wbbd_state[0] ;
 wire \wbbd_state[1] ;
 wire \wbbd_state[2] ;
 wire \wbbd_state[3] ;
 wire \wbbd_state[4] ;
 wire \wbbd_state[5] ;
 wire \wbbd_state[6] ;
 wire \wbbd_state[7] ;
 wire \wbbd_state[8] ;
 wire \wbbd_state[9] ;
 wire wbbd_write;
 wire \xfer_count[0] ;
 wire \xfer_count[1] ;
 wire \xfer_count[2] ;
 wire \xfer_count[3] ;
 wire \xfer_state[0] ;
 wire \xfer_state[1] ;
 wire \xfer_state[2] ;
 wire \xfer_state[3] ;
 wire net99;
 wire net98;
 wire net97;
 wire net96;
 wire net95;
 wire net94;
 wire net93;
 wire net92;
 wire net91;
 wire net90;
 wire net89;
 wire net88;
 wire net87;
 wire net86;
 wire net85;
 wire net84;
 wire net83;
 wire net82;
 wire net81;
 wire net80;
 wire net79;
 wire net78;
 wire net77;
 wire net76;
 wire net75;
 wire net74;
 wire net73;
 wire net72;
 wire net71;
 wire net70;
 wire net69;
 wire net68;
 wire net67;
 wire net66;
 wire net65;
 wire net64;
 wire net63;
 wire net62;
 wire net61;
 wire net60;
 wire net59;
 wire net58;
 wire net57;
 wire net56;
 wire net55;
 wire net54;
 wire net53;
 wire net52;
 wire net51;
 wire net50;
 wire net49;
 wire net48;
 wire net47;
 wire net46;
 wire net45;
 wire net44;
 wire net43;
 wire net42;
 wire net41;
 wire net40;
 wire net39;
 wire net38;
 wire net37;
 wire net36;
 wire net35;
 wire net34;
 wire net33;
 wire net32;
 wire net31;
 wire net30;
 wire net29;
 wire net28;
 wire net27;
 wire net26;
 wire net25;
 wire net24;
 wire net23;
 wire net22;
 wire net21;
 wire net20;
 wire net19;
 wire net18;
 wire net17;
 wire net16;
 wire net15;
 wire net14;
 wire net13;
 wire net12;
 wire net11;
 wire net10;
 wire net9;
 wire net8;
 wire net7;
 wire net6;
 wire net5;
 wire net4;
 wire net3;
 wire net2;
 wire net1;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net506;
 wire clknet_1_0_0_wb_clk_i;
 wire clknet_1_0_1_wb_clk_i;
 wire clknet_1_1_0_wb_clk_i;
 wire clknet_1_1_1_wb_clk_i;
 wire clknet_2_0_0_wb_clk_i;
 wire clknet_2_1_0_wb_clk_i;
 wire clknet_2_2_0_wb_clk_i;
 wire clknet_2_3_0_wb_clk_i;
 wire clknet_3_0_0_wb_clk_i;
 wire clknet_3_1_0_wb_clk_i;
 wire clknet_3_2_0_wb_clk_i;
 wire clknet_3_3_0_wb_clk_i;
 wire clknet_3_4_0_wb_clk_i;
 wire clknet_3_5_0_wb_clk_i;
 wire clknet_3_6_0_wb_clk_i;
 wire clknet_3_7_0_wb_clk_i;
 wire clknet_leaf_0_csclk;
 wire clknet_leaf_1_csclk;
 wire clknet_leaf_2_csclk;
 wire clknet_leaf_3_csclk;
 wire clknet_leaf_4_csclk;
 wire clknet_leaf_5_csclk;
 wire clknet_leaf_6_csclk;
 wire clknet_leaf_7_csclk;
 wire clknet_leaf_9_csclk;
 wire clknet_leaf_10_csclk;
 wire clknet_leaf_11_csclk;
 wire clknet_leaf_12_csclk;
 wire clknet_leaf_13_csclk;
 wire clknet_leaf_14_csclk;
 wire clknet_leaf_16_csclk;
 wire clknet_leaf_17_csclk;
 wire clknet_leaf_18_csclk;
 wire clknet_leaf_19_csclk;
 wire clknet_leaf_20_csclk;
 wire clknet_leaf_21_csclk;
 wire clknet_leaf_23_csclk;
 wire clknet_leaf_24_csclk;
 wire clknet_leaf_25_csclk;
 wire clknet_leaf_26_csclk;
 wire clknet_leaf_27_csclk;
 wire clknet_leaf_28_csclk;
 wire clknet_leaf_29_csclk;
 wire clknet_leaf_30_csclk;
 wire clknet_leaf_31_csclk;
 wire clknet_leaf_32_csclk;
 wire clknet_leaf_33_csclk;
 wire clknet_leaf_34_csclk;
 wire clknet_leaf_35_csclk;
 wire clknet_leaf_36_csclk;
 wire clknet_leaf_37_csclk;
 wire clknet_leaf_38_csclk;
 wire clknet_leaf_39_csclk;
 wire clknet_leaf_40_csclk;
 wire clknet_leaf_41_csclk;
 wire clknet_leaf_42_csclk;
 wire clknet_leaf_43_csclk;
 wire clknet_leaf_45_csclk;
 wire clknet_leaf_46_csclk;
 wire clknet_leaf_47_csclk;
 wire clknet_leaf_48_csclk;
 wire clknet_leaf_49_csclk;
 wire clknet_leaf_50_csclk;
 wire clknet_leaf_52_csclk;
 wire clknet_leaf_53_csclk;
 wire clknet_leaf_55_csclk;
 wire clknet_leaf_56_csclk;
 wire clknet_leaf_57_csclk;
 wire clknet_leaf_58_csclk;
 wire clknet_leaf_59_csclk;
 wire clknet_leaf_60_csclk;
 wire clknet_leaf_61_csclk;
 wire clknet_leaf_62_csclk;
 wire clknet_leaf_63_csclk;
 wire clknet_leaf_64_csclk;
 wire clknet_leaf_65_csclk;
 wire clknet_leaf_66_csclk;
 wire clknet_leaf_67_csclk;
 wire clknet_leaf_68_csclk;
 wire clknet_leaf_69_csclk;
 wire clknet_leaf_70_csclk;
 wire clknet_leaf_71_csclk;
 wire clknet_leaf_72_csclk;
 wire clknet_leaf_73_csclk;
 wire clknet_leaf_74_csclk;
 wire clknet_leaf_75_csclk;
 wire clknet_leaf_76_csclk;
 wire clknet_leaf_77_csclk;
 wire clknet_leaf_78_csclk;
 wire clknet_leaf_79_csclk;
 wire clknet_leaf_80_csclk;
 wire clknet_leaf_81_csclk;
 wire clknet_leaf_82_csclk;
 wire clknet_leaf_83_csclk;
 wire clknet_leaf_84_csclk;
 wire clknet_leaf_85_csclk;
 wire clknet_leaf_86_csclk;
 wire clknet_0_csclk;
 wire clknet_1_0_0_csclk;
 wire clknet_1_0_1_csclk;
 wire clknet_1_1_0_csclk;
 wire clknet_1_1_1_csclk;
 wire clknet_2_0_0_csclk;
 wire clknet_2_1_0_csclk;
 wire clknet_2_2_0_csclk;
 wire clknet_2_3_0_csclk;
 wire clknet_3_0_0_csclk;
 wire clknet_3_1_0_csclk;
 wire clknet_3_2_0_csclk;
 wire clknet_3_3_0_csclk;
 wire clknet_3_4_0_csclk;
 wire clknet_3_5_0_csclk;
 wire clknet_3_6_0_csclk;
 wire clknet_3_7_0_csclk;
 wire clknet_opt_1_0_csclk;
 wire clknet_opt_2_0_csclk;
 wire clknet_0__1160_;
 wire clknet_1_0__leaf__1160_;
 wire clknet_1_1__leaf__1160_;
 wire clknet_0_wbbd_sck;
 wire clknet_1_0__leaf_wbbd_sck;
 wire clknet_1_1__leaf_wbbd_sck;
 wire net507;
 wire net508;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net754;
 wire net755;
 wire net756;
 wire net757;
 wire net758;
 wire net759;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net770;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net778;
 wire net779;
 wire net780;
 wire net781;
 wire net782;
 wire net783;
 wire net784;
 wire net785;
 wire net786;
 wire net787;
 wire net788;
 wire net789;
 wire net790;
 wire net791;
 wire net792;
 wire net793;
 wire net794;
 wire net795;
 wire net796;
 wire net797;
 wire net798;
 wire net799;
 wire net800;
 wire net801;
 wire net802;
 wire net803;
 wire net804;
 wire net805;
 wire net806;
 wire net807;
 wire net808;
 wire net809;
 wire net810;
 wire net811;
 wire net812;
 wire net813;
 wire net814;
 wire net815;
 wire net816;
 wire net817;
 wire net818;
 wire net819;
 wire net820;
 wire net821;
 wire net822;
 wire net823;
 wire net824;
 wire net825;
 wire net826;
 wire net827;
 wire net828;
 wire net829;
 wire net830;
 wire net831;
 wire net832;
 wire net833;
 wire net834;
 wire net835;
 wire net836;
 wire net837;
 wire net838;
 wire net839;
 wire net840;
 wire net841;
 wire net842;
 wire net843;
 wire net844;
 wire net845;
 wire net846;
 wire net847;
 wire net848;
 wire net849;
 wire net850;
 wire net851;
 wire net852;
 wire net853;
 wire net854;
 wire net855;
 wire net856;
 wire net857;
 wire net858;
 wire net859;
 wire net860;
 wire net861;
 wire net862;
 wire net863;
 wire net864;
 wire net865;
 wire net866;
 wire net867;
 wire net868;
 wire net869;
 wire net870;
 wire net871;
 wire net872;
 wire net873;
 wire net874;
 wire net875;
 wire net876;
 wire net877;
 wire net878;
 wire net879;
 wire net880;
 wire net881;
 wire net882;
 wire net883;
 wire net884;
 wire net885;
 wire net886;
 wire net887;
 wire net888;
 wire net889;
 wire net890;
 wire net891;
 wire net892;
 wire net893;
 wire net894;
 wire net895;
 wire net896;
 wire net897;
 wire net898;
 wire net899;
 wire net900;
 wire net901;
 wire net902;
 wire net903;
 wire net904;
 wire net905;
 wire net906;
 wire net907;
 wire net908;
 wire net909;
 wire net910;
 wire net911;
 wire net912;
 wire net913;
 wire net914;
 wire net915;
 wire net916;
 wire net917;
 wire net918;
 wire net919;
 wire net920;
 wire net921;
 wire net922;
 wire net923;
 wire net924;
 wire net925;
 wire net926;
 wire net927;
 wire net928;
 wire net929;
 wire net930;
 wire net931;
 wire net932;
 wire net933;
 wire net934;
 wire net935;
 wire net936;
 wire net937;
 wire net938;
 wire net939;
 wire net940;
 wire net941;
 wire net942;
 wire net943;
 wire net944;
 wire net945;
 wire net946;
 wire net947;
 wire net948;
 wire net949;
 wire net950;
 wire net951;
 wire net952;
 wire net953;
 wire net954;
 wire net955;
 wire net956;
 wire net957;
 wire net958;
 wire net959;
 wire net960;
 wire net961;
 wire net962;
 wire net963;
 wire net964;
 wire net965;
 wire net966;
 wire net967;
 wire net968;
 wire net969;
 wire net970;
 wire net971;
 wire net972;
 wire net973;
 wire net974;
 wire net975;
 wire net976;
 wire net977;
 wire net978;
 wire net979;
 wire net980;
 wire net981;
 wire net982;
 wire net983;
 wire net984;
 wire net985;
 wire net986;
 wire net987;
 wire net988;
 wire net989;
 wire net990;
 wire net991;
 wire net992;
 wire net993;
 wire net994;
 wire net995;
 wire net996;
 wire net997;
 wire net998;
 wire net999;
 wire net1000;
 wire net1001;
 wire net1002;
 wire net1003;
 wire net1004;
 wire net1005;
 wire net1006;
 wire net1007;
 wire net1008;
 wire net1009;
 wire net1010;
 wire net1011;
 wire net1012;
 wire net1013;
 wire net1014;
 wire net1015;
 wire net1016;
 wire net1017;
 wire net1018;
 wire net1019;
 wire net1020;
 wire net1021;
 wire net1022;
 wire net1023;
 wire net1024;
 wire net1025;
 wire net1026;
 wire net1027;
 wire net1028;
 wire net1029;
 wire net1030;
 wire net1031;
 wire net1032;
 wire net1033;
 wire net1034;
 wire net1035;
 wire net1036;
 wire net1037;
 wire net1038;
 wire net1039;
 wire net1040;
 wire net1041;
 wire net1042;
 wire net1043;
 wire net1044;
 wire net1045;
 wire net1046;
 wire net1047;
 wire net1048;
 wire net1049;
 wire net1050;
 wire net1051;
 wire net1052;
 wire net1053;
 wire net1054;
 wire net1055;
 wire net1056;
 wire net1057;
 wire net1058;
 wire net1059;
 wire net1060;
 wire net1061;
 wire net1062;
 wire net1063;
 wire net1064;
 wire net1065;
 wire net1066;
 wire net1067;
 wire net1068;
 wire net1069;
 wire net1070;
 wire net1071;
 wire net1072;
 wire net1073;
 wire net1074;
 wire net1075;
 wire net1076;
 wire net1077;
 wire net1078;
 wire net1079;
 wire net1080;
 wire net1081;
 wire net1082;
 wire net1083;
 wire net1084;
 wire net1085;
 wire net1086;
 wire net1087;
 wire net1088;
 wire net1089;
 wire net1090;
 wire net1091;
 wire net1092;
 wire net1093;
 wire net1094;
 wire net1095;
 wire net1096;
 wire net1097;
 wire net1098;
 wire net1099;
 wire net1100;
 wire net1101;
 wire net1102;
 wire net1103;
 wire net1104;
 wire net1105;
 wire net1106;
 wire net1107;
 wire net1108;
 wire net1109;
 wire net1110;
 wire net1111;
 wire net1112;
 wire net1113;
 wire net1114;
 wire net1115;
 wire net1116;
 wire net1117;
 wire net1118;
 wire net1119;
 wire net1120;
 wire net1121;
 wire net1122;
 wire net1123;
 wire net1124;
 wire net1125;
 wire net1126;
 wire net1127;
 wire net1128;
 wire net1129;
 wire net1130;
 wire net1131;
 wire net1132;
 wire net1133;
 wire net1134;
 wire net1135;
 wire net1136;
 wire net1137;
 wire net1138;
 wire net1139;
 wire net1140;
 wire net1141;
 wire net1142;
 wire net1143;
 wire net1144;
 wire net1145;
 wire net1146;
 wire net1147;
 wire net1148;
 wire net1149;
 wire net1150;
 wire net1151;
 wire net1152;
 wire net1153;
 wire net1154;
 wire net1155;
 wire net1156;
 wire net1157;
 wire net1158;
 wire net1159;
 wire net1160;
 wire net1161;
 wire net1162;
 wire net1163;
 wire net1164;
 wire net1165;
 wire net1166;
 wire net1167;
 wire net1168;
 wire net1169;
 wire net1170;
 wire net1171;
 wire net1172;
 wire net1173;
 wire net1174;
 wire net1175;
 wire net1176;
 wire net1177;
 wire net1178;
 wire net1179;
 wire net1180;
 wire net1181;
 wire net1182;
 wire net1183;
 wire net1184;
 wire net1185;
 wire net1186;
 wire net1187;
 wire net1188;
 wire net1189;
 wire net1190;
 wire net1191;
 wire net1192;
 wire net1193;
 wire net1194;
 wire net1195;
 wire net1196;
 wire net1197;
 wire net1198;
 wire net1199;
 wire net1200;
 wire net1201;
 wire net1202;
 wire net1203;
 wire net1204;
 wire net1205;
 wire net1206;
 wire net1207;
 wire net1208;
 wire net1209;
 wire net1210;
 wire net1211;
 wire net1212;
 wire net1213;
 wire net1214;
 wire net1215;
 wire net1216;
 wire net1217;
 wire net1218;
 wire net1219;
 wire net1220;
 wire net1221;
 wire net1222;
 wire net1223;
 wire net1224;
 wire net1225;
 wire net1226;
 wire net1227;
 wire net1228;
 wire net1229;
 wire net1230;
 wire net1231;
 wire net1232;
 wire net1233;
 wire net1234;
 wire net1235;
 wire net1236;
 wire net1237;
 wire net1238;
 wire net1239;
 wire net1240;
 wire net1241;
 wire net1242;
 wire net1243;
 wire net1244;
 wire net1245;
 wire net1246;
 wire net1247;
 wire net1248;
 wire net1249;
 wire net1250;
 wire net1251;
 wire net1252;
 wire net1253;
 wire net1254;
 wire net1255;
 wire net1256;
 wire net1257;
 wire net1258;
 wire net1259;
 wire net1260;
 wire net1261;
 wire net1262;
 wire net1263;
 wire net1264;
 wire net1265;
 wire net1266;
 wire net1267;
 wire net1268;
 wire net1269;
 wire net1270;
 wire net1271;
 wire net1272;
 wire net1273;
 wire net1274;
 wire net1275;
 wire net1276;
 wire net1277;
 wire net1278;
 wire net1279;
 wire net1280;
 wire net1281;
 wire net1282;
 wire net1283;
 wire net1284;
 wire net1285;
 wire net1286;
 wire net1287;
 wire net1288;
 wire net1289;
 wire net1290;
 wire net1291;
 wire net1292;
 wire net1293;
 wire net1294;
 wire net1295;
 wire net1296;
 wire net1297;
 wire net1298;
 wire net1299;
 wire net1300;
 wire net1301;
 wire net1302;
 wire net1303;
 wire net1304;
 wire net1305;
 wire net1306;
 wire net1307;
 wire net1308;
 wire net1309;
 wire net1310;
 wire net1311;
 wire net1312;
 wire net1313;
 wire net1314;
 wire net1315;
 wire net1316;
 wire net1317;
 wire net1318;
 wire net1319;
 wire net1320;
 wire net1321;
 wire net1322;
 wire net1323;
 wire net1324;
 wire net1325;
 wire net1326;
 wire net1327;
 wire net1328;
 wire net1329;
 wire net1330;
 wire net1331;
 wire net1332;
 wire net1333;
 wire net1334;
 wire net1335;
 wire net1336;
 wire net1337;
 wire net1338;
 wire net1339;
 wire net1340;
 wire net1341;
 wire net1342;
 wire net1343;
 wire net1344;
 wire net1345;
 wire net1346;
 wire net1347;
 wire net1348;
 wire net1349;
 wire net1350;
 wire net1351;
 wire net1352;
 wire net1353;
 wire net1354;
 wire net1355;
 wire net1356;
 wire net1357;
 wire net1358;
 wire net1359;
 wire net1360;
 wire net1361;
 wire net1362;
 wire net1363;
 wire net1364;
 wire net1365;
 wire net1366;
 wire net1367;
 wire net1368;
 wire net1369;
 wire net1370;
 wire net1371;
 wire net1372;
 wire net1373;
 wire net1374;
 wire net1375;
 wire net1376;
 wire net1377;
 wire net1378;
 wire net1379;
 wire net1380;
 wire net1381;
 wire net1382;
 wire net1383;
 wire net1384;
 wire net1385;
 wire net1386;
 wire net1387;
 wire net1388;
 wire net1389;
 wire net1390;
 wire net1391;
 wire net1392;
 wire net1393;
 wire net1394;
 wire net1395;
 wire net1396;
 wire net1397;
 wire net1398;
 wire net1399;
 wire net1400;
 wire net1401;
 wire net1402;
 wire net1403;
 wire net1404;
 wire net1405;
 wire net1406;
 wire net1407;
 wire net1408;
 wire net1409;
 wire net1410;
 wire net1411;
 wire net1412;
 wire net1413;
 wire net1414;
 wire net1415;
 wire net1416;
 wire net1417;
 wire net1418;
 wire net1419;
 wire net1420;
 wire net1421;
 wire net1422;
 wire net1423;
 wire net1424;
 wire net1425;
 wire net1426;
 wire net1427;
 wire net1428;
 wire net1429;
 wire net1430;
 wire net1431;
 wire net1432;
 wire net1433;
 wire net1434;
 wire net1435;
 wire net1436;
 wire net1437;
 wire net1438;
 wire net1439;
 wire net1440;
 wire net1441;
 wire net1442;
 wire net1443;
 wire net1444;
 wire net1445;
 wire net1446;
 wire net1447;
 wire net1448;
 wire net1449;
 wire net1450;
 wire net1451;
 wire net1452;
 wire net1453;
 wire net1454;
 wire net1455;
 wire net1456;
 wire net1457;
 wire net1458;
 wire net1459;
 wire net1460;
 wire net1461;
 wire net1462;
 wire net1463;
 wire net1464;
 wire net1465;
 wire net1466;
 wire net1467;
 wire net1468;
 wire net1469;
 wire net1470;
 wire net1471;
 wire net1472;
 wire net1473;
 wire net1474;
 wire net1475;
 wire net1476;
 wire net1477;
 wire net1478;
 wire net1479;
 wire net1480;
 wire net1481;
 wire net1482;
 wire net1483;
 wire net1484;
 wire net1485;
 wire net1486;
 wire net1487;
 wire net1488;
 wire net1489;
 wire net1490;
 wire net1491;
 wire net1492;
 wire net1493;
 wire net1494;
 wire net1495;
 wire net1496;
 wire net1497;
 wire net1498;
 wire net1499;
 wire net1500;
 wire net1501;
 wire net1502;
 wire net1503;
 wire net1504;
 wire net1505;
 wire net1506;
 wire net1507;
 wire net1508;
 wire net1509;
 wire net1510;
 wire net1511;
 wire net1512;
 wire net1513;
 wire net1514;
 wire net1515;
 wire net1516;
 wire net1517;
 wire net1518;
 wire net1519;
 wire net1520;
 wire net1521;
 wire net1522;
 wire net1523;
 wire net1524;
 wire net1525;
 wire net1526;
 wire net1527;
 wire net1528;
 wire net1529;
 wire net1530;
 wire net1531;
 wire net1532;
 wire net1533;
 wire net1534;
 wire net1535;
 wire net1536;
 wire net1537;
 wire net1538;
 wire net1539;
 wire net1540;
 wire net1541;
 wire net1542;
 wire net1543;
 wire net1544;
 wire net1545;
 wire net1546;
 wire net1547;
 wire net1548;
 wire net1549;
 wire net1550;
 wire net1551;
 wire net1552;
 wire net1553;
 wire net1554;
 wire net1555;
 wire net1556;
 wire net1557;
 wire net1558;
 wire net1559;
 wire net1560;
 wire net1561;
 wire net1562;
 wire net1563;
 wire net1564;
 wire net509;
 wire net1565;
 wire net1566;
 wire net1567;
 wire net1568;
 wire net1569;
 wire net1570;
 wire net1571;
 wire net1572;
 wire net1573;
 wire net1574;
 wire net1575;
 wire net1576;
 wire net1577;
 wire net1578;
 wire net1579;
 wire net1580;
 wire net1581;
 wire net1582;
 wire net1583;
 wire net1584;
 wire net1585;
 wire net1586;
 wire net1587;
 wire net1588;
 wire net1589;
 wire net1590;
 wire net1591;
 wire net1592;
 wire net1593;
 wire net1594;
 wire net1595;
 wire net1596;
 wire net1597;
 wire net1598;
 wire net1599;
 wire net1600;
 wire net1601;
 wire net1602;
 wire net1603;
 wire net1604;
 wire net1605;
 wire net1606;
 wire net1607;
 wire net1608;
 wire net1609;
 wire net1610;
 wire net1611;
 wire net1612;
 wire net1613;
 wire net1614;
 wire net1615;
 wire net1616;
 wire net1617;
 wire net1618;
 wire net1619;
 wire net1620;
 wire net1621;
 wire net1622;
 wire net1623;
 wire net1624;
 wire net1625;
 wire net1626;
 wire net1627;
 wire net1628;
 wire net1629;
 wire net1630;
 wire net1631;
 wire net1632;
 wire net1633;
 wire net1634;
 wire net1635;
 wire net1636;
 wire net1637;
 wire net1638;
 wire net1639;
 wire net1640;
 wire net1641;
 wire net1642;
 wire net1643;
 wire net1644;
 wire net1645;
 wire net1646;
 wire net1647;
 wire net1648;
 wire net1649;
 wire net1650;
 wire net1651;
 wire net1652;
 wire net1653;
 wire net1654;
 wire net1655;
 wire net1656;
 wire net1657;
 wire net1658;
 wire net1659;
 wire net1660;
 wire net1661;
 wire net1662;
 wire net1663;
 wire net1664;
 wire net1665;
 wire net1666;
 wire net1667;
 wire net1668;
 wire net1669;
 wire net1670;
 wire net1671;
 wire net1672;
 wire net1673;
 wire net1674;
 wire net1675;
 wire net1676;
 wire net1677;
 wire net1678;
 wire net1679;
 wire net1680;
 wire net1681;
 wire net1682;
 wire net1683;
 wire net1684;
 wire net1685;
 wire net1686;
 wire net1687;
 wire net1688;
 wire net1689;
 wire net1690;
 wire net1691;
 wire net1692;
 wire net1693;
 wire net1694;
 wire net1695;
 wire net1696;
 wire net1697;
 wire net1698;
 wire net1699;
 wire net1700;
 wire net1701;
 wire net1702;
 wire net1703;
 wire net1704;
 wire net1705;
 wire net1706;
 wire net1707;
 wire net1708;
 wire net1709;
 wire net1710;
 wire net1711;
 wire net1712;
 wire net1713;
 wire net1714;
 wire net1715;
 wire net1716;
 wire net1717;
 wire net1718;
 wire net1719;
 wire net1720;
 wire net1721;
 wire net1722;
 wire net1723;
 wire net1724;
 wire net1725;
 wire net1726;
 wire net1727;
 wire net1728;
 wire net1729;
 wire net1730;
 wire net1731;
 wire net1732;
 wire net1733;
 wire net1734;
 wire net1735;
 wire net1736;
 wire net1737;
 wire net1738;
 wire net1739;
 wire net1740;
 wire net1741;
 wire net1742;
 wire net1743;
 wire net1744;
 wire net1745;
 wire net1746;
 wire net1747;
 wire net1748;
 wire net1749;
 wire net1750;
 wire net1751;
 wire net1752;
 wire net1753;
 wire net1754;
 wire net1755;
 wire net1756;
 wire net1757;
 wire net1758;
 wire net1759;
 wire net1760;
 wire net1761;
 wire net1762;
 wire net1763;
 wire net1764;
 wire net1765;
 wire net1766;
 wire net1767;
 wire net1768;
 wire net1769;
 wire net1770;
 wire net1771;
 wire net1772;
 wire net1773;
 wire net1774;
 wire net1775;
 wire net1776;
 wire net1777;
 wire net1778;
 wire net1779;
 wire net1780;
 wire net1781;
 wire net1782;
 wire net1783;
 wire net1784;
 wire net1785;
 wire net1786;
 wire net1787;
 wire net1788;
 wire net1789;
 wire net1790;
 wire net1791;
 wire [4:0] clknet_0_mgmt_gpio_in;
 wire [4:0] clknet_1_0_0_mgmt_gpio_in;
 wire [4:0] clknet_1_1_0_mgmt_gpio_in;
 wire [4:0] clknet_2_0_0_mgmt_gpio_in;
 wire [4:0] clknet_2_1_0_mgmt_gpio_in;
 wire [4:0] clknet_2_2_0_mgmt_gpio_in;
 wire [4:0] clknet_2_3_0_mgmt_gpio_in;

 sky130_fd_sc_hd__buf_6 _4349_ (.A(net579),
    .X(_0824_));
 sky130_fd_sc_hd__clkinv_2 _4350_ (.A(net528),
    .Y(_0825_));
 sky130_fd_sc_hd__and2_1 _4351_ (.A(\hkspi.addr[7] ),
    .B(_0825_),
    .X(_0826_));
 sky130_fd_sc_hd__a21oi_1 _4352_ (.A1(net535),
    .A2(net528),
    .B1(_0826_),
    .Y(_0827_));
 sky130_fd_sc_hd__and2_1 _4353_ (.A(net561),
    .B(net528),
    .X(_0828_));
 sky130_fd_sc_hd__or2b_1 _4354_ (.A(\wbbd_addr[6] ),
    .B_N(wbbd_busy),
    .X(_0829_));
 sky130_fd_sc_hd__o31a_1 _4355_ (.A1(net535),
    .A2(wbbd_busy),
    .A3(net562),
    .B1(_0829_),
    .X(_0830_));
 sky130_fd_sc_hd__o21bai_1 _4356_ (.A1(_0824_),
    .A2(net536),
    .B1_N(net563),
    .Y(_0831_));
 sky130_fd_sc_hd__nand2_1 _4357_ (.A(net561),
    .B(_0825_),
    .Y(_0832_));
 sky130_fd_sc_hd__a21bo_1 _4358_ (.A1(net586),
    .A2(net528),
    .B1_N(_0832_),
    .X(_0833_));
 sky130_fd_sc_hd__mux2_1 _4359_ (.A0(net587),
    .A1(net1280),
    .S(net579),
    .X(_0834_));
 sky130_fd_sc_hd__nand2_1 _4360_ (.A(\hkspi.addr[4] ),
    .B(_0825_),
    .Y(_0835_));
 sky130_fd_sc_hd__a21bo_1 _4361_ (.A1(net555),
    .A2(net528),
    .B1_N(_0835_),
    .X(_0836_));
 sky130_fd_sc_hd__mux2_1 _4362_ (.A0(net556),
    .A1(net1363),
    .S(net579),
    .X(_0837_));
 sky130_fd_sc_hd__or3b_1 _4363_ (.A(net564),
    .B(net588),
    .C_N(net557),
    .X(_0838_));
 sky130_fd_sc_hd__buf_8 _4364_ (.A(net1281),
    .X(_0839_));
 sky130_fd_sc_hd__mux2_1 _4365_ (.A0(net555),
    .A1(net545),
    .S(net528),
    .X(_0840_));
 sky130_fd_sc_hd__mux2_4 _4366_ (.A0(_0840_),
    .A1(net568),
    .S(_0824_),
    .X(_0841_));
 sky130_fd_sc_hd__mux2_1 _4367_ (.A0(net545),
    .A1(net514),
    .S(net528),
    .X(_0842_));
 sky130_fd_sc_hd__mux2_4 _4368_ (.A0(net546),
    .A1(net869),
    .S(net579),
    .X(_0843_));
 sky130_fd_sc_hd__nor2b_4 _4369_ (.A(net569),
    .B_N(net547),
    .Y(_0844_));
 sky130_fd_sc_hd__mux2_1 _4370_ (.A0(net514),
    .A1(net513),
    .S(net600),
    .X(_0845_));
 sky130_fd_sc_hd__mux2_4 _4371_ (.A0(net515),
    .A1(net604),
    .S(_0824_),
    .X(_0846_));
 sky130_fd_sc_hd__mux2_1 _4372_ (.A0(net583),
    .A1(net58),
    .S(net528),
    .X(_0847_));
 sky130_fd_sc_hd__mux2_4 _4373_ (.A0(_0847_),
    .A1(net541),
    .S(net580),
    .X(_0848_));
 sky130_fd_sc_hd__nor2b_4 _4374_ (.A(net516),
    .B_N(_0848_),
    .Y(_0849_));
 sky130_fd_sc_hd__nand2_8 _4375_ (.A(net400),
    .B(net399),
    .Y(_0850_));
 sky130_fd_sc_hd__nor2_8 _4376_ (.A(_0839_),
    .B(_0850_),
    .Y(_0851_));
 sky130_fd_sc_hd__nor2_8 _4377_ (.A(net516),
    .B(_0848_),
    .Y(_0852_));
 sky130_fd_sc_hd__nand2_8 _4378_ (.A(_0844_),
    .B(_0852_),
    .Y(_0853_));
 sky130_fd_sc_hd__or2b_1 _4379_ (.A(net557),
    .B_N(net588),
    .X(_0854_));
 sky130_fd_sc_hd__or2_1 _4380_ (.A(net564),
    .B(_0854_),
    .X(_0855_));
 sky130_fd_sc_hd__buf_8 _4381_ (.A(_0855_),
    .X(_0856_));
 sky130_fd_sc_hd__nor2_8 _4382_ (.A(_0853_),
    .B(_0856_),
    .Y(_0857_));
 sky130_fd_sc_hd__nor2b_4 _4383_ (.A(_0848_),
    .B_N(net516),
    .Y(_0858_));
 sky130_fd_sc_hd__nor2_8 _4384_ (.A(net569),
    .B(net547),
    .Y(_0859_));
 sky130_fd_sc_hd__nand2_8 _4385_ (.A(net398),
    .B(_0859_),
    .Y(_0860_));
 sky130_fd_sc_hd__o21ai_1 _4386_ (.A1(_0824_),
    .A2(net536),
    .B1(net563),
    .Y(_0861_));
 sky130_fd_sc_hd__or3b_1 _4387_ (.A(net537),
    .B(net588),
    .C_N(net557),
    .X(_0862_));
 sky130_fd_sc_hd__buf_6 _4388_ (.A(net589),
    .X(_0863_));
 sky130_fd_sc_hd__nor2_2 _4389_ (.A(_0860_),
    .B(_0863_),
    .Y(_0864_));
 sky130_fd_sc_hd__nand2_1 _4390_ (.A(_0834_),
    .B(net557),
    .Y(_0865_));
 sky130_fd_sc_hd__or2_1 _4391_ (.A(net564),
    .B(_0865_),
    .X(_0866_));
 sky130_fd_sc_hd__buf_8 _4392_ (.A(net565),
    .X(_0867_));
 sky130_fd_sc_hd__buf_12 _4393_ (.A(net566),
    .X(_0868_));
 sky130_fd_sc_hd__nand2_1 _4394_ (.A(net569),
    .B(net547),
    .Y(_0869_));
 sky130_fd_sc_hd__inv_4 _4395_ (.A(net570),
    .Y(_0870_));
 sky130_fd_sc_hd__nand2_8 _4396_ (.A(net398),
    .B(_0870_),
    .Y(_0871_));
 sky130_fd_sc_hd__nor2_8 _4397_ (.A(_0868_),
    .B(_0871_),
    .Y(_0872_));
 sky130_fd_sc_hd__a22o_1 _4398_ (.A1(\gpio_configure[26][7] ),
    .A2(net392),
    .B1(_0872_),
    .B2(\gpio_configure[16][7] ),
    .X(_0873_));
 sky130_fd_sc_hd__a221o_1 _4399_ (.A1(net323),
    .A2(_0851_),
    .B1(_0857_),
    .B2(\gpio_configure[3][7] ),
    .C1(_0873_),
    .X(_0874_));
 sky130_fd_sc_hd__nand2_8 _4400_ (.A(_0852_),
    .B(_0870_),
    .Y(_0875_));
 sky130_fd_sc_hd__nor2_8 _4401_ (.A(_0868_),
    .B(_0875_),
    .Y(_0876_));
 sky130_fd_sc_hd__nand2_8 _4402_ (.A(_0858_),
    .B(_0844_),
    .Y(_0877_));
 sky130_fd_sc_hd__or2_1 _4403_ (.A(net588),
    .B(net557),
    .X(_0878_));
 sky130_fd_sc_hd__or2_1 _4404_ (.A(net564),
    .B(net558),
    .X(_0879_));
 sky130_fd_sc_hd__clkbuf_16 _4405_ (.A(_0879_),
    .X(_0880_));
 sky130_fd_sc_hd__nor2_4 _4406_ (.A(_0877_),
    .B(_0880_),
    .Y(_0881_));
 sky130_fd_sc_hd__nor2_1 _4407_ (.A(net566),
    .B(_0877_),
    .Y(_0882_));
 sky130_fd_sc_hd__nand2_8 _4408_ (.A(_0859_),
    .B(_0852_),
    .Y(_0883_));
 sky130_fd_sc_hd__nor2_2 _4409_ (.A(_0868_),
    .B(_0883_),
    .Y(_0884_));
 sky130_fd_sc_hd__a22o_2 _4410_ (.A1(\gpio_configure[12][7] ),
    .A2(net387),
    .B1(net366),
    .B2(\gpio_configure[9][7] ),
    .X(_0885_));
 sky130_fd_sc_hd__a221o_1 _4411_ (.A1(\gpio_configure[15][7] ),
    .A2(_0876_),
    .B1(_0881_),
    .B2(net10),
    .C1(_0885_),
    .X(_0886_));
 sky130_fd_sc_hd__or2_1 _4412_ (.A(net537),
    .B(net558),
    .X(_0887_));
 sky130_fd_sc_hd__buf_8 _4413_ (.A(net559),
    .X(_0888_));
 sky130_fd_sc_hd__nor2_8 _4414_ (.A(_0888_),
    .B(_0853_),
    .Y(_0889_));
 sky130_fd_sc_hd__nor2_8 _4415_ (.A(_0888_),
    .B(_0871_),
    .Y(_0890_));
 sky130_fd_sc_hd__nor2_2 _4416_ (.A(_0860_),
    .B(_0856_),
    .Y(_0891_));
 sky130_fd_sc_hd__nor2b_4 _4417_ (.A(net547),
    .B_N(net569),
    .Y(_0892_));
 sky130_fd_sc_hd__nand2_8 _4418_ (.A(_0858_),
    .B(net548),
    .Y(_0893_));
 sky130_fd_sc_hd__nor2_1 _4419_ (.A(_0893_),
    .B(_0888_),
    .Y(_0894_));
 sky130_fd_sc_hd__a22o_1 _4420_ (.A1(\gpio_configure[2][7] ),
    .A2(net385),
    .B1(net384),
    .B2(\gpio_configure[22][7] ),
    .X(_0895_));
 sky130_fd_sc_hd__a221o_1 _4421_ (.A1(\gpio_configure[19][7] ),
    .A2(_0889_),
    .B1(_0890_),
    .B2(\gpio_configure[24][7] ),
    .C1(_0895_),
    .X(_0896_));
 sky130_fd_sc_hd__buf_12 _4422_ (.A(_0863_),
    .X(_0897_));
 sky130_fd_sc_hd__nor2_8 _4423_ (.A(_0897_),
    .B(_0871_),
    .Y(_0898_));
 sky130_fd_sc_hd__nor2_2 _4424_ (.A(_0883_),
    .B(_0856_),
    .Y(_0899_));
 sky130_fd_sc_hd__nand2_8 _4425_ (.A(net548),
    .B(_0852_),
    .Y(_0900_));
 sky130_fd_sc_hd__buf_12 _4426_ (.A(_0888_),
    .X(_0901_));
 sky130_fd_sc_hd__nor2_4 _4427_ (.A(_0900_),
    .B(_0901_),
    .Y(_0902_));
 sky130_fd_sc_hd__nor2_2 _4428_ (.A(_0893_),
    .B(_0856_),
    .Y(_0903_));
 sky130_fd_sc_hd__a22o_1 _4429_ (.A1(\gpio_configure[21][7] ),
    .A2(net365),
    .B1(net382),
    .B2(\gpio_configure[6][7] ),
    .X(_0904_));
 sky130_fd_sc_hd__a221o_1 _4430_ (.A1(\gpio_configure[32][7] ),
    .A2(_0898_),
    .B1(_0899_),
    .B2(\gpio_configure[1][7] ),
    .C1(_0904_),
    .X(_0905_));
 sky130_fd_sc_hd__or4_1 _4431_ (.A(_0874_),
    .B(_0886_),
    .C(_0896_),
    .D(_0905_),
    .X(_0906_));
 sky130_fd_sc_hd__or2_1 _4432_ (.A(net537),
    .B(_0854_),
    .X(_0907_));
 sky130_fd_sc_hd__buf_12 _4433_ (.A(net538),
    .X(_0908_));
 sky130_fd_sc_hd__clkbuf_16 _4434_ (.A(net539),
    .X(_0909_));
 sky130_fd_sc_hd__nor2_8 _4435_ (.A(_0909_),
    .B(_0875_),
    .Y(_0910_));
 sky130_fd_sc_hd__buf_8 _4436_ (.A(_0910_),
    .X(_0911_));
 sky130_fd_sc_hd__nor2_4 _4437_ (.A(_0893_),
    .B(_0863_),
    .Y(_0912_));
 sky130_fd_sc_hd__nor2_2 _4438_ (.A(_0877_),
    .B(_0897_),
    .Y(_0913_));
 sky130_fd_sc_hd__nor2_2 _4439_ (.A(_0900_),
    .B(_0863_),
    .Y(_0914_));
 sky130_fd_sc_hd__a22o_1 _4440_ (.A1(\gpio_configure[28][7] ),
    .A2(net381),
    .B1(net390),
    .B2(\gpio_configure[29][7] ),
    .X(_0915_));
 sky130_fd_sc_hd__a221o_1 _4441_ (.A1(net42),
    .A2(_0911_),
    .B1(net391),
    .B2(\gpio_configure[30][7] ),
    .C1(_0915_),
    .X(_0916_));
 sky130_fd_sc_hd__buf_12 _4442_ (.A(_0839_),
    .X(_0917_));
 sky130_fd_sc_hd__nand2_8 _4443_ (.A(net397),
    .B(_0849_),
    .Y(_0918_));
 sky130_fd_sc_hd__nor2_8 _4444_ (.A(_0917_),
    .B(_0918_),
    .Y(_0919_));
 sky130_fd_sc_hd__nor2_4 _4445_ (.A(_0883_),
    .B(_0897_),
    .Y(_0920_));
 sky130_fd_sc_hd__a22o_1 _4446_ (.A1(net122),
    .A2(_0919_),
    .B1(net380),
    .B2(\gpio_configure[25][7] ),
    .X(_0921_));
 sky130_fd_sc_hd__nor2_1 _4447_ (.A(net539),
    .B(_0853_),
    .Y(_0922_));
 sky130_fd_sc_hd__nor2_8 _4448_ (.A(net566),
    .B(_0853_),
    .Y(_0923_));
 sky130_fd_sc_hd__nor2_8 _4449_ (.A(_0856_),
    .B(_0875_),
    .Y(_0924_));
 sky130_fd_sc_hd__nor2_2 _4450_ (.A(_0909_),
    .B(_0860_),
    .Y(_0925_));
 sky130_fd_sc_hd__a22o_1 _4451_ (.A1(\gpio_configure[7][7] ),
    .A2(net377),
    .B1(net364),
    .B2(\gpio_configure[34][7] ),
    .X(_0926_));
 sky130_fd_sc_hd__a221o_1 _4452_ (.A1(\gpio_configure[35][7] ),
    .A2(net379),
    .B1(_0923_),
    .B2(\gpio_configure[11][7] ),
    .C1(_0926_),
    .X(_0927_));
 sky130_fd_sc_hd__buf_12 _4453_ (.A(_0856_),
    .X(_0928_));
 sky130_fd_sc_hd__nor2_4 _4454_ (.A(_0900_),
    .B(_0928_),
    .Y(_0929_));
 sky130_fd_sc_hd__nor2_2 _4455_ (.A(_0883_),
    .B(_0888_),
    .Y(_0930_));
 sky130_fd_sc_hd__a22o_1 _4456_ (.A1(\gpio_configure[5][7] ),
    .A2(net363),
    .B1(_0930_),
    .B2(\gpio_configure[17][7] ),
    .X(_0931_));
 sky130_fd_sc_hd__nor2_2 _4457_ (.A(net566),
    .B(_0893_),
    .Y(_0932_));
 sky130_fd_sc_hd__nor2_4 _4458_ (.A(_0868_),
    .B(_0860_),
    .Y(_0933_));
 sky130_fd_sc_hd__nor2_4 _4459_ (.A(_0901_),
    .B(_0860_),
    .Y(_0934_));
 sky130_fd_sc_hd__nor2_8 _4460_ (.A(_0853_),
    .B(_0880_),
    .Y(_0935_));
 sky130_fd_sc_hd__a22o_1 _4461_ (.A1(\gpio_configure[18][7] ),
    .A2(net361),
    .B1(_0935_),
    .B2(net28),
    .X(_0936_));
 sky130_fd_sc_hd__a221o_1 _4462_ (.A1(\gpio_configure[14][7] ),
    .A2(net375),
    .B1(net362),
    .B2(\gpio_configure[10][7] ),
    .C1(_0936_),
    .X(_0937_));
 sky130_fd_sc_hd__or4_1 _4463_ (.A(_0921_),
    .B(_0927_),
    .C(_0931_),
    .D(_0937_),
    .X(_0938_));
 sky130_fd_sc_hd__nor2_4 _4464_ (.A(net539),
    .B(_0900_),
    .Y(_0939_));
 sky130_fd_sc_hd__nand2_8 _4465_ (.A(_0870_),
    .B(_0849_),
    .Y(_0940_));
 sky130_fd_sc_hd__nor2_8 _4466_ (.A(_0880_),
    .B(_0940_),
    .Y(_0941_));
 sky130_fd_sc_hd__nor2_8 _4467_ (.A(_0877_),
    .B(net539),
    .Y(_0942_));
 sky130_fd_sc_hd__nand2_1 _4468_ (.A(net516),
    .B(_0848_),
    .Y(_0943_));
 sky130_fd_sc_hd__or2_1 _4469_ (.A(_0943_),
    .B(_0869_),
    .X(_0944_));
 sky130_fd_sc_hd__buf_6 _4470_ (.A(_0944_),
    .X(_0945_));
 sky130_fd_sc_hd__nor2_8 _4471_ (.A(_0880_),
    .B(_0945_),
    .Y(_0946_));
 sky130_fd_sc_hd__a22o_1 _4472_ (.A1(\gpio_configure[36][7] ),
    .A2(_0942_),
    .B1(_0946_),
    .B2(net289),
    .X(_0947_));
 sky130_fd_sc_hd__a221o_1 _4473_ (.A1(\gpio_configure[37][7] ),
    .A2(_0939_),
    .B1(_0941_),
    .B2(net297),
    .C1(_0947_),
    .X(_0948_));
 sky130_fd_sc_hd__nor2_8 _4474_ (.A(_0863_),
    .B(_0875_),
    .Y(_0949_));
 sky130_fd_sc_hd__inv_4 _4475_ (.A(_0943_),
    .Y(_0950_));
 sky130_fd_sc_hd__nand2_8 _4476_ (.A(net400),
    .B(_0950_),
    .Y(_0951_));
 sky130_fd_sc_hd__nor2_8 _4477_ (.A(_0880_),
    .B(_0951_),
    .Y(_0952_));
 sky130_fd_sc_hd__nor2_1 _4478_ (.A(_0877_),
    .B(_0901_),
    .Y(_0953_));
 sky130_fd_sc_hd__nor2_8 _4479_ (.A(net539),
    .B(_0940_),
    .Y(_0954_));
 sky130_fd_sc_hd__a22o_1 _4480_ (.A1(\gpio_configure[20][7] ),
    .A2(net360),
    .B1(_0954_),
    .B2(net70),
    .X(_0955_));
 sky130_fd_sc_hd__a221o_1 _4481_ (.A1(\gpio_configure[31][7] ),
    .A2(_0949_),
    .B1(_0952_),
    .B2(net33),
    .C1(_0955_),
    .X(_0956_));
 sky130_fd_sc_hd__nor2_8 _4482_ (.A(_0909_),
    .B(_0883_),
    .Y(_0957_));
 sky130_fd_sc_hd__nor2_8 _4483_ (.A(_0877_),
    .B(_0917_),
    .Y(_0958_));
 sky130_fd_sc_hd__nor2_4 _4484_ (.A(_0853_),
    .B(_0863_),
    .Y(_0959_));
 sky130_fd_sc_hd__nor2_4 _4485_ (.A(_0888_),
    .B(_0875_),
    .Y(_0960_));
 sky130_fd_sc_hd__a22o_1 _4486_ (.A1(\gpio_configure[27][7] ),
    .A2(net388),
    .B1(_0960_),
    .B2(\gpio_configure[23][7] ),
    .X(_0961_));
 sky130_fd_sc_hd__a221o_1 _4487_ (.A1(\gpio_configure[33][7] ),
    .A2(_0957_),
    .B1(_0958_),
    .B2(net117),
    .C1(_0961_),
    .X(_0962_));
 sky130_fd_sc_hd__nor2_4 _4488_ (.A(_0900_),
    .B(_0917_),
    .Y(_0963_));
 sky130_fd_sc_hd__nand2_8 _4489_ (.A(net397),
    .B(_0950_),
    .Y(_0964_));
 sky130_fd_sc_hd__nor2_8 _4490_ (.A(_0909_),
    .B(_0964_),
    .Y(_0965_));
 sky130_fd_sc_hd__nor2_2 _4491_ (.A(_0893_),
    .B(net539),
    .Y(_0966_));
 sky130_fd_sc_hd__nor2_8 _4492_ (.A(_0877_),
    .B(_0856_),
    .Y(_0967_));
 sky130_fd_sc_hd__a22o_1 _4493_ (.A1(net60),
    .A2(net372),
    .B1(_0967_),
    .B2(\gpio_configure[4][7] ),
    .X(_0968_));
 sky130_fd_sc_hd__a221o_1 _4494_ (.A1(net99),
    .A2(_0963_),
    .B1(_0965_),
    .B2(net51),
    .C1(_0968_),
    .X(_0969_));
 sky130_fd_sc_hd__or4_1 _4495_ (.A(_0948_),
    .B(_0956_),
    .C(_0962_),
    .D(_0969_),
    .X(_0970_));
 sky130_fd_sc_hd__nor2_8 _4496_ (.A(_0917_),
    .B(_0871_),
    .Y(_0971_));
 sky130_fd_sc_hd__nor2_8 _4497_ (.A(_0871_),
    .B(_0880_),
    .Y(_0972_));
 sky130_fd_sc_hd__nor2_8 _4498_ (.A(_0871_),
    .B(_0928_),
    .Y(_0973_));
 sky130_fd_sc_hd__buf_6 _4499_ (.A(_0880_),
    .X(_0974_));
 sky130_fd_sc_hd__nor2_8 _4500_ (.A(_0974_),
    .B(_0850_),
    .Y(_0975_));
 sky130_fd_sc_hd__nor2_1 _4501_ (.A(net566),
    .B(_0900_),
    .Y(_0976_));
 sky130_fd_sc_hd__nor2_8 _4502_ (.A(_0839_),
    .B(_0951_),
    .Y(_0977_));
 sky130_fd_sc_hd__a22o_1 _4503_ (.A1(\gpio_configure[13][7] ),
    .A2(net371),
    .B1(_0977_),
    .B2(net108),
    .X(_0978_));
 sky130_fd_sc_hd__a221o_1 _4504_ (.A1(\gpio_configure[8][7] ),
    .A2(_0973_),
    .B1(_0975_),
    .B2(net19),
    .C1(_0978_),
    .X(_0979_));
 sky130_fd_sc_hd__a221o_1 _4505_ (.A1(\gpio_configure[0][7] ),
    .A2(_0971_),
    .B1(_0972_),
    .B2(net280),
    .C1(_0979_),
    .X(_0980_));
 sky130_fd_sc_hd__or4_1 _4506_ (.A(_0916_),
    .B(_0938_),
    .C(_0970_),
    .D(_0980_),
    .X(_0981_));
 sky130_fd_sc_hd__or2_4 _4507_ (.A(_0906_),
    .B(_0981_),
    .X(_0982_));
 sky130_fd_sc_hd__nor3_2 _4508_ (.A(\hkspi.count[2] ),
    .B(\hkspi.count[1] ),
    .C(\hkspi.count[0] ),
    .Y(_0983_));
 sky130_fd_sc_hd__mux2_1 _4509_ (.A0(net1469),
    .A1(_0982_),
    .S(net402),
    .X(_0984_));
 sky130_fd_sc_hd__nand2_4 _4510_ (.A(\hkspi.readmode ),
    .B(\hkspi.state[2] ),
    .Y(_0985_));
 sky130_fd_sc_hd__mux2_1 _4511_ (.A0(_0984_),
    .A1(net1490),
    .S(_0985_),
    .X(_0986_));
 sky130_fd_sc_hd__clkbuf_1 _4512_ (.A(_0986_),
    .X(_0391_));
 sky130_fd_sc_hd__a22o_1 _4513_ (.A1(\gpio_configure[4][6] ),
    .A2(_0967_),
    .B1(_0942_),
    .B2(\gpio_configure[36][6] ),
    .X(_0987_));
 sky130_fd_sc_hd__a221o_1 _4514_ (.A1(net121),
    .A2(_0919_),
    .B1(net362),
    .B2(\gpio_configure[10][6] ),
    .C1(_0987_),
    .X(_0988_));
 sky130_fd_sc_hd__a22o_1 _4515_ (.A1(\gpio_configure[20][6] ),
    .A2(net360),
    .B1(_0851_),
    .B2(net322),
    .X(_0989_));
 sky130_fd_sc_hd__a221o_1 _4516_ (.A1(net116),
    .A2(_0958_),
    .B1(net385),
    .B2(\gpio_configure[2][6] ),
    .C1(_0989_),
    .X(_0990_));
 sky130_fd_sc_hd__a22o_1 _4517_ (.A1(\gpio_configure[32][6] ),
    .A2(_0898_),
    .B1(_0949_),
    .B2(\gpio_configure[31][6] ),
    .X(_0991_));
 sky130_fd_sc_hd__a221o_1 _4518_ (.A1(net59),
    .A2(net372),
    .B1(_0884_),
    .B2(\gpio_configure[9][6] ),
    .C1(_0991_),
    .X(_0992_));
 sky130_fd_sc_hd__a22o_1 _4519_ (.A1(net279),
    .A2(_0972_),
    .B1(_0857_),
    .B2(\gpio_configure[3][6] ),
    .X(_0993_));
 sky130_fd_sc_hd__a221o_1 _4520_ (.A1(\gpio_configure[5][6] ),
    .A2(net363),
    .B1(_0890_),
    .B2(\gpio_configure[24][6] ),
    .C1(_0993_),
    .X(_0994_));
 sky130_fd_sc_hd__or4_1 _4521_ (.A(_0988_),
    .B(_0990_),
    .C(_0992_),
    .D(_0994_),
    .X(_0995_));
 sky130_fd_sc_hd__a22o_1 _4522_ (.A1(\gpio_configure[7][6] ),
    .A2(_0924_),
    .B1(_0910_),
    .B2(net41),
    .X(_0996_));
 sky130_fd_sc_hd__a221o_1 _4523_ (.A1(\gpio_configure[1][6] ),
    .A2(_0899_),
    .B1(_0941_),
    .B2(net296),
    .C1(_0996_),
    .X(_0997_));
 sky130_fd_sc_hd__a22o_1 _4524_ (.A1(\gpio_configure[29][6] ),
    .A2(_0914_),
    .B1(_0946_),
    .B2(net288),
    .X(_0998_));
 sky130_fd_sc_hd__a221o_1 _4525_ (.A1(net50),
    .A2(_0965_),
    .B1(net365),
    .B2(\gpio_configure[21][6] ),
    .C1(_0998_),
    .X(_0999_));
 sky130_fd_sc_hd__a22o_1 _4526_ (.A1(\gpio_configure[12][6] ),
    .A2(_0882_),
    .B1(net381),
    .B2(\gpio_configure[28][6] ),
    .X(_1000_));
 sky130_fd_sc_hd__a221o_1 _4527_ (.A1(net98),
    .A2(_0963_),
    .B1(_0975_),
    .B2(net18),
    .C1(_1000_),
    .X(_1001_));
 sky130_fd_sc_hd__a22o_1 _4528_ (.A1(\gpio_configure[35][6] ),
    .A2(_0922_),
    .B1(_0957_),
    .B2(\gpio_configure[33][6] ),
    .X(_1002_));
 sky130_fd_sc_hd__a221o_1 _4529_ (.A1(net107),
    .A2(_0977_),
    .B1(net364),
    .B2(\gpio_configure[34][6] ),
    .C1(_1002_),
    .X(_1003_));
 sky130_fd_sc_hd__or4_1 _4530_ (.A(_0997_),
    .B(_0999_),
    .C(_1001_),
    .D(_1003_),
    .X(_1004_));
 sky130_fd_sc_hd__nor2_4 _4531_ (.A(_0860_),
    .B(_0974_),
    .Y(_1005_));
 sky130_fd_sc_hd__a22o_1 _4532_ (.A1(\gpio_configure[37][6] ),
    .A2(_0939_),
    .B1(_0930_),
    .B2(\gpio_configure[17][6] ),
    .X(_1006_));
 sky130_fd_sc_hd__a22o_1 _4533_ (.A1(\gpio_configure[14][6] ),
    .A2(_0932_),
    .B1(net382),
    .B2(\gpio_configure[6][6] ),
    .X(_1007_));
 sky130_fd_sc_hd__a221o_1 _4534_ (.A1(\gpio_configure[13][6] ),
    .A2(net371),
    .B1(_0971_),
    .B2(\gpio_configure[0][6] ),
    .C1(_1007_),
    .X(_1008_));
 sky130_fd_sc_hd__a2111o_1 _4535_ (.A1(\gpio_configure[26][6] ),
    .A2(net392),
    .B1(_1005_),
    .C1(_1006_),
    .D1(_1008_),
    .X(_1009_));
 sky130_fd_sc_hd__nand2_8 _4536_ (.A(_0859_),
    .B(_0950_),
    .Y(_1010_));
 sky130_fd_sc_hd__nor2_8 _4537_ (.A(_0917_),
    .B(_1010_),
    .Y(_1011_));
 sky130_fd_sc_hd__mux2_1 _4538_ (.A0(\serial_data_staging_2[12] ),
    .A1(serial_bb_data_2),
    .S(serial_bb_enable),
    .X(_1012_));
 sky130_fd_sc_hd__clkbuf_4 _4539_ (.A(_1012_),
    .X(net308));
 sky130_fd_sc_hd__a22o_1 _4540_ (.A1(\gpio_configure[23][6] ),
    .A2(net373),
    .B1(_1011_),
    .B2(net308),
    .X(_1013_));
 sky130_fd_sc_hd__a221o_1 _4541_ (.A1(\gpio_configure[19][6] ),
    .A2(_0889_),
    .B1(net378),
    .B2(\gpio_configure[11][6] ),
    .C1(_1013_),
    .X(_1014_));
 sky130_fd_sc_hd__a22o_1 _4542_ (.A1(net27),
    .A2(_0935_),
    .B1(_0952_),
    .B2(net32),
    .X(_1015_));
 sky130_fd_sc_hd__a221o_1 _4543_ (.A1(net69),
    .A2(_0954_),
    .B1(net384),
    .B2(\gpio_configure[22][6] ),
    .C1(_1015_),
    .X(_1016_));
 sky130_fd_sc_hd__a22o_1 _4544_ (.A1(\gpio_configure[18][6] ),
    .A2(net361),
    .B1(net388),
    .B2(\gpio_configure[27][6] ),
    .X(_1017_));
 sky130_fd_sc_hd__a221o_1 _4545_ (.A1(\gpio_configure[16][6] ),
    .A2(_0872_),
    .B1(_0973_),
    .B2(\gpio_configure[8][6] ),
    .C1(_1017_),
    .X(_1018_));
 sky130_fd_sc_hd__a22o_1 _4546_ (.A1(\gpio_configure[30][6] ),
    .A2(net391),
    .B1(_0881_),
    .B2(net9),
    .X(_1019_));
 sky130_fd_sc_hd__a221o_1 _4547_ (.A1(\gpio_configure[15][6] ),
    .A2(_0876_),
    .B1(net380),
    .B2(\gpio_configure[25][6] ),
    .C1(_1019_),
    .X(_1020_));
 sky130_fd_sc_hd__or4_1 _4548_ (.A(_1014_),
    .B(_1016_),
    .C(_1018_),
    .D(_1020_),
    .X(_1021_));
 sky130_fd_sc_hd__or4_4 _4549_ (.A(_0995_),
    .B(_1004_),
    .C(_1009_),
    .D(_1021_),
    .X(_1022_));
 sky130_fd_sc_hd__mux2_1 _4550_ (.A0(\hkspi.ldata[5] ),
    .A1(_1022_),
    .S(_0983_),
    .X(_1023_));
 sky130_fd_sc_hd__mux2_1 _4551_ (.A0(_1023_),
    .A1(net1469),
    .S(_0985_),
    .X(_1024_));
 sky130_fd_sc_hd__clkbuf_1 _4552_ (.A(net1470),
    .X(_0390_));
 sky130_fd_sc_hd__a22o_1 _4553_ (.A1(\gpio_configure[37][5] ),
    .A2(_0939_),
    .B1(_0967_),
    .B2(\gpio_configure[4][5] ),
    .X(_1025_));
 sky130_fd_sc_hd__a221o_1 _4554_ (.A1(\gpio_configure[23][5] ),
    .A2(_0960_),
    .B1(net380),
    .B2(\gpio_configure[25][5] ),
    .C1(_1025_),
    .X(_1026_));
 sky130_fd_sc_hd__nand2_8 _4555_ (.A(_0859_),
    .B(net399),
    .Y(_1027_));
 sky130_fd_sc_hd__nor2_4 _4556_ (.A(_0839_),
    .B(_1027_),
    .Y(_1028_));
 sky130_fd_sc_hd__a22o_2 _4557_ (.A1(\gpio_configure[32][5] ),
    .A2(_0898_),
    .B1(_1028_),
    .B2(net262),
    .X(_1029_));
 sky130_fd_sc_hd__a221o_2 _4558_ (.A1(\gpio_configure[11][5] ),
    .A2(_0923_),
    .B1(net381),
    .B2(\gpio_configure[28][5] ),
    .C1(_1029_),
    .X(_1030_));
 sky130_fd_sc_hd__a22o_1 _4559_ (.A1(net25),
    .A2(_0935_),
    .B1(_0894_),
    .B2(\gpio_configure[22][5] ),
    .X(_1031_));
 sky130_fd_sc_hd__a221o_1 _4560_ (.A1(\gpio_configure[30][5] ),
    .A2(_0912_),
    .B1(_0942_),
    .B2(\gpio_configure[36][5] ),
    .C1(_1031_),
    .X(_1032_));
 sky130_fd_sc_hd__mux2_1 _4561_ (.A0(\serial_data_staging_1[12] ),
    .A1(serial_bb_data_1),
    .S(serial_bb_enable),
    .X(_1033_));
 sky130_fd_sc_hd__buf_2 _4562_ (.A(_1033_),
    .X(net307));
 sky130_fd_sc_hd__a22o_1 _4563_ (.A1(\gpio_configure[7][5] ),
    .A2(_0924_),
    .B1(_0946_),
    .B2(net287),
    .X(_1034_));
 sky130_fd_sc_hd__a221o_1 _4564_ (.A1(\gpio_configure[9][5] ),
    .A2(_0884_),
    .B1(_1011_),
    .B2(net307),
    .C1(_1034_),
    .X(_1035_));
 sky130_fd_sc_hd__a22o_2 _4565_ (.A1(\gpio_configure[29][5] ),
    .A2(net390),
    .B1(_0876_),
    .B2(\gpio_configure[15][5] ),
    .X(_1036_));
 sky130_fd_sc_hd__a221o_1 _4566_ (.A1(\gpio_configure[0][5] ),
    .A2(_0971_),
    .B1(_0952_),
    .B2(net31),
    .C1(_1036_),
    .X(_1037_));
 sky130_fd_sc_hd__a22o_1 _4567_ (.A1(\gpio_configure[12][5] ),
    .A2(net387),
    .B1(net376),
    .B2(\gpio_configure[17][5] ),
    .X(_1038_));
 sky130_fd_sc_hd__a221o_2 _4568_ (.A1(\gpio_configure[13][5] ),
    .A2(net371),
    .B1(net359),
    .B2(\gpio_configure[33][5] ),
    .C1(_1038_),
    .X(_1039_));
 sky130_fd_sc_hd__or4_1 _4569_ (.A(_1032_),
    .B(_1035_),
    .C(_1037_),
    .D(_1039_),
    .X(_1040_));
 sky130_fd_sc_hd__a22o_2 _4570_ (.A1(\gpio_configure[21][5] ),
    .A2(net365),
    .B1(net382),
    .B2(\gpio_configure[6][5] ),
    .X(_1041_));
 sky130_fd_sc_hd__a221o_1 _4571_ (.A1(net8),
    .A2(_0881_),
    .B1(_0941_),
    .B2(net295),
    .C1(_1041_),
    .X(_1042_));
 sky130_fd_sc_hd__a221o_1 _4572_ (.A1(\gpio_configure[16][5] ),
    .A2(_0872_),
    .B1(_0851_),
    .B2(net321),
    .C1(_1042_),
    .X(_1043_));
 sky130_fd_sc_hd__or4_1 _4573_ (.A(_1026_),
    .B(_1030_),
    .C(_1040_),
    .D(_1043_),
    .X(_1044_));
 sky130_fd_sc_hd__a22o_1 _4574_ (.A1(net97),
    .A2(_0963_),
    .B1(_0949_),
    .B2(\gpio_configure[31][5] ),
    .X(_1045_));
 sky130_fd_sc_hd__a221o_1 _4575_ (.A1(\gpio_configure[8][5] ),
    .A2(_0973_),
    .B1(_0958_),
    .B2(net114),
    .C1(_1045_),
    .X(_1046_));
 sky130_fd_sc_hd__a22o_1 _4576_ (.A1(\gpio_configure[1][5] ),
    .A2(net383),
    .B1(net362),
    .B2(\gpio_configure[10][5] ),
    .X(_1047_));
 sky130_fd_sc_hd__a221o_2 _4577_ (.A1(net57),
    .A2(net372),
    .B1(net363),
    .B2(\gpio_configure[5][5] ),
    .C1(_1047_),
    .X(_1048_));
 sky130_fd_sc_hd__a211o_1 _4578_ (.A1(net17),
    .A2(_0975_),
    .B1(_1046_),
    .C1(_1048_),
    .X(_1049_));
 sky130_fd_sc_hd__a221o_1 _4579_ (.A1(net106),
    .A2(_0977_),
    .B1(_0857_),
    .B2(\gpio_configure[3][5] ),
    .C1(_1049_),
    .X(_1050_));
 sky130_fd_sc_hd__a22o_1 _4580_ (.A1(net68),
    .A2(_0954_),
    .B1(net385),
    .B2(\gpio_configure[2][5] ),
    .X(_1051_));
 sky130_fd_sc_hd__a221o_1 _4581_ (.A1(\gpio_configure[27][5] ),
    .A2(net388),
    .B1(net364),
    .B2(\gpio_configure[34][5] ),
    .C1(_1051_),
    .X(_1052_));
 sky130_fd_sc_hd__buf_6 _4582_ (.A(_0965_),
    .X(_1053_));
 sky130_fd_sc_hd__a22o_1 _4583_ (.A1(\gpio_configure[18][5] ),
    .A2(net361),
    .B1(_0890_),
    .B2(\gpio_configure[24][5] ),
    .X(_1054_));
 sky130_fd_sc_hd__a221o_1 _4584_ (.A1(\gpio_configure[14][5] ),
    .A2(net375),
    .B1(_1053_),
    .B2(net49),
    .C1(_1054_),
    .X(_1055_));
 sky130_fd_sc_hd__nor2_2 _4585_ (.A(net539),
    .B(_0918_),
    .Y(_1056_));
 sky130_fd_sc_hd__a22o_1 _4586_ (.A1(\gpio_configure[20][5] ),
    .A2(net360),
    .B1(net370),
    .B2(net66),
    .X(_1057_));
 sky130_fd_sc_hd__a221o_1 _4587_ (.A1(\gpio_configure[35][5] ),
    .A2(net379),
    .B1(net386),
    .B2(\gpio_configure[19][5] ),
    .C1(_1057_),
    .X(_1058_));
 sky130_fd_sc_hd__a22o_1 _4588_ (.A1(\gpio_configure[26][5] ),
    .A2(net392),
    .B1(_0910_),
    .B2(net40),
    .X(_1059_));
 sky130_fd_sc_hd__a221o_2 _4589_ (.A1(net120),
    .A2(_0919_),
    .B1(_0972_),
    .B2(net278),
    .C1(_1059_),
    .X(_1060_));
 sky130_fd_sc_hd__or4_1 _4590_ (.A(_1052_),
    .B(_1055_),
    .C(_1058_),
    .D(_1060_),
    .X(_1061_));
 sky130_fd_sc_hd__or3_4 _4591_ (.A(_1044_),
    .B(_1050_),
    .C(_1061_),
    .X(_1062_));
 sky130_fd_sc_hd__mux2_1 _4592_ (.A0(\hkspi.ldata[4] ),
    .A1(_1062_),
    .S(net402),
    .X(_1063_));
 sky130_fd_sc_hd__mux2_1 _4593_ (.A0(_1063_),
    .A1(net1478),
    .S(_0985_),
    .X(_1064_));
 sky130_fd_sc_hd__clkbuf_1 _4594_ (.A(net1479),
    .X(_0389_));
 sky130_fd_sc_hd__nor2_8 _4595_ (.A(_0897_),
    .B(_0918_),
    .Y(_1065_));
 sky130_fd_sc_hd__nor2_4 _4596_ (.A(_0928_),
    .B(_0945_),
    .Y(_1066_));
 sky130_fd_sc_hd__a22o_1 _4597_ (.A1(\gpio_configure[6][4] ),
    .A2(net382),
    .B1(_1066_),
    .B2(\gpio_configure[9][12] ),
    .X(_1067_));
 sky130_fd_sc_hd__a221o_1 _4598_ (.A1(\gpio_configure[20][4] ),
    .A2(_0953_),
    .B1(_0946_),
    .B2(net286),
    .C1(_1067_),
    .X(_1068_));
 sky130_fd_sc_hd__a22o_1 _4599_ (.A1(net24),
    .A2(_0935_),
    .B1(_0933_),
    .B2(\gpio_configure[10][4] ),
    .X(_1069_));
 sky130_fd_sc_hd__a221o_1 _4600_ (.A1(net39),
    .A2(_0910_),
    .B1(_0975_),
    .B2(net16),
    .C1(_1069_),
    .X(_1070_));
 sky130_fd_sc_hd__a211o_1 _4601_ (.A1(net119),
    .A2(_0919_),
    .B1(_1068_),
    .C1(_1070_),
    .X(_1071_));
 sky130_fd_sc_hd__a221o_1 _4602_ (.A1(\gpio_configure[28][4] ),
    .A2(_0913_),
    .B1(_1065_),
    .B2(\gpio_configure[30][12] ),
    .C1(_1071_),
    .X(_1072_));
 sky130_fd_sc_hd__nor2_4 _4603_ (.A(_0839_),
    .B(_0945_),
    .Y(_1073_));
 sky130_fd_sc_hd__a22o_1 _4604_ (.A1(\gpio_configure[21][4] ),
    .A2(_0902_),
    .B1(_1073_),
    .B2(\gpio_configure[1][12] ),
    .X(_1074_));
 sky130_fd_sc_hd__a221o_1 _4605_ (.A1(\gpio_configure[15][4] ),
    .A2(_0876_),
    .B1(_1011_),
    .B2(serial_bb_clock),
    .C1(_1074_),
    .X(_1075_));
 sky130_fd_sc_hd__nor2_8 _4606_ (.A(_0868_),
    .B(_0945_),
    .Y(_1076_));
 sky130_fd_sc_hd__nor2_8 _4607_ (.A(_0897_),
    .B(_1010_),
    .Y(_1077_));
 sky130_fd_sc_hd__nor2_2 _4608_ (.A(_0901_),
    .B(_0945_),
    .Y(_1078_));
 sky130_fd_sc_hd__a22o_1 _4609_ (.A1(net320),
    .A2(_0851_),
    .B1(_1078_),
    .B2(\gpio_configure[25][12] ),
    .X(_1079_));
 sky130_fd_sc_hd__a221o_1 _4610_ (.A1(\gpio_configure[17][12] ),
    .A2(_1076_),
    .B1(_1077_),
    .B2(\gpio_configure[27][12] ),
    .C1(_1079_),
    .X(_1080_));
 sky130_fd_sc_hd__nor2_2 _4611_ (.A(_0897_),
    .B(_0940_),
    .Y(_1081_));
 sky130_fd_sc_hd__a22o_1 _4612_ (.A1(\gpio_configure[5][4] ),
    .A2(_0929_),
    .B1(_1081_),
    .B2(\gpio_configure[32][12] ),
    .X(_1082_));
 sky130_fd_sc_hd__a221o_2 _4613_ (.A1(clknet_2_1_0_mgmt_gpio_in[4]),
    .A2(_0954_),
    .B1(_0952_),
    .B2(net30),
    .C1(_1082_),
    .X(_1083_));
 sky130_fd_sc_hd__nor2_8 _4614_ (.A(_0868_),
    .B(_0850_),
    .Y(_1084_));
 sky130_fd_sc_hd__a22o_1 _4615_ (.A1(\gpio_configure[32][4] ),
    .A2(_0898_),
    .B1(_1084_),
    .B2(\gpio_configure[12][12] ),
    .X(_1085_));
 sky130_fd_sc_hd__a221o_1 _4616_ (.A1(\gpio_configure[11][4] ),
    .A2(net378),
    .B1(_0958_),
    .B2(net113),
    .C1(_1085_),
    .X(_1086_));
 sky130_fd_sc_hd__or4_2 _4617_ (.A(_1075_),
    .B(_1080_),
    .C(_1083_),
    .D(_1086_),
    .X(_1087_));
 sky130_fd_sc_hd__nor2_8 _4618_ (.A(_0901_),
    .B(_0850_),
    .Y(_1088_));
 sky130_fd_sc_hd__a22o_1 _4619_ (.A1(net48),
    .A2(_0965_),
    .B1(_1088_),
    .B2(\gpio_configure[20][12] ),
    .X(_1089_));
 sky130_fd_sc_hd__a221o_1 _4620_ (.A1(\gpio_configure[35][4] ),
    .A2(net379),
    .B1(_0977_),
    .B2(net105),
    .C1(_1089_),
    .X(_1090_));
 sky130_fd_sc_hd__nor2_8 _4621_ (.A(_0897_),
    .B(_1027_),
    .Y(_1091_));
 sky130_fd_sc_hd__nor2_4 _4622_ (.A(_0901_),
    .B(_0964_),
    .Y(_1092_));
 sky130_fd_sc_hd__a22o_1 _4623_ (.A1(\gpio_configure[25][4] ),
    .A2(_0920_),
    .B1(_1092_),
    .B2(\gpio_configure[23][12] ),
    .X(_1093_));
 sky130_fd_sc_hd__a221o_1 _4624_ (.A1(net294),
    .A2(_0941_),
    .B1(_1091_),
    .B2(\gpio_configure[26][12] ),
    .C1(_1093_),
    .X(_1094_));
 sky130_fd_sc_hd__nor2_4 _4625_ (.A(_0897_),
    .B(_0945_),
    .Y(_1095_));
 sky130_fd_sc_hd__nor2_8 _4626_ (.A(_0928_),
    .B(_0918_),
    .Y(_1096_));
 sky130_fd_sc_hd__a22o_1 _4627_ (.A1(net7),
    .A2(_0881_),
    .B1(_1096_),
    .B2(\gpio_configure[6][12] ),
    .X(_1097_));
 sky130_fd_sc_hd__a221o_1 _4628_ (.A1(\gpio_configure[2][4] ),
    .A2(_0891_),
    .B1(_1095_),
    .B2(\gpio_configure[33][12] ),
    .C1(_1097_),
    .X(_1098_));
 sky130_fd_sc_hd__nor2_8 _4629_ (.A(_0897_),
    .B(_0951_),
    .Y(_1099_));
 sky130_fd_sc_hd__nor2_8 _4630_ (.A(_0868_),
    .B(_0951_),
    .Y(_1100_));
 sky130_fd_sc_hd__a22o_1 _4631_ (.A1(\gpio_configure[0][4] ),
    .A2(_0971_),
    .B1(_1100_),
    .B2(\gpio_configure[13][12] ),
    .X(_1101_));
 sky130_fd_sc_hd__a221o_1 _4632_ (.A1(\gpio_configure[33][4] ),
    .A2(net359),
    .B1(_1099_),
    .B2(\gpio_configure[29][12] ),
    .C1(_1101_),
    .X(_1102_));
 sky130_fd_sc_hd__or4_1 _4633_ (.A(_1090_),
    .B(_1094_),
    .C(_1098_),
    .D(_1102_),
    .X(_1103_));
 sky130_fd_sc_hd__nor2_8 _4634_ (.A(_0868_),
    .B(_0918_),
    .Y(_1104_));
 sky130_fd_sc_hd__nor2_8 _4635_ (.A(_0897_),
    .B(_0850_),
    .Y(_1105_));
 sky130_fd_sc_hd__a22o_1 _4636_ (.A1(\gpio_configure[14][4] ),
    .A2(net375),
    .B1(_1105_),
    .B2(\gpio_configure[28][12] ),
    .X(_1106_));
 sky130_fd_sc_hd__a221o_1 _4637_ (.A1(\gpio_configure[37][4] ),
    .A2(net374),
    .B1(_1104_),
    .B2(\gpio_configure[14][12] ),
    .C1(_1106_),
    .X(_1107_));
 sky130_fd_sc_hd__a22o_1 _4638_ (.A1(\gpio_configure[29][4] ),
    .A2(net390),
    .B1(_0890_),
    .B2(\gpio_configure[24][4] ),
    .X(_1108_));
 sky130_fd_sc_hd__a221o_1 _4639_ (.A1(\gpio_configure[7][4] ),
    .A2(_0924_),
    .B1(net364),
    .B2(\gpio_configure[34][4] ),
    .C1(_1108_),
    .X(_1109_));
 sky130_fd_sc_hd__nor2_8 _4640_ (.A(_0928_),
    .B(_0850_),
    .Y(_1110_));
 sky130_fd_sc_hd__nor2_4 _4641_ (.A(_0928_),
    .B(_1010_),
    .Y(_1111_));
 sky130_fd_sc_hd__nor2_8 _4642_ (.A(_0901_),
    .B(_0940_),
    .Y(_1112_));
 sky130_fd_sc_hd__a22o_1 _4643_ (.A1(\gpio_configure[4][4] ),
    .A2(_0967_),
    .B1(_1112_),
    .B2(\gpio_configure[24][12] ),
    .X(_1113_));
 sky130_fd_sc_hd__a221o_1 _4644_ (.A1(\gpio_configure[4][12] ),
    .A2(_1110_),
    .B1(_1111_),
    .B2(\gpio_configure[3][12] ),
    .C1(_1113_),
    .X(_1114_));
 sky130_fd_sc_hd__nor2_8 _4645_ (.A(_0901_),
    .B(_0918_),
    .Y(_1115_));
 sky130_fd_sc_hd__nor2_4 _4646_ (.A(_0928_),
    .B(_0940_),
    .Y(_1116_));
 sky130_fd_sc_hd__a22o_1 _4647_ (.A1(\gpio_configure[27][4] ),
    .A2(net388),
    .B1(net370),
    .B2(net65),
    .X(_1117_));
 sky130_fd_sc_hd__a221o_1 _4648_ (.A1(\gpio_configure[22][12] ),
    .A2(_1115_),
    .B1(_1116_),
    .B2(\gpio_configure[8][12] ),
    .C1(_1117_),
    .X(_1118_));
 sky130_fd_sc_hd__or4_1 _4649_ (.A(_1107_),
    .B(_1109_),
    .C(_1114_),
    .D(_1118_),
    .X(_1119_));
 sky130_fd_sc_hd__nor2_4 _4650_ (.A(_0974_),
    .B(_1010_),
    .Y(_1120_));
 sky130_fd_sc_hd__nor2_8 _4651_ (.A(_0868_),
    .B(_1027_),
    .Y(_1121_));
 sky130_fd_sc_hd__nor2_8 _4652_ (.A(_0901_),
    .B(_0951_),
    .Y(_1122_));
 sky130_fd_sc_hd__a22o_1 _4653_ (.A1(\gpio_configure[18][4] ),
    .A2(net361),
    .B1(_1122_),
    .B2(\gpio_configure[21][12] ),
    .X(_1123_));
 sky130_fd_sc_hd__a221o_1 _4654_ (.A1(\gpio_configure[30][4] ),
    .A2(net391),
    .B1(_1121_),
    .B2(\gpio_configure[10][12] ),
    .C1(_1123_),
    .X(_1124_));
 sky130_fd_sc_hd__a2111o_1 _4655_ (.A1(\gpio_configure[1][4] ),
    .A2(net383),
    .B1(_1005_),
    .C1(_1120_),
    .D1(_1124_),
    .X(_1125_));
 sky130_fd_sc_hd__nor2_4 _4656_ (.A(_0868_),
    .B(_0964_),
    .Y(_1126_));
 sky130_fd_sc_hd__a22o_1 _4657_ (.A1(\gpio_configure[3][4] ),
    .A2(_0857_),
    .B1(_1126_),
    .B2(\gpio_configure[15][12] ),
    .X(_1127_));
 sky130_fd_sc_hd__a221o_1 _4658_ (.A1(\gpio_configure[22][4] ),
    .A2(net384),
    .B1(_1028_),
    .B2(net261),
    .C1(_1127_),
    .X(_1128_));
 sky130_fd_sc_hd__nor2_4 _4659_ (.A(_0909_),
    .B(_1010_),
    .Y(_1129_));
 sky130_fd_sc_hd__nor2_4 _4660_ (.A(_0917_),
    .B(_0940_),
    .Y(_1130_));
 sky130_fd_sc_hd__nor2_8 _4661_ (.A(net539),
    .B(_0951_),
    .Y(_1131_));
 sky130_fd_sc_hd__a22o_1 _4662_ (.A1(net277),
    .A2(_0972_),
    .B1(_1131_),
    .B2(\gpio_configure[37][12] ),
    .X(_1132_));
 sky130_fd_sc_hd__a221o_1 _4663_ (.A1(\gpio_configure[35][12] ),
    .A2(_1129_),
    .B1(_1130_),
    .B2(\gpio_configure[0][12] ),
    .C1(_1132_),
    .X(_1133_));
 sky130_fd_sc_hd__nor2_4 _4664_ (.A(_0928_),
    .B(_1027_),
    .Y(_1134_));
 sky130_fd_sc_hd__nor2_8 _4665_ (.A(_0901_),
    .B(_1027_),
    .Y(_1135_));
 sky130_fd_sc_hd__nor2_8 _4666_ (.A(_0964_),
    .B(_0928_),
    .Y(_1136_));
 sky130_fd_sc_hd__nor2_4 _4667_ (.A(_0928_),
    .B(_0951_),
    .Y(_1137_));
 sky130_fd_sc_hd__a22o_1 _4668_ (.A1(\gpio_configure[7][12] ),
    .A2(_1136_),
    .B1(_1137_),
    .B2(\gpio_configure[5][12] ),
    .X(_1138_));
 sky130_fd_sc_hd__a221o_1 _4669_ (.A1(\gpio_configure[2][12] ),
    .A2(_1134_),
    .B1(_1135_),
    .B2(\gpio_configure[18][12] ),
    .C1(_1138_),
    .X(_1139_));
 sky130_fd_sc_hd__nor2_4 _4670_ (.A(_0839_),
    .B(_0860_),
    .Y(_1140_));
 sky130_fd_sc_hd__a22o_1 _4671_ (.A1(\gpio_configure[36][4] ),
    .A2(_0942_),
    .B1(_1140_),
    .B2(net269),
    .X(_1141_));
 sky130_fd_sc_hd__a221o_1 _4672_ (.A1(net96),
    .A2(_0963_),
    .B1(_0889_),
    .B2(\gpio_configure[19][4] ),
    .C1(_1141_),
    .X(_1142_));
 sky130_fd_sc_hd__or4_2 _4673_ (.A(_1128_),
    .B(_1133_),
    .C(_1139_),
    .D(_1142_),
    .X(_1143_));
 sky130_fd_sc_hd__nor2_8 _4674_ (.A(_0888_),
    .B(_1010_),
    .Y(_1144_));
 sky130_fd_sc_hd__nor2_4 _4675_ (.A(_0964_),
    .B(_0863_),
    .Y(_1145_));
 sky130_fd_sc_hd__a22o_2 _4676_ (.A1(\gpio_configure[19][12] ),
    .A2(_1144_),
    .B1(_1145_),
    .B2(\gpio_configure[31][12] ),
    .X(_1146_));
 sky130_fd_sc_hd__a221o_1 _4677_ (.A1(\gpio_configure[12][4] ),
    .A2(net387),
    .B1(_0872_),
    .B2(\gpio_configure[16][4] ),
    .C1(_1146_),
    .X(_1147_));
 sky130_fd_sc_hd__nor2_8 _4678_ (.A(net566),
    .B(_0940_),
    .Y(_1148_));
 sky130_fd_sc_hd__a22o_1 _4679_ (.A1(\gpio_configure[13][4] ),
    .A2(net371),
    .B1(_1148_),
    .B2(\gpio_configure[16][12] ),
    .X(_1149_));
 sky130_fd_sc_hd__a221o_1 _4680_ (.A1(\gpio_configure[9][4] ),
    .A2(net366),
    .B1(net389),
    .B2(\gpio_configure[31][4] ),
    .C1(_1149_),
    .X(_1150_));
 sky130_fd_sc_hd__nor2_8 _4681_ (.A(net566),
    .B(_1010_),
    .Y(_1151_));
 sky130_fd_sc_hd__a22o_1 _4682_ (.A1(net56),
    .A2(net372),
    .B1(_1151_),
    .B2(\gpio_configure[11][12] ),
    .X(_1152_));
 sky130_fd_sc_hd__a221o_1 _4683_ (.A1(\gpio_configure[26][4] ),
    .A2(net392),
    .B1(_0973_),
    .B2(\gpio_configure[8][4] ),
    .C1(_1152_),
    .X(_1153_));
 sky130_fd_sc_hd__nor2_8 _4684_ (.A(net539),
    .B(_1027_),
    .Y(_1154_));
 sky130_fd_sc_hd__nor2_8 _4685_ (.A(net539),
    .B(_0850_),
    .Y(_1155_));
 sky130_fd_sc_hd__a22o_1 _4686_ (.A1(\gpio_configure[17][4] ),
    .A2(net376),
    .B1(_1155_),
    .B2(\gpio_configure[36][12] ),
    .X(_1156_));
 sky130_fd_sc_hd__a221o_1 _4687_ (.A1(\gpio_configure[23][4] ),
    .A2(net373),
    .B1(_1154_),
    .B2(\gpio_configure[34][12] ),
    .C1(_1156_),
    .X(_1157_));
 sky130_fd_sc_hd__or4_1 _4688_ (.A(_1147_),
    .B(_1150_),
    .C(_1153_),
    .D(_1157_),
    .X(_1158_));
 sky130_fd_sc_hd__or4_1 _4689_ (.A(_1119_),
    .B(_1125_),
    .C(_1143_),
    .D(_1158_),
    .X(_1159_));
 sky130_fd_sc_hd__or4_2 _4690_ (.A(_1072_),
    .B(_1087_),
    .C(_1103_),
    .D(_1159_),
    .X(_1160_));
 sky130_fd_sc_hd__mux2_2 _4691_ (.A0(\hkspi.ldata[3] ),
    .A1(clknet_1_0__leaf__1160_),
    .S(net402),
    .X(_1161_));
 sky130_fd_sc_hd__mux2_2 _4692_ (.A0(_1161_),
    .A1(\hkspi.ldata[4] ),
    .S(_0985_),
    .X(_1162_));
 sky130_fd_sc_hd__buf_1 _4693_ (.A(_1162_),
    .X(_0388_));
 sky130_fd_sc_hd__a22o_1 _4694_ (.A1(\gpio_configure[7][3] ),
    .A2(_0924_),
    .B1(_1148_),
    .B2(\gpio_configure[16][11] ),
    .X(_1163_));
 sky130_fd_sc_hd__a221o_1 _4695_ (.A1(net112),
    .A2(_0958_),
    .B1(_0890_),
    .B2(\gpio_configure[24][3] ),
    .C1(_1163_),
    .X(_1164_));
 sky130_fd_sc_hd__a22o_1 _4696_ (.A1(\gpio_configure[3][3] ),
    .A2(_0857_),
    .B1(_1111_),
    .B2(\gpio_configure[3][11] ),
    .X(_1165_));
 sky130_fd_sc_hd__a221o_1 _4697_ (.A1(\gpio_configure[6][3] ),
    .A2(net382),
    .B1(_1099_),
    .B2(\gpio_configure[29][11] ),
    .C1(_1165_),
    .X(_1166_));
 sky130_fd_sc_hd__a22o_1 _4698_ (.A1(net67),
    .A2(_0954_),
    .B1(_0891_),
    .B2(\gpio_configure[2][3] ),
    .X(_1167_));
 sky130_fd_sc_hd__a221o_1 _4699_ (.A1(\gpio_configure[4][11] ),
    .A2(_1110_),
    .B1(_1155_),
    .B2(\gpio_configure[36][11] ),
    .C1(_1167_),
    .X(_1168_));
 sky130_fd_sc_hd__a22o_1 _4700_ (.A1(\gpio_configure[19][3] ),
    .A2(net386),
    .B1(net391),
    .B2(\gpio_configure[30][3] ),
    .X(_1169_));
 sky130_fd_sc_hd__a221o_2 _4701_ (.A1(\gpio_configure[37][3] ),
    .A2(net374),
    .B1(net381),
    .B2(\gpio_configure[28][3] ),
    .C1(_1169_),
    .X(_1170_));
 sky130_fd_sc_hd__or4_1 _4702_ (.A(_1164_),
    .B(_1166_),
    .C(_1168_),
    .D(_1170_),
    .X(_1171_));
 sky130_fd_sc_hd__a22o_2 _4703_ (.A1(\gpio_configure[12][3] ),
    .A2(net387),
    .B1(_1151_),
    .B2(\gpio_configure[11][11] ),
    .X(_1172_));
 sky130_fd_sc_hd__a221o_1 _4704_ (.A1(net103),
    .A2(_0977_),
    .B1(_0972_),
    .B2(net276),
    .C1(_1172_),
    .X(_1173_));
 sky130_fd_sc_hd__a22o_1 _4705_ (.A1(\gpio_configure[35][3] ),
    .A2(net379),
    .B1(net384),
    .B2(\gpio_configure[22][3] ),
    .X(_1174_));
 sky130_fd_sc_hd__a221o_1 _4706_ (.A1(\gpio_configure[9][3] ),
    .A2(net366),
    .B1(_0952_),
    .B2(net29),
    .C1(_1174_),
    .X(_1175_));
 sky130_fd_sc_hd__a22o_1 _4707_ (.A1(\gpio_configure[26][3] ),
    .A2(net392),
    .B1(net383),
    .B2(\gpio_configure[1][3] ),
    .X(_1176_));
 sky130_fd_sc_hd__a221o_1 _4708_ (.A1(\gpio_configure[20][11] ),
    .A2(_1088_),
    .B1(_1131_),
    .B2(\gpio_configure[37][11] ),
    .C1(_1176_),
    .X(_1177_));
 sky130_fd_sc_hd__a22o_1 _4709_ (.A1(\gpio_configure[31][11] ),
    .A2(_1145_),
    .B1(_1134_),
    .B2(\gpio_configure[2][11] ),
    .X(_1178_));
 sky130_fd_sc_hd__a221o_1 _4710_ (.A1(\gpio_configure[15][3] ),
    .A2(_0876_),
    .B1(net364),
    .B2(\gpio_configure[34][3] ),
    .C1(_1178_),
    .X(_1179_));
 sky130_fd_sc_hd__or4_1 _4711_ (.A(_1173_),
    .B(_1175_),
    .C(_1177_),
    .D(_1179_),
    .X(_1180_));
 sky130_fd_sc_hd__a22o_1 _4712_ (.A1(\gpio_configure[8][3] ),
    .A2(_0973_),
    .B1(_1073_),
    .B2(\gpio_configure[1][11] ),
    .X(_1181_));
 sky130_fd_sc_hd__a221o_1 _4713_ (.A1(\gpio_configure[15][11] ),
    .A2(_1126_),
    .B1(_1066_),
    .B2(\gpio_configure[9][11] ),
    .C1(_1181_),
    .X(_1182_));
 sky130_fd_sc_hd__a221o_1 _4714_ (.A1(\gpio_configure[33][11] ),
    .A2(_1095_),
    .B1(_1121_),
    .B2(\gpio_configure[10][11] ),
    .C1(_1182_),
    .X(_1183_));
 sky130_fd_sc_hd__a22o_2 _4715_ (.A1(net55),
    .A2(net372),
    .B1(net373),
    .B2(\gpio_configure[23][3] ),
    .X(_1184_));
 sky130_fd_sc_hd__a221o_1 _4716_ (.A1(\gpio_configure[14][11] ),
    .A2(_1104_),
    .B1(_1140_),
    .B2(net268),
    .C1(_1184_),
    .X(_1185_));
 sky130_fd_sc_hd__a22o_1 _4717_ (.A1(net260),
    .A2(_1028_),
    .B1(_1092_),
    .B2(\gpio_configure[23][11] ),
    .X(_1186_));
 sky130_fd_sc_hd__a221o_1 _4718_ (.A1(\gpio_configure[16][3] ),
    .A2(_0872_),
    .B1(_0851_),
    .B2(net319),
    .C1(_1186_),
    .X(_1187_));
 sky130_fd_sc_hd__a22o_1 _4719_ (.A1(\gpio_configure[8][11] ),
    .A2(_1116_),
    .B1(_1096_),
    .B2(\gpio_configure[6][11] ),
    .X(_1188_));
 sky130_fd_sc_hd__a221o_1 _4720_ (.A1(\gpio_configure[4][3] ),
    .A2(_0967_),
    .B1(_1077_),
    .B2(\gpio_configure[27][11] ),
    .C1(_1188_),
    .X(_1189_));
 sky130_fd_sc_hd__a22o_1 _4721_ (.A1(\gpio_configure[25][11] ),
    .A2(_1078_),
    .B1(_1154_),
    .B2(\gpio_configure[34][11] ),
    .X(_1190_));
 sky130_fd_sc_hd__a221o_1 _4722_ (.A1(\gpio_configure[25][3] ),
    .A2(_0920_),
    .B1(_1115_),
    .B2(\gpio_configure[22][11] ),
    .C1(_1190_),
    .X(_1191_));
 sky130_fd_sc_hd__or4_1 _4723_ (.A(_1185_),
    .B(_1187_),
    .C(_1189_),
    .D(_1191_),
    .X(_1192_));
 sky130_fd_sc_hd__or4_1 _4724_ (.A(_1171_),
    .B(_1180_),
    .C(_1183_),
    .D(_1192_),
    .X(_1193_));
 sky130_fd_sc_hd__a22o_2 _4725_ (.A1(\gpio_configure[27][3] ),
    .A2(net388),
    .B1(_1105_),
    .B2(\gpio_configure[28][11] ),
    .X(_1194_));
 sky130_fd_sc_hd__a221o_1 _4726_ (.A1(net23),
    .A2(_0935_),
    .B1(_0975_),
    .B2(net14),
    .C1(_1194_),
    .X(_1195_));
 sky130_fd_sc_hd__a22o_1 _4727_ (.A1(net95),
    .A2(_0963_),
    .B1(_1091_),
    .B2(\gpio_configure[26][11] ),
    .X(_1196_));
 sky130_fd_sc_hd__a22o_1 _4728_ (.A1(net46),
    .A2(_0965_),
    .B1(net363),
    .B2(\gpio_configure[5][3] ),
    .X(_1197_));
 sky130_fd_sc_hd__a221o_1 _4729_ (.A1(\gpio_configure[29][3] ),
    .A2(net390),
    .B1(_1130_),
    .B2(\gpio_configure[0][11] ),
    .C1(_1197_),
    .X(_1198_));
 sky130_fd_sc_hd__a22o_1 _4730_ (.A1(serial_bb_load),
    .A2(_1011_),
    .B1(_1056_),
    .B2(net64),
    .X(_1199_));
 sky130_fd_sc_hd__or4_1 _4731_ (.A(_1195_),
    .B(_1196_),
    .C(_1198_),
    .D(_1199_),
    .X(_1200_));
 sky130_fd_sc_hd__a22o_1 _4732_ (.A1(\gpio_configure[33][3] ),
    .A2(net359),
    .B1(_0946_),
    .B2(net284),
    .X(_1201_));
 sky130_fd_sc_hd__a221o_1 _4733_ (.A1(\gpio_configure[7][11] ),
    .A2(_1136_),
    .B1(_1065_),
    .B2(\gpio_configure[30][11] ),
    .C1(_1201_),
    .X(_1202_));
 sky130_fd_sc_hd__nor2_4 _4734_ (.A(_0893_),
    .B(_0839_),
    .Y(_1203_));
 sky130_fd_sc_hd__a22o_2 _4735_ (.A1(\gpio_configure[5][11] ),
    .A2(_1137_),
    .B1(_1081_),
    .B2(\gpio_configure[32][11] ),
    .X(_1204_));
 sky130_fd_sc_hd__a221o_2 _4736_ (.A1(\gpio_configure[14][3] ),
    .A2(net375),
    .B1(_1203_),
    .B2(net127),
    .C1(_1204_),
    .X(_1205_));
 sky130_fd_sc_hd__a22o_1 _4737_ (.A1(\gpio_configure[32][3] ),
    .A2(_0898_),
    .B1(_1084_),
    .B2(\gpio_configure[12][11] ),
    .X(_1206_));
 sky130_fd_sc_hd__a221o_2 _4738_ (.A1(\gpio_configure[18][3] ),
    .A2(net361),
    .B1(net376),
    .B2(\gpio_configure[17][3] ),
    .C1(_1206_),
    .X(_1207_));
 sky130_fd_sc_hd__a22o_1 _4739_ (.A1(net118),
    .A2(_0919_),
    .B1(_0881_),
    .B2(net6),
    .X(_1208_));
 sky130_fd_sc_hd__a221o_1 _4740_ (.A1(net38),
    .A2(_0910_),
    .B1(_1112_),
    .B2(\gpio_configure[24][11] ),
    .C1(_1208_),
    .X(_1209_));
 sky130_fd_sc_hd__or4_1 _4741_ (.A(_1202_),
    .B(_1205_),
    .C(_1207_),
    .D(_1209_),
    .X(_1210_));
 sky130_fd_sc_hd__a22o_1 _4742_ (.A1(\gpio_configure[21][11] ),
    .A2(_1122_),
    .B1(_1135_),
    .B2(\gpio_configure[18][11] ),
    .X(_1211_));
 sky130_fd_sc_hd__a221o_2 _4743_ (.A1(net293),
    .A2(_0941_),
    .B1(_1129_),
    .B2(\gpio_configure[35][11] ),
    .C1(_1211_),
    .X(_1212_));
 sky130_fd_sc_hd__a22o_1 _4744_ (.A1(\gpio_configure[11][3] ),
    .A2(net378),
    .B1(_1100_),
    .B2(\gpio_configure[13][11] ),
    .X(_1213_));
 sky130_fd_sc_hd__a221o_1 _4745_ (.A1(\gpio_configure[20][3] ),
    .A2(net360),
    .B1(_0971_),
    .B2(\gpio_configure[0][3] ),
    .C1(_1213_),
    .X(_1214_));
 sky130_fd_sc_hd__a22o_1 _4746_ (.A1(\gpio_configure[21][3] ),
    .A2(net365),
    .B1(_1144_),
    .B2(\gpio_configure[19][11] ),
    .X(_1215_));
 sky130_fd_sc_hd__a221o_1 _4747_ (.A1(\gpio_configure[10][3] ),
    .A2(_0933_),
    .B1(_1076_),
    .B2(\gpio_configure[17][11] ),
    .C1(_1215_),
    .X(_1216_));
 sky130_fd_sc_hd__nor2_4 _4748_ (.A(_0909_),
    .B(_0871_),
    .Y(_1217_));
 sky130_fd_sc_hd__a22o_2 _4749_ (.A1(\gpio_configure[36][3] ),
    .A2(_0942_),
    .B1(_1217_),
    .B2(net303),
    .X(_1218_));
 sky130_fd_sc_hd__a221o_1 _4750_ (.A1(\gpio_configure[31][3] ),
    .A2(net389),
    .B1(net371),
    .B2(\gpio_configure[13][3] ),
    .C1(_1218_),
    .X(_1219_));
 sky130_fd_sc_hd__or4_2 _4751_ (.A(_1212_),
    .B(_1214_),
    .C(_1216_),
    .D(_1219_),
    .X(_1220_));
 sky130_fd_sc_hd__or4_4 _4752_ (.A(_1193_),
    .B(_1200_),
    .C(_1210_),
    .D(_1220_),
    .X(_1221_));
 sky130_fd_sc_hd__mux2_1 _4753_ (.A0(\hkspi.ldata[2] ),
    .A1(_1221_),
    .S(net402),
    .X(_1222_));
 sky130_fd_sc_hd__mux2_1 _4754_ (.A0(_1222_),
    .A1(net1462),
    .S(_0985_),
    .X(_1223_));
 sky130_fd_sc_hd__clkbuf_1 _4755_ (.A(net1463),
    .X(_0387_));
 sky130_fd_sc_hd__a22o_1 _4756_ (.A1(\gpio_configure[13][2] ),
    .A2(net371),
    .B1(_1092_),
    .B2(\gpio_configure[23][10] ),
    .X(_1224_));
 sky130_fd_sc_hd__a221o_1 _4757_ (.A1(\gpio_configure[11][2] ),
    .A2(net378),
    .B1(_0890_),
    .B2(\gpio_configure[24][2] ),
    .C1(_1224_),
    .X(_1225_));
 sky130_fd_sc_hd__nor2_4 _4758_ (.A(_0839_),
    .B(_0964_),
    .Y(_1226_));
 sky130_fd_sc_hd__a22o_1 _4759_ (.A1(net102),
    .A2(_0977_),
    .B1(_1226_),
    .B2(clk1_output_dest),
    .X(_1227_));
 sky130_fd_sc_hd__a22o_2 _4760_ (.A1(\gpio_configure[16][2] ),
    .A2(_0872_),
    .B1(_1028_),
    .B2(net273),
    .X(_1228_));
 sky130_fd_sc_hd__a22o_1 _4761_ (.A1(\gpio_configure[6][2] ),
    .A2(net382),
    .B1(_1091_),
    .B2(\gpio_configure[26][10] ),
    .X(_1229_));
 sky130_fd_sc_hd__a221o_1 _4762_ (.A1(net37),
    .A2(_0910_),
    .B1(_1136_),
    .B2(\gpio_configure[7][10] ),
    .C1(_1229_),
    .X(_1230_));
 sky130_fd_sc_hd__or4_1 _4763_ (.A(_1225_),
    .B(_1227_),
    .C(_1228_),
    .D(_1230_),
    .X(_1231_));
 sky130_fd_sc_hd__a22o_1 _4764_ (.A1(net5),
    .A2(_0881_),
    .B1(_1081_),
    .B2(\gpio_configure[32][10] ),
    .X(_1232_));
 sky130_fd_sc_hd__a221o_4 _4765_ (.A1(net22),
    .A2(_0935_),
    .B1(_0942_),
    .B2(\gpio_configure[36][2] ),
    .C1(_1232_),
    .X(_1233_));
 sky130_fd_sc_hd__a22o_1 _4766_ (.A1(\gpio_configure[12][2] ),
    .A2(net387),
    .B1(_1077_),
    .B2(\gpio_configure[27][10] ),
    .X(_1234_));
 sky130_fd_sc_hd__a221o_1 _4767_ (.A1(\gpio_configure[19][2] ),
    .A2(net386),
    .B1(net362),
    .B2(\gpio_configure[10][2] ),
    .C1(_1234_),
    .X(_1235_));
 sky130_fd_sc_hd__a22o_1 _4768_ (.A1(\gpio_configure[29][2] ),
    .A2(net390),
    .B1(net391),
    .B2(\gpio_configure[30][2] ),
    .X(_1236_));
 sky130_fd_sc_hd__a221o_1 _4769_ (.A1(\gpio_configure[23][2] ),
    .A2(net373),
    .B1(net385),
    .B2(\gpio_configure[2][2] ),
    .C1(_1236_),
    .X(_1237_));
 sky130_fd_sc_hd__a22o_1 _4770_ (.A1(\gpio_configure[37][10] ),
    .A2(_1131_),
    .B1(_1116_),
    .B2(\gpio_configure[8][10] ),
    .X(_1238_));
 sky130_fd_sc_hd__a221o_1 _4771_ (.A1(\gpio_configure[9][2] ),
    .A2(net366),
    .B1(net370),
    .B2(net63),
    .C1(_1238_),
    .X(_1239_));
 sky130_fd_sc_hd__or4_2 _4772_ (.A(_1233_),
    .B(_1235_),
    .C(_1237_),
    .D(_1239_),
    .X(_1240_));
 sky130_fd_sc_hd__a22o_2 _4773_ (.A1(net26),
    .A2(_0952_),
    .B1(_1078_),
    .B2(\gpio_configure[25][10] ),
    .X(_1241_));
 sky130_fd_sc_hd__a221o_1 _4774_ (.A1(\gpio_configure[20][2] ),
    .A2(net360),
    .B1(_0973_),
    .B2(\gpio_configure[8][2] ),
    .C1(_1241_),
    .X(_1242_));
 sky130_fd_sc_hd__a22o_1 _4775_ (.A1(\gpio_configure[3][2] ),
    .A2(_0857_),
    .B1(_1115_),
    .B2(\gpio_configure[22][10] ),
    .X(_1243_));
 sky130_fd_sc_hd__a221o_1 _4776_ (.A1(net54),
    .A2(net372),
    .B1(_1155_),
    .B2(\gpio_configure[36][10] ),
    .C1(_1243_),
    .X(_1244_));
 sky130_fd_sc_hd__a22o_1 _4777_ (.A1(\gpio_configure[15][10] ),
    .A2(_1126_),
    .B1(_1099_),
    .B2(\gpio_configure[29][10] ),
    .X(_1245_));
 sky130_fd_sc_hd__a221o_1 _4778_ (.A1(\gpio_configure[14][2] ),
    .A2(net375),
    .B1(net376),
    .B2(\gpio_configure[17][2] ),
    .C1(_1245_),
    .X(_1246_));
 sky130_fd_sc_hd__a22o_1 _4779_ (.A1(net292),
    .A2(_0941_),
    .B1(_1129_),
    .B2(\gpio_configure[35][10] ),
    .X(_1247_));
 sky130_fd_sc_hd__a221o_1 _4780_ (.A1(\gpio_configure[5][2] ),
    .A2(_0929_),
    .B1(_0958_),
    .B2(net111),
    .C1(_1247_),
    .X(_1248_));
 sky130_fd_sc_hd__or4_1 _4781_ (.A(_1242_),
    .B(_1244_),
    .C(_1246_),
    .D(_1248_),
    .X(_1249_));
 sky130_fd_sc_hd__or3_1 _4782_ (.A(_1231_),
    .B(_1240_),
    .C(_1249_),
    .X(_1250_));
 sky130_fd_sc_hd__a22o_1 _4783_ (.A1(\gpio_configure[24][10] ),
    .A2(_1112_),
    .B1(_1135_),
    .B2(\gpio_configure[18][10] ),
    .X(_1251_));
 sky130_fd_sc_hd__a221o_4 _4784_ (.A1(\gpio_configure[27][2] ),
    .A2(net388),
    .B1(_1151_),
    .B2(\gpio_configure[11][10] ),
    .C1(_1251_),
    .X(_1252_));
 sky130_fd_sc_hd__a22o_1 _4785_ (.A1(\gpio_configure[33][10] ),
    .A2(_1095_),
    .B1(_1217_),
    .B2(net302),
    .X(_1253_));
 sky130_fd_sc_hd__a221o_1 _4786_ (.A1(\gpio_configure[25][2] ),
    .A2(_0920_),
    .B1(_1203_),
    .B2(net129),
    .C1(_1253_),
    .X(_1254_));
 sky130_fd_sc_hd__a22o_1 _4787_ (.A1(\gpio_configure[37][2] ),
    .A2(net374),
    .B1(_0975_),
    .B2(net13),
    .X(_1255_));
 sky130_fd_sc_hd__a221o_1 _4788_ (.A1(\gpio_configure[20][10] ),
    .A2(_1088_),
    .B1(_1140_),
    .B2(net267),
    .C1(_1255_),
    .X(_1256_));
 sky130_fd_sc_hd__a22o_2 _4789_ (.A1(\gpio_configure[12][10] ),
    .A2(_1084_),
    .B1(_1065_),
    .B2(\gpio_configure[30][10] ),
    .X(_1257_));
 sky130_fd_sc_hd__a221o_1 _4790_ (.A1(\gpio_configure[32][2] ),
    .A2(_0898_),
    .B1(_1096_),
    .B2(\gpio_configure[6][10] ),
    .C1(_1257_),
    .X(_1258_));
 sky130_fd_sc_hd__or4_1 _4791_ (.A(_1252_),
    .B(_1254_),
    .C(_1256_),
    .D(_1258_),
    .X(_1259_));
 sky130_fd_sc_hd__a22o_1 _4792_ (.A1(\gpio_configure[33][2] ),
    .A2(net359),
    .B1(_1145_),
    .B2(\gpio_configure[31][10] ),
    .X(_1260_));
 sky130_fd_sc_hd__a221o_1 _4793_ (.A1(net115),
    .A2(_0919_),
    .B1(_0925_),
    .B2(\gpio_configure[34][2] ),
    .C1(_1260_),
    .X(_1261_));
 sky130_fd_sc_hd__nor2_1 _4794_ (.A(_0974_),
    .B(_1027_),
    .Y(_1262_));
 sky130_fd_sc_hd__a211o_1 _4795_ (.A1(net318),
    .A2(_0851_),
    .B1(_1005_),
    .C1(_1262_),
    .X(_1263_));
 sky130_fd_sc_hd__a221o_1 _4796_ (.A1(\gpio_configure[4][2] ),
    .A2(_0967_),
    .B1(net384),
    .B2(\gpio_configure[22][2] ),
    .C1(_1263_),
    .X(_1264_));
 sky130_fd_sc_hd__or3_1 _4797_ (.A(_1259_),
    .B(_1261_),
    .C(_1264_),
    .X(_1265_));
 sky130_fd_sc_hd__a22o_1 _4798_ (.A1(\gpio_configure[19][10] ),
    .A2(_1144_),
    .B1(_1134_),
    .B2(\gpio_configure[2][10] ),
    .X(_1266_));
 sky130_fd_sc_hd__a221o_1 _4799_ (.A1(\gpio_configure[18][2] ),
    .A2(_0934_),
    .B1(_1110_),
    .B2(\gpio_configure[4][10] ),
    .C1(_1266_),
    .X(_1267_));
 sky130_fd_sc_hd__a22o_1 _4800_ (.A1(net283),
    .A2(_0946_),
    .B1(_1154_),
    .B2(\gpio_configure[34][10] ),
    .X(_1268_));
 sky130_fd_sc_hd__a221o_1 _4801_ (.A1(\gpio_configure[31][2] ),
    .A2(net389),
    .B1(_1130_),
    .B2(\gpio_configure[0][10] ),
    .C1(_1268_),
    .X(_1269_));
 sky130_fd_sc_hd__a22o_1 _4802_ (.A1(\gpio_configure[21][10] ),
    .A2(_1122_),
    .B1(_1066_),
    .B2(\gpio_configure[9][10] ),
    .X(_1270_));
 sky130_fd_sc_hd__a221o_1 _4803_ (.A1(net45),
    .A2(_0965_),
    .B1(_1121_),
    .B2(\gpio_configure[10][10] ),
    .C1(_1270_),
    .X(_1271_));
 sky130_fd_sc_hd__a22o_1 _4804_ (.A1(\gpio_configure[16][10] ),
    .A2(_1148_),
    .B1(_1076_),
    .B2(\gpio_configure[17][10] ),
    .X(_1272_));
 sky130_fd_sc_hd__a221o_1 _4805_ (.A1(serial_bb_resetn),
    .A2(_1011_),
    .B1(_1111_),
    .B2(\gpio_configure[3][10] ),
    .C1(_1272_),
    .X(_1273_));
 sky130_fd_sc_hd__or4_1 _4806_ (.A(_1267_),
    .B(_1269_),
    .C(_1271_),
    .D(_1273_),
    .X(_1274_));
 sky130_fd_sc_hd__a22o_1 _4807_ (.A1(\gpio_configure[28][2] ),
    .A2(net381),
    .B1(_1105_),
    .B2(\gpio_configure[28][10] ),
    .X(_1275_));
 sky130_fd_sc_hd__a221o_1 _4808_ (.A1(\gpio_configure[0][2] ),
    .A2(_0971_),
    .B1(_0876_),
    .B2(\gpio_configure[15][2] ),
    .C1(_1275_),
    .X(_1276_));
 sky130_fd_sc_hd__a22o_1 _4809_ (.A1(\gpio_configure[26][2] ),
    .A2(_0864_),
    .B1(_1137_),
    .B2(\gpio_configure[5][10] ),
    .X(_1277_));
 sky130_fd_sc_hd__a221o_1 _4810_ (.A1(net275),
    .A2(_0972_),
    .B1(net383),
    .B2(\gpio_configure[1][2] ),
    .C1(_1277_),
    .X(_1278_));
 sky130_fd_sc_hd__buf_8 _4811_ (.A(_0954_),
    .X(_1279_));
 sky130_fd_sc_hd__a22o_1 _4812_ (.A1(net94),
    .A2(_0963_),
    .B1(_0924_),
    .B2(\gpio_configure[7][2] ),
    .X(_1280_));
 sky130_fd_sc_hd__a221o_1 _4813_ (.A1(net58),
    .A2(_1279_),
    .B1(_1073_),
    .B2(\gpio_configure[1][10] ),
    .C1(_1280_),
    .X(_1281_));
 sky130_fd_sc_hd__a22o_1 _4814_ (.A1(\gpio_configure[13][10] ),
    .A2(_1100_),
    .B1(_1104_),
    .B2(\gpio_configure[14][10] ),
    .X(_1282_));
 sky130_fd_sc_hd__a221o_1 _4815_ (.A1(\gpio_configure[35][2] ),
    .A2(net379),
    .B1(net365),
    .B2(\gpio_configure[21][2] ),
    .C1(_1282_),
    .X(_1283_));
 sky130_fd_sc_hd__or4_1 _4816_ (.A(_1276_),
    .B(_1278_),
    .C(_1281_),
    .D(_1283_),
    .X(_1284_));
 sky130_fd_sc_hd__or4_4 _4817_ (.A(_1250_),
    .B(_1265_),
    .C(_1274_),
    .D(_1284_),
    .X(_1285_));
 sky130_fd_sc_hd__mux2_1 _4818_ (.A0(\hkspi.ldata[1] ),
    .A1(_1285_),
    .S(net402),
    .X(_1286_));
 sky130_fd_sc_hd__mux2_1 _4819_ (.A0(_1286_),
    .A1(net1467),
    .S(_0985_),
    .X(_1287_));
 sky130_fd_sc_hd__clkbuf_1 _4820_ (.A(net1468),
    .X(_0386_));
 sky130_fd_sc_hd__a22o_1 _4821_ (.A1(net124),
    .A2(_0963_),
    .B1(_1078_),
    .B2(\gpio_configure[25][9] ),
    .X(_1288_));
 sky130_fd_sc_hd__a221o_1 _4822_ (.A1(\gpio_configure[4][1] ),
    .A2(_0967_),
    .B1(_1076_),
    .B2(\gpio_configure[17][9] ),
    .C1(_1288_),
    .X(_1289_));
 sky130_fd_sc_hd__a22o_1 _4823_ (.A1(net272),
    .A2(_1028_),
    .B1(_1137_),
    .B2(\gpio_configure[5][9] ),
    .X(_1290_));
 sky130_fd_sc_hd__a221o_1 _4824_ (.A1(net299),
    .A2(_0972_),
    .B1(_1011_),
    .B2(serial_bb_enable),
    .C1(_1290_),
    .X(_1291_));
 sky130_fd_sc_hd__a22o_1 _4825_ (.A1(net53),
    .A2(_0966_),
    .B1(net374),
    .B2(\gpio_configure[37][1] ),
    .X(_1292_));
 sky130_fd_sc_hd__a221o_1 _4826_ (.A1(net266),
    .A2(_1140_),
    .B1(_1111_),
    .B2(\gpio_configure[3][9] ),
    .C1(_1292_),
    .X(_1293_));
 sky130_fd_sc_hd__a22o_1 _4827_ (.A1(\gpio_configure[24][9] ),
    .A2(_1112_),
    .B1(_1066_),
    .B2(\gpio_configure[9][9] ),
    .X(_1294_));
 sky130_fd_sc_hd__a221o_1 _4828_ (.A1(\gpio_configure[10][1] ),
    .A2(_0933_),
    .B1(_1110_),
    .B2(\gpio_configure[4][9] ),
    .C1(_1294_),
    .X(_1295_));
 sky130_fd_sc_hd__or4_2 _4829_ (.A(_1289_),
    .B(_1291_),
    .C(_1293_),
    .D(_1295_),
    .X(_1296_));
 sky130_fd_sc_hd__nor2_4 _4830_ (.A(_0917_),
    .B(_0875_),
    .Y(_1297_));
 sky130_fd_sc_hd__a22o_1 _4831_ (.A1(\gpio_configure[15][1] ),
    .A2(_0876_),
    .B1(_1297_),
    .B2(irq_2_inputsrc),
    .X(_1298_));
 sky130_fd_sc_hd__a221o_1 _4832_ (.A1(\gpio_configure[19][1] ),
    .A2(_0889_),
    .B1(_1100_),
    .B2(\gpio_configure[13][9] ),
    .C1(_1298_),
    .X(_1299_));
 sky130_fd_sc_hd__a22o_1 _4833_ (.A1(\gpio_configure[10][9] ),
    .A2(_1121_),
    .B1(_1105_),
    .B2(\gpio_configure[28][9] ),
    .X(_1300_));
 sky130_fd_sc_hd__a221o_1 _4834_ (.A1(net104),
    .A2(_0919_),
    .B1(_0924_),
    .B2(\gpio_configure[7][1] ),
    .C1(_1300_),
    .X(_1301_));
 sky130_fd_sc_hd__a22o_1 _4835_ (.A1(\gpio_configure[11][1] ),
    .A2(net378),
    .B1(_0857_),
    .B2(\gpio_configure[3][1] ),
    .X(_1302_));
 sky130_fd_sc_hd__a221o_1 _4836_ (.A1(\gpio_configure[33][1] ),
    .A2(net359),
    .B1(_1073_),
    .B2(\gpio_configure[1][9] ),
    .C1(_1302_),
    .X(_1303_));
 sky130_fd_sc_hd__a22o_1 _4837_ (.A1(\gpio_configure[33][9] ),
    .A2(_1095_),
    .B1(_1091_),
    .B2(\gpio_configure[26][9] ),
    .X(_1304_));
 sky130_fd_sc_hd__a221o_1 _4838_ (.A1(\gpio_configure[8][1] ),
    .A2(_0973_),
    .B1(_1151_),
    .B2(\gpio_configure[11][9] ),
    .C1(_1304_),
    .X(_1305_));
 sky130_fd_sc_hd__a22o_1 _4839_ (.A1(\gpio_configure[35][1] ),
    .A2(net379),
    .B1(net363),
    .B2(\gpio_configure[5][1] ),
    .X(_1306_));
 sky130_fd_sc_hd__a221o_1 _4840_ (.A1(net72),
    .A2(_0910_),
    .B1(_1144_),
    .B2(\gpio_configure[19][9] ),
    .C1(_1306_),
    .X(_1307_));
 sky130_fd_sc_hd__or4_1 _4841_ (.A(_1301_),
    .B(_1303_),
    .C(_1305_),
    .D(_1307_),
    .X(_1308_));
 sky130_fd_sc_hd__a22o_1 _4842_ (.A1(\gpio_configure[27][1] ),
    .A2(_0959_),
    .B1(_0942_),
    .B2(\gpio_configure[36][1] ),
    .X(_1309_));
 sky130_fd_sc_hd__a22o_1 _4843_ (.A1(\gpio_configure[32][1] ),
    .A2(_0898_),
    .B1(_1092_),
    .B2(\gpio_configure[23][9] ),
    .X(_1310_));
 sky130_fd_sc_hd__a221o_1 _4844_ (.A1(\gpio_configure[21][1] ),
    .A2(_0902_),
    .B1(_0881_),
    .B2(net35),
    .C1(_1310_),
    .X(_1311_));
 sky130_fd_sc_hd__a2111o_1 _4845_ (.A1(\gpio_configure[28][1] ),
    .A2(_0913_),
    .B1(_1005_),
    .C1(_1309_),
    .D1(_1311_),
    .X(_1312_));
 sky130_fd_sc_hd__a22o_1 _4846_ (.A1(\gpio_configure[20][9] ),
    .A2(_1088_),
    .B1(_1130_),
    .B2(\gpio_configure[0][9] ),
    .X(_1313_));
 sky130_fd_sc_hd__a22o_1 _4847_ (.A1(\gpio_configure[6][1] ),
    .A2(net382),
    .B1(_0890_),
    .B2(\gpio_configure[24][1] ),
    .X(_1314_));
 sky130_fd_sc_hd__a221o_1 _4848_ (.A1(\gpio_configure[14][1] ),
    .A2(net375),
    .B1(net383),
    .B2(\gpio_configure[1][1] ),
    .C1(_1314_),
    .X(_1315_));
 sky130_fd_sc_hd__a22o_1 _4849_ (.A1(\gpio_configure[7][9] ),
    .A2(_1136_),
    .B1(_1116_),
    .B2(\gpio_configure[8][9] ),
    .X(_1316_));
 sky130_fd_sc_hd__a22o_2 _4850_ (.A1(net285),
    .A2(_0941_),
    .B1(_1155_),
    .B2(\gpio_configure[36][9] ),
    .X(_1317_));
 sky130_fd_sc_hd__a221o_1 _4851_ (.A1(\gpio_configure[29][9] ),
    .A2(_1099_),
    .B1(_1135_),
    .B2(\gpio_configure[18][9] ),
    .C1(_1317_),
    .X(_1318_));
 sky130_fd_sc_hd__or4_1 _4852_ (.A(_1313_),
    .B(_1315_),
    .C(_1316_),
    .D(_1318_),
    .X(_1319_));
 sky130_fd_sc_hd__or4_1 _4853_ (.A(_1299_),
    .B(_1308_),
    .C(_1312_),
    .D(_1319_),
    .X(_1320_));
 sky130_fd_sc_hd__a22o_1 _4854_ (.A1(\gpio_configure[0][1] ),
    .A2(_0971_),
    .B1(_1081_),
    .B2(\gpio_configure[32][9] ),
    .X(_1321_));
 sky130_fd_sc_hd__a221o_1 _4855_ (.A1(\gpio_configure[12][1] ),
    .A2(net387),
    .B1(_1065_),
    .B2(\gpio_configure[30][9] ),
    .C1(_1321_),
    .X(_1322_));
 sky130_fd_sc_hd__a22o_2 _4856_ (.A1(\gpio_configure[2][1] ),
    .A2(net385),
    .B1(_1104_),
    .B2(\gpio_configure[14][9] ),
    .X(_1323_));
 sky130_fd_sc_hd__a221o_1 _4857_ (.A1(net110),
    .A2(_0958_),
    .B1(_0925_),
    .B2(\gpio_configure[34][1] ),
    .C1(_1323_),
    .X(_1324_));
 sky130_fd_sc_hd__nor2_2 _4858_ (.A(_0917_),
    .B(_0853_),
    .Y(_1325_));
 sky130_fd_sc_hd__a22o_2 _4859_ (.A1(\gpio_configure[26][1] ),
    .A2(net392),
    .B1(net380),
    .B2(\gpio_configure[25][1] ),
    .X(_1326_));
 sky130_fd_sc_hd__a221o_1 _4860_ (.A1(\gpio_configure[30][1] ),
    .A2(_0912_),
    .B1(_1325_),
    .B2(net324),
    .C1(_1326_),
    .X(_1327_));
 sky130_fd_sc_hd__nor2_1 _4861_ (.A(_0883_),
    .B(_0917_),
    .Y(_1328_));
 sky130_fd_sc_hd__a22o_1 _4862_ (.A1(net12),
    .A2(_0975_),
    .B1(_1096_),
    .B2(\gpio_configure[6][9] ),
    .X(_1329_));
 sky130_fd_sc_hd__a221o_1 _4863_ (.A1(net282),
    .A2(_0946_),
    .B1(_1328_),
    .B2(net291),
    .C1(_1329_),
    .X(_1330_));
 sky130_fd_sc_hd__or3_2 _4864_ (.A(_1324_),
    .B(_1327_),
    .C(_1330_),
    .X(_1331_));
 sky130_fd_sc_hd__a22o_1 _4865_ (.A1(\gpio_configure[13][1] ),
    .A2(net371),
    .B1(_0952_),
    .B2(net15),
    .X(_1332_));
 sky130_fd_sc_hd__a221o_1 _4866_ (.A1(\gpio_configure[16][1] ),
    .A2(_0872_),
    .B1(_1148_),
    .B2(\gpio_configure[16][9] ),
    .C1(_1332_),
    .X(_1333_));
 sky130_fd_sc_hd__a22o_2 _4867_ (.A1(net317),
    .A2(_0851_),
    .B1(_1145_),
    .B2(\gpio_configure[31][9] ),
    .X(_1334_));
 sky130_fd_sc_hd__a221o_1 _4868_ (.A1(\gpio_configure[9][1] ),
    .A2(net366),
    .B1(_1134_),
    .B2(\gpio_configure[2][9] ),
    .C1(_1334_),
    .X(_1335_));
 sky130_fd_sc_hd__a22o_1 _4869_ (.A1(\gpio_configure[21][9] ),
    .A2(_1122_),
    .B1(_1077_),
    .B2(\gpio_configure[27][9] ),
    .X(_1336_));
 sky130_fd_sc_hd__a221o_1 _4870_ (.A1(net44),
    .A2(_0965_),
    .B1(_1115_),
    .B2(\gpio_configure[22][9] ),
    .C1(_1336_),
    .X(_1337_));
 sky130_fd_sc_hd__a22o_1 _4871_ (.A1(net21),
    .A2(_0935_),
    .B1(_1203_),
    .B2(net128),
    .X(_1338_));
 sky130_fd_sc_hd__a221o_1 _4872_ (.A1(\gpio_configure[29][1] ),
    .A2(net390),
    .B1(net376),
    .B2(\gpio_configure[17][1] ),
    .C1(_1338_),
    .X(_1339_));
 sky130_fd_sc_hd__or4_1 _4873_ (.A(_1333_),
    .B(_1335_),
    .C(_1337_),
    .D(_1339_),
    .X(_1340_));
 sky130_fd_sc_hd__a22o_1 _4874_ (.A1(\gpio_configure[34][9] ),
    .A2(_1154_),
    .B1(_1226_),
    .B2(clk2_output_dest),
    .X(_1341_));
 sky130_fd_sc_hd__a221o_1 _4875_ (.A1(\gpio_configure[20][1] ),
    .A2(net360),
    .B1(net384),
    .B2(\gpio_configure[22][1] ),
    .C1(_1341_),
    .X(_1342_));
 sky130_fd_sc_hd__a22o_1 _4876_ (.A1(net62),
    .A2(net370),
    .B1(_1131_),
    .B2(\gpio_configure[37][9] ),
    .X(_1343_));
 sky130_fd_sc_hd__a221o_1 _4877_ (.A1(\gpio_configure[18][1] ),
    .A2(net361),
    .B1(_1084_),
    .B2(\gpio_configure[12][9] ),
    .C1(_1343_),
    .X(_1344_));
 sky130_fd_sc_hd__nor2_2 _4878_ (.A(_0900_),
    .B(_0974_),
    .Y(_1345_));
 sky130_fd_sc_hd__a22o_1 _4879_ (.A1(\gpio_configure[31][1] ),
    .A2(_0949_),
    .B1(_1345_),
    .B2(net264),
    .X(_1346_));
 sky130_fd_sc_hd__a221o_4 _4880_ (.A1(net47),
    .A2(_0954_),
    .B1(_0977_),
    .B2(net101),
    .C1(_1346_),
    .X(_1347_));
 sky130_fd_sc_hd__a22o_2 _4881_ (.A1(\gpio_configure[35][9] ),
    .A2(_1129_),
    .B1(_1217_),
    .B2(net301),
    .X(_1348_));
 sky130_fd_sc_hd__a221o_1 _4882_ (.A1(\gpio_configure[23][1] ),
    .A2(net373),
    .B1(_1126_),
    .B2(\gpio_configure[15][9] ),
    .C1(_1348_),
    .X(_1349_));
 sky130_fd_sc_hd__or4_1 _4883_ (.A(_1342_),
    .B(_1344_),
    .C(_1347_),
    .D(_1349_),
    .X(_1350_));
 sky130_fd_sc_hd__or4_1 _4884_ (.A(_1322_),
    .B(_1331_),
    .C(_1340_),
    .D(_1350_),
    .X(_1351_));
 sky130_fd_sc_hd__or3_4 _4885_ (.A(_1296_),
    .B(_1320_),
    .C(_1351_),
    .X(_1352_));
 sky130_fd_sc_hd__mux2_1 _4886_ (.A0(\hkspi.ldata[0] ),
    .A1(_1352_),
    .S(net402),
    .X(_1353_));
 sky130_fd_sc_hd__mux2_1 _4887_ (.A0(_1353_),
    .A1(net1486),
    .S(_0985_),
    .X(_1354_));
 sky130_fd_sc_hd__clkbuf_1 _4888_ (.A(_1354_),
    .X(_0385_));
 sky130_fd_sc_hd__inv_2 _4889_ (.A(_0875_),
    .Y(_1355_));
 sky130_fd_sc_hd__inv_2 _4890_ (.A(_0974_),
    .Y(_1356_));
 sky130_fd_sc_hd__nor2_2 _4891_ (.A(_0909_),
    .B(_0945_),
    .Y(_1357_));
 sky130_fd_sc_hd__a32o_1 _4892_ (.A1(net125),
    .A2(_1355_),
    .A3(_1356_),
    .B1(_1357_),
    .B2(hkspi_disable),
    .X(_1358_));
 sky130_fd_sc_hd__a22o_1 _4893_ (.A1(\gpio_configure[14][0] ),
    .A2(net375),
    .B1(_1099_),
    .B2(\gpio_configure[29][8] ),
    .X(_1359_));
 sky130_fd_sc_hd__a22o_1 _4894_ (.A1(\gpio_configure[10][0] ),
    .A2(net362),
    .B1(_1100_),
    .B2(\gpio_configure[13][8] ),
    .X(_1360_));
 sky130_fd_sc_hd__a22o_1 _4895_ (.A1(\gpio_configure[1][0] ),
    .A2(net383),
    .B1(net384),
    .B2(\gpio_configure[22][0] ),
    .X(_1361_));
 sky130_fd_sc_hd__or4_1 _4896_ (.A(_1358_),
    .B(_1359_),
    .C(_1360_),
    .D(_1361_),
    .X(_1362_));
 sky130_fd_sc_hd__a22o_1 _4897_ (.A1(\gpio_configure[5][8] ),
    .A2(_1137_),
    .B1(_1297_),
    .B2(irq_1_inputsrc),
    .X(_1363_));
 sky130_fd_sc_hd__a22o_1 _4898_ (.A1(\gpio_configure[37][0] ),
    .A2(net374),
    .B1(_1112_),
    .B2(\gpio_configure[24][8] ),
    .X(_1364_));
 sky130_fd_sc_hd__a221o_1 _4899_ (.A1(\gpio_configure[30][0] ),
    .A2(_0912_),
    .B1(_1122_),
    .B2(\gpio_configure[21][8] ),
    .C1(_1364_),
    .X(_1365_));
 sky130_fd_sc_hd__a211o_1 _4900_ (.A1(\gpio_configure[15][8] ),
    .A2(_1126_),
    .B1(_1363_),
    .C1(_1365_),
    .X(_1366_));
 sky130_fd_sc_hd__a22o_1 _4901_ (.A1(\gpio_configure[18][0] ),
    .A2(_0934_),
    .B1(_0857_),
    .B2(\gpio_configure[3][0] ),
    .X(_1367_));
 sky130_fd_sc_hd__a221o_1 _4902_ (.A1(\gpio_configure[8][0] ),
    .A2(_0973_),
    .B1(_1151_),
    .B2(\gpio_configure[11][8] ),
    .C1(_1367_),
    .X(_1368_));
 sky130_fd_sc_hd__a22o_1 _4903_ (.A1(\gpio_configure[31][8] ),
    .A2(_1145_),
    .B1(_1091_),
    .B2(\gpio_configure[26][8] ),
    .X(_1369_));
 sky130_fd_sc_hd__a221o_1 _4904_ (.A1(net123),
    .A2(_0963_),
    .B1(net380),
    .B2(\gpio_configure[25][0] ),
    .C1(_1369_),
    .X(_1370_));
 sky130_fd_sc_hd__a22o_1 _4905_ (.A1(\gpio_configure[17][8] ),
    .A2(_1076_),
    .B1(_1134_),
    .B2(\gpio_configure[2][8] ),
    .X(_1371_));
 sky130_fd_sc_hd__a221o_1 _4906_ (.A1(\gpio_configure[31][0] ),
    .A2(net389),
    .B1(_1096_),
    .B2(\gpio_configure[6][8] ),
    .C1(_1371_),
    .X(_1372_));
 sky130_fd_sc_hd__a22o_1 _4907_ (.A1(\gpio_configure[16][0] ),
    .A2(_0872_),
    .B1(_1104_),
    .B2(\gpio_configure[14][8] ),
    .X(_1373_));
 sky130_fd_sc_hd__a221o_1 _4908_ (.A1(net316),
    .A2(_0851_),
    .B1(_1148_),
    .B2(\gpio_configure[16][8] ),
    .C1(_1373_),
    .X(_1374_));
 sky130_fd_sc_hd__or4_1 _4909_ (.A(_1368_),
    .B(_1370_),
    .C(_1372_),
    .D(_1374_),
    .X(_1375_));
 sky130_fd_sc_hd__a22o_1 _4910_ (.A1(\gpio_configure[2][0] ),
    .A2(net385),
    .B1(_1115_),
    .B2(\gpio_configure[22][8] ),
    .X(_1376_));
 sky130_fd_sc_hd__a221o_1 _4911_ (.A1(\gpio_configure[27][0] ),
    .A2(_0959_),
    .B1(_1028_),
    .B2(net271),
    .C1(_1376_),
    .X(_1377_));
 sky130_fd_sc_hd__a22o_1 _4912_ (.A1(\gpio_configure[35][0] ),
    .A2(net379),
    .B1(net381),
    .B2(\gpio_configure[28][0] ),
    .X(_1378_));
 sky130_fd_sc_hd__a221o_1 _4913_ (.A1(net71),
    .A2(_0910_),
    .B1(_1077_),
    .B2(\gpio_configure[27][8] ),
    .C1(_1378_),
    .X(_1379_));
 sky130_fd_sc_hd__or3_1 _4914_ (.A(\hkspi.pass_thru_mgmt_delay ),
    .B(\hkspi.pre_pass_thru_mgmt ),
    .C(reset_reg),
    .X(_1380_));
 sky130_fd_sc_hd__clkbuf_2 _4915_ (.A(_1380_),
    .X(net304));
 sky130_fd_sc_hd__nor2_1 _4916_ (.A(_0964_),
    .B(_0974_),
    .Y(_1381_));
 sky130_fd_sc_hd__a22o_1 _4917_ (.A1(\gpio_configure[7][0] ),
    .A2(net377),
    .B1(net304),
    .B2(_1381_),
    .X(_1382_));
 sky130_fd_sc_hd__a221o_1 _4918_ (.A1(net100),
    .A2(_0977_),
    .B1(_1325_),
    .B2(net325),
    .C1(_1382_),
    .X(_1383_));
 sky130_fd_sc_hd__a22o_1 _4919_ (.A1(\gpio_configure[36][0] ),
    .A2(_0942_),
    .B1(_0941_),
    .B2(net274),
    .X(_1384_));
 sky130_fd_sc_hd__a221o_1 _4920_ (.A1(\gpio_configure[6][0] ),
    .A2(_0903_),
    .B1(_1130_),
    .B2(\gpio_configure[0][8] ),
    .C1(_1384_),
    .X(_1385_));
 sky130_fd_sc_hd__or4_1 _4921_ (.A(_1377_),
    .B(_1379_),
    .C(_1383_),
    .D(_1385_),
    .X(_1386_));
 sky130_fd_sc_hd__or4_1 _4922_ (.A(_1362_),
    .B(_1366_),
    .C(_1375_),
    .D(_1386_),
    .X(_1387_));
 sky130_fd_sc_hd__a22o_1 _4923_ (.A1(\gpio_configure[37][8] ),
    .A2(_1131_),
    .B1(_1092_),
    .B2(\gpio_configure[23][8] ),
    .X(_1388_));
 sky130_fd_sc_hd__a221o_1 _4924_ (.A1(net298),
    .A2(_0972_),
    .B1(_1140_),
    .B2(net265),
    .C1(_1388_),
    .X(_1389_));
 sky130_fd_sc_hd__a22o_1 _4925_ (.A1(\gpio_configure[21][0] ),
    .A2(_0902_),
    .B1(_1066_),
    .B2(\gpio_configure[9][8] ),
    .X(_1390_));
 sky130_fd_sc_hd__a221o_1 _4926_ (.A1(net4),
    .A2(_0952_),
    .B1(_1095_),
    .B2(\gpio_configure[33][8] ),
    .C1(_1390_),
    .X(_1391_));
 sky130_fd_sc_hd__a22o_1 _4927_ (.A1(\gpio_configure[5][0] ),
    .A2(_0929_),
    .B1(net376),
    .B2(\gpio_configure[17][0] ),
    .X(_1392_));
 sky130_fd_sc_hd__a221o_1 _4928_ (.A1(\gpio_configure[28][8] ),
    .A2(_1105_),
    .B1(_1217_),
    .B2(net300),
    .C1(_1392_),
    .X(_1393_));
 sky130_fd_sc_hd__a22o_1 _4929_ (.A1(\gpio_configure[24][0] ),
    .A2(_0890_),
    .B1(_1110_),
    .B2(\gpio_configure[4][8] ),
    .X(_1394_));
 sky130_fd_sc_hd__a221o_1 _4930_ (.A1(net93),
    .A2(_0919_),
    .B1(_0976_),
    .B2(\gpio_configure[13][0] ),
    .C1(_1394_),
    .X(_1395_));
 sky130_fd_sc_hd__or4_1 _4931_ (.A(_1389_),
    .B(_1391_),
    .C(_1393_),
    .D(_1395_),
    .X(_1396_));
 sky130_fd_sc_hd__a22o_1 _4932_ (.A1(\gpio_configure[12][8] ),
    .A2(_1084_),
    .B1(_1065_),
    .B2(\gpio_configure[30][8] ),
    .X(_1397_));
 sky130_fd_sc_hd__a221o_1 _4933_ (.A1(\gpio_configure[10][8] ),
    .A2(_1121_),
    .B1(_1226_),
    .B2(trap_output_dest),
    .C1(_1397_),
    .X(_1398_));
 sky130_fd_sc_hd__a211o_2 _4934_ (.A1(\gpio_configure[12][0] ),
    .A2(net387),
    .B1(_1120_),
    .C1(_1398_),
    .X(_1399_));
 sky130_fd_sc_hd__a22o_1 _4935_ (.A1(\gpio_configure[19][8] ),
    .A2(_1144_),
    .B1(_1088_),
    .B2(\gpio_configure[20][8] ),
    .X(_1400_));
 sky130_fd_sc_hd__a221o_1 _4936_ (.A1(net281),
    .A2(_0946_),
    .B1(_1136_),
    .B2(\gpio_configure[7][8] ),
    .C1(_1400_),
    .X(_1401_));
 sky130_fd_sc_hd__a22o_1 _4937_ (.A1(\gpio_configure[32][0] ),
    .A2(_0898_),
    .B1(_0889_),
    .B2(\gpio_configure[19][0] ),
    .X(_1402_));
 sky130_fd_sc_hd__a221o_1 _4938_ (.A1(\gpio_configure[11][0] ),
    .A2(net378),
    .B1(net364),
    .B2(\gpio_configure[34][0] ),
    .C1(_1402_),
    .X(_1403_));
 sky130_fd_sc_hd__or4_1 _4939_ (.A(_1396_),
    .B(_1399_),
    .C(_1401_),
    .D(_1403_),
    .X(_1404_));
 sky130_fd_sc_hd__a22o_1 _4940_ (.A1(\gpio_configure[33][0] ),
    .A2(_0957_),
    .B1(_0881_),
    .B2(net34),
    .X(_1405_));
 sky130_fd_sc_hd__a221o_1 _4941_ (.A1(net36),
    .A2(_0954_),
    .B1(_1203_),
    .B2(net130),
    .C1(_1405_),
    .X(_1406_));
 sky130_fd_sc_hd__a22o_1 _4942_ (.A1(\gpio_configure[23][0] ),
    .A2(net373),
    .B1(_1111_),
    .B2(\gpio_configure[3][8] ),
    .X(_1407_));
 sky130_fd_sc_hd__a221o_1 _4943_ (.A1(net43),
    .A2(_0965_),
    .B1(_1155_),
    .B2(\gpio_configure[36][8] ),
    .C1(_1407_),
    .X(_1408_));
 sky130_fd_sc_hd__nor2_1 _4944_ (.A(_0893_),
    .B(_0974_),
    .Y(_1409_));
 sky130_fd_sc_hd__a22o_1 _4945_ (.A1(net20),
    .A2(_0935_),
    .B1(_1409_),
    .B2(net204),
    .X(_1410_));
 sky130_fd_sc_hd__a221o_1 _4946_ (.A1(net11),
    .A2(_0975_),
    .B1(_1011_),
    .B2(serial_busy),
    .C1(_1410_),
    .X(_1411_));
 sky130_fd_sc_hd__a22o_1 _4947_ (.A1(net52),
    .A2(net372),
    .B1(_1135_),
    .B2(\gpio_configure[18][8] ),
    .X(_1412_));
 sky130_fd_sc_hd__a221o_2 _4948_ (.A1(\gpio_configure[9][0] ),
    .A2(net366),
    .B1(net370),
    .B2(net61),
    .C1(_1412_),
    .X(_1413_));
 sky130_fd_sc_hd__or4_1 _4949_ (.A(_1406_),
    .B(_1408_),
    .C(_1411_),
    .D(_1413_),
    .X(_1414_));
 sky130_fd_sc_hd__a22o_1 _4950_ (.A1(\gpio_configure[25][8] ),
    .A2(_1078_),
    .B1(_1116_),
    .B2(\gpio_configure[8][8] ),
    .X(_1415_));
 sky130_fd_sc_hd__a221o_1 _4951_ (.A1(\gpio_configure[20][0] ),
    .A2(net360),
    .B1(_0958_),
    .B2(net109),
    .C1(_1415_),
    .X(_1416_));
 sky130_fd_sc_hd__a22o_1 _4952_ (.A1(net290),
    .A2(_1328_),
    .B1(_1345_),
    .B2(net270),
    .X(_1417_));
 sky130_fd_sc_hd__a221o_1 _4953_ (.A1(\gpio_configure[26][0] ),
    .A2(_0864_),
    .B1(_1129_),
    .B2(\gpio_configure[35][8] ),
    .C1(_1417_),
    .X(_1418_));
 sky130_fd_sc_hd__a22o_1 _4954_ (.A1(\gpio_configure[29][0] ),
    .A2(_0914_),
    .B1(_1081_),
    .B2(\gpio_configure[32][8] ),
    .X(_1419_));
 sky130_fd_sc_hd__a221o_1 _4955_ (.A1(\gpio_configure[4][0] ),
    .A2(_0967_),
    .B1(_0971_),
    .B2(\gpio_configure[0][0] ),
    .C1(_1419_),
    .X(_1420_));
 sky130_fd_sc_hd__nor2_1 _4956_ (.A(_0918_),
    .B(_0974_),
    .Y(_1421_));
 sky130_fd_sc_hd__a22o_1 _4957_ (.A1(\gpio_configure[34][8] ),
    .A2(_1154_),
    .B1(_1421_),
    .B2(net263),
    .X(_1422_));
 sky130_fd_sc_hd__a221o_1 _4958_ (.A1(\gpio_configure[15][0] ),
    .A2(_0876_),
    .B1(_1073_),
    .B2(\gpio_configure[1][8] ),
    .C1(_1422_),
    .X(_1423_));
 sky130_fd_sc_hd__or2_1 _4959_ (.A(_1420_),
    .B(_1423_),
    .X(_1424_));
 sky130_fd_sc_hd__or4_1 _4960_ (.A(_1414_),
    .B(_1416_),
    .C(_1418_),
    .D(_1424_),
    .X(_1425_));
 sky130_fd_sc_hd__or3_4 _4961_ (.A(_1387_),
    .B(_1404_),
    .C(_1425_),
    .X(_1426_));
 sky130_fd_sc_hd__buf_2 _4962_ (.A(\hkspi.count[0] ),
    .X(_1427_));
 sky130_fd_sc_hd__or3_1 _4963_ (.A(\hkspi.count[2] ),
    .B(\hkspi.count[1] ),
    .C(_1427_),
    .X(_1428_));
 sky130_fd_sc_hd__nor2_1 _4964_ (.A(_1428_),
    .B(_0985_),
    .Y(_1429_));
 sky130_fd_sc_hd__a22o_1 _4965_ (.A1(net1449),
    .A2(_0985_),
    .B1(_1426_),
    .B2(_1429_),
    .X(_0384_));
 sky130_fd_sc_hd__buf_2 _4966_ (.A(\hkspi.state[3] ),
    .X(_1430_));
 sky130_fd_sc_hd__or3_2 _4967_ (.A(\hkspi.state[0] ),
    .B(_1430_),
    .C(\hkspi.state[2] ),
    .X(_1431_));
 sky130_fd_sc_hd__and3_1 _4968_ (.A(\hkspi.count[1] ),
    .B(_1427_),
    .C(_1431_),
    .X(_1432_));
 sky130_fd_sc_hd__xor2_1 _4969_ (.A(net1509),
    .B(_1432_),
    .X(_0100_));
 sky130_fd_sc_hd__a21oi_1 _4970_ (.A1(_1427_),
    .A2(_1431_),
    .B1(net1528),
    .Y(_1433_));
 sky130_fd_sc_hd__nor2_1 _4971_ (.A(_1432_),
    .B(_1433_),
    .Y(_0099_));
 sky130_fd_sc_hd__xor2_1 _4972_ (.A(_1427_),
    .B(_1431_),
    .X(_0098_));
 sky130_fd_sc_hd__clkinv_2 _4973_ (.A(\hkspi.state[0] ),
    .Y(_1434_));
 sky130_fd_sc_hd__and3_1 _4974_ (.A(\hkspi.count[2] ),
    .B(\hkspi.count[1] ),
    .C(\hkspi.count[0] ),
    .X(_1435_));
 sky130_fd_sc_hd__clkbuf_2 _4975_ (.A(_1435_),
    .X(_1436_));
 sky130_fd_sc_hd__nor2_1 _4976_ (.A(\hkspi.fixed[2] ),
    .B(\hkspi.fixed[1] ),
    .Y(_1437_));
 sky130_fd_sc_hd__nand2_1 _4977_ (.A(\hkspi.fixed[0] ),
    .B(_1437_),
    .Y(_1438_));
 sky130_fd_sc_hd__a31o_1 _4978_ (.A1(\hkspi.state[2] ),
    .A2(_1436_),
    .A3(_1438_),
    .B1(_1430_),
    .X(_1439_));
 sky130_fd_sc_hd__nand2_4 _4979_ (.A(_1434_),
    .B(_1439_),
    .Y(_1440_));
 sky130_fd_sc_hd__and3_1 _4980_ (.A(\hkspi.addr[2] ),
    .B(\hkspi.addr[1] ),
    .C(\hkspi.addr[0] ),
    .X(_1441_));
 sky130_fd_sc_hd__and2_1 _4981_ (.A(\hkspi.addr[3] ),
    .B(_1441_),
    .X(_1442_));
 sky130_fd_sc_hd__nand4_1 _4982_ (.A(\hkspi.addr[6] ),
    .B(\hkspi.addr[5] ),
    .C(\hkspi.addr[4] ),
    .D(_1442_),
    .Y(_1443_));
 sky130_fd_sc_hd__mux2_1 _4983_ (.A0(_0826_),
    .A1(_0827_),
    .S(_1443_),
    .X(_1444_));
 sky130_fd_sc_hd__nor2_1 _4984_ (.A(_1440_),
    .B(_1444_),
    .Y(_1445_));
 sky130_fd_sc_hd__a21o_1 _4985_ (.A1(net1450),
    .A2(_1440_),
    .B1(_1445_),
    .X(_0097_));
 sky130_fd_sc_hd__a31o_1 _4986_ (.A1(\hkspi.addr[5] ),
    .A2(\hkspi.addr[4] ),
    .A3(_1442_),
    .B1(\hkspi.addr[6] ),
    .X(_1446_));
 sky130_fd_sc_hd__a31o_1 _4987_ (.A1(_0825_),
    .A2(_1443_),
    .A3(_1446_),
    .B1(_0828_),
    .X(_1447_));
 sky130_fd_sc_hd__mux2_1 _4988_ (.A0(_1447_),
    .A1(\hkspi.addr[6] ),
    .S(_1440_),
    .X(_1448_));
 sky130_fd_sc_hd__clkbuf_1 _4989_ (.A(_1448_),
    .X(_0096_));
 sky130_fd_sc_hd__o21a_1 _4990_ (.A1(_1430_),
    .A2(_1442_),
    .B1(\hkspi.addr[4] ),
    .X(_1449_));
 sky130_fd_sc_hd__xnor2_1 _4991_ (.A(_0832_),
    .B(_1449_),
    .Y(_1450_));
 sky130_fd_sc_hd__mux2_1 _4992_ (.A0(_1450_),
    .A1(\hkspi.addr[5] ),
    .S(_1440_),
    .X(_1451_));
 sky130_fd_sc_hd__clkbuf_1 _4993_ (.A(_1451_),
    .X(_0095_));
 sky130_fd_sc_hd__mux2_1 _4994_ (.A0(_0836_),
    .A1(_0835_),
    .S(_1442_),
    .X(_1452_));
 sky130_fd_sc_hd__mux2_1 _4995_ (.A0(_1452_),
    .A1(\hkspi.addr[4] ),
    .S(_1440_),
    .X(_1453_));
 sky130_fd_sc_hd__clkbuf_1 _4996_ (.A(_1453_),
    .X(_0094_));
 sky130_fd_sc_hd__nor2_1 _4997_ (.A(_1430_),
    .B(_1442_),
    .Y(_1454_));
 sky130_fd_sc_hd__or2_1 _4998_ (.A(\hkspi.addr[3] ),
    .B(_1441_),
    .X(_1455_));
 sky130_fd_sc_hd__a22o_1 _4999_ (.A1(\hkspi.addr[2] ),
    .A2(_1430_),
    .B1(_1454_),
    .B2(_1455_),
    .X(_1456_));
 sky130_fd_sc_hd__mux2_1 _5000_ (.A0(_1456_),
    .A1(net1561),
    .S(_1440_),
    .X(_1457_));
 sky130_fd_sc_hd__clkbuf_1 _5001_ (.A(_1457_),
    .X(_0093_));
 sky130_fd_sc_hd__nor2_1 _5002_ (.A(_1430_),
    .B(_1441_),
    .Y(_1458_));
 sky130_fd_sc_hd__a21o_1 _5003_ (.A1(\hkspi.addr[1] ),
    .A2(\hkspi.addr[0] ),
    .B1(\hkspi.addr[2] ),
    .X(_1459_));
 sky130_fd_sc_hd__a22o_1 _5004_ (.A1(\hkspi.addr[1] ),
    .A2(_1430_),
    .B1(_1458_),
    .B2(_1459_),
    .X(_1460_));
 sky130_fd_sc_hd__mux2_1 _5005_ (.A0(_1460_),
    .A1(\hkspi.addr[2] ),
    .S(_1440_),
    .X(_1461_));
 sky130_fd_sc_hd__clkbuf_1 _5006_ (.A(_1461_),
    .X(_0092_));
 sky130_fd_sc_hd__buf_2 _5007_ (.A(\hkspi.state[0] ),
    .X(_1462_));
 sky130_fd_sc_hd__o21ai_1 _5008_ (.A1(_1462_),
    .A2(_0825_),
    .B1(\hkspi.addr[1] ),
    .Y(_1463_));
 sky130_fd_sc_hd__inv_2 _5009_ (.A(net1562),
    .Y(_1464_));
 sky130_fd_sc_hd__nor2_1 _5010_ (.A(_1464_),
    .B(_1440_),
    .Y(_1465_));
 sky130_fd_sc_hd__xnor2_1 _5011_ (.A(_1463_),
    .B(_1465_),
    .Y(_0091_));
 sky130_fd_sc_hd__buf_8 _5012_ (.A(net58),
    .X(_1466_));
 sky130_fd_sc_hd__mux2_1 _5013_ (.A0(_1464_),
    .A1(_1466_),
    .S(_1430_),
    .X(_1467_));
 sky130_fd_sc_hd__mux2_1 _5014_ (.A0(_1467_),
    .A1(\hkspi.addr[0] ),
    .S(_1440_),
    .X(_1468_));
 sky130_fd_sc_hd__clkbuf_1 _5015_ (.A(_1468_),
    .X(_0090_));
 sky130_fd_sc_hd__nand2_1 _5016_ (.A(_1462_),
    .B(_1436_),
    .Y(_1469_));
 sky130_fd_sc_hd__mux2_1 _5017_ (.A0(net1500),
    .A1(\hkspi.pass_thru_user_delay ),
    .S(_1469_),
    .X(_1470_));
 sky130_fd_sc_hd__clkbuf_1 _5018_ (.A(_1470_),
    .X(_0089_));
 sky130_fd_sc_hd__inv_2 _5019_ (.A(net1457),
    .Y(_1471_));
 sky130_fd_sc_hd__inv_2 _5020_ (.A(\hkspi.state[2] ),
    .Y(_1472_));
 sky130_fd_sc_hd__and3_1 _5021_ (.A(_1434_),
    .B(_0825_),
    .C(_1472_),
    .X(_1473_));
 sky130_fd_sc_hd__a31o_1 _5022_ (.A1(net1455),
    .A2(_1471_),
    .A3(_1473_),
    .B1(\hkspi.pass_thru_user ),
    .X(_0088_));
 sky130_fd_sc_hd__and2_1 _5023_ (.A(\hkspi.count[2] ),
    .B(\hkspi.count[1] ),
    .X(_1474_));
 sky130_fd_sc_hd__nand2_1 _5024_ (.A(_1462_),
    .B(_1474_),
    .Y(_1475_));
 sky130_fd_sc_hd__nor2_1 _5025_ (.A(_1427_),
    .B(_1475_),
    .Y(_1476_));
 sky130_fd_sc_hd__mux2_1 _5026_ (.A0(\hkspi.pass_thru_mgmt_delay ),
    .A1(net1505),
    .S(_1476_),
    .X(_1477_));
 sky130_fd_sc_hd__clkbuf_1 _5027_ (.A(_1477_),
    .X(_0087_));
 sky130_fd_sc_hd__a21o_1 _5028_ (.A1(net1457),
    .A2(_1473_),
    .B1(\hkspi.pass_thru_mgmt ),
    .X(_0086_));
 sky130_fd_sc_hd__a21oi_1 _5029_ (.A1(\hkspi.readmode ),
    .A2(_1431_),
    .B1(net1530),
    .Y(_1478_));
 sky130_fd_sc_hd__a21oi_1 _5030_ (.A1(_1434_),
    .A2(_1436_),
    .B1(_1473_),
    .Y(_1479_));
 sky130_fd_sc_hd__nor2_1 _5031_ (.A(_1478_),
    .B(_1479_),
    .Y(_0085_));
 sky130_fd_sc_hd__o21a_1 _5032_ (.A1(_1434_),
    .A2(_1428_),
    .B1(net1518),
    .X(_1480_));
 sky130_fd_sc_hd__a31o_1 _5033_ (.A1(_1466_),
    .A2(_1462_),
    .A3(_0983_),
    .B1(_1480_),
    .X(_0084_));
 sky130_fd_sc_hd__inv_2 _5034_ (.A(\hkspi.count[1] ),
    .Y(_1481_));
 sky130_fd_sc_hd__and4b_1 _5035_ (.A_N(\hkspi.count[2] ),
    .B(_1481_),
    .C(_1427_),
    .D(\hkspi.state[0] ),
    .X(_1482_));
 sky130_fd_sc_hd__mux2_1 _5036_ (.A0(\hkspi.readmode ),
    .A1(_1466_),
    .S(_1482_),
    .X(_1483_));
 sky130_fd_sc_hd__clkbuf_1 _5037_ (.A(_1483_),
    .X(_0083_));
 sky130_fd_sc_hd__a2111oi_2 _5038_ (.A1(_1481_),
    .A2(\hkspi.count[0] ),
    .B1(_1434_),
    .C1(_0983_),
    .D1(_1474_),
    .Y(_1484_));
 sky130_fd_sc_hd__nand2_1 _5039_ (.A(_1427_),
    .B(_1474_),
    .Y(_1485_));
 sky130_fd_sc_hd__or3_1 _5040_ (.A(\hkspi.state[0] ),
    .B(_1430_),
    .C(_1472_),
    .X(_1486_));
 sky130_fd_sc_hd__buf_6 _5041_ (.A(_1486_),
    .X(_1487_));
 sky130_fd_sc_hd__inv_2 _5042_ (.A(_1484_),
    .Y(_1488_));
 sky130_fd_sc_hd__o31a_1 _5043_ (.A1(_1485_),
    .A2(_1437_),
    .A3(_1487_),
    .B1(_1488_),
    .X(_1489_));
 sky130_fd_sc_hd__nor2_1 _5044_ (.A(\hkspi.fixed[0] ),
    .B(_1489_),
    .Y(_1490_));
 sky130_fd_sc_hd__nor2_1 _5045_ (.A(net401),
    .B(_1490_),
    .Y(_1491_));
 sky130_fd_sc_hd__o22a_1 _5046_ (.A1(\hkspi.fixed[2] ),
    .A2(net401),
    .B1(_1491_),
    .B2(net1471),
    .X(_0082_));
 sky130_fd_sc_hd__inv_2 _5047_ (.A(net1471),
    .Y(_1492_));
 sky130_fd_sc_hd__o21a_1 _5048_ (.A1(net1471),
    .A2(net401),
    .B1(_1490_),
    .X(_1493_));
 sky130_fd_sc_hd__a21oi_1 _5049_ (.A1(_1492_),
    .A2(_1491_),
    .B1(_1493_),
    .Y(_0081_));
 sky130_fd_sc_hd__and2_1 _5050_ (.A(net1506),
    .B(_1489_),
    .X(_1494_));
 sky130_fd_sc_hd__and3_1 _5051_ (.A(_1466_),
    .B(_1462_),
    .C(_1484_),
    .X(_1495_));
 sky130_fd_sc_hd__a211o_1 _5052_ (.A1(_1434_),
    .A2(_1490_),
    .B1(_1494_),
    .C1(_1495_),
    .X(_0080_));
 sky130_fd_sc_hd__mux2_1 _5053_ (.A0(net1534),
    .A1(net510),
    .S(_1487_),
    .X(_1496_));
 sky130_fd_sc_hd__clkbuf_1 _5054_ (.A(_1496_),
    .X(_0079_));
 sky130_fd_sc_hd__mux2_1 _5055_ (.A0(net1556),
    .A1(net1534),
    .S(_1487_),
    .X(_1497_));
 sky130_fd_sc_hd__clkbuf_1 _5056_ (.A(_1497_),
    .X(_0078_));
 sky130_fd_sc_hd__mux2_1 _5057_ (.A0(net1536),
    .A1(net1556),
    .S(_1487_),
    .X(_1498_));
 sky130_fd_sc_hd__clkbuf_1 _5058_ (.A(_1498_),
    .X(_0077_));
 sky130_fd_sc_hd__mux2_1 _5059_ (.A0(net550),
    .A1(net1536),
    .S(_1487_),
    .X(_1499_));
 sky130_fd_sc_hd__clkbuf_1 _5060_ (.A(_1499_),
    .X(_0076_));
 sky130_fd_sc_hd__mux2_1 _5061_ (.A0(net517),
    .A1(net550),
    .S(_1487_),
    .X(_1500_));
 sky130_fd_sc_hd__clkbuf_1 _5062_ (.A(_1500_),
    .X(_0075_));
 sky130_fd_sc_hd__mux2_1 _5063_ (.A0(net1535),
    .A1(net517),
    .S(_1487_),
    .X(_1501_));
 sky130_fd_sc_hd__clkbuf_1 _5064_ (.A(_1501_),
    .X(_0074_));
 sky130_fd_sc_hd__mux2_1 _5065_ (.A0(_1466_),
    .A1(net1535),
    .S(_1487_),
    .X(_1502_));
 sky130_fd_sc_hd__clkbuf_1 _5066_ (.A(_1502_),
    .X(_0073_));
 sky130_fd_sc_hd__and3_1 _5067_ (.A(\hkspi.count[2] ),
    .B(_1466_),
    .C(_1462_),
    .X(_1503_));
 sky130_fd_sc_hd__nand3_1 _5068_ (.A(\hkspi.count[2] ),
    .B(_1427_),
    .C(_1462_),
    .Y(_1504_));
 sky130_fd_sc_hd__a32o_1 _5069_ (.A1(_1481_),
    .A2(_1427_),
    .A3(_1503_),
    .B1(_1504_),
    .B2(net1505),
    .X(_0072_));
 sky130_fd_sc_hd__clkbuf_8 _5070_ (.A(net417),
    .X(_1505_));
 sky130_fd_sc_hd__nor3_1 _5071_ (.A(\gpio_configure[3][3] ),
    .B(hkspi_disable),
    .C(net67),
    .Y(_1506_));
 sky130_fd_sc_hd__buf_4 _5072_ (.A(_1506_),
    .X(_1507_));
 sky130_fd_sc_hd__buf_2 _5073_ (.A(_1507_),
    .X(_1508_));
 sky130_fd_sc_hd__buf_4 _5074_ (.A(_1508_),
    .X(_1509_));
 sky130_fd_sc_hd__and2_1 _5075_ (.A(_1505_),
    .B(_1509_),
    .X(_1510_));
 sky130_fd_sc_hd__clkbuf_1 _5076_ (.A(_1510_),
    .X(_0021_));
 sky130_fd_sc_hd__a21o_1 _5077_ (.A1(_1427_),
    .A2(\hkspi.pre_pass_thru_mgmt ),
    .B1(_1475_),
    .X(_1511_));
 sky130_fd_sc_hd__a22o_1 _5078_ (.A1(_1466_),
    .A2(_1476_),
    .B1(_1511_),
    .B2(net1500),
    .X(_0071_));
 sky130_fd_sc_hd__o211a_1 _5079_ (.A1(\hkspi.writemode ),
    .A2(net523),
    .B1(\hkspi.state[2] ),
    .C1(_1436_),
    .X(_0070_));
 sky130_fd_sc_hd__inv_2 _5080_ (.A(\gpio_configure[34][3] ),
    .Y(_4347_));
 sky130_fd_sc_hd__inv_2 _5081_ (.A(\gpio_configure[33][3] ),
    .Y(_4346_));
 sky130_fd_sc_hd__inv_2 _5082_ (.A(\gpio_configure[32][3] ),
    .Y(_4345_));
 sky130_fd_sc_hd__inv_2 _5083_ (.A(\gpio_configure[31][3] ),
    .Y(_4344_));
 sky130_fd_sc_hd__inv_2 _5084_ (.A(\gpio_configure[30][3] ),
    .Y(_4343_));
 sky130_fd_sc_hd__inv_2 _5085_ (.A(\gpio_configure[29][3] ),
    .Y(_4342_));
 sky130_fd_sc_hd__inv_2 _5086_ (.A(\gpio_configure[28][3] ),
    .Y(_4341_));
 sky130_fd_sc_hd__inv_2 _5087_ (.A(\gpio_configure[27][3] ),
    .Y(_4340_));
 sky130_fd_sc_hd__inv_2 _5088_ (.A(\gpio_configure[26][3] ),
    .Y(_4339_));
 sky130_fd_sc_hd__inv_2 _5089_ (.A(\gpio_configure[25][3] ),
    .Y(_4338_));
 sky130_fd_sc_hd__inv_2 _5090_ (.A(\gpio_configure[24][3] ),
    .Y(_4337_));
 sky130_fd_sc_hd__inv_2 _5091_ (.A(\gpio_configure[23][3] ),
    .Y(_4336_));
 sky130_fd_sc_hd__inv_2 _5092_ (.A(\gpio_configure[22][3] ),
    .Y(_4335_));
 sky130_fd_sc_hd__inv_2 _5093_ (.A(\gpio_configure[21][3] ),
    .Y(_4334_));
 sky130_fd_sc_hd__inv_2 _5094_ (.A(\gpio_configure[20][3] ),
    .Y(_4333_));
 sky130_fd_sc_hd__inv_2 _5095_ (.A(\gpio_configure[19][3] ),
    .Y(_4332_));
 sky130_fd_sc_hd__inv_2 _5096_ (.A(\gpio_configure[18][3] ),
    .Y(_4331_));
 sky130_fd_sc_hd__inv_2 _5097_ (.A(\gpio_configure[17][3] ),
    .Y(_4330_));
 sky130_fd_sc_hd__inv_2 _5098_ (.A(\gpio_configure[16][3] ),
    .Y(_4329_));
 sky130_fd_sc_hd__inv_2 _5099_ (.A(\gpio_configure[15][3] ),
    .Y(_4328_));
 sky130_fd_sc_hd__inv_2 _5100_ (.A(\gpio_configure[14][3] ),
    .Y(_4327_));
 sky130_fd_sc_hd__inv_2 _5101_ (.A(\gpio_configure[13][3] ),
    .Y(_4326_));
 sky130_fd_sc_hd__inv_2 _5102_ (.A(\gpio_configure[12][3] ),
    .Y(_4325_));
 sky130_fd_sc_hd__inv_2 _5103_ (.A(\gpio_configure[11][3] ),
    .Y(_4324_));
 sky130_fd_sc_hd__inv_2 _5104_ (.A(\gpio_configure[10][3] ),
    .Y(_4323_));
 sky130_fd_sc_hd__inv_2 _5105_ (.A(\gpio_configure[9][3] ),
    .Y(_4322_));
 sky130_fd_sc_hd__inv_2 _5106_ (.A(\gpio_configure[8][3] ),
    .Y(_4321_));
 sky130_fd_sc_hd__inv_2 _5107_ (.A(\gpio_configure[7][3] ),
    .Y(_4320_));
 sky130_fd_sc_hd__inv_2 _5108_ (.A(\gpio_configure[6][3] ),
    .Y(_4319_));
 sky130_fd_sc_hd__inv_2 _5109_ (.A(\gpio_configure[5][3] ),
    .Y(_4318_));
 sky130_fd_sc_hd__inv_2 _5110_ (.A(\gpio_configure[4][3] ),
    .Y(_4317_));
 sky130_fd_sc_hd__inv_2 _5111_ (.A(\gpio_configure[3][3] ),
    .Y(_4316_));
 sky130_fd_sc_hd__inv_2 _5112_ (.A(\gpio_configure[2][3] ),
    .Y(_4315_));
 sky130_fd_sc_hd__mux2_1 _5113_ (.A0(serial_clock_pre),
    .A1(serial_bb_clock),
    .S(serial_bb_enable),
    .X(_1512_));
 sky130_fd_sc_hd__clkbuf_2 _5114_ (.A(_1512_),
    .X(net306));
 sky130_fd_sc_hd__o21a_4 _5115_ (.A1(\hkspi.rdstb ),
    .A2(\hkspi.wrstb ),
    .B1(_1508_),
    .X(_1513_));
 sky130_fd_sc_hd__or2_1 _5116_ (.A(net162),
    .B(net161),
    .X(_1514_));
 sky130_fd_sc_hd__or4_1 _5117_ (.A(net133),
    .B(net132),
    .C(net135),
    .D(net134),
    .X(_1515_));
 sky130_fd_sc_hd__or4b_1 _5118_ (.A(net141),
    .B(net140),
    .C(net147),
    .D_N(net148),
    .X(_1516_));
 sky130_fd_sc_hd__or4_1 _5119_ (.A(net137),
    .B(net136),
    .C(net139),
    .D(net138),
    .X(_1517_));
 sky130_fd_sc_hd__or4_1 _5120_ (.A(_1514_),
    .B(_1515_),
    .C(_1516_),
    .D(_1517_),
    .X(_1518_));
 sky130_fd_sc_hd__buf_4 _5121_ (.A(net143),
    .X(_1519_));
 sky130_fd_sc_hd__a211o_2 _5122_ (.A1(net144),
    .A2(_1519_),
    .B1(net146),
    .C1(net145),
    .X(_1520_));
 sky130_fd_sc_hd__and4bb_1 _5123_ (.A_N(net155),
    .B_N(net154),
    .C(net163),
    .D(net201),
    .X(_1521_));
 sky130_fd_sc_hd__and4bb_1 _5124_ (.A_N(net150),
    .B_N(net151),
    .C(net152),
    .D(net149),
    .X(_1522_));
 sky130_fd_sc_hd__and4bb_2 _5125_ (.A_N(_1518_),
    .B_N(_1520_),
    .C(_1521_),
    .D(_1522_),
    .X(_1523_));
 sky130_fd_sc_hd__a22o_1 _5126_ (.A1(net1555),
    .A2(_1513_),
    .B1(_1523_),
    .B2(net1502),
    .X(_0010_));
 sky130_fd_sc_hd__nor2_1 _5127_ (.A(_1485_),
    .B(_1438_),
    .Y(_1524_));
 sky130_fd_sc_hd__a22o_1 _5128_ (.A1(_1462_),
    .A2(_1485_),
    .B1(_1524_),
    .B2(net1514),
    .X(_0004_));
 sky130_fd_sc_hd__clkbuf_4 _5129_ (.A(\xfer_state[1] ),
    .X(_1525_));
 sky130_fd_sc_hd__clkbuf_4 _5130_ (.A(_1525_),
    .X(_1526_));
 sky130_fd_sc_hd__nand2b_4 _5131_ (.A_N(\pad_count_2[4] ),
    .B(\pad_count_2[5] ),
    .Y(_1527_));
 sky130_fd_sc_hd__nor2b_2 _5132_ (.A(\pad_count_2[0] ),
    .B_N(\pad_count_2[1] ),
    .Y(_1528_));
 sky130_fd_sc_hd__nor2b_2 _5133_ (.A(\pad_count_2[3] ),
    .B_N(\pad_count_2[2] ),
    .Y(_1529_));
 sky130_fd_sc_hd__nand2_2 _5134_ (.A(_1528_),
    .B(_1529_),
    .Y(_1530_));
 sky130_fd_sc_hd__or2_2 _5135_ (.A(_1527_),
    .B(_1530_),
    .X(_1531_));
 sky130_fd_sc_hd__nor2_1 _5136_ (.A(\xfer_count[0] ),
    .B(\xfer_count[1] ),
    .Y(_1532_));
 sky130_fd_sc_hd__and4b_1 _5137_ (.A_N(net306),
    .B(_1532_),
    .C(\xfer_count[2] ),
    .D(\xfer_count[3] ),
    .X(_1533_));
 sky130_fd_sc_hd__a32o_1 _5138_ (.A1(_1526_),
    .A2(_1531_),
    .A3(_1533_),
    .B1(serial_xfer),
    .B2(\xfer_state[0] ),
    .X(_0016_));
 sky130_fd_sc_hd__nand2_1 _5139_ (.A(_1526_),
    .B(_1533_),
    .Y(_1534_));
 sky130_fd_sc_hd__or4b_1 _5140_ (.A(\xfer_count[0] ),
    .B(\xfer_count[2] ),
    .C(\xfer_count[3] ),
    .D_N(\xfer_count[1] ),
    .X(_1535_));
 sky130_fd_sc_hd__a2bb2o_1 _5141_ (.A1_N(_1531_),
    .A2_N(_1534_),
    .B1(_1535_),
    .B2(net1525),
    .X(_0017_));
 sky130_fd_sc_hd__buf_2 _5142_ (.A(\wbbd_state[7] ),
    .X(_1536_));
 sky130_fd_sc_hd__a21o_1 _5143_ (.A1(_1536_),
    .A2(_1513_),
    .B1(net1487),
    .X(_0011_));
 sky130_fd_sc_hd__buf_2 _5144_ (.A(\wbbd_state[8] ),
    .X(_1537_));
 sky130_fd_sc_hd__a21o_1 _5145_ (.A1(_1537_),
    .A2(_1513_),
    .B1(net1473),
    .X(_0012_));
 sky130_fd_sc_hd__buf_2 _5146_ (.A(\wbbd_state[9] ),
    .X(_1538_));
 sky130_fd_sc_hd__a21o_1 _5147_ (.A1(_1538_),
    .A2(_1513_),
    .B1(net1464),
    .X(_0013_));
 sky130_fd_sc_hd__inv_2 _5148_ (.A(net1502),
    .Y(_1539_));
 sky130_fd_sc_hd__inv_2 _5149_ (.A(net1498),
    .Y(_1540_));
 sky130_fd_sc_hd__o21ai_1 _5150_ (.A1(_1539_),
    .A2(_1523_),
    .B1(_1540_),
    .Y(_0009_));
 sky130_fd_sc_hd__inv_2 _5151_ (.A(\hkspi.pre_pass_thru_mgmt ),
    .Y(_1541_));
 sky130_fd_sc_hd__a41o_1 _5152_ (.A1(\hkspi.pre_pass_thru_user ),
    .A2(_1541_),
    .A3(_1462_),
    .A4(_1436_),
    .B1(net1455),
    .X(_0005_));
 sky130_fd_sc_hd__clkinv_2 _5153_ (.A(\xfer_state[0] ),
    .Y(_1542_));
 sky130_fd_sc_hd__inv_2 _5154_ (.A(\xfer_state[3] ),
    .Y(_1543_));
 sky130_fd_sc_hd__or2_1 _5155_ (.A(_1543_),
    .B(_1535_),
    .X(_1544_));
 sky130_fd_sc_hd__o21ai_1 _5156_ (.A1(serial_xfer),
    .A2(_1542_),
    .B1(_1544_),
    .Y(_0014_));
 sky130_fd_sc_hd__a31o_1 _5157_ (.A1(net1505),
    .A2(_1462_),
    .A3(_1436_),
    .B1(net1457),
    .X(_0008_));
 sky130_fd_sc_hd__buf_4 _5158_ (.A(\xfer_state[2] ),
    .X(_1545_));
 sky130_fd_sc_hd__inv_2 _5159_ (.A(\xfer_state[1] ),
    .Y(_1546_));
 sky130_fd_sc_hd__nor2_1 _5160_ (.A(_1546_),
    .B(_1533_),
    .Y(_1547_));
 sky130_fd_sc_hd__or2_1 _5161_ (.A(_1545_),
    .B(_1547_),
    .X(_1548_));
 sky130_fd_sc_hd__clkbuf_1 _5162_ (.A(_1548_),
    .X(_0015_));
 sky130_fd_sc_hd__o32ai_1 _5163_ (.A1(net1500),
    .A2(\hkspi.pre_pass_thru_mgmt ),
    .A3(_1469_),
    .B1(_1436_),
    .B2(_0825_),
    .Y(_0007_));
 sky130_fd_sc_hd__a2bb2o_1 _5164_ (.A1_N(_1472_),
    .A2_N(_1524_),
    .B1(_1436_),
    .B2(_1430_),
    .X(_0006_));
 sky130_fd_sc_hd__mux2_1 _5165_ (.A0(net84),
    .A1(net67),
    .S(\hkspi.pass_thru_mgmt_delay ),
    .X(_1549_));
 sky130_fd_sc_hd__clkbuf_1 _5166_ (.A(_1549_),
    .X(net252));
 sky130_fd_sc_hd__nor2_2 _5167_ (.A(\hkspi.pass_thru_mgmt_delay ),
    .B(_1505_),
    .Y(net253));
 sky130_fd_sc_hd__mux2_2 _5168_ (.A0(net83),
    .A1(clknet_2_1_0_mgmt_gpio_in[4]),
    .S(\hkspi.pass_thru_mgmt ),
    .X(_1550_));
 sky130_fd_sc_hd__buf_1 _5169_ (.A(_1550_),
    .X(net250));
 sky130_fd_sc_hd__nor2_2 _5170_ (.A(\hkspi.pass_thru_mgmt ),
    .B(_1505_),
    .Y(net251));
 sky130_fd_sc_hd__or2b_1 _5171_ (.A(\hkspi.pass_thru_mgmt_delay ),
    .B_N(net86),
    .X(_1551_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _5172_ (.A(_1551_),
    .X(net255));
 sky130_fd_sc_hd__inv_2 _5173_ (.A(net255),
    .Y(net256));
 sky130_fd_sc_hd__or2_1 _5174_ (.A(\hkspi.pass_thru_mgmt ),
    .B(net88),
    .X(_1552_));
 sky130_fd_sc_hd__clkbuf_2 _5175_ (.A(_1552_),
    .X(net259));
 sky130_fd_sc_hd__inv_2 _5176_ (.A(net259),
    .Y(net258));
 sky130_fd_sc_hd__mux2_1 _5177_ (.A0(net85),
    .A1(_1466_),
    .S(\hkspi.pass_thru_mgmt_delay ),
    .X(_1553_));
 sky130_fd_sc_hd__clkbuf_1 _5178_ (.A(_1553_),
    .X(net254));
 sky130_fd_sc_hd__and2b_1 _5179_ (.A_N(\hkspi.pass_thru_mgmt_delay ),
    .B(net73),
    .X(_1554_));
 sky130_fd_sc_hd__clkbuf_4 _5180_ (.A(_1554_),
    .X(net312));
 sky130_fd_sc_hd__and2b_1 _5181_ (.A_N(\hkspi.pass_thru_mgmt ),
    .B(net74),
    .X(_1555_));
 sky130_fd_sc_hd__clkbuf_4 _5182_ (.A(_1555_),
    .X(net313));
 sky130_fd_sc_hd__nor2_1 _5183_ (.A(\hkspi.state[1] ),
    .B(\hkspi.state[4] ),
    .Y(_1556_));
 sky130_fd_sc_hd__o21a_1 _5184_ (.A1(\hkspi.state[2] ),
    .A2(_1556_),
    .B1(_0985_),
    .X(_0018_));
 sky130_fd_sc_hd__inv_2 _5185_ (.A(\gpio_configure[26][3] ),
    .Y(net225));
 sky130_fd_sc_hd__mux2_2 _5186_ (.A0(\mgmt_gpio_data[37] ),
    .A1(net91),
    .S(net76),
    .X(_1557_));
 sky130_fd_sc_hd__clkbuf_1 _5187_ (.A(_1557_),
    .X(net249));
 sky130_fd_sc_hd__mux2_2 _5188_ (.A0(\mgmt_gpio_data[36] ),
    .A1(net89),
    .S(net76),
    .X(_1558_));
 sky130_fd_sc_hd__clkbuf_1 _5189_ (.A(_1558_),
    .X(net248));
 sky130_fd_sc_hd__clkinv_2 _5190_ (.A(\gpio_configure[37][3] ),
    .Y(_1559_));
 sky130_fd_sc_hd__mux2_1 _5191_ (.A0(_1559_),
    .A1(net92),
    .S(net76),
    .X(_1560_));
 sky130_fd_sc_hd__clkbuf_1 _5192_ (.A(_1560_),
    .X(net237));
 sky130_fd_sc_hd__clkinv_2 _5193_ (.A(\gpio_configure[36][3] ),
    .Y(_1561_));
 sky130_fd_sc_hd__mux2_1 _5194_ (.A0(_1561_),
    .A1(net90),
    .S(net76),
    .X(_1562_));
 sky130_fd_sc_hd__clkbuf_1 _5195_ (.A(_1562_),
    .X(net236));
 sky130_fd_sc_hd__inv_2 _5196_ (.A(\gpio_configure[35][3] ),
    .Y(_1563_));
 sky130_fd_sc_hd__mux2_8 _5197_ (.A0(_1563_),
    .A1(net82),
    .S(net79),
    .X(_1564_));
 sky130_fd_sc_hd__clkbuf_1 _5198_ (.A(_1564_),
    .X(net235));
 sky130_fd_sc_hd__mux2_4 _5199_ (.A0(\mgmt_gpio_data[32] ),
    .A1(net80),
    .S(net79),
    .X(_1565_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _5200_ (.A(_1565_),
    .X(\mgmt_gpio_out_pre[32] ));
 sky130_fd_sc_hd__mux2_4 _5201_ (.A0(\mgmt_gpio_data[33] ),
    .A1(net78),
    .S(net79),
    .X(_1566_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _5202_ (.A(_1566_),
    .X(\mgmt_gpio_out_pre[33] ));
 sky130_fd_sc_hd__mux2_8 _5203_ (.A0(\mgmt_gpio_data[35] ),
    .A1(net81),
    .S(net79),
    .X(_1567_));
 sky130_fd_sc_hd__clkbuf_1 _5204_ (.A(_1567_),
    .X(net247));
 sky130_fd_sc_hd__mux2_1 _5205_ (.A0(\mgmt_gpio_data[10] ),
    .A1(_1466_),
    .S(\hkspi.pass_thru_user_delay ),
    .X(_1568_));
 sky130_fd_sc_hd__clkbuf_1 _5206_ (.A(_1568_),
    .X(\mgmt_gpio_out_pre[10] ));
 sky130_fd_sc_hd__mux2_2 _5207_ (.A0(\mgmt_gpio_data[9] ),
    .A1(clknet_2_3_0_mgmt_gpio_in[4]),
    .S(\hkspi.pass_thru_user ),
    .X(_1569_));
 sky130_fd_sc_hd__buf_1 _5208_ (.A(_1569_),
    .X(\mgmt_gpio_out_pre[9] ));
 sky130_fd_sc_hd__mux2_1 _5209_ (.A0(\mgmt_gpio_data[8] ),
    .A1(net67),
    .S(\hkspi.pass_thru_user_delay ),
    .X(_1570_));
 sky130_fd_sc_hd__clkbuf_1 _5210_ (.A(_1570_),
    .X(\mgmt_gpio_out_pre[8] ));
 sky130_fd_sc_hd__mux2_1 _5211_ (.A0(\mgmt_gpio_data[6] ),
    .A1(net77),
    .S(net126),
    .X(_1571_));
 sky130_fd_sc_hd__buf_2 _5212_ (.A(_1571_),
    .X(\mgmt_gpio_out_pre[6] ));
 sky130_fd_sc_hd__mux2_1 _5213_ (.A0(\mgmt_gpio_data[1] ),
    .A1(\hkspi.SDO ),
    .S(_1507_),
    .X(_1572_));
 sky130_fd_sc_hd__mux2_1 _5214_ (.A0(_1572_),
    .A1(net38),
    .S(\hkspi.pass_thru_user ),
    .X(_1573_));
 sky130_fd_sc_hd__mux2_4 _5215_ (.A0(_1573_),
    .A1(net74),
    .S(\hkspi.pass_thru_mgmt ),
    .X(_1574_));
 sky130_fd_sc_hd__clkbuf_1 _5216_ (.A(_1574_),
    .X(net246));
 sky130_fd_sc_hd__mux2_4 _5217_ (.A0(\mgmt_gpio_data[0] ),
    .A1(net3),
    .S(net1),
    .X(_1575_));
 sky130_fd_sc_hd__clkbuf_1 _5218_ (.A(_1575_),
    .X(net245));
 sky130_fd_sc_hd__inv_2 _5219_ (.A(\gpio_configure[0][3] ),
    .Y(_1576_));
 sky130_fd_sc_hd__mux2_4 _5220_ (.A0(_1576_),
    .A1(\hkspi.sdoenb ),
    .S(_1508_),
    .X(_1577_));
 sky130_fd_sc_hd__clkbuf_1 _5221_ (.A(_1577_),
    .X(net218));
 sky130_fd_sc_hd__mux2_4 _5222_ (.A0(_1576_),
    .A1(net2),
    .S(net1),
    .X(_1578_));
 sky130_fd_sc_hd__clkbuf_1 _5223_ (.A(_1578_),
    .X(net207));
 sky130_fd_sc_hd__mux2_2 _5224_ (.A0(\mgmt_gpio_data[15] ),
    .A1(user_clock),
    .S(clk2_output_dest),
    .X(_1579_));
 sky130_fd_sc_hd__buf_1 _5225_ (.A(_1579_),
    .X(\mgmt_gpio_out_pre[15] ));
 sky130_fd_sc_hd__mux2_4 _5226_ (.A0(\mgmt_gpio_data[14] ),
    .A1(clknet_3_6_0_wb_clk_i),
    .S(clk1_output_dest),
    .X(_1580_));
 sky130_fd_sc_hd__buf_1 _5227_ (.A(_1580_),
    .X(\mgmt_gpio_out_pre[14] ));
 sky130_fd_sc_hd__mux2_1 _5228_ (.A0(\mgmt_gpio_data[13] ),
    .A1(net125),
    .S(trap_output_dest),
    .X(_1581_));
 sky130_fd_sc_hd__clkbuf_1 _5229_ (.A(_1581_),
    .X(\mgmt_gpio_out_pre[13] ));
 sky130_fd_sc_hd__mux2_1 _5230_ (.A0(serial_resetn_pre),
    .A1(serial_bb_resetn),
    .S(serial_bb_enable),
    .X(_1582_));
 sky130_fd_sc_hd__clkbuf_1 _5231_ (.A(_1582_),
    .X(net310));
 sky130_fd_sc_hd__mux2_1 _5232_ (.A0(serial_load_pre),
    .A1(serial_bb_load),
    .S(serial_bb_enable),
    .X(_1583_));
 sky130_fd_sc_hd__clkbuf_1 _5233_ (.A(_1583_),
    .X(net309));
 sky130_fd_sc_hd__buf_6 _5234_ (.A(net580),
    .X(_1584_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_wb_clk_i (.A(wb_clk_i),
    .X(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__nor2_2 _5236_ (.A(_1584_),
    .B(net506),
    .Y(_1585_));
 sky130_fd_sc_hd__a22o_2 _5237_ (.A1(_1584_),
    .A2(clknet_1_0__leaf_wbbd_sck),
    .B1(_1509_),
    .B2(_1585_),
    .X(csclk));
 sky130_fd_sc_hd__inv_2 _5238_ (.A(\gpio_configure[3][3] ),
    .Y(net238));
 sky130_fd_sc_hd__inv_2 _5239_ (.A(\gpio_configure[2][3] ),
    .Y(net229));
 sky130_fd_sc_hd__inv_2 _5240_ (.A(\gpio_configure[4][3] ),
    .Y(net239));
 sky130_fd_sc_hd__inv_2 _5241_ (.A(\gpio_configure[5][3] ),
    .Y(net240));
 sky130_fd_sc_hd__inv_2 _5242_ (.A(\gpio_configure[6][3] ),
    .Y(net241));
 sky130_fd_sc_hd__inv_2 _5243_ (.A(\gpio_configure[7][3] ),
    .Y(net242));
 sky130_fd_sc_hd__inv_2 _5244_ (.A(\gpio_configure[8][3] ),
    .Y(net243));
 sky130_fd_sc_hd__inv_2 _5245_ (.A(\gpio_configure[9][3] ),
    .Y(net244));
 sky130_fd_sc_hd__inv_2 _5246_ (.A(\gpio_configure[10][3] ),
    .Y(net208));
 sky130_fd_sc_hd__inv_2 _5247_ (.A(\gpio_configure[11][3] ),
    .Y(net209));
 sky130_fd_sc_hd__inv_2 _5248_ (.A(\gpio_configure[12][3] ),
    .Y(net210));
 sky130_fd_sc_hd__inv_2 _5249_ (.A(\gpio_configure[13][3] ),
    .Y(net211));
 sky130_fd_sc_hd__inv_2 _5250_ (.A(\gpio_configure[14][3] ),
    .Y(net212));
 sky130_fd_sc_hd__inv_2 _5251_ (.A(\gpio_configure[15][3] ),
    .Y(net213));
 sky130_fd_sc_hd__inv_2 _5252_ (.A(\gpio_configure[16][3] ),
    .Y(net214));
 sky130_fd_sc_hd__inv_2 _5253_ (.A(\gpio_configure[17][3] ),
    .Y(net215));
 sky130_fd_sc_hd__inv_2 _5254_ (.A(\gpio_configure[18][3] ),
    .Y(net216));
 sky130_fd_sc_hd__inv_2 _5255_ (.A(\gpio_configure[19][3] ),
    .Y(net217));
 sky130_fd_sc_hd__inv_2 _5256_ (.A(\gpio_configure[20][3] ),
    .Y(net219));
 sky130_fd_sc_hd__inv_2 _5257_ (.A(\gpio_configure[21][3] ),
    .Y(net220));
 sky130_fd_sc_hd__inv_2 _5258_ (.A(\gpio_configure[22][3] ),
    .Y(net221));
 sky130_fd_sc_hd__inv_2 _5259_ (.A(\gpio_configure[23][3] ),
    .Y(net222));
 sky130_fd_sc_hd__inv_2 _5260_ (.A(\gpio_configure[24][3] ),
    .Y(net223));
 sky130_fd_sc_hd__inv_2 _5261_ (.A(\gpio_configure[25][3] ),
    .Y(net224));
 sky130_fd_sc_hd__inv_2 _5262_ (.A(\gpio_configure[27][3] ),
    .Y(net226));
 sky130_fd_sc_hd__inv_2 _5263_ (.A(\gpio_configure[28][3] ),
    .Y(net227));
 sky130_fd_sc_hd__inv_2 _5264_ (.A(\gpio_configure[29][3] ),
    .Y(net228));
 sky130_fd_sc_hd__inv_2 _5265_ (.A(\gpio_configure[30][3] ),
    .Y(net230));
 sky130_fd_sc_hd__inv_2 _5266_ (.A(\gpio_configure[31][3] ),
    .Y(net231));
 sky130_fd_sc_hd__inv_2 _5267_ (.A(\gpio_configure[32][3] ),
    .Y(net232));
 sky130_fd_sc_hd__inv_2 _5268_ (.A(\gpio_configure[33][3] ),
    .Y(net233));
 sky130_fd_sc_hd__inv_2 _5269_ (.A(\gpio_configure[34][3] ),
    .Y(net234));
 sky130_fd_sc_hd__o21ai_1 _5270_ (.A1(\hkspi.rdstb ),
    .A2(net403),
    .B1(_1508_),
    .Y(_1586_));
 sky130_fd_sc_hd__and2_1 _5271_ (.A(_1536_),
    .B(net396),
    .X(_1587_));
 sky130_fd_sc_hd__clkbuf_1 _5272_ (.A(_1587_),
    .X(_0003_));
 sky130_fd_sc_hd__and2_1 _5273_ (.A(\wbbd_state[5] ),
    .B(net396),
    .X(_1588_));
 sky130_fd_sc_hd__clkbuf_1 _5274_ (.A(_1588_),
    .X(_0002_));
 sky130_fd_sc_hd__and2_1 _5275_ (.A(_1537_),
    .B(net396),
    .X(_1589_));
 sky130_fd_sc_hd__clkbuf_1 _5276_ (.A(_1589_),
    .X(_0001_));
 sky130_fd_sc_hd__and2_1 _5277_ (.A(net68),
    .B(net126),
    .X(_1590_));
 sky130_fd_sc_hd__clkbuf_1 _5278_ (.A(_1590_),
    .X(net305));
 sky130_fd_sc_hd__and2_1 _5279_ (.A(net63),
    .B(net79),
    .X(_1591_));
 sky130_fd_sc_hd__clkbuf_1 _5280_ (.A(_1591_),
    .X(net311));
 sky130_fd_sc_hd__and2_1 _5281_ (.A(net36),
    .B(net1),
    .X(_1592_));
 sky130_fd_sc_hd__clkbuf_1 _5282_ (.A(_1592_),
    .X(net203));
 sky130_fd_sc_hd__and2_1 _5283_ (.A(irq_1_inputsrc),
    .B(net70),
    .X(_1593_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _5284_ (.A(_1593_),
    .X(net205));
 sky130_fd_sc_hd__and2_1 _5285_ (.A(irq_2_inputsrc),
    .B(net39),
    .X(_1594_));
 sky130_fd_sc_hd__clkbuf_1 _5286_ (.A(_1594_),
    .X(net206));
 sky130_fd_sc_hd__and2_1 _5287_ (.A(_1538_),
    .B(net396),
    .X(_1595_));
 sky130_fd_sc_hd__clkbuf_1 _5288_ (.A(_1595_),
    .X(_0000_));
 sky130_fd_sc_hd__mux2_1 _5289_ (.A0(_1466_),
    .A1(net937),
    .S(_1584_),
    .X(_1596_));
 sky130_fd_sc_hd__buf_6 _5290_ (.A(net938),
    .X(_1597_));
 sky130_fd_sc_hd__buf_6 _5291_ (.A(_1597_),
    .X(_1598_));
 sky130_fd_sc_hd__or2b_1 _5292_ (.A(net609),
    .B_N(net580),
    .X(_1599_));
 sky130_fd_sc_hd__o21a_4 _5293_ (.A1(net524),
    .A2(_0824_),
    .B1(_1599_),
    .X(_1600_));
 sky130_fd_sc_hd__buf_8 _5294_ (.A(net525),
    .X(_1601_));
 sky130_fd_sc_hd__buf_4 _5295_ (.A(net526),
    .X(_1602_));
 sky130_fd_sc_hd__nand2_4 _5296_ (.A(_1091_),
    .B(_1602_),
    .Y(_1603_));
 sky130_fd_sc_hd__mux2_1 _5297_ (.A0(_1598_),
    .A1(net1326),
    .S(_1603_),
    .X(_1604_));
 sky130_fd_sc_hd__clkbuf_1 _5298_ (.A(net1694),
    .X(_0065_));
 sky130_fd_sc_hd__mux2_8 _5299_ (.A0(net542),
    .A1(net574),
    .S(_1584_),
    .X(_1605_));
 sky130_fd_sc_hd__buf_6 _5300_ (.A(net543),
    .X(_1606_));
 sky130_fd_sc_hd__buf_6 _5301_ (.A(_1606_),
    .X(_1607_));
 sky130_fd_sc_hd__mux2_1 _5302_ (.A0(_1607_),
    .A1(net968),
    .S(_1603_),
    .X(_1608_));
 sky130_fd_sc_hd__clkbuf_1 _5303_ (.A(net1750),
    .X(_0066_));
 sky130_fd_sc_hd__mux2_2 _5304_ (.A0(net517),
    .A1(net1063),
    .S(_0824_),
    .X(_1609_));
 sky130_fd_sc_hd__buf_6 _5305_ (.A(net518),
    .X(_1610_));
 sky130_fd_sc_hd__clkbuf_8 _5306_ (.A(_1610_),
    .X(_1611_));
 sky130_fd_sc_hd__mux2_1 _5307_ (.A0(_1611_),
    .A1(net1020),
    .S(_1603_),
    .X(_1612_));
 sky130_fd_sc_hd__clkbuf_1 _5308_ (.A(net1021),
    .X(_0067_));
 sky130_fd_sc_hd__mux2_1 _5309_ (.A0(net550),
    .A1(net703),
    .S(_0824_),
    .X(_1613_));
 sky130_fd_sc_hd__buf_4 _5310_ (.A(net551),
    .X(_1614_));
 sky130_fd_sc_hd__clkbuf_8 _5311_ (.A(_1614_),
    .X(_1615_));
 sky130_fd_sc_hd__mux2_1 _5312_ (.A0(_1615_),
    .A1(net903),
    .S(_1603_),
    .X(_1616_));
 sky130_fd_sc_hd__clkbuf_1 _5313_ (.A(_1616_),
    .X(_0068_));
 sky130_fd_sc_hd__mux2_8 _5314_ (.A0(net529),
    .A1(net618),
    .S(_1584_),
    .X(_1617_));
 sky130_fd_sc_hd__buf_6 _5315_ (.A(net530),
    .X(_1618_));
 sky130_fd_sc_hd__mux2_1 _5316_ (.A0(_1618_),
    .A1(net637),
    .S(_1603_),
    .X(_1619_));
 sky130_fd_sc_hd__clkbuf_1 _5317_ (.A(net638),
    .X(_0069_));
 sky130_fd_sc_hd__and2_1 _5318_ (.A(_1505_),
    .B(_1509_),
    .X(_1620_));
 sky130_fd_sc_hd__clkbuf_1 _5319_ (.A(_1620_),
    .X(_0019_));
 sky130_fd_sc_hd__and2_1 _5320_ (.A(_1505_),
    .B(_1509_),
    .X(_1621_));
 sky130_fd_sc_hd__clkbuf_1 _5321_ (.A(_1621_),
    .X(_0020_));
 sky130_fd_sc_hd__and2_1 _5322_ (.A(_1505_),
    .B(_1509_),
    .X(_1622_));
 sky130_fd_sc_hd__clkbuf_1 _5323_ (.A(_1622_),
    .X(_0023_));
 sky130_fd_sc_hd__and2_1 _5324_ (.A(_1505_),
    .B(_1509_),
    .X(_1623_));
 sky130_fd_sc_hd__clkbuf_1 _5325_ (.A(_1623_),
    .X(_0024_));
 sky130_fd_sc_hd__and2_1 _5326_ (.A(_1505_),
    .B(_1509_),
    .X(_1624_));
 sky130_fd_sc_hd__clkbuf_1 _5327_ (.A(_1624_),
    .X(_0025_));
 sky130_fd_sc_hd__and2_1 _5328_ (.A(_1505_),
    .B(_1509_),
    .X(_1625_));
 sky130_fd_sc_hd__clkbuf_1 _5329_ (.A(_1625_),
    .X(_0026_));
 sky130_fd_sc_hd__and2_1 _5330_ (.A(_1505_),
    .B(_1509_),
    .X(_1626_));
 sky130_fd_sc_hd__clkbuf_1 _5331_ (.A(_1626_),
    .X(_0027_));
 sky130_fd_sc_hd__clkbuf_2 _5332_ (.A(net418),
    .X(_1627_));
 sky130_fd_sc_hd__buf_4 _5333_ (.A(_1627_),
    .X(_1628_));
 sky130_fd_sc_hd__and2_1 _5334_ (.A(_1628_),
    .B(_1509_),
    .X(_1629_));
 sky130_fd_sc_hd__clkbuf_1 _5335_ (.A(_1629_),
    .X(_0028_));
 sky130_fd_sc_hd__buf_4 _5336_ (.A(_1507_),
    .X(_1630_));
 sky130_fd_sc_hd__and2_1 _5337_ (.A(_1628_),
    .B(_1630_),
    .X(_1631_));
 sky130_fd_sc_hd__clkbuf_1 _5338_ (.A(_1631_),
    .X(_0029_));
 sky130_fd_sc_hd__and2_1 _5339_ (.A(_1628_),
    .B(_1630_),
    .X(_1632_));
 sky130_fd_sc_hd__clkbuf_1 _5340_ (.A(_1632_),
    .X(_0030_));
 sky130_fd_sc_hd__and2_1 _5341_ (.A(_1628_),
    .B(_1630_),
    .X(_1633_));
 sky130_fd_sc_hd__clkbuf_1 _5342_ (.A(_1633_),
    .X(_0031_));
 sky130_fd_sc_hd__and2_1 _5343_ (.A(_1628_),
    .B(_1630_),
    .X(_1634_));
 sky130_fd_sc_hd__clkbuf_1 _5344_ (.A(_1634_),
    .X(_0032_));
 sky130_fd_sc_hd__and2_1 _5345_ (.A(_1628_),
    .B(_1630_),
    .X(_1635_));
 sky130_fd_sc_hd__clkbuf_1 _5346_ (.A(_1635_),
    .X(_0033_));
 sky130_fd_sc_hd__and2_1 _5347_ (.A(_1628_),
    .B(_1630_),
    .X(_1636_));
 sky130_fd_sc_hd__clkbuf_1 _5348_ (.A(_1636_),
    .X(_0034_));
 sky130_fd_sc_hd__and2_1 _5349_ (.A(_1628_),
    .B(_1630_),
    .X(_1637_));
 sky130_fd_sc_hd__clkbuf_1 _5350_ (.A(_1637_),
    .X(_0035_));
 sky130_fd_sc_hd__and2_1 _5351_ (.A(_1628_),
    .B(_1630_),
    .X(_1638_));
 sky130_fd_sc_hd__clkbuf_1 _5352_ (.A(_1638_),
    .X(_0036_));
 sky130_fd_sc_hd__and2_1 _5353_ (.A(_1628_),
    .B(_1630_),
    .X(_1639_));
 sky130_fd_sc_hd__clkbuf_1 _5354_ (.A(_1639_),
    .X(_0037_));
 sky130_fd_sc_hd__clkbuf_2 _5355_ (.A(_1627_),
    .X(_1640_));
 sky130_fd_sc_hd__and2_1 _5356_ (.A(_1640_),
    .B(_1630_),
    .X(_1641_));
 sky130_fd_sc_hd__clkbuf_1 _5357_ (.A(_1641_),
    .X(_0038_));
 sky130_fd_sc_hd__buf_2 _5358_ (.A(_1507_),
    .X(_1642_));
 sky130_fd_sc_hd__and2_1 _5359_ (.A(_1640_),
    .B(_1642_),
    .X(_1643_));
 sky130_fd_sc_hd__clkbuf_1 _5360_ (.A(_1643_),
    .X(_0039_));
 sky130_fd_sc_hd__and2_1 _5361_ (.A(_1640_),
    .B(_1642_),
    .X(_1644_));
 sky130_fd_sc_hd__clkbuf_1 _5362_ (.A(_1644_),
    .X(_0040_));
 sky130_fd_sc_hd__and2_1 _5363_ (.A(_1640_),
    .B(_1642_),
    .X(_1645_));
 sky130_fd_sc_hd__clkbuf_1 _5364_ (.A(_1645_),
    .X(_0041_));
 sky130_fd_sc_hd__and2_1 _5365_ (.A(_1640_),
    .B(_1642_),
    .X(_1646_));
 sky130_fd_sc_hd__clkbuf_1 _5366_ (.A(_1646_),
    .X(_0042_));
 sky130_fd_sc_hd__and2_1 _5367_ (.A(_1640_),
    .B(_1642_),
    .X(_1647_));
 sky130_fd_sc_hd__clkbuf_1 _5368_ (.A(_1647_),
    .X(_0043_));
 sky130_fd_sc_hd__and2_1 _5369_ (.A(_1640_),
    .B(_1642_),
    .X(_1648_));
 sky130_fd_sc_hd__clkbuf_1 _5370_ (.A(_1648_),
    .X(_0044_));
 sky130_fd_sc_hd__and2_1 _5371_ (.A(_1640_),
    .B(_1642_),
    .X(_1649_));
 sky130_fd_sc_hd__clkbuf_1 _5372_ (.A(_1649_),
    .X(_0045_));
 sky130_fd_sc_hd__and2_1 _5373_ (.A(_1640_),
    .B(_1642_),
    .X(_1650_));
 sky130_fd_sc_hd__clkbuf_1 _5374_ (.A(_1650_),
    .X(_0046_));
 sky130_fd_sc_hd__and2_1 _5375_ (.A(_1640_),
    .B(_1642_),
    .X(_1651_));
 sky130_fd_sc_hd__clkbuf_1 _5376_ (.A(_1651_),
    .X(_0047_));
 sky130_fd_sc_hd__clkbuf_2 _5377_ (.A(_1627_),
    .X(_1652_));
 sky130_fd_sc_hd__and2_1 _5378_ (.A(_1652_),
    .B(_1642_),
    .X(_1653_));
 sky130_fd_sc_hd__clkbuf_1 _5379_ (.A(_1653_),
    .X(_0048_));
 sky130_fd_sc_hd__buf_2 _5380_ (.A(_1507_),
    .X(_1654_));
 sky130_fd_sc_hd__and2_1 _5381_ (.A(_1652_),
    .B(_1654_),
    .X(_1655_));
 sky130_fd_sc_hd__clkbuf_1 _5382_ (.A(_1655_),
    .X(_0049_));
 sky130_fd_sc_hd__and2_1 _5383_ (.A(_1652_),
    .B(_1654_),
    .X(_1656_));
 sky130_fd_sc_hd__clkbuf_1 _5384_ (.A(_1656_),
    .X(_0050_));
 sky130_fd_sc_hd__and2_1 _5385_ (.A(_1652_),
    .B(_1654_),
    .X(_1657_));
 sky130_fd_sc_hd__clkbuf_1 _5386_ (.A(_1657_),
    .X(_0051_));
 sky130_fd_sc_hd__buf_6 _5387_ (.A(_1597_),
    .X(_1658_));
 sky130_fd_sc_hd__and2_1 _5388_ (.A(_0972_),
    .B(_1601_),
    .X(_1659_));
 sky130_fd_sc_hd__clkbuf_4 _5389_ (.A(_1659_),
    .X(_1660_));
 sky130_fd_sc_hd__mux2_1 _5390_ (.A0(net298),
    .A1(_1658_),
    .S(_1660_),
    .X(_1661_));
 sky130_fd_sc_hd__clkbuf_1 _5391_ (.A(net1443),
    .X(_0101_));
 sky130_fd_sc_hd__buf_6 _5392_ (.A(_1606_),
    .X(_1662_));
 sky130_fd_sc_hd__mux2_1 _5393_ (.A0(net299),
    .A1(_1662_),
    .S(_1660_),
    .X(_1663_));
 sky130_fd_sc_hd__clkbuf_1 _5394_ (.A(net958),
    .X(_0102_));
 sky130_fd_sc_hd__clkbuf_4 _5395_ (.A(_1610_),
    .X(_1664_));
 sky130_fd_sc_hd__mux2_1 _5396_ (.A0(net275),
    .A1(_1664_),
    .S(_1660_),
    .X(_1665_));
 sky130_fd_sc_hd__clkbuf_1 _5397_ (.A(net1129),
    .X(_0103_));
 sky130_fd_sc_hd__buf_6 _5398_ (.A(_1614_),
    .X(_1666_));
 sky130_fd_sc_hd__mux2_1 _5399_ (.A0(net276),
    .A1(_1666_),
    .S(_1660_),
    .X(_1667_));
 sky130_fd_sc_hd__clkbuf_1 _5400_ (.A(net949),
    .X(_0104_));
 sky130_fd_sc_hd__buf_6 _5401_ (.A(net530),
    .X(_1668_));
 sky130_fd_sc_hd__clkbuf_4 _5402_ (.A(_1668_),
    .X(_1669_));
 sky130_fd_sc_hd__mux2_1 _5403_ (.A0(net277),
    .A1(_1669_),
    .S(_1660_),
    .X(_1670_));
 sky130_fd_sc_hd__clkbuf_1 _5404_ (.A(net1082),
    .X(_0105_));
 sky130_fd_sc_hd__mux2_8 _5405_ (.A0(net520),
    .A1(net1553),
    .S(_1584_),
    .X(_1671_));
 sky130_fd_sc_hd__buf_4 _5406_ (.A(net521),
    .X(_1672_));
 sky130_fd_sc_hd__mux2_1 _5407_ (.A0(net278),
    .A1(_1672_),
    .S(_1660_),
    .X(_1673_));
 sky130_fd_sc_hd__clkbuf_1 _5408_ (.A(net844),
    .X(_0106_));
 sky130_fd_sc_hd__mux2_8 _5409_ (.A0(net532),
    .A1(net1533),
    .S(_1584_),
    .X(_1674_));
 sky130_fd_sc_hd__buf_4 _5410_ (.A(net533),
    .X(_1675_));
 sky130_fd_sc_hd__mux2_1 _5411_ (.A0(net279),
    .A1(_1675_),
    .S(_1660_),
    .X(_1676_));
 sky130_fd_sc_hd__clkbuf_1 _5412_ (.A(net819),
    .X(_0107_));
 sky130_fd_sc_hd__mux2_4 _5413_ (.A0(net510),
    .A1(net1541),
    .S(_1584_),
    .X(_1677_));
 sky130_fd_sc_hd__buf_6 _5414_ (.A(net511),
    .X(_1678_));
 sky130_fd_sc_hd__clkbuf_4 _5415_ (.A(_1678_),
    .X(_1679_));
 sky130_fd_sc_hd__mux2_1 _5416_ (.A0(net280),
    .A1(_1679_),
    .S(_1660_),
    .X(_1680_));
 sky130_fd_sc_hd__clkbuf_1 _5417_ (.A(net1235),
    .X(_0108_));
 sky130_fd_sc_hd__and2_1 _5418_ (.A(_0941_),
    .B(net525),
    .X(_1681_));
 sky130_fd_sc_hd__clkbuf_4 _5419_ (.A(_1681_),
    .X(_1682_));
 sky130_fd_sc_hd__mux2_1 _5420_ (.A0(net274),
    .A1(_1658_),
    .S(_1682_),
    .X(_1683_));
 sky130_fd_sc_hd__clkbuf_1 _5421_ (.A(net1366),
    .X(_0109_));
 sky130_fd_sc_hd__mux2_1 _5422_ (.A0(net285),
    .A1(_1662_),
    .S(_1682_),
    .X(_1684_));
 sky130_fd_sc_hd__clkbuf_1 _5423_ (.A(net953),
    .X(_0110_));
 sky130_fd_sc_hd__mux2_1 _5424_ (.A0(net292),
    .A1(_1664_),
    .S(_1682_),
    .X(_1685_));
 sky130_fd_sc_hd__clkbuf_1 _5425_ (.A(net1124),
    .X(_0111_));
 sky130_fd_sc_hd__mux2_1 _5426_ (.A0(net293),
    .A1(_1666_),
    .S(_1682_),
    .X(_1686_));
 sky130_fd_sc_hd__clkbuf_1 _5427_ (.A(net934),
    .X(_0112_));
 sky130_fd_sc_hd__mux2_1 _5428_ (.A0(net294),
    .A1(_1669_),
    .S(_1682_),
    .X(_1687_));
 sky130_fd_sc_hd__clkbuf_1 _5429_ (.A(net1087),
    .X(_0113_));
 sky130_fd_sc_hd__mux2_1 _5430_ (.A0(net295),
    .A1(_1672_),
    .S(_1682_),
    .X(_1688_));
 sky130_fd_sc_hd__clkbuf_1 _5431_ (.A(net875),
    .X(_0114_));
 sky130_fd_sc_hd__buf_4 _5432_ (.A(net533),
    .X(_1689_));
 sky130_fd_sc_hd__mux2_1 _5433_ (.A0(net296),
    .A1(_1689_),
    .S(_1682_),
    .X(_1690_));
 sky130_fd_sc_hd__clkbuf_1 _5434_ (.A(net883),
    .X(_0115_));
 sky130_fd_sc_hd__mux2_1 _5435_ (.A0(net297),
    .A1(_1679_),
    .S(_1682_),
    .X(_1691_));
 sky130_fd_sc_hd__clkbuf_1 _5436_ (.A(net1267),
    .X(_0116_));
 sky130_fd_sc_hd__nand2_1 _5437_ (.A(_1328_),
    .B(_1602_),
    .Y(_1692_));
 sky130_fd_sc_hd__mux2_1 _5438_ (.A0(_1598_),
    .A1(net290),
    .S(_1692_),
    .X(_1693_));
 sky130_fd_sc_hd__clkbuf_1 _5439_ (.A(net1303),
    .X(_0117_));
 sky130_fd_sc_hd__mux2_1 _5440_ (.A0(_1607_),
    .A1(net291),
    .S(_1692_),
    .X(_1694_));
 sky130_fd_sc_hd__clkbuf_1 _5441_ (.A(net1081),
    .X(_0118_));
 sky130_fd_sc_hd__and2_1 _5442_ (.A(_1652_),
    .B(_1654_),
    .X(_1695_));
 sky130_fd_sc_hd__clkbuf_1 _5443_ (.A(_1695_),
    .X(_0052_));
 sky130_fd_sc_hd__and2_1 _5444_ (.A(_1652_),
    .B(_1654_),
    .X(_1696_));
 sky130_fd_sc_hd__clkbuf_1 _5445_ (.A(_1696_),
    .X(_0053_));
 sky130_fd_sc_hd__and2_1 _5446_ (.A(_1652_),
    .B(_1654_),
    .X(_1697_));
 sky130_fd_sc_hd__clkbuf_1 _5447_ (.A(_1697_),
    .X(_0054_));
 sky130_fd_sc_hd__and2_1 _5448_ (.A(_1652_),
    .B(_1654_),
    .X(_1698_));
 sky130_fd_sc_hd__clkbuf_1 _5449_ (.A(_1698_),
    .X(_0055_));
 sky130_fd_sc_hd__and2_1 _5450_ (.A(_1652_),
    .B(_1654_),
    .X(_1699_));
 sky130_fd_sc_hd__clkbuf_1 _5451_ (.A(_1699_),
    .X(_0056_));
 sky130_fd_sc_hd__o21ai_1 _5452_ (.A1(net524),
    .A2(_1584_),
    .B1(net610),
    .Y(_1700_));
 sky130_fd_sc_hd__or4_2 _5453_ (.A(_0909_),
    .B(_0964_),
    .C(_1507_),
    .D(net611),
    .X(_1701_));
 sky130_fd_sc_hd__buf_4 _5454_ (.A(_1701_),
    .X(_1702_));
 sky130_fd_sc_hd__mux2_1 _5455_ (.A0(_1598_),
    .A1(net1334),
    .S(_1702_),
    .X(_1703_));
 sky130_fd_sc_hd__clkbuf_1 _5456_ (.A(net1335),
    .X(_0119_));
 sky130_fd_sc_hd__mux2_1 _5457_ (.A0(_1607_),
    .A1(net977),
    .S(_1702_),
    .X(_1704_));
 sky130_fd_sc_hd__clkbuf_1 _5458_ (.A(net978),
    .X(_0120_));
 sky130_fd_sc_hd__mux2_1 _5459_ (.A0(_1611_),
    .A1(net962),
    .S(_1702_),
    .X(_1705_));
 sky130_fd_sc_hd__clkbuf_1 _5460_ (.A(net963),
    .X(_0121_));
 sky130_fd_sc_hd__mux2_1 _5461_ (.A0(_1615_),
    .A1(net889),
    .S(_1702_),
    .X(_1706_));
 sky130_fd_sc_hd__clkbuf_1 _5462_ (.A(net890),
    .X(_0122_));
 sky130_fd_sc_hd__mux2_1 _5463_ (.A0(_1618_),
    .A1(net616),
    .S(_1702_),
    .X(_1707_));
 sky130_fd_sc_hd__clkbuf_1 _5464_ (.A(net617),
    .X(_0123_));
 sky130_fd_sc_hd__clkbuf_16 _5465_ (.A(_1672_),
    .X(_1708_));
 sky130_fd_sc_hd__mux2_1 _5466_ (.A0(_1708_),
    .A1(net1322),
    .S(_1702_),
    .X(_1709_));
 sky130_fd_sc_hd__clkbuf_1 _5467_ (.A(net1323),
    .X(_0124_));
 sky130_fd_sc_hd__buf_12 _5468_ (.A(_1689_),
    .X(_1710_));
 sky130_fd_sc_hd__mux2_1 _5469_ (.A0(_1710_),
    .A1(net1327),
    .S(_1702_),
    .X(_1711_));
 sky130_fd_sc_hd__clkbuf_1 _5470_ (.A(net1328),
    .X(_0125_));
 sky130_fd_sc_hd__buf_6 _5471_ (.A(_1678_),
    .X(_1712_));
 sky130_fd_sc_hd__mux2_1 _5472_ (.A0(_1712_),
    .A1(net956),
    .S(_1702_),
    .X(_1713_));
 sky130_fd_sc_hd__clkbuf_1 _5473_ (.A(net957),
    .X(_0126_));
 sky130_fd_sc_hd__or4_4 _5474_ (.A(_0909_),
    .B(_0875_),
    .C(_1506_),
    .D(net611),
    .X(_1714_));
 sky130_fd_sc_hd__clkbuf_4 _5475_ (.A(_1714_),
    .X(_1715_));
 sky130_fd_sc_hd__mux2_1 _5476_ (.A0(_1598_),
    .A1(net1344),
    .S(_1715_),
    .X(_1716_));
 sky130_fd_sc_hd__clkbuf_1 _5477_ (.A(net1345),
    .X(_0127_));
 sky130_fd_sc_hd__mux2_1 _5478_ (.A0(_1607_),
    .A1(net1024),
    .S(_1715_),
    .X(_1717_));
 sky130_fd_sc_hd__clkbuf_1 _5479_ (.A(net1025),
    .X(_0128_));
 sky130_fd_sc_hd__mux2_1 _5480_ (.A0(_1611_),
    .A1(net1012),
    .S(_1715_),
    .X(_1718_));
 sky130_fd_sc_hd__clkbuf_1 _5481_ (.A(net1013),
    .X(_0129_));
 sky130_fd_sc_hd__mux2_1 _5482_ (.A0(_1615_),
    .A1(net873),
    .S(_1715_),
    .X(_1719_));
 sky130_fd_sc_hd__clkbuf_1 _5483_ (.A(net874),
    .X(_0130_));
 sky130_fd_sc_hd__mux2_1 _5484_ (.A0(_1618_),
    .A1(net643),
    .S(_1715_),
    .X(_1720_));
 sky130_fd_sc_hd__clkbuf_1 _5485_ (.A(net644),
    .X(_0131_));
 sky130_fd_sc_hd__mux2_1 _5486_ (.A0(_1708_),
    .A1(net1119),
    .S(_1715_),
    .X(_1721_));
 sky130_fd_sc_hd__clkbuf_1 _5487_ (.A(net1120),
    .X(_0132_));
 sky130_fd_sc_hd__mux2_1 _5488_ (.A0(_1710_),
    .A1(net1117),
    .S(_1715_),
    .X(_1722_));
 sky130_fd_sc_hd__clkbuf_1 _5489_ (.A(net1118),
    .X(_0133_));
 sky130_fd_sc_hd__mux2_1 _5490_ (.A0(_1712_),
    .A1(net975),
    .S(_1715_),
    .X(_1723_));
 sky130_fd_sc_hd__clkbuf_1 _5491_ (.A(net976),
    .X(_0134_));
 sky130_fd_sc_hd__buf_2 _5492_ (.A(_1601_),
    .X(_1724_));
 sky130_fd_sc_hd__and2_2 _5493_ (.A(_1130_),
    .B(_1724_),
    .X(_1725_));
 sky130_fd_sc_hd__mux2_1 _5494_ (.A0(net1446),
    .A1(_1658_),
    .S(_1725_),
    .X(_1726_));
 sky130_fd_sc_hd__clkbuf_1 _5495_ (.A(_1726_),
    .X(_0135_));
 sky130_fd_sc_hd__mux2_1 _5496_ (.A0(net983),
    .A1(_1662_),
    .S(_1725_),
    .X(_1727_));
 sky130_fd_sc_hd__clkbuf_1 _5497_ (.A(net984),
    .X(_0136_));
 sky130_fd_sc_hd__mux2_1 _5498_ (.A0(net1098),
    .A1(_1664_),
    .S(_1725_),
    .X(_1728_));
 sky130_fd_sc_hd__clkbuf_1 _5499_ (.A(net1099),
    .X(_0137_));
 sky130_fd_sc_hd__mux2_1 _5500_ (.A0(net925),
    .A1(_1666_),
    .S(_1725_),
    .X(_1729_));
 sky130_fd_sc_hd__clkbuf_1 _5501_ (.A(net926),
    .X(_0138_));
 sky130_fd_sc_hd__mux2_1 _5502_ (.A0(net1329),
    .A1(_1669_),
    .S(_1725_),
    .X(_1730_));
 sky130_fd_sc_hd__clkbuf_1 _5503_ (.A(_1730_),
    .X(_0139_));
 sky130_fd_sc_hd__buf_8 _5504_ (.A(net938),
    .X(_1731_));
 sky130_fd_sc_hd__clkbuf_4 _5505_ (.A(_1731_),
    .X(_1732_));
 sky130_fd_sc_hd__and2_2 _5506_ (.A(_1073_),
    .B(_1724_),
    .X(_1733_));
 sky130_fd_sc_hd__mux2_1 _5507_ (.A0(net1423),
    .A1(_1732_),
    .S(_1733_),
    .X(_1734_));
 sky130_fd_sc_hd__clkbuf_1 _5508_ (.A(_1734_),
    .X(_0140_));
 sky130_fd_sc_hd__mux2_1 _5509_ (.A0(net985),
    .A1(_1662_),
    .S(_1733_),
    .X(_1735_));
 sky130_fd_sc_hd__clkbuf_1 _5510_ (.A(net986),
    .X(_0141_));
 sky130_fd_sc_hd__mux2_1 _5511_ (.A0(net1107),
    .A1(_1664_),
    .S(_1733_),
    .X(_1736_));
 sky130_fd_sc_hd__clkbuf_1 _5512_ (.A(net1108),
    .X(_0142_));
 sky130_fd_sc_hd__mux2_1 _5513_ (.A0(net943),
    .A1(_1666_),
    .S(_1733_),
    .X(_1737_));
 sky130_fd_sc_hd__clkbuf_1 _5514_ (.A(net944),
    .X(_0143_));
 sky130_fd_sc_hd__mux2_1 _5515_ (.A0(net1113),
    .A1(_1669_),
    .S(_1733_),
    .X(_1738_));
 sky130_fd_sc_hd__clkbuf_1 _5516_ (.A(net1114),
    .X(_0144_));
 sky130_fd_sc_hd__buf_8 _5517_ (.A(net526),
    .X(_1739_));
 sky130_fd_sc_hd__nand2_2 _5518_ (.A(_1110_),
    .B(_1739_),
    .Y(_1740_));
 sky130_fd_sc_hd__mux2_1 _5519_ (.A0(_1598_),
    .A1(net1397),
    .S(_1740_),
    .X(_1741_));
 sky130_fd_sc_hd__clkbuf_1 _5520_ (.A(_1741_),
    .X(_0145_));
 sky130_fd_sc_hd__mux2_1 _5521_ (.A0(_1607_),
    .A1(net969),
    .S(_1740_),
    .X(_1742_));
 sky130_fd_sc_hd__clkbuf_1 _5522_ (.A(net970),
    .X(_0146_));
 sky130_fd_sc_hd__mux2_1 _5523_ (.A0(_1611_),
    .A1(net1014),
    .S(_1740_),
    .X(_1743_));
 sky130_fd_sc_hd__clkbuf_1 _5524_ (.A(net1015),
    .X(_0147_));
 sky130_fd_sc_hd__mux2_1 _5525_ (.A0(_1615_),
    .A1(net906),
    .S(_1740_),
    .X(_1744_));
 sky130_fd_sc_hd__clkbuf_1 _5526_ (.A(net907),
    .X(_0148_));
 sky130_fd_sc_hd__mux2_1 _5527_ (.A0(_1618_),
    .A1(net692),
    .S(_1740_),
    .X(_1745_));
 sky130_fd_sc_hd__clkbuf_1 _5528_ (.A(net693),
    .X(_0149_));
 sky130_fd_sc_hd__nand2_4 _5529_ (.A(_1121_),
    .B(_1739_),
    .Y(_1746_));
 sky130_fd_sc_hd__mux2_1 _5530_ (.A0(_1598_),
    .A1(net1387),
    .S(_1746_),
    .X(_1747_));
 sky130_fd_sc_hd__clkbuf_1 _5531_ (.A(_1747_),
    .X(_0150_));
 sky130_fd_sc_hd__mux2_1 _5532_ (.A0(_1607_),
    .A1(net1001),
    .S(_1746_),
    .X(_1748_));
 sky130_fd_sc_hd__clkbuf_1 _5533_ (.A(_1748_),
    .X(_0151_));
 sky130_fd_sc_hd__mux2_1 _5534_ (.A0(_1611_),
    .A1(net979),
    .S(_1746_),
    .X(_1749_));
 sky130_fd_sc_hd__clkbuf_1 _5535_ (.A(net980),
    .X(_0152_));
 sky130_fd_sc_hd__mux2_1 _5536_ (.A0(_1615_),
    .A1(net928),
    .S(_1746_),
    .X(_1750_));
 sky130_fd_sc_hd__clkbuf_1 _5537_ (.A(_1750_),
    .X(_0153_));
 sky130_fd_sc_hd__mux2_1 _5538_ (.A0(_1618_),
    .A1(net1766),
    .S(_1746_),
    .X(_1751_));
 sky130_fd_sc_hd__clkbuf_1 _5539_ (.A(net619),
    .X(_0154_));
 sky130_fd_sc_hd__nand2_2 _5540_ (.A(_1151_),
    .B(_1739_),
    .Y(_1752_));
 sky130_fd_sc_hd__mux2_1 _5541_ (.A0(_1598_),
    .A1(net1412),
    .S(_1752_),
    .X(_1753_));
 sky130_fd_sc_hd__clkbuf_1 _5542_ (.A(_1753_),
    .X(_0155_));
 sky130_fd_sc_hd__mux2_1 _5543_ (.A0(_1607_),
    .A1(net1038),
    .S(_1752_),
    .X(_1754_));
 sky130_fd_sc_hd__clkbuf_1 _5544_ (.A(_1754_),
    .X(_0156_));
 sky130_fd_sc_hd__mux2_1 _5545_ (.A0(_1611_),
    .A1(net997),
    .S(_1752_),
    .X(_1755_));
 sky130_fd_sc_hd__clkbuf_1 _5546_ (.A(net998),
    .X(_0157_));
 sky130_fd_sc_hd__mux2_1 _5547_ (.A0(_1615_),
    .A1(net893),
    .S(_1752_),
    .X(_1756_));
 sky130_fd_sc_hd__clkbuf_1 _5548_ (.A(_1756_),
    .X(_0158_));
 sky130_fd_sc_hd__mux2_1 _5549_ (.A0(_1618_),
    .A1(net647),
    .S(_1752_),
    .X(_1757_));
 sky130_fd_sc_hd__clkbuf_1 _5550_ (.A(net648),
    .X(_0159_));
 sky130_fd_sc_hd__nand2_2 _5551_ (.A(_1084_),
    .B(_1739_),
    .Y(_1758_));
 sky130_fd_sc_hd__mux2_1 _5552_ (.A0(_1598_),
    .A1(net1405),
    .S(_1758_),
    .X(_1759_));
 sky130_fd_sc_hd__clkbuf_1 _5553_ (.A(_1759_),
    .X(_0160_));
 sky130_fd_sc_hd__mux2_1 _5554_ (.A0(_1607_),
    .A1(net1100),
    .S(_1758_),
    .X(_1760_));
 sky130_fd_sc_hd__clkbuf_1 _5555_ (.A(_1760_),
    .X(_0161_));
 sky130_fd_sc_hd__mux2_1 _5556_ (.A0(_1611_),
    .A1(net1046),
    .S(_1758_),
    .X(_1761_));
 sky130_fd_sc_hd__clkbuf_1 _5557_ (.A(net1047),
    .X(_0162_));
 sky130_fd_sc_hd__mux2_1 _5558_ (.A0(_1615_),
    .A1(net959),
    .S(_1758_),
    .X(_1762_));
 sky130_fd_sc_hd__clkbuf_1 _5559_ (.A(_1762_),
    .X(_0163_));
 sky130_fd_sc_hd__mux2_1 _5560_ (.A0(_1618_),
    .A1(net655),
    .S(_1758_),
    .X(_1763_));
 sky130_fd_sc_hd__clkbuf_1 _5561_ (.A(net656),
    .X(_0164_));
 sky130_fd_sc_hd__and2_2 _5562_ (.A(_1100_),
    .B(_1724_),
    .X(_1764_));
 sky130_fd_sc_hd__mux2_1 _5563_ (.A0(net1438),
    .A1(_1732_),
    .S(_1764_),
    .X(_1765_));
 sky130_fd_sc_hd__clkbuf_1 _5564_ (.A(_1765_),
    .X(_0165_));
 sky130_fd_sc_hd__mux2_1 _5565_ (.A0(net965),
    .A1(_1662_),
    .S(_1764_),
    .X(_1766_));
 sky130_fd_sc_hd__clkbuf_1 _5566_ (.A(_1766_),
    .X(_0166_));
 sky130_fd_sc_hd__mux2_1 _5567_ (.A0(net1294),
    .A1(_1664_),
    .S(_1764_),
    .X(_1767_));
 sky130_fd_sc_hd__clkbuf_1 _5568_ (.A(_1767_),
    .X(_0167_));
 sky130_fd_sc_hd__mux2_1 _5569_ (.A0(net916),
    .A1(_1666_),
    .S(_1764_),
    .X(_1768_));
 sky130_fd_sc_hd__clkbuf_1 _5570_ (.A(_1768_),
    .X(_0168_));
 sky130_fd_sc_hd__mux2_1 _5571_ (.A0(net1170),
    .A1(_1669_),
    .S(_1764_),
    .X(_1769_));
 sky130_fd_sc_hd__clkbuf_1 _5572_ (.A(_1769_),
    .X(_0169_));
 sky130_fd_sc_hd__nand2_2 _5573_ (.A(_1104_),
    .B(_1739_),
    .Y(_1770_));
 sky130_fd_sc_hd__mux2_1 _5574_ (.A0(_1598_),
    .A1(net1352),
    .S(_1770_),
    .X(_1771_));
 sky130_fd_sc_hd__clkbuf_1 _5575_ (.A(_1771_),
    .X(_0170_));
 sky130_fd_sc_hd__mux2_1 _5576_ (.A0(_1607_),
    .A1(net1035),
    .S(_1770_),
    .X(_1772_));
 sky130_fd_sc_hd__clkbuf_1 _5577_ (.A(_1772_),
    .X(_0171_));
 sky130_fd_sc_hd__mux2_1 _5578_ (.A0(_1611_),
    .A1(net1048),
    .S(_1770_),
    .X(_1773_));
 sky130_fd_sc_hd__clkbuf_1 _5579_ (.A(net1049),
    .X(_0172_));
 sky130_fd_sc_hd__mux2_1 _5580_ (.A0(_1615_),
    .A1(net929),
    .S(_1770_),
    .X(_1774_));
 sky130_fd_sc_hd__clkbuf_1 _5581_ (.A(_1774_),
    .X(_0173_));
 sky130_fd_sc_hd__mux2_1 _5582_ (.A0(_1618_),
    .A1(net663),
    .S(_1770_),
    .X(_1775_));
 sky130_fd_sc_hd__clkbuf_1 _5583_ (.A(net664),
    .X(_0174_));
 sky130_fd_sc_hd__and2_2 _5584_ (.A(_1126_),
    .B(_1724_),
    .X(_1776_));
 sky130_fd_sc_hd__mux2_1 _5585_ (.A0(net1445),
    .A1(_1732_),
    .S(_1776_),
    .X(_1777_));
 sky130_fd_sc_hd__clkbuf_1 _5586_ (.A(_1777_),
    .X(_0175_));
 sky130_fd_sc_hd__buf_4 _5587_ (.A(_1606_),
    .X(_1778_));
 sky130_fd_sc_hd__mux2_1 _5588_ (.A0(net1255),
    .A1(_1778_),
    .S(_1776_),
    .X(_1779_));
 sky130_fd_sc_hd__clkbuf_1 _5589_ (.A(_1779_),
    .X(_0176_));
 sky130_fd_sc_hd__mux2_1 _5590_ (.A0(net1290),
    .A1(_1664_),
    .S(_1776_),
    .X(_1780_));
 sky130_fd_sc_hd__clkbuf_1 _5591_ (.A(_1780_),
    .X(_0177_));
 sky130_fd_sc_hd__mux2_1 _5592_ (.A0(net1173),
    .A1(_1666_),
    .S(_1776_),
    .X(_1781_));
 sky130_fd_sc_hd__clkbuf_1 _5593_ (.A(_1781_),
    .X(_0178_));
 sky130_fd_sc_hd__mux2_1 _5594_ (.A0(net1310),
    .A1(_1669_),
    .S(_1776_),
    .X(_1782_));
 sky130_fd_sc_hd__clkbuf_1 _5595_ (.A(_1782_),
    .X(_0179_));
 sky130_fd_sc_hd__and2_2 _5596_ (.A(_1131_),
    .B(_1724_),
    .X(_1783_));
 sky130_fd_sc_hd__mux2_1 _5597_ (.A0(net1419),
    .A1(_1732_),
    .S(_1783_),
    .X(_1784_));
 sky130_fd_sc_hd__clkbuf_1 _5598_ (.A(_1784_),
    .X(_0180_));
 sky130_fd_sc_hd__mux2_1 _5599_ (.A0(net1028),
    .A1(_1778_),
    .S(_1783_),
    .X(_1785_));
 sky130_fd_sc_hd__clkbuf_1 _5600_ (.A(_1785_),
    .X(_0181_));
 sky130_fd_sc_hd__mux2_1 _5601_ (.A0(net1144),
    .A1(_1664_),
    .S(_1783_),
    .X(_1786_));
 sky130_fd_sc_hd__clkbuf_1 _5602_ (.A(_1786_),
    .X(_0182_));
 sky130_fd_sc_hd__mux2_1 _5603_ (.A0(net955),
    .A1(_1666_),
    .S(_1783_),
    .X(_1787_));
 sky130_fd_sc_hd__clkbuf_1 _5604_ (.A(_1787_),
    .X(_0183_));
 sky130_fd_sc_hd__mux2_1 _5605_ (.A0(net1126),
    .A1(_1669_),
    .S(_1783_),
    .X(_1788_));
 sky130_fd_sc_hd__clkbuf_1 _5606_ (.A(_1788_),
    .X(_0184_));
 sky130_fd_sc_hd__nand2_2 _5607_ (.A(_1129_),
    .B(_1739_),
    .Y(_1789_));
 sky130_fd_sc_hd__mux2_1 _5608_ (.A0(_1598_),
    .A1(net1351),
    .S(_1789_),
    .X(_1790_));
 sky130_fd_sc_hd__clkbuf_1 _5609_ (.A(_1790_),
    .X(_0185_));
 sky130_fd_sc_hd__mux2_1 _5610_ (.A0(_1607_),
    .A1(net1000),
    .S(_1789_),
    .X(_1791_));
 sky130_fd_sc_hd__clkbuf_1 _5611_ (.A(_1791_),
    .X(_0186_));
 sky130_fd_sc_hd__mux2_1 _5612_ (.A0(_1611_),
    .A1(net1041),
    .S(_1789_),
    .X(_1792_));
 sky130_fd_sc_hd__clkbuf_1 _5613_ (.A(net1042),
    .X(_0187_));
 sky130_fd_sc_hd__mux2_1 _5614_ (.A0(_1615_),
    .A1(net905),
    .S(_1789_),
    .X(_1793_));
 sky130_fd_sc_hd__clkbuf_1 _5615_ (.A(_1793_),
    .X(_0188_));
 sky130_fd_sc_hd__mux2_1 _5616_ (.A0(_1618_),
    .A1(net675),
    .S(_1789_),
    .X(_1794_));
 sky130_fd_sc_hd__clkbuf_1 _5617_ (.A(net676),
    .X(_0189_));
 sky130_fd_sc_hd__and2_2 _5618_ (.A(_1076_),
    .B(_1724_),
    .X(_1795_));
 sky130_fd_sc_hd__mux2_1 _5619_ (.A0(net1429),
    .A1(_1732_),
    .S(_1795_),
    .X(_1796_));
 sky130_fd_sc_hd__clkbuf_1 _5620_ (.A(_1796_),
    .X(_0190_));
 sky130_fd_sc_hd__mux2_1 _5621_ (.A0(net1031),
    .A1(_1778_),
    .S(_1795_),
    .X(_1797_));
 sky130_fd_sc_hd__clkbuf_1 _5622_ (.A(_1797_),
    .X(_0191_));
 sky130_fd_sc_hd__mux2_1 _5623_ (.A0(net1116),
    .A1(_1664_),
    .S(_1795_),
    .X(_1798_));
 sky130_fd_sc_hd__clkbuf_1 _5624_ (.A(_1798_),
    .X(_0192_));
 sky130_fd_sc_hd__mux2_1 _5625_ (.A0(net941),
    .A1(_1666_),
    .S(_1795_),
    .X(_1799_));
 sky130_fd_sc_hd__clkbuf_1 _5626_ (.A(_1799_),
    .X(_0193_));
 sky130_fd_sc_hd__mux2_1 _5627_ (.A0(net1128),
    .A1(_1669_),
    .S(_1795_),
    .X(_1800_));
 sky130_fd_sc_hd__clkbuf_1 _5628_ (.A(_1800_),
    .X(_0194_));
 sky130_fd_sc_hd__buf_4 _5629_ (.A(_1597_),
    .X(_1801_));
 sky130_fd_sc_hd__nand2_4 _5630_ (.A(_1154_),
    .B(_1739_),
    .Y(_1802_));
 sky130_fd_sc_hd__mux2_1 _5631_ (.A0(_1801_),
    .A1(net1355),
    .S(_1802_),
    .X(_1803_));
 sky130_fd_sc_hd__clkbuf_1 _5632_ (.A(_1803_),
    .X(_0195_));
 sky130_fd_sc_hd__buf_4 _5633_ (.A(_1606_),
    .X(_1804_));
 sky130_fd_sc_hd__mux2_1 _5634_ (.A0(_1804_),
    .A1(net1234),
    .S(_1802_),
    .X(_1805_));
 sky130_fd_sc_hd__clkbuf_1 _5635_ (.A(_1805_),
    .X(_0196_));
 sky130_fd_sc_hd__mux2_1 _5636_ (.A0(_1611_),
    .A1(net1007),
    .S(_1802_),
    .X(_1806_));
 sky130_fd_sc_hd__clkbuf_1 _5637_ (.A(net1008),
    .X(_0197_));
 sky130_fd_sc_hd__mux2_1 _5638_ (.A0(_1615_),
    .A1(net1178),
    .S(_1802_),
    .X(_1807_));
 sky130_fd_sc_hd__clkbuf_1 _5639_ (.A(net1179),
    .X(_0198_));
 sky130_fd_sc_hd__mux2_1 _5640_ (.A0(_1618_),
    .A1(net834),
    .S(_1802_),
    .X(_1808_));
 sky130_fd_sc_hd__clkbuf_1 _5641_ (.A(net835),
    .X(_0199_));
 sky130_fd_sc_hd__nand2_4 _5642_ (.A(_1135_),
    .B(_1739_),
    .Y(_1809_));
 sky130_fd_sc_hd__mux2_1 _5643_ (.A0(_1801_),
    .A1(net1336),
    .S(_1809_),
    .X(_1810_));
 sky130_fd_sc_hd__clkbuf_1 _5644_ (.A(_1810_),
    .X(_0200_));
 sky130_fd_sc_hd__mux2_1 _5645_ (.A0(_1804_),
    .A1(net945),
    .S(_1809_),
    .X(_1811_));
 sky130_fd_sc_hd__clkbuf_1 _5646_ (.A(_1811_),
    .X(_0201_));
 sky130_fd_sc_hd__buf_4 _5647_ (.A(_1610_),
    .X(_1812_));
 sky130_fd_sc_hd__mux2_1 _5648_ (.A0(_1812_),
    .A1(net1078),
    .S(_1809_),
    .X(_1813_));
 sky130_fd_sc_hd__clkbuf_1 _5649_ (.A(_1813_),
    .X(_0202_));
 sky130_fd_sc_hd__buf_4 _5650_ (.A(_1614_),
    .X(_1814_));
 sky130_fd_sc_hd__mux2_1 _5651_ (.A0(_1814_),
    .A1(net894),
    .S(_1809_),
    .X(_1815_));
 sky130_fd_sc_hd__clkbuf_1 _5652_ (.A(_1815_),
    .X(_0203_));
 sky130_fd_sc_hd__buf_4 _5653_ (.A(net530),
    .X(_1816_));
 sky130_fd_sc_hd__mux2_1 _5654_ (.A0(_1816_),
    .A1(net668),
    .S(_1809_),
    .X(_1817_));
 sky130_fd_sc_hd__clkbuf_1 _5655_ (.A(net669),
    .X(_0204_));
 sky130_fd_sc_hd__and2_2 _5656_ (.A(_1095_),
    .B(_1724_),
    .X(_1818_));
 sky130_fd_sc_hd__mux2_1 _5657_ (.A0(net1436),
    .A1(_1732_),
    .S(_1818_),
    .X(_1819_));
 sky130_fd_sc_hd__clkbuf_1 _5658_ (.A(_1819_),
    .X(_0205_));
 sky130_fd_sc_hd__mux2_1 _5659_ (.A0(net1248),
    .A1(_1778_),
    .S(_1818_),
    .X(_1820_));
 sky130_fd_sc_hd__clkbuf_1 _5660_ (.A(_1820_),
    .X(_0206_));
 sky130_fd_sc_hd__mux2_1 _5661_ (.A0(net1123),
    .A1(_1664_),
    .S(_1818_),
    .X(_1821_));
 sky130_fd_sc_hd__clkbuf_1 _5662_ (.A(_1821_),
    .X(_0207_));
 sky130_fd_sc_hd__mux2_1 _5663_ (.A0(net927),
    .A1(_1666_),
    .S(_1818_),
    .X(_1822_));
 sky130_fd_sc_hd__clkbuf_1 _5664_ (.A(_1822_),
    .X(_0208_));
 sky130_fd_sc_hd__mux2_1 _5665_ (.A0(net1168),
    .A1(_1669_),
    .S(_1818_),
    .X(_1823_));
 sky130_fd_sc_hd__clkbuf_1 _5666_ (.A(_1823_),
    .X(_0209_));
 sky130_fd_sc_hd__nand2_2 _5667_ (.A(_1144_),
    .B(_1739_),
    .Y(_1824_));
 sky130_fd_sc_hd__mux2_1 _5668_ (.A0(_1801_),
    .A1(net1353),
    .S(_1824_),
    .X(_1825_));
 sky130_fd_sc_hd__clkbuf_1 _5669_ (.A(_1825_),
    .X(_0210_));
 sky130_fd_sc_hd__mux2_1 _5670_ (.A0(_1804_),
    .A1(net950),
    .S(_1824_),
    .X(_1826_));
 sky130_fd_sc_hd__clkbuf_1 _5671_ (.A(_1826_),
    .X(_0211_));
 sky130_fd_sc_hd__mux2_1 _5672_ (.A0(_1812_),
    .A1(net1083),
    .S(_1824_),
    .X(_1827_));
 sky130_fd_sc_hd__clkbuf_1 _5673_ (.A(_1827_),
    .X(_0212_));
 sky130_fd_sc_hd__mux2_1 _5674_ (.A0(_1814_),
    .A1(net901),
    .S(_1824_),
    .X(_1828_));
 sky130_fd_sc_hd__clkbuf_1 _5675_ (.A(_1828_),
    .X(_0213_));
 sky130_fd_sc_hd__mux2_1 _5676_ (.A0(_1816_),
    .A1(net627),
    .S(_1824_),
    .X(_1829_));
 sky130_fd_sc_hd__clkbuf_1 _5677_ (.A(net628),
    .X(_0214_));
 sky130_fd_sc_hd__and2_2 _5678_ (.A(_1081_),
    .B(_1724_),
    .X(_1830_));
 sky130_fd_sc_hd__mux2_1 _5679_ (.A0(net1424),
    .A1(_1732_),
    .S(_1830_),
    .X(_1831_));
 sky130_fd_sc_hd__clkbuf_1 _5680_ (.A(_1831_),
    .X(_0215_));
 sky130_fd_sc_hd__mux2_1 _5681_ (.A0(net1094),
    .A1(_1778_),
    .S(_1830_),
    .X(_1832_));
 sky130_fd_sc_hd__clkbuf_1 _5682_ (.A(_1832_),
    .X(_0216_));
 sky130_fd_sc_hd__clkbuf_4 _5683_ (.A(_1610_),
    .X(_1833_));
 sky130_fd_sc_hd__mux2_1 _5684_ (.A0(net1111),
    .A1(_1833_),
    .S(_1830_),
    .X(_1834_));
 sky130_fd_sc_hd__clkbuf_1 _5685_ (.A(_1834_),
    .X(_0217_));
 sky130_fd_sc_hd__buf_6 _5686_ (.A(net551),
    .X(_1835_));
 sky130_fd_sc_hd__clkbuf_4 _5687_ (.A(net552),
    .X(_1836_));
 sky130_fd_sc_hd__mux2_1 _5688_ (.A0(net911),
    .A1(_1836_),
    .S(_1830_),
    .X(_1837_));
 sky130_fd_sc_hd__clkbuf_1 _5689_ (.A(_1837_),
    .X(_0218_));
 sky130_fd_sc_hd__buf_4 _5690_ (.A(_1668_),
    .X(_1838_));
 sky130_fd_sc_hd__mux2_1 _5691_ (.A0(net1022),
    .A1(_1838_),
    .S(_1830_),
    .X(_1839_));
 sky130_fd_sc_hd__clkbuf_1 _5692_ (.A(_1839_),
    .X(_0219_));
 sky130_fd_sc_hd__nand2_4 _5693_ (.A(_1088_),
    .B(_1739_),
    .Y(_1840_));
 sky130_fd_sc_hd__mux2_1 _5694_ (.A0(_1801_),
    .A1(net1378),
    .S(_1840_),
    .X(_1841_));
 sky130_fd_sc_hd__clkbuf_1 _5695_ (.A(_1841_),
    .X(_0220_));
 sky130_fd_sc_hd__mux2_1 _5696_ (.A0(_1804_),
    .A1(net972),
    .S(_1840_),
    .X(_1842_));
 sky130_fd_sc_hd__clkbuf_1 _5697_ (.A(_1842_),
    .X(_0221_));
 sky130_fd_sc_hd__mux2_1 _5698_ (.A0(_1812_),
    .A1(net1084),
    .S(_1840_),
    .X(_1843_));
 sky130_fd_sc_hd__clkbuf_1 _5699_ (.A(_1843_),
    .X(_0222_));
 sky130_fd_sc_hd__mux2_1 _5700_ (.A0(_1814_),
    .A1(net902),
    .S(_1840_),
    .X(_1844_));
 sky130_fd_sc_hd__clkbuf_1 _5701_ (.A(_1844_),
    .X(_0223_));
 sky130_fd_sc_hd__mux2_1 _5702_ (.A0(_1816_),
    .A1(net677),
    .S(_1840_),
    .X(_1845_));
 sky130_fd_sc_hd__clkbuf_1 _5703_ (.A(net678),
    .X(_0224_));
 sky130_fd_sc_hd__and2_2 _5704_ (.A(_1145_),
    .B(_1724_),
    .X(_1846_));
 sky130_fd_sc_hd__mux2_1 _5705_ (.A0(net1409),
    .A1(_1732_),
    .S(_1846_),
    .X(_1847_));
 sky130_fd_sc_hd__clkbuf_1 _5706_ (.A(_1847_),
    .X(_0225_));
 sky130_fd_sc_hd__mux2_1 _5707_ (.A0(net1089),
    .A1(_1778_),
    .S(_1846_),
    .X(_1848_));
 sky130_fd_sc_hd__clkbuf_1 _5708_ (.A(_1848_),
    .X(_0226_));
 sky130_fd_sc_hd__mux2_1 _5709_ (.A0(net1169),
    .A1(_1833_),
    .S(_1846_),
    .X(_1849_));
 sky130_fd_sc_hd__clkbuf_1 _5710_ (.A(_1849_),
    .X(_0227_));
 sky130_fd_sc_hd__mux2_1 _5711_ (.A0(net1011),
    .A1(_1836_),
    .S(_1846_),
    .X(_1850_));
 sky130_fd_sc_hd__clkbuf_1 _5712_ (.A(_1850_),
    .X(_0228_));
 sky130_fd_sc_hd__mux2_1 _5713_ (.A0(net1122),
    .A1(_1838_),
    .S(_1846_),
    .X(_1851_));
 sky130_fd_sc_hd__clkbuf_1 _5714_ (.A(_1851_),
    .X(_0229_));
 sky130_fd_sc_hd__and2_2 _5715_ (.A(_1122_),
    .B(_1724_),
    .X(_1852_));
 sky130_fd_sc_hd__mux2_1 _5716_ (.A0(net1447),
    .A1(_1732_),
    .S(_1852_),
    .X(_1853_));
 sky130_fd_sc_hd__clkbuf_1 _5717_ (.A(_1853_),
    .X(_0230_));
 sky130_fd_sc_hd__mux2_1 _5718_ (.A0(net1302),
    .A1(_1778_),
    .S(_1852_),
    .X(_1854_));
 sky130_fd_sc_hd__clkbuf_1 _5719_ (.A(_1854_),
    .X(_0231_));
 sky130_fd_sc_hd__mux2_1 _5720_ (.A0(net1044),
    .A1(_1833_),
    .S(_1852_),
    .X(_1855_));
 sky130_fd_sc_hd__clkbuf_1 _5721_ (.A(net1045),
    .X(_0232_));
 sky130_fd_sc_hd__mux2_1 _5722_ (.A0(net1184),
    .A1(_1836_),
    .S(_1852_),
    .X(_1856_));
 sky130_fd_sc_hd__clkbuf_1 _5723_ (.A(_1856_),
    .X(_0233_));
 sky130_fd_sc_hd__mux2_1 _5724_ (.A0(net991),
    .A1(_1838_),
    .S(_1852_),
    .X(_1857_));
 sky130_fd_sc_hd__clkbuf_1 _5725_ (.A(_1857_),
    .X(_0234_));
 sky130_fd_sc_hd__buf_12 _5726_ (.A(net526),
    .X(_1858_));
 sky130_fd_sc_hd__nand2_4 _5727_ (.A(_1065_),
    .B(_1858_),
    .Y(_1859_));
 sky130_fd_sc_hd__mux2_1 _5728_ (.A0(_1801_),
    .A1(net1337),
    .S(_1859_),
    .X(_1860_));
 sky130_fd_sc_hd__clkbuf_1 _5729_ (.A(_1860_),
    .X(_0235_));
 sky130_fd_sc_hd__mux2_1 _5730_ (.A0(_1804_),
    .A1(net961),
    .S(_1859_),
    .X(_1861_));
 sky130_fd_sc_hd__clkbuf_1 _5731_ (.A(_1861_),
    .X(_0236_));
 sky130_fd_sc_hd__mux2_1 _5732_ (.A0(_1812_),
    .A1(net1103),
    .S(_1859_),
    .X(_1862_));
 sky130_fd_sc_hd__clkbuf_1 _5733_ (.A(_1862_),
    .X(_0237_));
 sky130_fd_sc_hd__mux2_1 _5734_ (.A0(_1814_),
    .A1(net896),
    .S(_1859_),
    .X(_1863_));
 sky130_fd_sc_hd__clkbuf_1 _5735_ (.A(_1863_),
    .X(_0238_));
 sky130_fd_sc_hd__mux2_1 _5736_ (.A0(_1816_),
    .A1(net629),
    .S(_1859_),
    .X(_1864_));
 sky130_fd_sc_hd__clkbuf_1 _5737_ (.A(net630),
    .X(_0239_));
 sky130_fd_sc_hd__nand2_4 _5738_ (.A(_1115_),
    .B(_1858_),
    .Y(_1865_));
 sky130_fd_sc_hd__mux2_1 _5739_ (.A0(_1801_),
    .A1(net1375),
    .S(_1865_),
    .X(_1866_));
 sky130_fd_sc_hd__clkbuf_1 _5740_ (.A(_1866_),
    .X(_0240_));
 sky130_fd_sc_hd__mux2_1 _5741_ (.A0(_1804_),
    .A1(net1356),
    .S(_1865_),
    .X(_1867_));
 sky130_fd_sc_hd__clkbuf_1 _5742_ (.A(_1867_),
    .X(_0241_));
 sky130_fd_sc_hd__mux2_1 _5743_ (.A0(_1812_),
    .A1(net1317),
    .S(_1865_),
    .X(_1868_));
 sky130_fd_sc_hd__clkbuf_1 _5744_ (.A(_1868_),
    .X(_0242_));
 sky130_fd_sc_hd__mux2_1 _5745_ (.A0(_1814_),
    .A1(net1216),
    .S(_1865_),
    .X(_1869_));
 sky130_fd_sc_hd__clkbuf_1 _5746_ (.A(_1869_),
    .X(_0243_));
 sky130_fd_sc_hd__mux2_1 _5747_ (.A0(_1816_),
    .A1(net842),
    .S(_1865_),
    .X(_1870_));
 sky130_fd_sc_hd__clkbuf_1 _5748_ (.A(net1666),
    .X(_0244_));
 sky130_fd_sc_hd__buf_4 _5749_ (.A(net525),
    .X(_1871_));
 sky130_fd_sc_hd__and2_4 _5750_ (.A(_1099_),
    .B(_1871_),
    .X(_1872_));
 sky130_fd_sc_hd__mux2_1 _5751_ (.A0(net1376),
    .A1(_1732_),
    .S(_1872_),
    .X(_1873_));
 sky130_fd_sc_hd__clkbuf_1 _5752_ (.A(_1873_),
    .X(_0245_));
 sky130_fd_sc_hd__mux2_1 _5753_ (.A0(net973),
    .A1(_1778_),
    .S(_1872_),
    .X(_1874_));
 sky130_fd_sc_hd__clkbuf_1 _5754_ (.A(_1874_),
    .X(_0246_));
 sky130_fd_sc_hd__mux2_1 _5755_ (.A0(net1075),
    .A1(_1833_),
    .S(_1872_),
    .X(_1875_));
 sky130_fd_sc_hd__clkbuf_1 _5756_ (.A(_1875_),
    .X(_0247_));
 sky130_fd_sc_hd__mux2_1 _5757_ (.A0(net919),
    .A1(_1836_),
    .S(_1872_),
    .X(_1876_));
 sky130_fd_sc_hd__clkbuf_1 _5758_ (.A(_1876_),
    .X(_0248_));
 sky130_fd_sc_hd__mux2_1 _5759_ (.A0(net1148),
    .A1(_1838_),
    .S(_1872_),
    .X(_1877_));
 sky130_fd_sc_hd__clkbuf_1 _5760_ (.A(_1877_),
    .X(_0249_));
 sky130_fd_sc_hd__buf_4 _5761_ (.A(_1731_),
    .X(_1878_));
 sky130_fd_sc_hd__and2_2 _5762_ (.A(_1092_),
    .B(_1871_),
    .X(_1879_));
 sky130_fd_sc_hd__mux2_1 _5763_ (.A0(net1398),
    .A1(_1878_),
    .S(_1879_),
    .X(_1880_));
 sky130_fd_sc_hd__clkbuf_1 _5764_ (.A(_1880_),
    .X(_0250_));
 sky130_fd_sc_hd__mux2_1 _5765_ (.A0(net1059),
    .A1(_1778_),
    .S(_1879_),
    .X(_1881_));
 sky130_fd_sc_hd__clkbuf_1 _5766_ (.A(_1881_),
    .X(_0251_));
 sky130_fd_sc_hd__mux2_1 _5767_ (.A0(net1125),
    .A1(_1833_),
    .S(_1879_),
    .X(_1882_));
 sky130_fd_sc_hd__clkbuf_1 _5768_ (.A(_1882_),
    .X(_0252_));
 sky130_fd_sc_hd__mux2_1 _5769_ (.A0(net913),
    .A1(_1836_),
    .S(_1879_),
    .X(_1883_));
 sky130_fd_sc_hd__clkbuf_1 _5770_ (.A(_1883_),
    .X(_0253_));
 sky130_fd_sc_hd__mux2_1 _5771_ (.A0(net1141),
    .A1(_1838_),
    .S(_1879_),
    .X(_1884_));
 sky130_fd_sc_hd__clkbuf_1 _5772_ (.A(_1884_),
    .X(_0254_));
 sky130_fd_sc_hd__nand2_4 _5773_ (.A(_1105_),
    .B(_1858_),
    .Y(_1885_));
 sky130_fd_sc_hd__mux2_1 _5774_ (.A0(_1801_),
    .A1(net1386),
    .S(_1885_),
    .X(_1886_));
 sky130_fd_sc_hd__clkbuf_1 _5775_ (.A(_1886_),
    .X(_0255_));
 sky130_fd_sc_hd__mux2_1 _5776_ (.A0(_1804_),
    .A1(net964),
    .S(_1885_),
    .X(_1887_));
 sky130_fd_sc_hd__clkbuf_1 _5777_ (.A(_1887_),
    .X(_0256_));
 sky130_fd_sc_hd__mux2_1 _5778_ (.A0(_1812_),
    .A1(net1121),
    .S(_1885_),
    .X(_1888_));
 sky130_fd_sc_hd__clkbuf_1 _5779_ (.A(_1888_),
    .X(_0257_));
 sky130_fd_sc_hd__mux2_1 _5780_ (.A0(_1814_),
    .A1(net910),
    .S(_1885_),
    .X(_1889_));
 sky130_fd_sc_hd__clkbuf_1 _5781_ (.A(_1889_),
    .X(_0258_));
 sky130_fd_sc_hd__mux2_1 _5782_ (.A0(_1816_),
    .A1(net635),
    .S(_1885_),
    .X(_1890_));
 sky130_fd_sc_hd__clkbuf_1 _5783_ (.A(net636),
    .X(_0259_));
 sky130_fd_sc_hd__and2_2 _5784_ (.A(_1112_),
    .B(_1871_),
    .X(_1891_));
 sky130_fd_sc_hd__mux2_1 _5785_ (.A0(net1421),
    .A1(_1878_),
    .S(_1891_),
    .X(_1892_));
 sky130_fd_sc_hd__clkbuf_1 _5786_ (.A(_1892_),
    .X(_0260_));
 sky130_fd_sc_hd__mux2_1 _5787_ (.A0(net1274),
    .A1(_1778_),
    .S(_1891_),
    .X(_1893_));
 sky130_fd_sc_hd__clkbuf_1 _5788_ (.A(_1893_),
    .X(_0261_));
 sky130_fd_sc_hd__mux2_1 _5789_ (.A0(net1315),
    .A1(_1833_),
    .S(_1891_),
    .X(_1894_));
 sky130_fd_sc_hd__clkbuf_1 _5790_ (.A(_1894_),
    .X(_0262_));
 sky130_fd_sc_hd__mux2_1 _5791_ (.A0(net1218),
    .A1(_1836_),
    .S(_1891_),
    .X(_1895_));
 sky130_fd_sc_hd__clkbuf_1 _5792_ (.A(_1895_),
    .X(_0263_));
 sky130_fd_sc_hd__mux2_1 _5793_ (.A0(net1147),
    .A1(_1838_),
    .S(_1891_),
    .X(_1896_));
 sky130_fd_sc_hd__clkbuf_1 _5794_ (.A(_1896_),
    .X(_0264_));
 sky130_fd_sc_hd__nand2_4 _5795_ (.A(_1077_),
    .B(_1858_),
    .Y(_1897_));
 sky130_fd_sc_hd__mux2_1 _5796_ (.A0(_1801_),
    .A1(net1388),
    .S(_1897_),
    .X(_1898_));
 sky130_fd_sc_hd__clkbuf_1 _5797_ (.A(_1898_),
    .X(_0265_));
 sky130_fd_sc_hd__mux2_1 _5798_ (.A0(_1804_),
    .A1(net960),
    .S(_1897_),
    .X(_1899_));
 sky130_fd_sc_hd__clkbuf_1 _5799_ (.A(_1899_),
    .X(_0266_));
 sky130_fd_sc_hd__mux2_1 _5800_ (.A0(_1812_),
    .A1(net1088),
    .S(_1897_),
    .X(_1900_));
 sky130_fd_sc_hd__clkbuf_1 _5801_ (.A(_1900_),
    .X(_0267_));
 sky130_fd_sc_hd__mux2_1 _5802_ (.A0(_1814_),
    .A1(net912),
    .S(_1897_),
    .X(_1901_));
 sky130_fd_sc_hd__clkbuf_1 _5803_ (.A(_1901_),
    .X(_0268_));
 sky130_fd_sc_hd__mux2_1 _5804_ (.A0(_1816_),
    .A1(net679),
    .S(_1897_),
    .X(_1902_));
 sky130_fd_sc_hd__clkbuf_1 _5805_ (.A(net680),
    .X(_0269_));
 sky130_fd_sc_hd__and2_2 _5806_ (.A(_1078_),
    .B(_1871_),
    .X(_1903_));
 sky130_fd_sc_hd__mux2_1 _5807_ (.A0(net1401),
    .A1(_1878_),
    .S(_1903_),
    .X(_1904_));
 sky130_fd_sc_hd__clkbuf_1 _5808_ (.A(_1904_),
    .X(_0270_));
 sky130_fd_sc_hd__buf_6 _5809_ (.A(_1606_),
    .X(_1905_));
 sky130_fd_sc_hd__mux2_1 _5810_ (.A0(net1032),
    .A1(_1905_),
    .S(_1903_),
    .X(_1906_));
 sky130_fd_sc_hd__clkbuf_1 _5811_ (.A(_1906_),
    .X(_0271_));
 sky130_fd_sc_hd__mux2_1 _5812_ (.A0(net1112),
    .A1(_1833_),
    .S(_1903_),
    .X(_1907_));
 sky130_fd_sc_hd__clkbuf_1 _5813_ (.A(_1907_),
    .X(_0272_));
 sky130_fd_sc_hd__mux2_1 _5814_ (.A0(net942),
    .A1(_1836_),
    .S(_1903_),
    .X(_1908_));
 sky130_fd_sc_hd__clkbuf_1 _5815_ (.A(_1908_),
    .X(_0273_));
 sky130_fd_sc_hd__mux2_1 _5816_ (.A0(net1154),
    .A1(_1838_),
    .S(_1903_),
    .X(_1909_));
 sky130_fd_sc_hd__clkbuf_1 _5817_ (.A(_1909_),
    .X(_0274_));
 sky130_fd_sc_hd__mux2_1 _5818_ (.A0(net1334),
    .A1(_1597_),
    .S(_1053_),
    .X(_1910_));
 sky130_fd_sc_hd__and2b_1 _5819_ (.A_N(_1507_),
    .B(net372),
    .X(_1911_));
 sky130_fd_sc_hd__buf_12 _5820_ (.A(_1601_),
    .X(_1912_));
 sky130_fd_sc_hd__o221a_4 _5821_ (.A1(_0964_),
    .A2(_1507_),
    .B1(_1911_),
    .B2(_1053_),
    .C1(_1912_),
    .X(_1913_));
 sky130_fd_sc_hd__mux2_1 _5822_ (.A0(\mgmt_gpio_data[16] ),
    .A1(_1910_),
    .S(net549),
    .X(_1914_));
 sky130_fd_sc_hd__clkbuf_1 _5823_ (.A(net1569),
    .X(_0275_));
 sky130_fd_sc_hd__mux2_1 _5824_ (.A0(net977),
    .A1(net543),
    .S(_1053_),
    .X(_1915_));
 sky130_fd_sc_hd__mux2_1 _5825_ (.A0(\mgmt_gpio_data[17] ),
    .A1(_1915_),
    .S(net549),
    .X(_1916_));
 sky130_fd_sc_hd__clkbuf_1 _5826_ (.A(net1567),
    .X(_0276_));
 sky130_fd_sc_hd__mux2_1 _5827_ (.A0(net962),
    .A1(_1610_),
    .S(_1053_),
    .X(_1917_));
 sky130_fd_sc_hd__mux2_1 _5828_ (.A0(\mgmt_gpio_data[18] ),
    .A1(_1917_),
    .S(net549),
    .X(_1918_));
 sky130_fd_sc_hd__clkbuf_1 _5829_ (.A(net1565),
    .X(_0277_));
 sky130_fd_sc_hd__mux2_1 _5830_ (.A0(net889),
    .A1(_1614_),
    .S(_1053_),
    .X(_1919_));
 sky130_fd_sc_hd__mux2_1 _5831_ (.A0(\mgmt_gpio_data[19] ),
    .A1(_1919_),
    .S(net549),
    .X(_1920_));
 sky130_fd_sc_hd__clkbuf_1 _5832_ (.A(net1587),
    .X(_0278_));
 sky130_fd_sc_hd__mux2_1 _5833_ (.A0(\mgmt_gpio_data_buf[20] ),
    .A1(net530),
    .S(_1053_),
    .X(_1921_));
 sky130_fd_sc_hd__mux2_1 _5834_ (.A0(\mgmt_gpio_data[20] ),
    .A1(net531),
    .S(net549),
    .X(_1922_));
 sky130_fd_sc_hd__clkbuf_1 _5835_ (.A(net1585),
    .X(_0279_));
 sky130_fd_sc_hd__mux2_1 _5836_ (.A0(net1322),
    .A1(net521),
    .S(_1053_),
    .X(_1923_));
 sky130_fd_sc_hd__mux2_1 _5837_ (.A0(\mgmt_gpio_data[21] ),
    .A1(_1923_),
    .S(net549),
    .X(_1924_));
 sky130_fd_sc_hd__clkbuf_1 _5838_ (.A(net1583),
    .X(_0280_));
 sky130_fd_sc_hd__mux2_1 _5839_ (.A0(net1327),
    .A1(net533),
    .S(_1053_),
    .X(_1925_));
 sky130_fd_sc_hd__mux2_1 _5840_ (.A0(\mgmt_gpio_data[22] ),
    .A1(_1925_),
    .S(net549),
    .X(_1926_));
 sky130_fd_sc_hd__clkbuf_1 _5841_ (.A(net1571),
    .X(_0281_));
 sky130_fd_sc_hd__mux2_1 _5842_ (.A0(\mgmt_gpio_data_buf[23] ),
    .A1(net511),
    .S(_1053_),
    .X(_1927_));
 sky130_fd_sc_hd__mux2_1 _5843_ (.A0(\mgmt_gpio_data[23] ),
    .A1(net512),
    .S(net549),
    .X(_1928_));
 sky130_fd_sc_hd__clkbuf_1 _5844_ (.A(net1589),
    .X(_0282_));
 sky130_fd_sc_hd__mux2_1 _5845_ (.A0(net1344),
    .A1(_1597_),
    .S(_0911_),
    .X(_1929_));
 sky130_fd_sc_hd__o221a_4 _5846_ (.A1(_0875_),
    .A2(_1507_),
    .B1(_1911_),
    .B2(_0911_),
    .C1(_1912_),
    .X(_1930_));
 sky130_fd_sc_hd__mux2_1 _5847_ (.A0(\mgmt_gpio_data[8] ),
    .A1(_1929_),
    .S(_1930_),
    .X(_1931_));
 sky130_fd_sc_hd__clkbuf_1 _5848_ (.A(net1383),
    .X(_0283_));
 sky130_fd_sc_hd__mux2_1 _5849_ (.A0(\mgmt_gpio_data_buf[9] ),
    .A1(net543),
    .S(_0911_),
    .X(_1932_));
 sky130_fd_sc_hd__mux2_1 _5850_ (.A0(\mgmt_gpio_data[9] ),
    .A1(net544),
    .S(_1930_),
    .X(_1933_));
 sky130_fd_sc_hd__clkbuf_1 _5851_ (.A(net1581),
    .X(_0284_));
 sky130_fd_sc_hd__mux2_1 _5852_ (.A0(net1012),
    .A1(net518),
    .S(_0911_),
    .X(_1934_));
 sky130_fd_sc_hd__mux2_1 _5853_ (.A0(\mgmt_gpio_data[10] ),
    .A1(_1934_),
    .S(_1930_),
    .X(_1935_));
 sky130_fd_sc_hd__clkbuf_1 _5854_ (.A(net1546),
    .X(_0285_));
 sky130_fd_sc_hd__mux2_1 _5855_ (.A0(\mgmt_gpio_data_buf[11] ),
    .A1(_1614_),
    .S(_0911_),
    .X(_1936_));
 sky130_fd_sc_hd__mux2_1 _5856_ (.A0(\mgmt_gpio_data[11] ),
    .A1(_1936_),
    .S(_1930_),
    .X(_1937_));
 sky130_fd_sc_hd__clkbuf_1 _5857_ (.A(net717),
    .X(_0286_));
 sky130_fd_sc_hd__mux2_1 _5858_ (.A0(net643),
    .A1(net530),
    .S(_0911_),
    .X(_1938_));
 sky130_fd_sc_hd__mux2_1 _5859_ (.A0(\mgmt_gpio_data[12] ),
    .A1(_1938_),
    .S(_1930_),
    .X(_1939_));
 sky130_fd_sc_hd__clkbuf_1 _5860_ (.A(net1544),
    .X(_0287_));
 sky130_fd_sc_hd__mux2_1 _5861_ (.A0(\mgmt_gpio_data_buf[13] ),
    .A1(net521),
    .S(_0911_),
    .X(_1940_));
 sky130_fd_sc_hd__mux2_1 _5862_ (.A0(\mgmt_gpio_data[13] ),
    .A1(net522),
    .S(_1930_),
    .X(_1941_));
 sky130_fd_sc_hd__clkbuf_1 _5863_ (.A(net1575),
    .X(_0288_));
 sky130_fd_sc_hd__mux2_1 _5864_ (.A0(\mgmt_gpio_data_buf[14] ),
    .A1(net533),
    .S(_0911_),
    .X(_1942_));
 sky130_fd_sc_hd__mux2_1 _5865_ (.A0(\mgmt_gpio_data[14] ),
    .A1(net534),
    .S(_1930_),
    .X(_1943_));
 sky130_fd_sc_hd__clkbuf_1 _5866_ (.A(net1577),
    .X(_0289_));
 sky130_fd_sc_hd__mux2_1 _5867_ (.A0(net975),
    .A1(net511),
    .S(_0911_),
    .X(_1944_));
 sky130_fd_sc_hd__mux2_1 _5868_ (.A0(\mgmt_gpio_data[15] ),
    .A1(_1944_),
    .S(_1930_),
    .X(_1945_));
 sky130_fd_sc_hd__clkbuf_1 _5869_ (.A(net1539),
    .X(_0290_));
 sky130_fd_sc_hd__or4_1 _5870_ (.A(net1448),
    .B(net1487),
    .C(net1464),
    .D(net1473),
    .X(_1946_));
 sky130_fd_sc_hd__or3_4 _5871_ (.A(net1521),
    .B(net1538),
    .C(\wbbd_state[9] ),
    .X(_1947_));
 sky130_fd_sc_hd__or2_1 _5872_ (.A(\wbbd_state[5] ),
    .B(_1947_),
    .X(_1948_));
 sky130_fd_sc_hd__clkbuf_4 _5873_ (.A(_1948_),
    .X(_1949_));
 sky130_fd_sc_hd__a2111o_4 _5874_ (.A1(_1584_),
    .A2(_1539_),
    .B1(net1498),
    .C1(_1946_),
    .D1(_1949_),
    .X(_0291_));
 sky130_fd_sc_hd__mux2_1 _5875_ (.A0(net1320),
    .A1(_1597_),
    .S(_1279_),
    .X(_1950_));
 sky130_fd_sc_hd__o221a_4 _5876_ (.A1(_0940_),
    .A2(_1507_),
    .B1(_1911_),
    .B2(_1279_),
    .C1(_1912_),
    .X(_1951_));
 sky130_fd_sc_hd__mux2_1 _5877_ (.A0(\mgmt_gpio_data[0] ),
    .A1(_1950_),
    .S(_1951_),
    .X(_1952_));
 sky130_fd_sc_hd__clkbuf_1 _5878_ (.A(net1402),
    .X(_0292_));
 sky130_fd_sc_hd__mux2_1 _5879_ (.A0(\mgmt_gpio_data_buf[1] ),
    .A1(net543),
    .S(_1279_),
    .X(_1953_));
 sky130_fd_sc_hd__mux2_1 _5880_ (.A0(\mgmt_gpio_data[1] ),
    .A1(net576),
    .S(_1951_),
    .X(_1954_));
 sky130_fd_sc_hd__clkbuf_1 _5881_ (.A(net1573),
    .X(_0293_));
 sky130_fd_sc_hd__mux2_1 _5882_ (.A0(\mgmt_gpio_data_buf[2] ),
    .A1(net518),
    .S(_1279_),
    .X(_1955_));
 sky130_fd_sc_hd__mux2_1 _5883_ (.A0(\mgmt_gpio_data[2] ),
    .A1(net519),
    .S(_1951_),
    .X(_1956_));
 sky130_fd_sc_hd__clkbuf_1 _5884_ (.A(net1548),
    .X(_0294_));
 sky130_fd_sc_hd__mux2_1 _5885_ (.A0(\mgmt_gpio_data_buf[3] ),
    .A1(_1614_),
    .S(_1279_),
    .X(_1957_));
 sky130_fd_sc_hd__mux2_1 _5886_ (.A0(\mgmt_gpio_data[3] ),
    .A1(net705),
    .S(_1951_),
    .X(_1958_));
 sky130_fd_sc_hd__clkbuf_1 _5887_ (.A(net706),
    .X(_0295_));
 sky130_fd_sc_hd__mux2_1 _5888_ (.A0(\mgmt_gpio_data_buf[4] ),
    .A1(net530),
    .S(_1279_),
    .X(_1959_));
 sky130_fd_sc_hd__mux2_1 _5889_ (.A0(\mgmt_gpio_data[4] ),
    .A1(net540),
    .S(_1951_),
    .X(_1960_));
 sky130_fd_sc_hd__clkbuf_1 _5890_ (.A(net1545),
    .X(_0296_));
 sky130_fd_sc_hd__mux2_1 _5891_ (.A0(net1145),
    .A1(net521),
    .S(_1279_),
    .X(_1961_));
 sky130_fd_sc_hd__mux2_1 _5892_ (.A0(\mgmt_gpio_data[5] ),
    .A1(_1961_),
    .S(_1951_),
    .X(_1962_));
 sky130_fd_sc_hd__clkbuf_1 _5893_ (.A(net1547),
    .X(_0297_));
 sky130_fd_sc_hd__mux2_1 _5894_ (.A0(\mgmt_gpio_data_buf[6] ),
    .A1(net533),
    .S(_1279_),
    .X(_1963_));
 sky130_fd_sc_hd__mux2_1 _5895_ (.A0(\mgmt_gpio_data[6] ),
    .A1(_1963_),
    .S(_1951_),
    .X(_1964_));
 sky130_fd_sc_hd__clkbuf_1 _5896_ (.A(net607),
    .X(_0298_));
 sky130_fd_sc_hd__mux2_1 _5897_ (.A0(net1073),
    .A1(net511),
    .S(_1279_),
    .X(_1965_));
 sky130_fd_sc_hd__mux2_1 _5898_ (.A0(\mgmt_gpio_data[7] ),
    .A1(_1965_),
    .S(_1951_),
    .X(_1966_));
 sky130_fd_sc_hd__clkbuf_1 _5899_ (.A(net1543),
    .X(_0299_));
 sky130_fd_sc_hd__buf_12 _5900_ (.A(_1601_),
    .X(_1967_));
 sky130_fd_sc_hd__nand2_4 _5901_ (.A(net372),
    .B(_1967_),
    .Y(_1968_));
 sky130_fd_sc_hd__mux2_1 _5902_ (.A0(_1801_),
    .A1(\mgmt_gpio_data[24] ),
    .S(_1968_),
    .X(_1969_));
 sky130_fd_sc_hd__clkbuf_1 _5903_ (.A(net1392),
    .X(_0300_));
 sky130_fd_sc_hd__mux2_1 _5904_ (.A0(_1804_),
    .A1(\mgmt_gpio_data[25] ),
    .S(_1968_),
    .X(_1970_));
 sky130_fd_sc_hd__clkbuf_1 _5905_ (.A(net947),
    .X(_0301_));
 sky130_fd_sc_hd__mux2_1 _5906_ (.A0(_1812_),
    .A1(\mgmt_gpio_data[26] ),
    .S(_1968_),
    .X(_1971_));
 sky130_fd_sc_hd__clkbuf_1 _5907_ (.A(net1029),
    .X(_0302_));
 sky130_fd_sc_hd__mux2_1 _5908_ (.A0(_1814_),
    .A1(\mgmt_gpio_data[27] ),
    .S(_1968_),
    .X(_1972_));
 sky130_fd_sc_hd__clkbuf_1 _5909_ (.A(net897),
    .X(_0303_));
 sky130_fd_sc_hd__mux2_1 _5910_ (.A0(_1816_),
    .A1(\mgmt_gpio_data[28] ),
    .S(_1968_),
    .X(_1973_));
 sky130_fd_sc_hd__clkbuf_1 _5911_ (.A(net659),
    .X(_0304_));
 sky130_fd_sc_hd__mux2_1 _5912_ (.A0(_1708_),
    .A1(\mgmt_gpio_data[29] ),
    .S(_1968_),
    .X(_1974_));
 sky130_fd_sc_hd__clkbuf_1 _5913_ (.A(net1166),
    .X(_0305_));
 sky130_fd_sc_hd__mux2_1 _5914_ (.A0(_1710_),
    .A1(\mgmt_gpio_data[30] ),
    .S(_1968_),
    .X(_1975_));
 sky130_fd_sc_hd__clkbuf_1 _5915_ (.A(net1164),
    .X(_0306_));
 sky130_fd_sc_hd__mux2_1 _5916_ (.A0(_1712_),
    .A1(\mgmt_gpio_data[31] ),
    .S(_1968_),
    .X(_1976_));
 sky130_fd_sc_hd__clkbuf_1 _5917_ (.A(net987),
    .X(_0307_));
 sky130_fd_sc_hd__nand2_4 _5918_ (.A(_1134_),
    .B(_1858_),
    .Y(_1977_));
 sky130_fd_sc_hd__mux2_1 _5919_ (.A0(_1801_),
    .A1(net1396),
    .S(_1977_),
    .X(_1978_));
 sky130_fd_sc_hd__clkbuf_1 _5920_ (.A(_1978_),
    .X(_0308_));
 sky130_fd_sc_hd__mux2_1 _5921_ (.A0(_1804_),
    .A1(net1213),
    .S(_1977_),
    .X(_1979_));
 sky130_fd_sc_hd__clkbuf_1 _5922_ (.A(net1214),
    .X(_0309_));
 sky130_fd_sc_hd__mux2_1 _5923_ (.A0(_1812_),
    .A1(net1318),
    .S(_1977_),
    .X(_1980_));
 sky130_fd_sc_hd__clkbuf_1 _5924_ (.A(net1319),
    .X(_0310_));
 sky130_fd_sc_hd__mux2_1 _5925_ (.A0(_1814_),
    .A1(net1357),
    .S(_1977_),
    .X(_1981_));
 sky130_fd_sc_hd__clkbuf_1 _5926_ (.A(_1981_),
    .X(_0311_));
 sky130_fd_sc_hd__mux2_1 _5927_ (.A0(_1816_),
    .A1(net866),
    .S(_1977_),
    .X(_1982_));
 sky130_fd_sc_hd__clkbuf_1 _5928_ (.A(net867),
    .X(_0312_));
 sky130_fd_sc_hd__and2_1 _5929_ (.A(\wbbd_state[4] ),
    .B(net502),
    .X(_1983_));
 sky130_fd_sc_hd__clkbuf_4 _5930_ (.A(_1983_),
    .X(_1984_));
 sky130_fd_sc_hd__mux2_1 _5931_ (.A0(net334),
    .A1(_1426_),
    .S(_1984_),
    .X(_1985_));
 sky130_fd_sc_hd__clkbuf_1 _5932_ (.A(_1985_),
    .X(_0313_));
 sky130_fd_sc_hd__mux2_1 _5933_ (.A0(net335),
    .A1(_1352_),
    .S(_1984_),
    .X(_1986_));
 sky130_fd_sc_hd__clkbuf_1 _5934_ (.A(_1986_),
    .X(_0314_));
 sky130_fd_sc_hd__mux2_1 _5935_ (.A0(net336),
    .A1(_1285_),
    .S(_1984_),
    .X(_1987_));
 sky130_fd_sc_hd__clkbuf_1 _5936_ (.A(_1987_),
    .X(_0315_));
 sky130_fd_sc_hd__mux2_1 _5937_ (.A0(net337),
    .A1(_1221_),
    .S(_1984_),
    .X(_1988_));
 sky130_fd_sc_hd__clkbuf_1 _5938_ (.A(_1988_),
    .X(_0316_));
 sky130_fd_sc_hd__mux2_2 _5939_ (.A0(net339),
    .A1(clknet_1_1__leaf__1160_),
    .S(_1984_),
    .X(_1989_));
 sky130_fd_sc_hd__buf_1 _5940_ (.A(_1989_),
    .X(_0317_));
 sky130_fd_sc_hd__mux2_1 _5941_ (.A0(net340),
    .A1(_1062_),
    .S(_1984_),
    .X(_1990_));
 sky130_fd_sc_hd__clkbuf_1 _5942_ (.A(_1990_),
    .X(_0318_));
 sky130_fd_sc_hd__mux2_1 _5943_ (.A0(net341),
    .A1(_1022_),
    .S(_1984_),
    .X(_1991_));
 sky130_fd_sc_hd__clkbuf_1 _5944_ (.A(_1991_),
    .X(_0319_));
 sky130_fd_sc_hd__mux2_1 _5945_ (.A0(net342),
    .A1(_0982_),
    .S(_1984_),
    .X(_1992_));
 sky130_fd_sc_hd__clkbuf_1 _5946_ (.A(_1992_),
    .X(_0320_));
 sky130_fd_sc_hd__clkbuf_4 _5947_ (.A(_1597_),
    .X(_1993_));
 sky130_fd_sc_hd__nand2_4 _5948_ (.A(_1111_),
    .B(_1858_),
    .Y(_1994_));
 sky130_fd_sc_hd__mux2_1 _5949_ (.A0(_1993_),
    .A1(net1361),
    .S(_1994_),
    .X(_1995_));
 sky130_fd_sc_hd__clkbuf_1 _5950_ (.A(net1362),
    .X(_0321_));
 sky130_fd_sc_hd__buf_4 _5951_ (.A(_1606_),
    .X(_1996_));
 sky130_fd_sc_hd__mux2_1 _5952_ (.A0(_1996_),
    .A1(net1050),
    .S(_1994_),
    .X(_1997_));
 sky130_fd_sc_hd__clkbuf_1 _5953_ (.A(net1051),
    .X(_0322_));
 sky130_fd_sc_hd__mux2_1 _5954_ (.A0(_1812_),
    .A1(net1085),
    .S(_1994_),
    .X(_1998_));
 sky130_fd_sc_hd__clkbuf_1 _5955_ (.A(net1086),
    .X(_0323_));
 sky130_fd_sc_hd__mux2_1 _5956_ (.A0(_1814_),
    .A1(net1180),
    .S(_1994_),
    .X(_1999_));
 sky130_fd_sc_hd__clkbuf_1 _5957_ (.A(net1181),
    .X(_0324_));
 sky130_fd_sc_hd__mux2_1 _5958_ (.A0(_1816_),
    .A1(net862),
    .S(_1994_),
    .X(_2000_));
 sky130_fd_sc_hd__clkbuf_1 _5959_ (.A(net863),
    .X(_0325_));
 sky130_fd_sc_hd__and2_1 _5960_ (.A(\wbbd_state[2] ),
    .B(net501),
    .X(_2001_));
 sky130_fd_sc_hd__clkbuf_4 _5961_ (.A(_2001_),
    .X(_2002_));
 sky130_fd_sc_hd__mux2_1 _5962_ (.A0(net357),
    .A1(_1426_),
    .S(_2002_),
    .X(_2003_));
 sky130_fd_sc_hd__clkbuf_1 _5963_ (.A(_2003_),
    .X(_0326_));
 sky130_fd_sc_hd__mux2_1 _5964_ (.A0(net358),
    .A1(_1352_),
    .S(_2002_),
    .X(_2004_));
 sky130_fd_sc_hd__clkbuf_1 _5965_ (.A(_2004_),
    .X(_0327_));
 sky130_fd_sc_hd__mux2_1 _5966_ (.A0(net328),
    .A1(_1285_),
    .S(_2002_),
    .X(_2005_));
 sky130_fd_sc_hd__clkbuf_1 _5967_ (.A(_2005_),
    .X(_0328_));
 sky130_fd_sc_hd__mux2_1 _5968_ (.A0(net329),
    .A1(_1221_),
    .S(_2002_),
    .X(_2006_));
 sky130_fd_sc_hd__clkbuf_1 _5969_ (.A(_2006_),
    .X(_0329_));
 sky130_fd_sc_hd__mux2_2 _5970_ (.A0(net330),
    .A1(clknet_1_1__leaf__1160_),
    .S(_2002_),
    .X(_2007_));
 sky130_fd_sc_hd__buf_1 _5971_ (.A(_2007_),
    .X(_0330_));
 sky130_fd_sc_hd__mux2_1 _5972_ (.A0(net331),
    .A1(_1062_),
    .S(_2002_),
    .X(_2008_));
 sky130_fd_sc_hd__clkbuf_1 _5973_ (.A(_2008_),
    .X(_0331_));
 sky130_fd_sc_hd__mux2_1 _5974_ (.A0(net332),
    .A1(_1022_),
    .S(_2002_),
    .X(_2009_));
 sky130_fd_sc_hd__clkbuf_1 _5975_ (.A(_2009_),
    .X(_0332_));
 sky130_fd_sc_hd__mux2_1 _5976_ (.A0(net333),
    .A1(_0982_),
    .S(_2002_),
    .X(_2010_));
 sky130_fd_sc_hd__clkbuf_1 _5977_ (.A(_2010_),
    .X(_0333_));
 sky130_fd_sc_hd__and2_2 _5978_ (.A(\wbbd_state[3] ),
    .B(net501),
    .X(_2011_));
 sky130_fd_sc_hd__buf_2 _5979_ (.A(_2011_),
    .X(_2012_));
 sky130_fd_sc_hd__mux2_1 _5980_ (.A0(net327),
    .A1(_1426_),
    .S(_2012_),
    .X(_2013_));
 sky130_fd_sc_hd__clkbuf_1 _5981_ (.A(_2013_),
    .X(_0334_));
 sky130_fd_sc_hd__mux2_1 _5982_ (.A0(net338),
    .A1(_1352_),
    .S(_2012_),
    .X(_2014_));
 sky130_fd_sc_hd__clkbuf_1 _5983_ (.A(_2014_),
    .X(_0335_));
 sky130_fd_sc_hd__mux2_1 _5984_ (.A0(net349),
    .A1(_1285_),
    .S(_2012_),
    .X(_2015_));
 sky130_fd_sc_hd__clkbuf_1 _5985_ (.A(_2015_),
    .X(_0336_));
 sky130_fd_sc_hd__mux2_1 _5986_ (.A0(net352),
    .A1(_1221_),
    .S(_2012_),
    .X(_2016_));
 sky130_fd_sc_hd__clkbuf_1 _5987_ (.A(_2016_),
    .X(_0337_));
 sky130_fd_sc_hd__mux2_2 _5988_ (.A0(net353),
    .A1(clknet_1_0__leaf__1160_),
    .S(_2012_),
    .X(_2017_));
 sky130_fd_sc_hd__buf_1 _5989_ (.A(_2017_),
    .X(_0338_));
 sky130_fd_sc_hd__mux2_1 _5990_ (.A0(net354),
    .A1(_1062_),
    .S(_2012_),
    .X(_2018_));
 sky130_fd_sc_hd__clkbuf_1 _5991_ (.A(_2018_),
    .X(_0339_));
 sky130_fd_sc_hd__mux2_1 _5992_ (.A0(net355),
    .A1(_1022_),
    .S(_2012_),
    .X(_2019_));
 sky130_fd_sc_hd__clkbuf_1 _5993_ (.A(_2019_),
    .X(_0340_));
 sky130_fd_sc_hd__mux2_1 _5994_ (.A0(net356),
    .A1(_0982_),
    .S(_2012_),
    .X(_2020_));
 sky130_fd_sc_hd__clkbuf_1 _5995_ (.A(_2020_),
    .X(_0341_));
 sky130_fd_sc_hd__and2_2 _5996_ (.A(_1137_),
    .B(_1871_),
    .X(_2021_));
 sky130_fd_sc_hd__mux2_1 _5997_ (.A0(net1407),
    .A1(_1878_),
    .S(_2021_),
    .X(_2022_));
 sky130_fd_sc_hd__clkbuf_1 _5998_ (.A(_2022_),
    .X(_0342_));
 sky130_fd_sc_hd__mux2_1 _5999_ (.A0(net1052),
    .A1(_1905_),
    .S(_2021_),
    .X(_2023_));
 sky130_fd_sc_hd__clkbuf_1 _6000_ (.A(_2023_),
    .X(_0343_));
 sky130_fd_sc_hd__mux2_1 _6001_ (.A0(net1151),
    .A1(_1833_),
    .S(_2021_),
    .X(_2024_));
 sky130_fd_sc_hd__clkbuf_1 _6002_ (.A(_2024_),
    .X(_0344_));
 sky130_fd_sc_hd__mux2_1 _6003_ (.A0(net954),
    .A1(_1836_),
    .S(_2021_),
    .X(_2025_));
 sky130_fd_sc_hd__clkbuf_1 _6004_ (.A(_2025_),
    .X(_0345_));
 sky130_fd_sc_hd__mux2_1 _6005_ (.A0(net1115),
    .A1(_1838_),
    .S(_2021_),
    .X(_2026_));
 sky130_fd_sc_hd__clkbuf_1 _6006_ (.A(_2026_),
    .X(_0346_));
 sky130_fd_sc_hd__nand2_2 _6007_ (.A(_1096_),
    .B(_1858_),
    .Y(_2027_));
 sky130_fd_sc_hd__mux2_1 _6008_ (.A0(_1993_),
    .A1(net1349),
    .S(_2027_),
    .X(_2028_));
 sky130_fd_sc_hd__clkbuf_1 _6009_ (.A(net1350),
    .X(_0347_));
 sky130_fd_sc_hd__mux2_1 _6010_ (.A0(_1996_),
    .A1(net1060),
    .S(_2027_),
    .X(_2029_));
 sky130_fd_sc_hd__clkbuf_1 _6011_ (.A(net1061),
    .X(_0348_));
 sky130_fd_sc_hd__buf_8 _6012_ (.A(_1610_),
    .X(_2030_));
 sky130_fd_sc_hd__mux2_1 _6013_ (.A0(_2030_),
    .A1(\gpio_configure[6][10] ),
    .S(_2027_),
    .X(_2031_));
 sky130_fd_sc_hd__clkbuf_1 _6014_ (.A(net1065),
    .X(_0349_));
 sky130_fd_sc_hd__clkbuf_16 _6015_ (.A(_1614_),
    .X(_2032_));
 sky130_fd_sc_hd__mux2_1 _6016_ (.A0(_2032_),
    .A1(net951),
    .S(_2027_),
    .X(_2033_));
 sky130_fd_sc_hd__clkbuf_1 _6017_ (.A(net952),
    .X(_0350_));
 sky130_fd_sc_hd__clkbuf_16 _6018_ (.A(net530),
    .X(_2034_));
 sky130_fd_sc_hd__mux2_1 _6019_ (.A0(_2034_),
    .A1(net645),
    .S(_2027_),
    .X(_2035_));
 sky130_fd_sc_hd__clkbuf_1 _6020_ (.A(net646),
    .X(_0351_));
 sky130_fd_sc_hd__and2_2 _6021_ (.A(_1136_),
    .B(_1871_),
    .X(_2036_));
 sky130_fd_sc_hd__mux2_1 _6022_ (.A0(net1390),
    .A1(_1878_),
    .S(_2036_),
    .X(_2037_));
 sky130_fd_sc_hd__clkbuf_1 _6023_ (.A(_2037_),
    .X(_0352_));
 sky130_fd_sc_hd__mux2_1 _6024_ (.A0(net989),
    .A1(_1905_),
    .S(_2036_),
    .X(_2038_));
 sky130_fd_sc_hd__clkbuf_1 _6025_ (.A(net990),
    .X(_0353_));
 sky130_fd_sc_hd__mux2_1 _6026_ (.A0(net1157),
    .A1(_1833_),
    .S(_2036_),
    .X(_2039_));
 sky130_fd_sc_hd__clkbuf_1 _6027_ (.A(net1158),
    .X(_0354_));
 sky130_fd_sc_hd__mux2_1 _6028_ (.A0(net917),
    .A1(_1836_),
    .S(_2036_),
    .X(_2040_));
 sky130_fd_sc_hd__clkbuf_1 _6029_ (.A(net918),
    .X(_0355_));
 sky130_fd_sc_hd__mux2_1 _6030_ (.A0(net1053),
    .A1(_1838_),
    .S(_2036_),
    .X(_2041_));
 sky130_fd_sc_hd__clkbuf_1 _6031_ (.A(net1054),
    .X(_0356_));
 sky130_fd_sc_hd__and2_2 _6032_ (.A(_1116_),
    .B(_1871_),
    .X(_2042_));
 sky130_fd_sc_hd__mux2_1 _6033_ (.A0(net1404),
    .A1(_1878_),
    .S(_2042_),
    .X(_2043_));
 sky130_fd_sc_hd__clkbuf_1 _6034_ (.A(_2043_),
    .X(_0357_));
 sky130_fd_sc_hd__mux2_1 _6035_ (.A0(net974),
    .A1(_1905_),
    .S(_2042_),
    .X(_2044_));
 sky130_fd_sc_hd__clkbuf_1 _6036_ (.A(_2044_),
    .X(_0358_));
 sky130_fd_sc_hd__mux2_1 _6037_ (.A0(net1057),
    .A1(_1833_),
    .S(_2042_),
    .X(_2045_));
 sky130_fd_sc_hd__clkbuf_1 _6038_ (.A(net1058),
    .X(_0359_));
 sky130_fd_sc_hd__mux2_1 _6039_ (.A0(net1006),
    .A1(_1836_),
    .S(_2042_),
    .X(_2046_));
 sky130_fd_sc_hd__clkbuf_1 _6040_ (.A(_2046_),
    .X(_0360_));
 sky130_fd_sc_hd__mux2_1 _6041_ (.A0(net1004),
    .A1(_1838_),
    .S(_2042_),
    .X(_2047_));
 sky130_fd_sc_hd__clkbuf_1 _6042_ (.A(_2047_),
    .X(_0361_));
 sky130_fd_sc_hd__and2_4 _6043_ (.A(_1066_),
    .B(_1871_),
    .X(_2048_));
 sky130_fd_sc_hd__mux2_1 _6044_ (.A0(net1389),
    .A1(_1878_),
    .S(_2048_),
    .X(_2049_));
 sky130_fd_sc_hd__clkbuf_1 _6045_ (.A(_2049_),
    .X(_0362_));
 sky130_fd_sc_hd__mux2_1 _6046_ (.A0(net1372),
    .A1(_1905_),
    .S(_2048_),
    .X(_2050_));
 sky130_fd_sc_hd__clkbuf_1 _6047_ (.A(_2050_),
    .X(_0363_));
 sky130_fd_sc_hd__buf_8 _6048_ (.A(_1610_),
    .X(_2051_));
 sky130_fd_sc_hd__mux2_1 _6049_ (.A0(net1259),
    .A1(_2051_),
    .S(_2048_),
    .X(_2052_));
 sky130_fd_sc_hd__clkbuf_1 _6050_ (.A(_2052_),
    .X(_0364_));
 sky130_fd_sc_hd__mux2_1 _6051_ (.A0(net710),
    .A1(net552),
    .S(_2048_),
    .X(_2053_));
 sky130_fd_sc_hd__clkbuf_1 _6052_ (.A(_2053_),
    .X(_0365_));
 sky130_fd_sc_hd__mux2_1 _6053_ (.A0(net843),
    .A1(_1668_),
    .S(_2048_),
    .X(_2054_));
 sky130_fd_sc_hd__clkbuf_1 _6054_ (.A(net1620),
    .X(_0366_));
 sky130_fd_sc_hd__nand2_2 _6055_ (.A(_1155_),
    .B(_1858_),
    .Y(_2055_));
 sky130_fd_sc_hd__mux2_1 _6056_ (.A0(_1993_),
    .A1(net1368),
    .S(_2055_),
    .X(_2056_));
 sky130_fd_sc_hd__clkbuf_1 _6057_ (.A(_2056_),
    .X(_0367_));
 sky130_fd_sc_hd__mux2_1 _6058_ (.A0(_1996_),
    .A1(net1136),
    .S(_2055_),
    .X(_2057_));
 sky130_fd_sc_hd__clkbuf_1 _6059_ (.A(_2057_),
    .X(_0368_));
 sky130_fd_sc_hd__mux2_1 _6060_ (.A0(_2030_),
    .A1(net1106),
    .S(_2055_),
    .X(_2058_));
 sky130_fd_sc_hd__clkbuf_1 _6061_ (.A(_2058_),
    .X(_0369_));
 sky130_fd_sc_hd__mux2_1 _6062_ (.A0(_2032_),
    .A1(net996),
    .S(_2055_),
    .X(_2059_));
 sky130_fd_sc_hd__clkbuf_1 _6063_ (.A(_2059_),
    .X(_0370_));
 sky130_fd_sc_hd__mux2_1 _6064_ (.A0(_2034_),
    .A1(net661),
    .S(_2055_),
    .X(_2060_));
 sky130_fd_sc_hd__clkbuf_1 _6065_ (.A(net662),
    .X(_0371_));
 sky130_fd_sc_hd__and2_2 _6066_ (.A(_1148_),
    .B(_1871_),
    .X(_2061_));
 sky130_fd_sc_hd__mux2_1 _6067_ (.A0(net1400),
    .A1(_1878_),
    .S(_2061_),
    .X(_2062_));
 sky130_fd_sc_hd__clkbuf_1 _6068_ (.A(_2062_),
    .X(_0372_));
 sky130_fd_sc_hd__mux2_1 _6069_ (.A0(net1062),
    .A1(_1905_),
    .S(_2061_),
    .X(_2063_));
 sky130_fd_sc_hd__clkbuf_1 _6070_ (.A(_2063_),
    .X(_0373_));
 sky130_fd_sc_hd__mux2_1 _6071_ (.A0(net1018),
    .A1(_2051_),
    .S(_2061_),
    .X(_2064_));
 sky130_fd_sc_hd__clkbuf_1 _6072_ (.A(net1019),
    .X(_0374_));
 sky130_fd_sc_hd__mux2_1 _6073_ (.A0(net577),
    .A1(net552),
    .S(_2061_),
    .X(_2065_));
 sky130_fd_sc_hd__clkbuf_1 _6074_ (.A(net578),
    .X(_0375_));
 sky130_fd_sc_hd__mux2_1 _6075_ (.A0(net665),
    .A1(_1668_),
    .S(_2061_),
    .X(_2066_));
 sky130_fd_sc_hd__clkbuf_1 _6076_ (.A(net666),
    .X(_0376_));
 sky130_fd_sc_hd__or2_4 _6077_ (.A(net144),
    .B(_1520_),
    .X(_2067_));
 sky130_fd_sc_hd__and4_1 _6078_ (.A(net139),
    .B(net138),
    .C(net141),
    .D(net140),
    .X(_2068_));
 sky130_fd_sc_hd__and4_1 _6079_ (.A(net135),
    .B(net134),
    .C(net137),
    .D(net136),
    .X(_2069_));
 sky130_fd_sc_hd__and4_1 _6080_ (.A(net162),
    .B(net161),
    .C(net133),
    .D(net132),
    .X(_2070_));
 sky130_fd_sc_hd__and3_1 _6081_ (.A(_2068_),
    .B(_2069_),
    .C(_2070_),
    .X(_2071_));
 sky130_fd_sc_hd__clkbuf_4 _6082_ (.A(net159),
    .X(_2072_));
 sky130_fd_sc_hd__and2_1 _6083_ (.A(net157),
    .B(net158),
    .X(_2073_));
 sky130_fd_sc_hd__clkbuf_2 _6084_ (.A(_2073_),
    .X(_2074_));
 sky130_fd_sc_hd__buf_4 _6085_ (.A(net142),
    .X(_2075_));
 sky130_fd_sc_hd__o211a_1 _6086_ (.A1(_2075_),
    .A2(net131),
    .B1(net156),
    .C1(net153),
    .X(_2076_));
 sky130_fd_sc_hd__and3_1 _6087_ (.A(_2072_),
    .B(_2074_),
    .C(_2076_),
    .X(_2077_));
 sky130_fd_sc_hd__and3_1 _6088_ (.A(net160),
    .B(_2071_),
    .C(_2077_),
    .X(_2078_));
 sky130_fd_sc_hd__xnor2_1 _6089_ (.A(_1519_),
    .B(_2078_),
    .Y(_2079_));
 sky130_fd_sc_hd__or2_1 _6090_ (.A(_2067_),
    .B(_2079_),
    .X(_2080_));
 sky130_fd_sc_hd__a21oi_1 _6091_ (.A1(_2074_),
    .A2(_2076_),
    .B1(_2072_),
    .Y(_2081_));
 sky130_fd_sc_hd__or2_2 _6092_ (.A(_2077_),
    .B(_2081_),
    .X(_2082_));
 sky130_fd_sc_hd__xnor2_2 _6093_ (.A(net160),
    .B(_2077_),
    .Y(_2083_));
 sky130_fd_sc_hd__nand2_2 _6094_ (.A(_2082_),
    .B(_2083_),
    .Y(_2084_));
 sky130_fd_sc_hd__xor2_2 _6095_ (.A(net157),
    .B(_2076_),
    .X(_2085_));
 sky130_fd_sc_hd__buf_2 _6096_ (.A(net158),
    .X(_2086_));
 sky130_fd_sc_hd__a21oi_1 _6097_ (.A1(net157),
    .A2(_2076_),
    .B1(_2086_),
    .Y(_2087_));
 sky130_fd_sc_hd__a21oi_1 _6098_ (.A1(_2074_),
    .A2(_2076_),
    .B1(_2087_),
    .Y(_2088_));
 sky130_fd_sc_hd__or3_2 _6099_ (.A(_2084_),
    .B(_2085_),
    .C(_2088_),
    .X(_2089_));
 sky130_fd_sc_hd__or2_1 _6100_ (.A(_2080_),
    .B(_2089_),
    .X(_2090_));
 sky130_fd_sc_hd__clkbuf_4 _6101_ (.A(_2090_),
    .X(_2091_));
 sky130_fd_sc_hd__buf_4 _6102_ (.A(net153),
    .X(_2092_));
 sky130_fd_sc_hd__or2_1 _6103_ (.A(net156),
    .B(_2092_),
    .X(_2093_));
 sky130_fd_sc_hd__buf_4 _6104_ (.A(_2093_),
    .X(_2094_));
 sky130_fd_sc_hd__nand2_8 _6105_ (.A(_2075_),
    .B(net131),
    .Y(_2095_));
 sky130_fd_sc_hd__or2_1 _6106_ (.A(_2094_),
    .B(_2095_),
    .X(_2096_));
 sky130_fd_sc_hd__buf_4 _6107_ (.A(_2096_),
    .X(_2097_));
 sky130_fd_sc_hd__nor2_1 _6108_ (.A(_2091_),
    .B(_2097_),
    .Y(_2098_));
 sky130_fd_sc_hd__buf_4 _6109_ (.A(net160),
    .X(_2099_));
 sky130_fd_sc_hd__or2_4 _6110_ (.A(net157),
    .B(_2086_),
    .X(_2100_));
 sky130_fd_sc_hd__or3_4 _6111_ (.A(_2072_),
    .B(_2099_),
    .C(_2100_),
    .X(_2101_));
 sky130_fd_sc_hd__clkbuf_4 _6112_ (.A(net156),
    .X(_2102_));
 sky130_fd_sc_hd__inv_2 _6113_ (.A(_2092_),
    .Y(_2103_));
 sky130_fd_sc_hd__clkinv_4 _6114_ (.A(net142),
    .Y(_2104_));
 sky130_fd_sc_hd__buf_4 _6115_ (.A(net131),
    .X(_2105_));
 sky130_fd_sc_hd__nand2_8 _6116_ (.A(_2104_),
    .B(_2105_),
    .Y(_2106_));
 sky130_fd_sc_hd__or3_1 _6117_ (.A(_2102_),
    .B(_2103_),
    .C(_2106_),
    .X(_2107_));
 sky130_fd_sc_hd__clkbuf_4 _6118_ (.A(_2107_),
    .X(_2108_));
 sky130_fd_sc_hd__nor2_2 _6119_ (.A(net144),
    .B(_1520_),
    .Y(_2109_));
 sky130_fd_sc_hd__nand2_4 _6120_ (.A(_1519_),
    .B(_2109_),
    .Y(_2110_));
 sky130_fd_sc_hd__nor3_2 _6121_ (.A(_2101_),
    .B(_2108_),
    .C(_2110_),
    .Y(_2111_));
 sky130_fd_sc_hd__and2_1 _6122_ (.A(_2104_),
    .B(_2105_),
    .X(_2112_));
 sky130_fd_sc_hd__inv_2 _6123_ (.A(_2094_),
    .Y(_2113_));
 sky130_fd_sc_hd__nand2_1 _6124_ (.A(_2112_),
    .B(_2113_),
    .Y(_2114_));
 sky130_fd_sc_hd__buf_6 _6125_ (.A(_2114_),
    .X(_2115_));
 sky130_fd_sc_hd__nor2_1 _6126_ (.A(_2091_),
    .B(_2115_),
    .Y(_2116_));
 sky130_fd_sc_hd__clkinv_2 _6127_ (.A(_2086_),
    .Y(_2117_));
 sky130_fd_sc_hd__and2_2 _6128_ (.A(_2117_),
    .B(_2085_),
    .X(_2118_));
 sky130_fd_sc_hd__or3b_1 _6129_ (.A(_2080_),
    .B(_2084_),
    .C_N(_2118_),
    .X(_2119_));
 sky130_fd_sc_hd__buf_4 _6130_ (.A(_2119_),
    .X(_2120_));
 sky130_fd_sc_hd__inv_2 _6131_ (.A(_2120_),
    .Y(_2121_));
 sky130_fd_sc_hd__nor2_8 _6132_ (.A(net156),
    .B(_2095_),
    .Y(_2122_));
 sky130_fd_sc_hd__nand2_4 _6133_ (.A(_2092_),
    .B(_2122_),
    .Y(_2123_));
 sky130_fd_sc_hd__nor2_1 _6134_ (.A(_2091_),
    .B(_2123_),
    .Y(_2124_));
 sky130_fd_sc_hd__nand2b_4 _6135_ (.A_N(net153),
    .B(net156),
    .Y(_2125_));
 sky130_fd_sc_hd__nor2_1 _6136_ (.A(_2104_),
    .B(_2125_),
    .Y(_2126_));
 sky130_fd_sc_hd__nand2_2 _6137_ (.A(_2105_),
    .B(_2126_),
    .Y(_2127_));
 sky130_fd_sc_hd__clkbuf_4 _6138_ (.A(_2127_),
    .X(_2128_));
 sky130_fd_sc_hd__nor2_1 _6139_ (.A(_2128_),
    .B(_2120_),
    .Y(_2129_));
 sky130_fd_sc_hd__or2b_1 _6140_ (.A(_2085_),
    .B_N(_2088_),
    .X(_2130_));
 sky130_fd_sc_hd__or3_1 _6141_ (.A(_2080_),
    .B(_2084_),
    .C(_2130_),
    .X(_2131_));
 sky130_fd_sc_hd__clkbuf_4 _6142_ (.A(_2131_),
    .X(_2132_));
 sky130_fd_sc_hd__or2_1 _6143_ (.A(_2106_),
    .B(_2125_),
    .X(_2133_));
 sky130_fd_sc_hd__buf_4 _6144_ (.A(_2133_),
    .X(_2134_));
 sky130_fd_sc_hd__nor2_1 _6145_ (.A(_2132_),
    .B(_2134_),
    .Y(_2135_));
 sky130_fd_sc_hd__nor2_1 _6146_ (.A(_2128_),
    .B(_2132_),
    .Y(_2136_));
 sky130_fd_sc_hd__nand2_1 _6147_ (.A(net156),
    .B(net153),
    .Y(_2137_));
 sky130_fd_sc_hd__clkbuf_8 _6148_ (.A(_2137_),
    .X(_2138_));
 sky130_fd_sc_hd__or2_1 _6149_ (.A(_2138_),
    .B(_2106_),
    .X(_2139_));
 sky130_fd_sc_hd__buf_4 _6150_ (.A(_2139_),
    .X(_2140_));
 sky130_fd_sc_hd__nand2_1 _6151_ (.A(net144),
    .B(_1519_),
    .Y(_2141_));
 sky130_fd_sc_hd__or2_1 _6152_ (.A(net144),
    .B(_1519_),
    .X(_2142_));
 sky130_fd_sc_hd__nand2_1 _6153_ (.A(net146),
    .B(net145),
    .Y(_2143_));
 sky130_fd_sc_hd__o21a_1 _6154_ (.A1(_2141_),
    .A2(_2143_),
    .B1(_1520_),
    .X(_2144_));
 sky130_fd_sc_hd__a21oi_1 _6155_ (.A1(_2141_),
    .A2(_2142_),
    .B1(_2144_),
    .Y(_2145_));
 sky130_fd_sc_hd__nand2_1 _6156_ (.A(_2079_),
    .B(_2145_),
    .Y(_2146_));
 sky130_fd_sc_hd__or2_2 _6157_ (.A(_2089_),
    .B(_2146_),
    .X(_2147_));
 sky130_fd_sc_hd__nor2_2 _6158_ (.A(_2140_),
    .B(_2147_),
    .Y(_2148_));
 sky130_fd_sc_hd__buf_4 _6159_ (.A(net157),
    .X(_2149_));
 sky130_fd_sc_hd__or2_4 _6160_ (.A(_2149_),
    .B(_2117_),
    .X(_2150_));
 sky130_fd_sc_hd__or3_4 _6161_ (.A(_2072_),
    .B(_2099_),
    .C(_2150_),
    .X(_2151_));
 sky130_fd_sc_hd__or2_1 _6162_ (.A(_2110_),
    .B(_2151_),
    .X(_2152_));
 sky130_fd_sc_hd__buf_2 _6163_ (.A(_2152_),
    .X(_2153_));
 sky130_fd_sc_hd__nor2_1 _6164_ (.A(_2140_),
    .B(_2153_),
    .Y(_2154_));
 sky130_fd_sc_hd__or3_1 _6165_ (.A(_2104_),
    .B(net131),
    .C(net156),
    .X(_2155_));
 sky130_fd_sc_hd__buf_4 _6166_ (.A(_2155_),
    .X(_2156_));
 sky130_fd_sc_hd__and3_1 _6167_ (.A(net142),
    .B(net156),
    .C(net153),
    .X(_2157_));
 sky130_fd_sc_hd__buf_2 _6168_ (.A(_2157_),
    .X(_2158_));
 sky130_fd_sc_hd__and3_1 _6169_ (.A(net159),
    .B(_2074_),
    .C(_2158_),
    .X(_2159_));
 sky130_fd_sc_hd__and4_1 _6170_ (.A(net160),
    .B(_2068_),
    .C(_2069_),
    .D(_2070_),
    .X(_2160_));
 sky130_fd_sc_hd__clkinv_2 _6171_ (.A(_1519_),
    .Y(_2161_));
 sky130_fd_sc_hd__a21oi_2 _6172_ (.A1(_2159_),
    .A2(_2160_),
    .B1(_2161_),
    .Y(_2162_));
 sky130_fd_sc_hd__and3_1 _6173_ (.A(_2161_),
    .B(_2159_),
    .C(_2160_),
    .X(_2163_));
 sky130_fd_sc_hd__nor3b_4 _6174_ (.A(_2162_),
    .B(_2163_),
    .C_N(_2145_),
    .Y(_2164_));
 sky130_fd_sc_hd__nand2_1 _6175_ (.A(_2074_),
    .B(_2158_),
    .Y(_2165_));
 sky130_fd_sc_hd__a21o_1 _6176_ (.A1(net157),
    .A2(_2158_),
    .B1(net158),
    .X(_2166_));
 sky130_fd_sc_hd__xnor2_1 _6177_ (.A(net157),
    .B(_2158_),
    .Y(_2167_));
 sky130_fd_sc_hd__and3_1 _6178_ (.A(_2165_),
    .B(_2166_),
    .C(_2167_),
    .X(_2168_));
 sky130_fd_sc_hd__nand2_2 _6179_ (.A(net395),
    .B(_2168_),
    .Y(_2169_));
 sky130_fd_sc_hd__inv_2 _6180_ (.A(net160),
    .Y(_2170_));
 sky130_fd_sc_hd__nand2_8 _6181_ (.A(net157),
    .B(net158),
    .Y(_2171_));
 sky130_fd_sc_hd__or2b_1 _6182_ (.A(net160),
    .B_N(net159),
    .X(_2172_));
 sky130_fd_sc_hd__buf_6 _6183_ (.A(_2172_),
    .X(_2173_));
 sky130_fd_sc_hd__nor2_8 _6184_ (.A(_2171_),
    .B(_2173_),
    .Y(_2174_));
 sky130_fd_sc_hd__a2bb2o_1 _6185_ (.A1_N(_2170_),
    .A2_N(_2159_),
    .B1(_2174_),
    .B2(_2158_),
    .X(_2175_));
 sky130_fd_sc_hd__a21oi_1 _6186_ (.A1(_2074_),
    .A2(_2158_),
    .B1(_2072_),
    .Y(_2176_));
 sky130_fd_sc_hd__or2_2 _6187_ (.A(_2159_),
    .B(_2176_),
    .X(_2177_));
 sky130_fd_sc_hd__nand2b_2 _6188_ (.A_N(_2175_),
    .B(_2177_),
    .Y(_2178_));
 sky130_fd_sc_hd__or2_1 _6189_ (.A(_2169_),
    .B(_2178_),
    .X(_2179_));
 sky130_fd_sc_hd__buf_2 _6190_ (.A(_2179_),
    .X(_2180_));
 sky130_fd_sc_hd__nor2_8 _6191_ (.A(_2106_),
    .B(_2094_),
    .Y(_2181_));
 sky130_fd_sc_hd__nor2_1 _6192_ (.A(net144),
    .B(_1519_),
    .Y(_2182_));
 sky130_fd_sc_hd__or3b_2 _6193_ (.A(_1520_),
    .B(_2182_),
    .C_N(_2079_),
    .X(_2183_));
 sky130_fd_sc_hd__nor2_2 _6194_ (.A(_2089_),
    .B(_2183_),
    .Y(_2184_));
 sky130_fd_sc_hd__nand2_1 _6195_ (.A(_2181_),
    .B(_2184_),
    .Y(_2185_));
 sky130_fd_sc_hd__nor2_1 _6196_ (.A(_2117_),
    .B(_2167_),
    .Y(_2186_));
 sky130_fd_sc_hd__nand2_1 _6197_ (.A(net395),
    .B(_2186_),
    .Y(_2187_));
 sky130_fd_sc_hd__or2_1 _6198_ (.A(_2187_),
    .B(_2178_),
    .X(_2188_));
 sky130_fd_sc_hd__buf_2 _6199_ (.A(_2188_),
    .X(_2189_));
 sky130_fd_sc_hd__or3_4 _6200_ (.A(_2104_),
    .B(_2105_),
    .C(_2138_),
    .X(_2190_));
 sky130_fd_sc_hd__buf_4 _6201_ (.A(_2190_),
    .X(_2191_));
 sky130_fd_sc_hd__or2_1 _6202_ (.A(_2191_),
    .B(_2189_),
    .X(_2192_));
 sky130_fd_sc_hd__or2_2 _6203_ (.A(_2099_),
    .B(_2177_),
    .X(_2193_));
 sky130_fd_sc_hd__or3b_2 _6204_ (.A(_2162_),
    .B(_2163_),
    .C_N(_2145_),
    .X(_2194_));
 sky130_fd_sc_hd__a21bo_1 _6205_ (.A1(_2165_),
    .A2(_2166_),
    .B1_N(_2167_),
    .X(_2195_));
 sky130_fd_sc_hd__or2_2 _6206_ (.A(_2194_),
    .B(_2195_),
    .X(_2196_));
 sky130_fd_sc_hd__or2_1 _6207_ (.A(_2193_),
    .B(_2196_),
    .X(_2197_));
 sky130_fd_sc_hd__buf_2 _6208_ (.A(_2197_),
    .X(_2198_));
 sky130_fd_sc_hd__or2_1 _6209_ (.A(_2191_),
    .B(_2198_),
    .X(_2199_));
 sky130_fd_sc_hd__nor2_1 _6210_ (.A(_2086_),
    .B(_2167_),
    .Y(_2200_));
 sky130_fd_sc_hd__nand2_2 _6211_ (.A(_2164_),
    .B(_2200_),
    .Y(_2201_));
 sky130_fd_sc_hd__or2_1 _6212_ (.A(_2201_),
    .B(_2193_),
    .X(_2202_));
 sky130_fd_sc_hd__clkbuf_4 _6213_ (.A(_2202_),
    .X(_2203_));
 sky130_fd_sc_hd__and2b_1 _6214_ (.A_N(_2105_),
    .B(_2158_),
    .X(_2204_));
 sky130_fd_sc_hd__clkbuf_4 _6215_ (.A(_2204_),
    .X(_2205_));
 sky130_fd_sc_hd__nor2_2 _6216_ (.A(_2201_),
    .B(_2193_),
    .Y(_2206_));
 sky130_fd_sc_hd__nand2_1 _6217_ (.A(_2205_),
    .B(_2206_),
    .Y(_2207_));
 sky130_fd_sc_hd__or2_1 _6218_ (.A(_2092_),
    .B(_2156_),
    .X(_2208_));
 sky130_fd_sc_hd__clkbuf_4 _6219_ (.A(_2208_),
    .X(_2209_));
 sky130_fd_sc_hd__nand2_4 _6220_ (.A(_2177_),
    .B(_2175_),
    .Y(_2210_));
 sky130_fd_sc_hd__or2_1 _6221_ (.A(_2210_),
    .B(_2196_),
    .X(_2211_));
 sky130_fd_sc_hd__buf_2 _6222_ (.A(_2211_),
    .X(_2212_));
 sky130_fd_sc_hd__a21oi_1 _6223_ (.A1(_2209_),
    .A2(_2190_),
    .B1(_2212_),
    .Y(_2213_));
 sky130_fd_sc_hd__clkbuf_4 _6224_ (.A(_2146_),
    .X(_2214_));
 sky130_fd_sc_hd__nor2_4 _6225_ (.A(_2138_),
    .B(_2106_),
    .Y(_2215_));
 sky130_fd_sc_hd__nor3_4 _6226_ (.A(_2072_),
    .B(_2099_),
    .C(_2100_),
    .Y(_2216_));
 sky130_fd_sc_hd__nand2_2 _6227_ (.A(_2215_),
    .B(_2216_),
    .Y(_2217_));
 sky130_fd_sc_hd__nor2_1 _6228_ (.A(_2089_),
    .B(_2214_),
    .Y(_2218_));
 sky130_fd_sc_hd__and2_1 _6229_ (.A(_2075_),
    .B(_2105_),
    .X(_2219_));
 sky130_fd_sc_hd__and3_2 _6230_ (.A(_2102_),
    .B(_2103_),
    .C(_2219_),
    .X(_2220_));
 sky130_fd_sc_hd__a2bb2o_1 _6231_ (.A1_N(_2214_),
    .A2_N(_2217_),
    .B1(_2218_),
    .B2(_2220_),
    .X(_2221_));
 sky130_fd_sc_hd__or4_1 _6232_ (.A(_2086_),
    .B(_2194_),
    .C(_2167_),
    .D(_2210_),
    .X(_2222_));
 sky130_fd_sc_hd__buf_4 _6233_ (.A(_2222_),
    .X(_2223_));
 sky130_fd_sc_hd__or2_1 _6234_ (.A(_2104_),
    .B(_2125_),
    .X(_2224_));
 sky130_fd_sc_hd__buf_2 _6235_ (.A(_2224_),
    .X(_2225_));
 sky130_fd_sc_hd__or2_1 _6236_ (.A(net131),
    .B(_2225_),
    .X(_2226_));
 sky130_fd_sc_hd__clkbuf_4 _6237_ (.A(_2226_),
    .X(_2227_));
 sky130_fd_sc_hd__nor2_1 _6238_ (.A(_2223_),
    .B(_2227_),
    .Y(_2228_));
 sky130_fd_sc_hd__or2_2 _6239_ (.A(_2210_),
    .B(_2169_),
    .X(_2229_));
 sky130_fd_sc_hd__nor2_1 _6240_ (.A(_2190_),
    .B(_2229_),
    .Y(_2230_));
 sky130_fd_sc_hd__nor2_1 _6241_ (.A(_2227_),
    .B(_2229_),
    .Y(_2231_));
 sky130_fd_sc_hd__o22a_1 _6242_ (.A1(_2217_),
    .A2(_2183_),
    .B1(_2133_),
    .B2(_2147_),
    .X(_2232_));
 sky130_fd_sc_hd__or2b_2 _6243_ (.A(_2083_),
    .B_N(_2082_),
    .X(_2233_));
 sky130_fd_sc_hd__or2_1 _6244_ (.A(_2233_),
    .B(_2130_),
    .X(_2234_));
 sky130_fd_sc_hd__nand2_1 _6245_ (.A(_2086_),
    .B(_2085_),
    .Y(_2235_));
 sky130_fd_sc_hd__or2_1 _6246_ (.A(_2233_),
    .B(_2235_),
    .X(_2236_));
 sky130_fd_sc_hd__a211o_1 _6247_ (.A1(_2234_),
    .A2(_2236_),
    .B1(_2102_),
    .C1(_2146_),
    .X(_2237_));
 sky130_fd_sc_hd__or3_1 _6248_ (.A(_2104_),
    .B(_2105_),
    .C(_2237_),
    .X(_2238_));
 sky130_fd_sc_hd__or3_1 _6249_ (.A(_2146_),
    .B(_2190_),
    .C(_2236_),
    .X(_2239_));
 sky130_fd_sc_hd__and4b_1 _6250_ (.A_N(_2231_),
    .B(_2232_),
    .C(_2238_),
    .D(_2239_),
    .X(_2240_));
 sky130_fd_sc_hd__or4b_2 _6251_ (.A(_2221_),
    .B(_2228_),
    .C(_2230_),
    .D_N(_2240_),
    .X(_2241_));
 sky130_fd_sc_hd__nor2_1 _6252_ (.A(_2156_),
    .B(_2223_),
    .Y(_2242_));
 sky130_fd_sc_hd__or2_1 _6253_ (.A(_2103_),
    .B(_2156_),
    .X(_2243_));
 sky130_fd_sc_hd__clkbuf_4 _6254_ (.A(_2243_),
    .X(_2244_));
 sky130_fd_sc_hd__or2_1 _6255_ (.A(_2212_),
    .B(_2244_),
    .X(_2245_));
 sky130_fd_sc_hd__o221a_1 _6256_ (.A1(_2223_),
    .A2(_2190_),
    .B1(_2227_),
    .B2(_2212_),
    .C1(_2245_),
    .X(_2246_));
 sky130_fd_sc_hd__or4b_1 _6257_ (.A(_2213_),
    .B(_2241_),
    .C(_2242_),
    .D_N(_2246_),
    .X(_2247_));
 sky130_fd_sc_hd__or2_1 _6258_ (.A(_2193_),
    .B(_2187_),
    .X(_2248_));
 sky130_fd_sc_hd__clkbuf_4 _6259_ (.A(_2248_),
    .X(_2249_));
 sky130_fd_sc_hd__nor2_1 _6260_ (.A(_2227_),
    .B(_2249_),
    .Y(_2250_));
 sky130_fd_sc_hd__nor2_1 _6261_ (.A(_2156_),
    .B(_2249_),
    .Y(_2251_));
 sky130_fd_sc_hd__or2_1 _6262_ (.A(_2193_),
    .B(_2169_),
    .X(_2252_));
 sky130_fd_sc_hd__buf_2 _6263_ (.A(_2252_),
    .X(_2253_));
 sky130_fd_sc_hd__nor2_1 _6264_ (.A(_2253_),
    .B(_2244_),
    .Y(_2254_));
 sky130_fd_sc_hd__nor2_1 _6265_ (.A(_2253_),
    .B(_2227_),
    .Y(_2255_));
 sky130_fd_sc_hd__or2_1 _6266_ (.A(_2190_),
    .B(_2249_),
    .X(_2256_));
 sky130_fd_sc_hd__or3b_1 _6267_ (.A(_2254_),
    .B(_2255_),
    .C_N(_2256_),
    .X(_2257_));
 sky130_fd_sc_hd__or4_1 _6268_ (.A(_2247_),
    .B(_2250_),
    .C(_2251_),
    .D(_2257_),
    .X(_2258_));
 sky130_fd_sc_hd__nor2_1 _6269_ (.A(_2227_),
    .B(_2203_),
    .Y(_2259_));
 sky130_fd_sc_hd__or2_1 _6270_ (.A(_2253_),
    .B(_2209_),
    .X(_2260_));
 sky130_fd_sc_hd__or2_1 _6271_ (.A(_2253_),
    .B(_2191_),
    .X(_2261_));
 sky130_fd_sc_hd__and4bb_1 _6272_ (.A_N(_2258_),
    .B_N(_2259_),
    .C(_2260_),
    .D(_2261_),
    .X(_2262_));
 sky130_fd_sc_hd__clkbuf_4 _6273_ (.A(_2227_),
    .X(_2263_));
 sky130_fd_sc_hd__or2_1 _6274_ (.A(_2263_),
    .B(_2198_),
    .X(_2264_));
 sky130_fd_sc_hd__o2111a_1 _6275_ (.A1(_2156_),
    .A2(_2203_),
    .B1(_2207_),
    .C1(_2262_),
    .D1(_2264_),
    .X(_2265_));
 sky130_fd_sc_hd__nor2_1 _6276_ (.A(_2263_),
    .B(_2189_),
    .Y(_2266_));
 sky130_fd_sc_hd__inv_2 _6277_ (.A(_2266_),
    .Y(_2267_));
 sky130_fd_sc_hd__o2111a_1 _6278_ (.A1(_2156_),
    .A2(_2198_),
    .B1(_2199_),
    .C1(_2265_),
    .D1(_2267_),
    .X(_2268_));
 sky130_fd_sc_hd__clkinv_2 _6279_ (.A(_2227_),
    .Y(_2269_));
 sky130_fd_sc_hd__nor2_2 _6280_ (.A(_2169_),
    .B(_2178_),
    .Y(_2270_));
 sky130_fd_sc_hd__nand2_1 _6281_ (.A(_2269_),
    .B(_2270_),
    .Y(_2271_));
 sky130_fd_sc_hd__o2111a_1 _6282_ (.A1(_2156_),
    .A2(_2189_),
    .B1(_2192_),
    .C1(_2268_),
    .D1(_2271_),
    .X(_2272_));
 sky130_fd_sc_hd__o211a_1 _6283_ (.A1(_2156_),
    .A2(_2180_),
    .B1(_2185_),
    .C1(_2272_),
    .X(_2273_));
 sky130_fd_sc_hd__or4b_1 _6284_ (.A(_2136_),
    .B(_2148_),
    .C(_2154_),
    .D_N(_2273_),
    .X(_2274_));
 sky130_fd_sc_hd__nor2_8 _6285_ (.A(_2106_),
    .B(_2125_),
    .Y(_2275_));
 sky130_fd_sc_hd__nand2_4 _6286_ (.A(_2149_),
    .B(_2117_),
    .Y(_2276_));
 sky130_fd_sc_hd__or3_2 _6287_ (.A(_2072_),
    .B(_2099_),
    .C(_2276_),
    .X(_2277_));
 sky130_fd_sc_hd__nor3_1 _6288_ (.A(_2140_),
    .B(_2110_),
    .C(_2277_),
    .Y(_2278_));
 sky130_fd_sc_hd__a21oi_1 _6289_ (.A1(_2121_),
    .A2(_2275_),
    .B1(_2278_),
    .Y(_2279_));
 sky130_fd_sc_hd__or4b_1 _6290_ (.A(_2129_),
    .B(_2135_),
    .C(_2274_),
    .D_N(_2279_),
    .X(_2280_));
 sky130_fd_sc_hd__a311o_1 _6291_ (.A1(_2092_),
    .A2(_2112_),
    .A3(_2121_),
    .B1(_2124_),
    .C1(_2280_),
    .X(_2281_));
 sky130_fd_sc_hd__o21a_1 _6292_ (.A1(_2091_),
    .A2(_2140_),
    .B1(\wbbd_state[9] ),
    .X(_2282_));
 sky130_fd_sc_hd__o41a_1 _6293_ (.A1(_2098_),
    .A2(_2111_),
    .A3(_2116_),
    .A4(_2281_),
    .B1(_2282_),
    .X(_2283_));
 sky130_fd_sc_hd__buf_4 _6294_ (.A(_2244_),
    .X(_2284_));
 sky130_fd_sc_hd__nor2_4 _6295_ (.A(_2091_),
    .B(_2284_),
    .Y(_2285_));
 sky130_fd_sc_hd__nor2_1 _6296_ (.A(_2091_),
    .B(_2209_),
    .Y(_2286_));
 sky130_fd_sc_hd__or2_1 _6297_ (.A(_2162_),
    .B(_2163_),
    .X(_2287_));
 sky130_fd_sc_hd__nor3b_1 _6298_ (.A(_2067_),
    .B(_2178_),
    .C_N(_2287_),
    .Y(_2288_));
 sky130_fd_sc_hd__nand2_1 _6299_ (.A(_2200_),
    .B(net394),
    .Y(_2289_));
 sky130_fd_sc_hd__nor2_2 _6300_ (.A(_2156_),
    .B(_2289_),
    .Y(_2290_));
 sky130_fd_sc_hd__nor2_1 _6301_ (.A(_2132_),
    .B(_2263_),
    .Y(_2291_));
 sky130_fd_sc_hd__or2_1 _6302_ (.A(_2075_),
    .B(net131),
    .X(_2292_));
 sky130_fd_sc_hd__buf_4 _6303_ (.A(_2292_),
    .X(_2293_));
 sky130_fd_sc_hd__or2_1 _6304_ (.A(_2138_),
    .B(_2293_),
    .X(_2294_));
 sky130_fd_sc_hd__buf_4 _6305_ (.A(_2294_),
    .X(_2295_));
 sky130_fd_sc_hd__nor2_2 _6306_ (.A(_2120_),
    .B(_2295_),
    .Y(_2296_));
 sky130_fd_sc_hd__nor2_1 _6307_ (.A(_2153_),
    .B(_2295_),
    .Y(_2297_));
 sky130_fd_sc_hd__nor2_1 _6308_ (.A(_2191_),
    .B(_2153_),
    .Y(_2298_));
 sky130_fd_sc_hd__nor2_1 _6309_ (.A(_2195_),
    .B(_2178_),
    .Y(_2299_));
 sky130_fd_sc_hd__and3_1 _6310_ (.A(net395),
    .B(_2205_),
    .C(_2299_),
    .X(_2300_));
 sky130_fd_sc_hd__nor2_4 _6311_ (.A(_2092_),
    .B(_2156_),
    .Y(_2301_));
 sky130_fd_sc_hd__or2_1 _6312_ (.A(_1520_),
    .B(_2182_),
    .X(_2302_));
 sky130_fd_sc_hd__nor2_2 _6313_ (.A(_2287_),
    .B(_2302_),
    .Y(_2303_));
 sky130_fd_sc_hd__and3_1 _6314_ (.A(_2301_),
    .B(_2303_),
    .C(_2299_),
    .X(_2304_));
 sky130_fd_sc_hd__inv_2 _6315_ (.A(_2189_),
    .Y(_2305_));
 sky130_fd_sc_hd__nor2_4 _6316_ (.A(_2137_),
    .B(_2095_),
    .Y(_2306_));
 sky130_fd_sc_hd__and2_1 _6317_ (.A(net131),
    .B(_2159_),
    .X(_2307_));
 sky130_fd_sc_hd__nand2_1 _6318_ (.A(_2160_),
    .B(_2307_),
    .Y(_2308_));
 sky130_fd_sc_hd__mux2_1 _6319_ (.A0(_2141_),
    .A1(_2142_),
    .S(_2308_),
    .X(_2309_));
 sky130_fd_sc_hd__nor2_4 _6320_ (.A(_2144_),
    .B(_2309_),
    .Y(_2310_));
 sky130_fd_sc_hd__and3b_1 _6321_ (.A_N(_2151_),
    .B(_2306_),
    .C(_2310_),
    .X(_2311_));
 sky130_fd_sc_hd__nor2_1 _6322_ (.A(_2128_),
    .B(_2180_),
    .Y(_2312_));
 sky130_fd_sc_hd__nor2_1 _6323_ (.A(_2128_),
    .B(_2189_),
    .Y(_2313_));
 sky130_fd_sc_hd__or2_1 _6324_ (.A(_2137_),
    .B(_2095_),
    .X(_2314_));
 sky130_fd_sc_hd__buf_2 _6325_ (.A(_2314_),
    .X(_2315_));
 sky130_fd_sc_hd__buf_4 _6326_ (.A(_2315_),
    .X(_2316_));
 sky130_fd_sc_hd__nor2_1 _6327_ (.A(_2198_),
    .B(_2316_),
    .Y(_2317_));
 sky130_fd_sc_hd__inv_2 _6328_ (.A(_2197_),
    .Y(_2318_));
 sky130_fd_sc_hd__nor2_1 _6329_ (.A(_2128_),
    .B(_2197_),
    .Y(_2319_));
 sky130_fd_sc_hd__nor2_1 _6330_ (.A(_2203_),
    .B(_2316_),
    .Y(_2320_));
 sky130_fd_sc_hd__inv_2 _6331_ (.A(_2253_),
    .Y(_2321_));
 sky130_fd_sc_hd__nor2_1 _6332_ (.A(_2253_),
    .B(_2316_),
    .Y(_2322_));
 sky130_fd_sc_hd__nor2_1 _6333_ (.A(_2128_),
    .B(_2203_),
    .Y(_2323_));
 sky130_fd_sc_hd__nor2_1 _6334_ (.A(_2253_),
    .B(_2128_),
    .Y(_2324_));
 sky130_fd_sc_hd__nor2_1 _6335_ (.A(_2249_),
    .B(_2315_),
    .Y(_2325_));
 sky130_fd_sc_hd__nor2_1 _6336_ (.A(_2249_),
    .B(_2097_),
    .Y(_2326_));
 sky130_fd_sc_hd__nor2_1 _6337_ (.A(_2127_),
    .B(_2248_),
    .Y(_2327_));
 sky130_fd_sc_hd__nor2_1 _6338_ (.A(_2248_),
    .B(_2123_),
    .Y(_2328_));
 sky130_fd_sc_hd__nor2_1 _6339_ (.A(_2212_),
    .B(_2315_),
    .Y(_2329_));
 sky130_fd_sc_hd__nor2_2 _6340_ (.A(_2210_),
    .B(_2196_),
    .Y(_2330_));
 sky130_fd_sc_hd__nor2_1 _6341_ (.A(_2127_),
    .B(_2212_),
    .Y(_2331_));
 sky130_fd_sc_hd__nor2_1 _6342_ (.A(_2223_),
    .B(_2123_),
    .Y(_2332_));
 sky130_fd_sc_hd__and3_1 _6343_ (.A(_2205_),
    .B(_2216_),
    .C(_2303_),
    .X(_2333_));
 sky130_fd_sc_hd__and2_1 _6344_ (.A(_2177_),
    .B(_2175_),
    .X(_2334_));
 sky130_fd_sc_hd__and3_2 _6345_ (.A(_2164_),
    .B(_2200_),
    .C(_2334_),
    .X(_2335_));
 sky130_fd_sc_hd__a31o_1 _6346_ (.A1(_2164_),
    .A2(_2334_),
    .A3(_2168_),
    .B1(_2125_),
    .X(_2336_));
 sky130_fd_sc_hd__o2111a_1 _6347_ (.A1(_2168_),
    .A2(_2186_),
    .B1(_2219_),
    .C1(_2164_),
    .D1(_2334_),
    .X(_2337_));
 sky130_fd_sc_hd__nor2_8 _6348_ (.A(_2138_),
    .B(_2293_),
    .Y(_2338_));
 sky130_fd_sc_hd__o311a_1 _6349_ (.A1(_2204_),
    .A2(_2269_),
    .A3(_2338_),
    .B1(_2216_),
    .C1(_2164_),
    .X(_2339_));
 sky130_fd_sc_hd__a221o_1 _6350_ (.A1(_2335_),
    .A2(_2220_),
    .B1(_2336_),
    .B2(_2337_),
    .C1(_2339_),
    .X(_2340_));
 sky130_fd_sc_hd__a21oi_1 _6351_ (.A1(_2097_),
    .A2(_2315_),
    .B1(_2223_),
    .Y(_2341_));
 sky130_fd_sc_hd__or4_1 _6352_ (.A(_2332_),
    .B(_2333_),
    .C(_2340_),
    .D(_2341_),
    .X(_2342_));
 sky130_fd_sc_hd__a211o_1 _6353_ (.A1(_2330_),
    .A2(_2122_),
    .B1(_2331_),
    .C1(_2342_),
    .X(_2343_));
 sky130_fd_sc_hd__or4_1 _6354_ (.A(_2327_),
    .B(_2328_),
    .C(_2329_),
    .D(_2343_),
    .X(_2344_));
 sky130_fd_sc_hd__or4_1 _6355_ (.A(_2324_),
    .B(_2325_),
    .C(_2326_),
    .D(_2344_),
    .X(_2345_));
 sky130_fd_sc_hd__a2111o_1 _6356_ (.A1(_2321_),
    .A2(_2122_),
    .B1(_2322_),
    .C1(_2323_),
    .D1(_2345_),
    .X(_2346_));
 sky130_fd_sc_hd__a211o_1 _6357_ (.A1(_2206_),
    .A2(_2122_),
    .B1(_2320_),
    .C1(_2346_),
    .X(_2347_));
 sky130_fd_sc_hd__a211o_1 _6358_ (.A1(_2318_),
    .A2(_2122_),
    .B1(_2319_),
    .C1(_2347_),
    .X(_2348_));
 sky130_fd_sc_hd__or3_1 _6359_ (.A(_2313_),
    .B(_2317_),
    .C(_2348_),
    .X(_2349_));
 sky130_fd_sc_hd__a2111o_1 _6360_ (.A1(_2305_),
    .A2(_2122_),
    .B1(_2311_),
    .C1(_2312_),
    .D1(_2349_),
    .X(_2350_));
 sky130_fd_sc_hd__a211o_1 _6361_ (.A1(_2270_),
    .A2(_2122_),
    .B1(_2304_),
    .C1(_2350_),
    .X(_2351_));
 sky130_fd_sc_hd__or4_1 _6362_ (.A(_2297_),
    .B(_2298_),
    .C(_2300_),
    .D(_2351_),
    .X(_2352_));
 sky130_fd_sc_hd__o32a_1 _6363_ (.A1(_2191_),
    .A2(_2110_),
    .A3(_2277_),
    .B1(_2263_),
    .B2(_2120_),
    .X(_2353_));
 sky130_fd_sc_hd__or4b_1 _6364_ (.A(_2291_),
    .B(_2296_),
    .C(_2352_),
    .D_N(_2353_),
    .X(_2354_));
 sky130_fd_sc_hd__nor2_1 _6365_ (.A(_2191_),
    .B(_2289_),
    .Y(_2355_));
 sky130_fd_sc_hd__or2_2 _6366_ (.A(_2293_),
    .B(_2125_),
    .X(_2356_));
 sky130_fd_sc_hd__buf_4 _6367_ (.A(_2356_),
    .X(_2357_));
 sky130_fd_sc_hd__nor2_1 _6368_ (.A(_2091_),
    .B(_2357_),
    .Y(_2358_));
 sky130_fd_sc_hd__a2111o_1 _6369_ (.A1(_2092_),
    .A2(_2290_),
    .B1(_2354_),
    .C1(_2355_),
    .D1(_2358_),
    .X(_2359_));
 sky130_fd_sc_hd__clkbuf_4 _6370_ (.A(_2216_),
    .X(_2360_));
 sky130_fd_sc_hd__nor2_2 _6371_ (.A(_2161_),
    .B(_2067_),
    .Y(_2361_));
 sky130_fd_sc_hd__or2_1 _6372_ (.A(_2102_),
    .B(_2293_),
    .X(_2362_));
 sky130_fd_sc_hd__clkbuf_4 _6373_ (.A(_2362_),
    .X(_2363_));
 sky130_fd_sc_hd__nor2_4 _6374_ (.A(_2103_),
    .B(_2363_),
    .Y(_2364_));
 sky130_fd_sc_hd__and3_1 _6375_ (.A(_2360_),
    .B(_2361_),
    .C(_2364_),
    .X(_2365_));
 sky130_fd_sc_hd__inv_2 _6376_ (.A(_2288_),
    .Y(_2366_));
 sky130_fd_sc_hd__o31a_1 _6377_ (.A1(_2171_),
    .A2(_2191_),
    .A3(_2366_),
    .B1(\wbbd_state[7] ),
    .X(_2367_));
 sky130_fd_sc_hd__o41a_1 _6378_ (.A1(_2285_),
    .A2(_2286_),
    .A3(_2359_),
    .A4(_2365_),
    .B1(_2367_),
    .X(_2368_));
 sky130_fd_sc_hd__nand2_1 _6379_ (.A(_2099_),
    .B(_2307_),
    .Y(_2369_));
 sky130_fd_sc_hd__xnor2_1 _6380_ (.A(_1519_),
    .B(_2308_),
    .Y(_2370_));
 sky130_fd_sc_hd__nand2_1 _6381_ (.A(_2109_),
    .B(_2370_),
    .Y(_2371_));
 sky130_fd_sc_hd__o21a_1 _6382_ (.A1(_2369_),
    .A2(_2371_),
    .B1(\wbbd_state[8] ),
    .X(_2372_));
 sky130_fd_sc_hd__nor2_4 _6383_ (.A(_2094_),
    .B(_2095_),
    .Y(_2373_));
 sky130_fd_sc_hd__a31o_1 _6384_ (.A1(net131),
    .A2(_2074_),
    .A3(_2158_),
    .B1(_2072_),
    .X(_2374_));
 sky130_fd_sc_hd__or2b_1 _6385_ (.A(_2307_),
    .B_N(_2374_),
    .X(_2375_));
 sky130_fd_sc_hd__xnor2_1 _6386_ (.A(_2099_),
    .B(_2307_),
    .Y(_2376_));
 sky130_fd_sc_hd__a21oi_1 _6387_ (.A1(_2149_),
    .A2(_2306_),
    .B1(_2086_),
    .Y(_2377_));
 sky130_fd_sc_hd__a31o_1 _6388_ (.A1(_2105_),
    .A2(_2074_),
    .A3(_2158_),
    .B1(_2377_),
    .X(_2378_));
 sky130_fd_sc_hd__xnor2_1 _6389_ (.A(_2149_),
    .B(_2306_),
    .Y(_2379_));
 sky130_fd_sc_hd__and4_1 _6390_ (.A(_2375_),
    .B(_2376_),
    .C(_2378_),
    .D(_2379_),
    .X(_2380_));
 sky130_fd_sc_hd__nor2_2 _6391_ (.A(_2302_),
    .B(_2370_),
    .Y(_2381_));
 sky130_fd_sc_hd__or2_2 _6392_ (.A(_2144_),
    .B(_2309_),
    .X(_2382_));
 sky130_fd_sc_hd__nor2_1 _6393_ (.A(_2369_),
    .B(_2382_),
    .Y(_2383_));
 sky130_fd_sc_hd__a31o_1 _6394_ (.A1(_2373_),
    .A2(_2380_),
    .A3(_2381_),
    .B1(_2383_),
    .X(_2384_));
 sky130_fd_sc_hd__nor2_1 _6395_ (.A(_2102_),
    .B(_2293_),
    .Y(_2385_));
 sky130_fd_sc_hd__nand2_1 _6396_ (.A(_2092_),
    .B(_2385_),
    .Y(_2386_));
 sky130_fd_sc_hd__clkbuf_4 _6397_ (.A(_2386_),
    .X(_2387_));
 sky130_fd_sc_hd__or2_4 _6398_ (.A(_2072_),
    .B(_2170_),
    .X(_2388_));
 sky130_fd_sc_hd__or2_2 _6399_ (.A(_2117_),
    .B(_2388_),
    .X(_2389_));
 sky130_fd_sc_hd__or2_1 _6400_ (.A(_2150_),
    .B(_2388_),
    .X(_2390_));
 sky130_fd_sc_hd__buf_4 _6401_ (.A(_2390_),
    .X(_2391_));
 sky130_fd_sc_hd__or2_1 _6402_ (.A(_2092_),
    .B(_2293_),
    .X(_2392_));
 sky130_fd_sc_hd__o221a_1 _6403_ (.A1(_2387_),
    .A2(_2389_),
    .B1(_2391_),
    .B2(_2392_),
    .C1(_2217_),
    .X(_2393_));
 sky130_fd_sc_hd__o21ai_1 _6404_ (.A1(_2128_),
    .A2(_2101_),
    .B1(_2393_),
    .Y(_2394_));
 sky130_fd_sc_hd__or2_1 _6405_ (.A(_2110_),
    .B(_2277_),
    .X(_2395_));
 sky130_fd_sc_hd__clkbuf_2 _6406_ (.A(_2395_),
    .X(_2396_));
 sky130_fd_sc_hd__nor2_1 _6407_ (.A(_2140_),
    .B(_2396_),
    .Y(_2397_));
 sky130_fd_sc_hd__or2_1 _6408_ (.A(_2138_),
    .B(_2153_),
    .X(_2398_));
 sky130_fd_sc_hd__nor2_1 _6409_ (.A(_2106_),
    .B(_2398_),
    .Y(_2399_));
 sky130_fd_sc_hd__nor2_8 _6410_ (.A(_1519_),
    .B(_2067_),
    .Y(_2400_));
 sky130_fd_sc_hd__clkbuf_4 _6411_ (.A(_2400_),
    .X(_2401_));
 sky130_fd_sc_hd__nor2_2 _6412_ (.A(_2173_),
    .B(_2100_),
    .Y(_2402_));
 sky130_fd_sc_hd__nand2_4 _6413_ (.A(_2401_),
    .B(_2402_),
    .Y(_2403_));
 sky130_fd_sc_hd__nor2_1 _6414_ (.A(_2295_),
    .B(_2403_),
    .Y(_2404_));
 sky130_fd_sc_hd__nand2_4 _6415_ (.A(_2161_),
    .B(_2109_),
    .Y(_2405_));
 sky130_fd_sc_hd__or2_2 _6416_ (.A(_2100_),
    .B(_2388_),
    .X(_2406_));
 sky130_fd_sc_hd__or2_4 _6417_ (.A(_2405_),
    .B(_2406_),
    .X(_2407_));
 sky130_fd_sc_hd__a21oi_1 _6418_ (.A1(_2356_),
    .A2(_2295_),
    .B1(_2407_),
    .Y(_2408_));
 sky130_fd_sc_hd__nand2_4 _6419_ (.A(_2174_),
    .B(_2401_),
    .Y(_2409_));
 sky130_fd_sc_hd__nor2_1 _6420_ (.A(_2293_),
    .B(_2125_),
    .Y(_2410_));
 sky130_fd_sc_hd__buf_4 _6421_ (.A(_2410_),
    .X(_2411_));
 sky130_fd_sc_hd__nor2_2 _6422_ (.A(_2411_),
    .B(_2364_),
    .Y(_2412_));
 sky130_fd_sc_hd__nor2_1 _6423_ (.A(_2409_),
    .B(_2412_),
    .Y(_2413_));
 sky130_fd_sc_hd__buf_2 _6424_ (.A(_2405_),
    .X(_2414_));
 sky130_fd_sc_hd__or2_1 _6425_ (.A(_2151_),
    .B(_2414_),
    .X(_2415_));
 sky130_fd_sc_hd__or2_1 _6426_ (.A(_2295_),
    .B(_2409_),
    .X(_2416_));
 sky130_fd_sc_hd__or2_4 _6427_ (.A(_2293_),
    .B(_2094_),
    .X(_2417_));
 sky130_fd_sc_hd__nor2_1 _6428_ (.A(_2173_),
    .B(_2150_),
    .Y(_2418_));
 sky130_fd_sc_hd__nand2_1 _6429_ (.A(_2400_),
    .B(_2418_),
    .Y(_2419_));
 sky130_fd_sc_hd__clkbuf_4 _6430_ (.A(_2419_),
    .X(_2420_));
 sky130_fd_sc_hd__o22a_1 _6431_ (.A1(_2152_),
    .A2(_2316_),
    .B1(_2417_),
    .B2(_2420_),
    .X(_2421_));
 sky130_fd_sc_hd__o211a_1 _6432_ (.A1(_2412_),
    .A2(_2415_),
    .B1(_2416_),
    .C1(_2421_),
    .X(_2422_));
 sky130_fd_sc_hd__or4b_1 _6433_ (.A(_2404_),
    .B(_2408_),
    .C(_2413_),
    .D_N(_2422_),
    .X(_2423_));
 sky130_fd_sc_hd__nor2_1 _6434_ (.A(_2409_),
    .B(_2417_),
    .Y(_2424_));
 sky130_fd_sc_hd__nor2_1 _6435_ (.A(_2295_),
    .B(_2420_),
    .Y(_2425_));
 sky130_fd_sc_hd__nand2_1 _6436_ (.A(_2392_),
    .B(_2363_),
    .Y(_2426_));
 sky130_fd_sc_hd__or3_1 _6437_ (.A(_2072_),
    .B(_2099_),
    .C(_2171_),
    .X(_2427_));
 sky130_fd_sc_hd__buf_4 _6438_ (.A(_2427_),
    .X(_2428_));
 sky130_fd_sc_hd__nor2_4 _6439_ (.A(_2405_),
    .B(_2428_),
    .Y(_2429_));
 sky130_fd_sc_hd__nor2_4 _6440_ (.A(_2293_),
    .B(_2094_),
    .Y(_2430_));
 sky130_fd_sc_hd__nand2_2 _6441_ (.A(_2400_),
    .B(_2430_),
    .Y(_2431_));
 sky130_fd_sc_hd__nor2_1 _6442_ (.A(_2406_),
    .B(_2431_),
    .Y(_2432_));
 sky130_fd_sc_hd__or2_1 _6443_ (.A(_2276_),
    .B(_2388_),
    .X(_2433_));
 sky130_fd_sc_hd__clkbuf_4 _6444_ (.A(_2433_),
    .X(_2434_));
 sky130_fd_sc_hd__nor2_2 _6445_ (.A(_2405_),
    .B(_2434_),
    .Y(_2435_));
 sky130_fd_sc_hd__and3_2 _6446_ (.A(_2216_),
    .B(_2306_),
    .C(_2400_),
    .X(_2436_));
 sky130_fd_sc_hd__a21o_1 _6447_ (.A1(_2426_),
    .A2(_2435_),
    .B1(_2436_),
    .X(_2437_));
 sky130_fd_sc_hd__a211o_1 _6448_ (.A1(_2426_),
    .A2(_2429_),
    .B1(_2432_),
    .C1(_2437_),
    .X(_2438_));
 sky130_fd_sc_hd__nor2_1 _6449_ (.A(_2386_),
    .B(_2407_),
    .Y(_2439_));
 sky130_fd_sc_hd__nand2_1 _6450_ (.A(_2338_),
    .B(_2400_),
    .Y(_2440_));
 sky130_fd_sc_hd__nor2_1 _6451_ (.A(_2434_),
    .B(_2440_),
    .Y(_2441_));
 sky130_fd_sc_hd__nor2_1 _6452_ (.A(_2391_),
    .B(_2440_),
    .Y(_2442_));
 sky130_fd_sc_hd__or2_1 _6453_ (.A(_2151_),
    .B(_2440_),
    .X(_2443_));
 sky130_fd_sc_hd__or4b_1 _6454_ (.A(_2439_),
    .B(_2441_),
    .C(_2442_),
    .D_N(_2443_),
    .X(_2444_));
 sky130_fd_sc_hd__or4_1 _6455_ (.A(_2424_),
    .B(_2425_),
    .C(_2438_),
    .D(_2444_),
    .X(_2445_));
 sky130_fd_sc_hd__a21oi_1 _6456_ (.A1(_2357_),
    .A2(_2386_),
    .B1(_2403_),
    .Y(_2446_));
 sky130_fd_sc_hd__or2_1 _6457_ (.A(_2403_),
    .B(_2417_),
    .X(_2447_));
 sky130_fd_sc_hd__o21ai_1 _6458_ (.A1(_2357_),
    .A2(_2420_),
    .B1(_2447_),
    .Y(_2448_));
 sky130_fd_sc_hd__nor2_2 _6459_ (.A(_2173_),
    .B(_2276_),
    .Y(_2449_));
 sky130_fd_sc_hd__nand2_2 _6460_ (.A(_2400_),
    .B(_2449_),
    .Y(_2450_));
 sky130_fd_sc_hd__or2_1 _6461_ (.A(_2294_),
    .B(_2450_),
    .X(_2451_));
 sky130_fd_sc_hd__nand2_1 _6462_ (.A(_2338_),
    .B(_2429_),
    .Y(_2452_));
 sky130_fd_sc_hd__nand2_1 _6463_ (.A(_2451_),
    .B(_2452_),
    .Y(_2453_));
 sky130_fd_sc_hd__a21oi_1 _6464_ (.A1(_2356_),
    .A2(_2363_),
    .B1(_2450_),
    .Y(_2454_));
 sky130_fd_sc_hd__nor2_2 _6465_ (.A(_2396_),
    .B(_2316_),
    .Y(_2455_));
 sky130_fd_sc_hd__nor2_1 _6466_ (.A(_2386_),
    .B(_2420_),
    .Y(_2456_));
 sky130_fd_sc_hd__or4_1 _6467_ (.A(_2453_),
    .B(_2454_),
    .C(_2455_),
    .D(_2456_),
    .X(_2457_));
 sky130_fd_sc_hd__or4_1 _6468_ (.A(_2445_),
    .B(_2446_),
    .C(_2448_),
    .D(_2457_),
    .X(_2458_));
 sky130_fd_sc_hd__or4_1 _6469_ (.A(_2397_),
    .B(_2399_),
    .C(_2423_),
    .D(_2458_),
    .X(_2459_));
 sky130_fd_sc_hd__nand2_1 _6470_ (.A(_2375_),
    .B(_2376_),
    .Y(_2460_));
 sky130_fd_sc_hd__or3_1 _6471_ (.A(_2086_),
    .B(_2460_),
    .C(_2379_),
    .X(_2461_));
 sky130_fd_sc_hd__or2_1 _6472_ (.A(_2371_),
    .B(_2461_),
    .X(_2462_));
 sky130_fd_sc_hd__nor3_1 _6473_ (.A(_2103_),
    .B(_2095_),
    .C(_2462_),
    .Y(_2463_));
 sky130_fd_sc_hd__a211o_1 _6474_ (.A1(_2310_),
    .A2(_2394_),
    .B1(_2459_),
    .C1(_2463_),
    .X(_2464_));
 sky130_fd_sc_hd__or4_1 _6475_ (.A(_2136_),
    .B(_2129_),
    .C(_2384_),
    .D(_2464_),
    .X(_2465_));
 sky130_fd_sc_hd__or3_1 _6476_ (.A(_2124_),
    .B(_2098_),
    .C(_2111_),
    .X(_2466_));
 sky130_fd_sc_hd__clkinv_2 _6477_ (.A(_2461_),
    .Y(_2467_));
 sky130_fd_sc_hd__and3_1 _6478_ (.A(_2306_),
    .B(_2381_),
    .C(_2467_),
    .X(_2468_));
 sky130_fd_sc_hd__nor2_1 _6479_ (.A(_2091_),
    .B(_2134_),
    .Y(_2469_));
 sky130_fd_sc_hd__nor2_1 _6480_ (.A(_2171_),
    .B(_2388_),
    .Y(_2470_));
 sky130_fd_sc_hd__nand2_1 _6481_ (.A(_2310_),
    .B(_2470_),
    .Y(_2471_));
 sky130_fd_sc_hd__nor2_1 _6482_ (.A(_2392_),
    .B(_2471_),
    .Y(_2472_));
 sky130_fd_sc_hd__or4_1 _6483_ (.A(_2466_),
    .B(_2468_),
    .C(_2469_),
    .D(_2472_),
    .X(_2473_));
 sky130_fd_sc_hd__or2_1 _6484_ (.A(_2465_),
    .B(_2473_),
    .X(_2474_));
 sky130_fd_sc_hd__a31o_1 _6485_ (.A1(_2360_),
    .A2(_2361_),
    .A3(_2430_),
    .B1(_1947_),
    .X(_2475_));
 sky130_fd_sc_hd__inv_2 _6486_ (.A(_2475_),
    .Y(_2476_));
 sky130_fd_sc_hd__o22a_1 _6487_ (.A1(_2120_),
    .A2(_2295_),
    .B1(_2417_),
    .B2(_2153_),
    .X(_2477_));
 sky130_fd_sc_hd__or2_1 _6488_ (.A(_2108_),
    .B(_2414_),
    .X(_2478_));
 sky130_fd_sc_hd__clkbuf_4 _6489_ (.A(_2478_),
    .X(_2479_));
 sky130_fd_sc_hd__nor2_1 _6490_ (.A(_2151_),
    .B(_2479_),
    .Y(_2480_));
 sky130_fd_sc_hd__nor2_1 _6491_ (.A(_2191_),
    .B(_2396_),
    .Y(_2481_));
 sky130_fd_sc_hd__nor2_2 _6492_ (.A(_2115_),
    .B(_2419_),
    .Y(_2482_));
 sky130_fd_sc_hd__or2_1 _6493_ (.A(_2101_),
    .B(_2263_),
    .X(_2483_));
 sky130_fd_sc_hd__nor2_1 _6494_ (.A(_2110_),
    .B(_2483_),
    .Y(_2484_));
 sky130_fd_sc_hd__nor2_1 _6495_ (.A(_2396_),
    .B(_2356_),
    .Y(_2485_));
 sky130_fd_sc_hd__or4_1 _6496_ (.A(_2481_),
    .B(_2482_),
    .C(_2484_),
    .D(_2485_),
    .X(_2486_));
 sky130_fd_sc_hd__nor2_2 _6497_ (.A(_2115_),
    .B(_2403_),
    .Y(_2487_));
 sky130_fd_sc_hd__nand2_1 _6498_ (.A(_2138_),
    .B(_2112_),
    .Y(_2488_));
 sky130_fd_sc_hd__or2_1 _6499_ (.A(_2113_),
    .B(_2488_),
    .X(_2489_));
 sky130_fd_sc_hd__buf_4 _6500_ (.A(_2489_),
    .X(_2490_));
 sky130_fd_sc_hd__o22a_1 _6501_ (.A1(_2108_),
    .A2(_2403_),
    .B1(_2420_),
    .B2(_2490_),
    .X(_2491_));
 sky130_fd_sc_hd__or4b_1 _6502_ (.A(_2480_),
    .B(_2486_),
    .C(_2487_),
    .D_N(_2491_),
    .X(_2492_));
 sky130_fd_sc_hd__clkbuf_4 _6503_ (.A(_2401_),
    .X(_2493_));
 sky130_fd_sc_hd__or4b_4 _6504_ (.A(_1519_),
    .B(net146),
    .C(net145),
    .D_N(net144),
    .X(_2494_));
 sky130_fd_sc_hd__or2_1 _6505_ (.A(_2277_),
    .B(_2417_),
    .X(_2495_));
 sky130_fd_sc_hd__nor2_1 _6506_ (.A(_2494_),
    .B(_2495_),
    .Y(_2496_));
 sky130_fd_sc_hd__nand2_1 _6507_ (.A(_2205_),
    .B(_2216_),
    .Y(_2497_));
 sky130_fd_sc_hd__nand2_1 _6508_ (.A(_2497_),
    .B(_2495_),
    .Y(_2498_));
 sky130_fd_sc_hd__a21o_1 _6509_ (.A1(_2391_),
    .A2(_2434_),
    .B1(_2140_),
    .X(_2499_));
 sky130_fd_sc_hd__nand2_2 _6510_ (.A(_2216_),
    .B(_2338_),
    .Y(_2500_));
 sky130_fd_sc_hd__o211ai_1 _6511_ (.A1(_2389_),
    .A2(_2488_),
    .B1(_2499_),
    .C1(_2500_),
    .Y(_2501_));
 sky130_fd_sc_hd__o22a_1 _6512_ (.A1(_2493_),
    .A2(_2496_),
    .B1(_2498_),
    .B2(_2501_),
    .X(_2502_));
 sky130_fd_sc_hd__nor2_1 _6513_ (.A(_2108_),
    .B(_2409_),
    .Y(_2503_));
 sky130_fd_sc_hd__inv_2 _6514_ (.A(_2403_),
    .Y(_2504_));
 sky130_fd_sc_hd__nor2_2 _6515_ (.A(_2115_),
    .B(_2409_),
    .Y(_2505_));
 sky130_fd_sc_hd__a21o_1 _6516_ (.A1(_2275_),
    .A2(_2504_),
    .B1(_2505_),
    .X(_2506_));
 sky130_fd_sc_hd__or4_1 _6517_ (.A(_2492_),
    .B(_2502_),
    .C(_2503_),
    .D(_2506_),
    .X(_2507_));
 sky130_fd_sc_hd__nor2_4 _6518_ (.A(_2405_),
    .B(_2406_),
    .Y(_2508_));
 sky130_fd_sc_hd__or2_1 _6519_ (.A(_2414_),
    .B(_2434_),
    .X(_2509_));
 sky130_fd_sc_hd__nor2_1 _6520_ (.A(_2509_),
    .B(_2490_),
    .Y(_2510_));
 sky130_fd_sc_hd__nand2_1 _6521_ (.A(_2181_),
    .B(_2493_),
    .Y(_2511_));
 sky130_fd_sc_hd__nor2_1 _6522_ (.A(_2434_),
    .B(_2511_),
    .Y(_2512_));
 sky130_fd_sc_hd__a211o_1 _6523_ (.A1(_2215_),
    .A2(_2508_),
    .B1(_2510_),
    .C1(_2512_),
    .X(_2513_));
 sky130_fd_sc_hd__or3_1 _6524_ (.A(_2110_),
    .B(_2277_),
    .C(_2417_),
    .X(_2514_));
 sky130_fd_sc_hd__o21a_1 _6525_ (.A1(_2105_),
    .A2(_2398_),
    .B1(_2514_),
    .X(_2515_));
 sky130_fd_sc_hd__or2_1 _6526_ (.A(_2101_),
    .B(_2431_),
    .X(_2516_));
 sky130_fd_sc_hd__or2_1 _6527_ (.A(_2406_),
    .B(_2511_),
    .X(_2517_));
 sky130_fd_sc_hd__or2_1 _6528_ (.A(_2428_),
    .B(_2511_),
    .X(_2518_));
 sky130_fd_sc_hd__or2_2 _6529_ (.A(_2115_),
    .B(_2450_),
    .X(_2519_));
 sky130_fd_sc_hd__and4_1 _6530_ (.A(_2516_),
    .B(_2517_),
    .C(_2518_),
    .D(_2519_),
    .X(_2520_));
 sky130_fd_sc_hd__or2_1 _6531_ (.A(_2414_),
    .B(_2428_),
    .X(_2521_));
 sky130_fd_sc_hd__o32a_1 _6532_ (.A1(_2106_),
    .A2(_2113_),
    .A3(_2521_),
    .B1(_2415_),
    .B2(_2140_),
    .X(_2522_));
 sky130_fd_sc_hd__o211ai_2 _6533_ (.A1(_2092_),
    .A2(_2149_),
    .B1(_2112_),
    .C1(_2102_),
    .Y(_2523_));
 sky130_fd_sc_hd__o32a_1 _6534_ (.A1(_2173_),
    .A2(_2414_),
    .A3(_2523_),
    .B1(_2490_),
    .B2(_2407_),
    .X(_2524_));
 sky130_fd_sc_hd__nor2_2 _6535_ (.A(_2151_),
    .B(_2414_),
    .Y(_2525_));
 sky130_fd_sc_hd__nand2_1 _6536_ (.A(_2275_),
    .B(_2525_),
    .Y(_2526_));
 sky130_fd_sc_hd__o32a_1 _6537_ (.A1(_2101_),
    .A2(_2387_),
    .A3(_2494_),
    .B1(_2450_),
    .B2(_2108_),
    .X(_2527_));
 sky130_fd_sc_hd__o311a_1 _6538_ (.A1(_2110_),
    .A2(_2417_),
    .A3(_2428_),
    .B1(_2526_),
    .C1(_2527_),
    .X(_2528_));
 sky130_fd_sc_hd__and4_1 _6539_ (.A(_2520_),
    .B(_2522_),
    .C(_2524_),
    .D(_2528_),
    .X(_2529_));
 sky130_fd_sc_hd__and4bb_1 _6540_ (.A_N(_2507_),
    .B_N(_2513_),
    .C(_2515_),
    .D(_2529_),
    .X(_2530_));
 sky130_fd_sc_hd__nand2_1 _6541_ (.A(_2477_),
    .B(_2530_),
    .Y(_2531_));
 sky130_fd_sc_hd__or4_1 _6542_ (.A(_2358_),
    .B(_2285_),
    .C(_2365_),
    .D(_2531_),
    .X(_2532_));
 sky130_fd_sc_hd__nor2_8 _6543_ (.A(net1537),
    .B(_1947_),
    .Y(_2533_));
 sky130_fd_sc_hd__a221o_1 _6544_ (.A1(_2372_),
    .A2(_2474_),
    .B1(_2476_),
    .B2(_2532_),
    .C1(_2533_),
    .X(_2534_));
 sky130_fd_sc_hd__o32a_1 _6545_ (.A1(_2283_),
    .A2(_2368_),
    .A3(_2534_),
    .B1(_1949_),
    .B2(net591),
    .X(_0377_));
 sky130_fd_sc_hd__or2_1 _6546_ (.A(_2129_),
    .B(_2296_),
    .X(_2535_));
 sky130_fd_sc_hd__nand2_1 _6547_ (.A(_2168_),
    .B(net394),
    .Y(_2536_));
 sky130_fd_sc_hd__nor2_1 _6548_ (.A(_2209_),
    .B(_2536_),
    .Y(_2537_));
 sky130_fd_sc_hd__or2_1 _6549_ (.A(_2075_),
    .B(_2138_),
    .X(_2538_));
 sky130_fd_sc_hd__nor2_1 _6550_ (.A(_2538_),
    .B(_2153_),
    .Y(_2539_));
 sky130_fd_sc_hd__nand2_2 _6551_ (.A(_2209_),
    .B(_2123_),
    .Y(_2540_));
 sky130_fd_sc_hd__nor2_1 _6552_ (.A(_2263_),
    .B(_2180_),
    .Y(_2541_));
 sky130_fd_sc_hd__or2_1 _6553_ (.A(_2541_),
    .B(_2311_),
    .X(_2542_));
 sky130_fd_sc_hd__a21o_1 _6554_ (.A1(_2269_),
    .A2(_2318_),
    .B1(_2320_),
    .X(_2543_));
 sky130_fd_sc_hd__or2_1 _6555_ (.A(_2259_),
    .B(_2322_),
    .X(_2544_));
 sky130_fd_sc_hd__nor2_2 _6556_ (.A(_2210_),
    .B(_2169_),
    .Y(_2545_));
 sky130_fd_sc_hd__a21oi_1 _6557_ (.A1(_2217_),
    .A2(_2500_),
    .B1(_2194_),
    .Y(_2546_));
 sky130_fd_sc_hd__or3_1 _6558_ (.A(_2209_),
    .B(_2196_),
    .C(_2178_),
    .X(_2547_));
 sky130_fd_sc_hd__inv_2 _6559_ (.A(_2547_),
    .Y(_2548_));
 sky130_fd_sc_hd__or2_1 _6560_ (.A(_2333_),
    .B(_2548_),
    .X(_2549_));
 sky130_fd_sc_hd__or2_1 _6561_ (.A(_2210_),
    .B(_2187_),
    .X(_2550_));
 sky130_fd_sc_hd__nor2_1 _6562_ (.A(_2210_),
    .B(_2187_),
    .Y(_2551_));
 sky130_fd_sc_hd__nor2_1 _6563_ (.A(_2545_),
    .B(_2551_),
    .Y(_2552_));
 sky130_fd_sc_hd__inv_2 _6564_ (.A(_2122_),
    .Y(_2553_));
 sky130_fd_sc_hd__nor2_2 _6565_ (.A(_2103_),
    .B(_2553_),
    .Y(_2554_));
 sky130_fd_sc_hd__nor2_2 _6566_ (.A(_2301_),
    .B(_2554_),
    .Y(_2555_));
 sky130_fd_sc_hd__o22a_1 _6567_ (.A1(_2316_),
    .A2(_2550_),
    .B1(_2552_),
    .B2(_2555_),
    .X(_2556_));
 sky130_fd_sc_hd__or4b_1 _6568_ (.A(_2231_),
    .B(_2546_),
    .C(_2549_),
    .D_N(_2556_),
    .X(_2557_));
 sky130_fd_sc_hd__a221o_1 _6569_ (.A1(_2545_),
    .A2(_2306_),
    .B1(_2540_),
    .B2(_2335_),
    .C1(_2557_),
    .X(_2558_));
 sky130_fd_sc_hd__or2_1 _6570_ (.A(_2250_),
    .B(_2329_),
    .X(_2559_));
 sky130_fd_sc_hd__a22o_1 _6571_ (.A1(_2330_),
    .A2(_2269_),
    .B1(_2306_),
    .B2(_2335_),
    .X(_2560_));
 sky130_fd_sc_hd__a211o_1 _6572_ (.A1(_2330_),
    .A2(_2540_),
    .B1(_2559_),
    .C1(_2560_),
    .X(_2561_));
 sky130_fd_sc_hd__or2_1 _6573_ (.A(_2255_),
    .B(_2325_),
    .X(_2562_));
 sky130_fd_sc_hd__nor2_1 _6574_ (.A(_2249_),
    .B(_2555_),
    .Y(_2563_));
 sky130_fd_sc_hd__a211o_1 _6575_ (.A1(_2321_),
    .A2(_2540_),
    .B1(_2562_),
    .C1(_2563_),
    .X(_2564_));
 sky130_fd_sc_hd__or4_1 _6576_ (.A(_2228_),
    .B(_2558_),
    .C(_2561_),
    .D(_2564_),
    .X(_2565_));
 sky130_fd_sc_hd__a211o_1 _6577_ (.A1(_2206_),
    .A2(_2540_),
    .B1(_2544_),
    .C1(_2565_),
    .X(_2566_));
 sky130_fd_sc_hd__a211o_1 _6578_ (.A1(_2318_),
    .A2(_2540_),
    .B1(_2543_),
    .C1(_2566_),
    .X(_2567_));
 sky130_fd_sc_hd__a2111o_1 _6579_ (.A1(_2305_),
    .A2(_2540_),
    .B1(_2567_),
    .C1(_2266_),
    .D1(_2317_),
    .X(_2568_));
 sky130_fd_sc_hd__a311o_1 _6580_ (.A1(_2205_),
    .A2(_2303_),
    .A3(_2299_),
    .B1(_2300_),
    .C1(_2304_),
    .X(_2569_));
 sky130_fd_sc_hd__a2111o_1 _6581_ (.A1(_2270_),
    .A2(_2540_),
    .B1(_2542_),
    .C1(_2568_),
    .D1(_2569_),
    .X(_2570_));
 sky130_fd_sc_hd__or4_1 _6582_ (.A(_2535_),
    .B(_2537_),
    .C(_2539_),
    .D(_2570_),
    .X(_2571_));
 sky130_fd_sc_hd__or4_1 _6583_ (.A(_2124_),
    .B(_2285_),
    .C(_2290_),
    .D(_2571_),
    .X(_2572_));
 sky130_fd_sc_hd__o31a_1 _6584_ (.A1(_2098_),
    .A2(_2286_),
    .A3(_2572_),
    .B1(_2367_),
    .X(_2573_));
 sky130_fd_sc_hd__or2_1 _6585_ (.A(_2116_),
    .B(_2286_),
    .X(_2574_));
 sky130_fd_sc_hd__or2_1 _6586_ (.A(_2111_),
    .B(_2285_),
    .X(_2575_));
 sky130_fd_sc_hd__nor2_1 _6587_ (.A(_2132_),
    .B(_2115_),
    .Y(_2576_));
 sky130_fd_sc_hd__or2_2 _6588_ (.A(_2136_),
    .B(_2297_),
    .X(_2577_));
 sky130_fd_sc_hd__and4_1 _6589_ (.A(_2075_),
    .B(_2102_),
    .C(_2103_),
    .D(_2121_),
    .X(_2578_));
 sky130_fd_sc_hd__o21a_1 _6590_ (.A1(_2215_),
    .A2(_2181_),
    .B1(_2184_),
    .X(_2579_));
 sky130_fd_sc_hd__nand2_1 _6591_ (.A(_2192_),
    .B(_2526_),
    .Y(_2580_));
 sky130_fd_sc_hd__nor2_1 _6592_ (.A(_2284_),
    .B(_2198_),
    .Y(_2581_));
 sky130_fd_sc_hd__o21ai_1 _6593_ (.A1(_2134_),
    .A2(_2521_),
    .B1(_2199_),
    .Y(_2582_));
 sky130_fd_sc_hd__o21ai_1 _6594_ (.A1(_2284_),
    .A2(_2203_),
    .B1(_2519_),
    .Y(_2583_));
 sky130_fd_sc_hd__a32o_1 _6595_ (.A1(_2275_),
    .A2(_2401_),
    .A3(_2402_),
    .B1(_2206_),
    .B2(_2205_),
    .X(_2584_));
 sky130_fd_sc_hd__or2_1 _6596_ (.A(_2173_),
    .B(_2276_),
    .X(_2585_));
 sky130_fd_sc_hd__nand2_2 _6597_ (.A(_2275_),
    .B(_2400_),
    .Y(_2586_));
 sky130_fd_sc_hd__o21ai_1 _6598_ (.A1(_2585_),
    .A2(_2586_),
    .B1(_2261_),
    .Y(_2587_));
 sky130_fd_sc_hd__a32o_1 _6599_ (.A1(_2174_),
    .A2(_2275_),
    .A3(_2400_),
    .B1(_2330_),
    .B2(_2205_),
    .X(_2588_));
 sky130_fd_sc_hd__nor2_1 _6600_ (.A(_2244_),
    .B(_2249_),
    .Y(_2589_));
 sky130_fd_sc_hd__a31o_1 _6601_ (.A1(_2174_),
    .A2(_2181_),
    .A3(_2400_),
    .B1(_2589_),
    .X(_2590_));
 sky130_fd_sc_hd__a22o_1 _6602_ (.A1(_2335_),
    .A2(_2205_),
    .B1(_2275_),
    .B2(_2508_),
    .X(_2591_));
 sky130_fd_sc_hd__nor2_1 _6603_ (.A(_2223_),
    .B(_2244_),
    .Y(_2592_));
 sky130_fd_sc_hd__a21o_1 _6604_ (.A1(_2181_),
    .A2(_2435_),
    .B1(_2592_),
    .X(_2593_));
 sky130_fd_sc_hd__o221a_1 _6605_ (.A1(_2127_),
    .A2(_2147_),
    .B1(_2391_),
    .B2(_2586_),
    .C1(_2239_),
    .X(_2594_));
 sky130_fd_sc_hd__o22a_1 _6606_ (.A1(_2234_),
    .A2(_2244_),
    .B1(_2114_),
    .B2(_2390_),
    .X(_2595_));
 sky130_fd_sc_hd__nor2_1 _6607_ (.A(_2214_),
    .B(_2595_),
    .Y(_2596_));
 sky130_fd_sc_hd__o22ai_1 _6608_ (.A1(_2147_),
    .A2(_2114_),
    .B1(_2183_),
    .B2(_2217_),
    .Y(_2597_));
 sky130_fd_sc_hd__nand2_1 _6609_ (.A(_2181_),
    .B(_2470_),
    .Y(_2598_));
 sky130_fd_sc_hd__or2_1 _6610_ (.A(_2244_),
    .B(_2236_),
    .X(_2599_));
 sky130_fd_sc_hd__a21oi_1 _6611_ (.A1(_2598_),
    .A2(_2599_),
    .B1(_2214_),
    .Y(_2600_));
 sky130_fd_sc_hd__a2111oi_1 _6612_ (.A1(_2218_),
    .A2(_2338_),
    .B1(_2596_),
    .C1(_2597_),
    .D1(_2600_),
    .Y(_2601_));
 sky130_fd_sc_hd__o211a_1 _6613_ (.A1(_2434_),
    .A2(_2586_),
    .B1(_2594_),
    .C1(net367),
    .X(_2602_));
 sky130_fd_sc_hd__or4b_1 _6614_ (.A(_2230_),
    .B(_2591_),
    .C(_2593_),
    .D_N(_2602_),
    .X(_2603_));
 sky130_fd_sc_hd__o21ai_1 _6615_ (.A1(_2115_),
    .A2(_2407_),
    .B1(_2245_),
    .Y(_2604_));
 sky130_fd_sc_hd__or4_1 _6616_ (.A(_2588_),
    .B(_2590_),
    .C(_2603_),
    .D(_2604_),
    .X(_2605_));
 sky130_fd_sc_hd__o31ai_1 _6617_ (.A1(_2173_),
    .A2(_2150_),
    .A3(_2586_),
    .B1(_2256_),
    .Y(_2606_));
 sky130_fd_sc_hd__or4_1 _6618_ (.A(_2254_),
    .B(_2482_),
    .C(_2605_),
    .D(_2606_),
    .X(_2607_));
 sky130_fd_sc_hd__or4_1 _6619_ (.A(_2583_),
    .B(_2584_),
    .C(_2587_),
    .D(_2607_),
    .X(_2608_));
 sky130_fd_sc_hd__or4_1 _6620_ (.A(_2581_),
    .B(_2487_),
    .C(_2582_),
    .D(_2608_),
    .X(_2609_));
 sky130_fd_sc_hd__nor2_1 _6621_ (.A(_2284_),
    .B(_2189_),
    .Y(_2610_));
 sky130_fd_sc_hd__a2111o_1 _6622_ (.A1(_2181_),
    .A2(_2429_),
    .B1(_2580_),
    .C1(_2609_),
    .D1(_2610_),
    .X(_2611_));
 sky130_fd_sc_hd__nor2_2 _6623_ (.A(_2130_),
    .B(_2214_),
    .Y(_2612_));
 sky130_fd_sc_hd__nor2_2 _6624_ (.A(_2284_),
    .B(_2180_),
    .Y(_2613_));
 sky130_fd_sc_hd__a41o_1 _6625_ (.A1(_2082_),
    .A2(_2083_),
    .A3(_2612_),
    .A4(_2181_),
    .B1(_2613_),
    .X(_2614_));
 sky130_fd_sc_hd__or4_1 _6626_ (.A(_2148_),
    .B(_2579_),
    .C(_2611_),
    .D(_2614_),
    .X(_2615_));
 sky130_fd_sc_hd__or4_1 _6627_ (.A(_2576_),
    .B(_2577_),
    .C(_2578_),
    .D(_2615_),
    .X(_2616_));
 sky130_fd_sc_hd__or3_1 _6628_ (.A(_2102_),
    .B(_2106_),
    .C(_2120_),
    .X(_2617_));
 sky130_fd_sc_hd__or4b_1 _6629_ (.A(_2574_),
    .B(_2575_),
    .C(_2616_),
    .D_N(_2617_),
    .X(_2618_));
 sky130_fd_sc_hd__or2_1 _6630_ (.A(_2358_),
    .B(_2469_),
    .X(_2619_));
 sky130_fd_sc_hd__nand2_1 _6631_ (.A(_2134_),
    .B(_2387_),
    .Y(_2620_));
 sky130_fd_sc_hd__a21oi_1 _6632_ (.A1(_2117_),
    .A2(_2338_),
    .B1(_2620_),
    .Y(_2621_));
 sky130_fd_sc_hd__nand2_1 _6633_ (.A(_2158_),
    .B(_2360_),
    .Y(_2622_));
 sky130_fd_sc_hd__o21ai_1 _6634_ (.A1(_2388_),
    .A2(_2621_),
    .B1(_2622_),
    .Y(_2623_));
 sky130_fd_sc_hd__nor2_2 _6635_ (.A(_2138_),
    .B(_2152_),
    .Y(_2624_));
 sky130_fd_sc_hd__o21ai_2 _6636_ (.A1(_2115_),
    .A2(_2420_),
    .B1(_2451_),
    .Y(_2625_));
 sky130_fd_sc_hd__a21o_1 _6637_ (.A1(_2075_),
    .A2(_2624_),
    .B1(_2625_),
    .X(_2626_));
 sky130_fd_sc_hd__or2_1 _6638_ (.A(_2397_),
    .B(_2481_),
    .X(_2627_));
 sky130_fd_sc_hd__o21ai_1 _6639_ (.A1(_2153_),
    .A2(_2387_),
    .B1(_2516_),
    .Y(_2628_));
 sky130_fd_sc_hd__nor2_1 _6640_ (.A(_2173_),
    .B(_2414_),
    .Y(_2629_));
 sky130_fd_sc_hd__a21o_1 _6641_ (.A1(_2171_),
    .A2(_2629_),
    .B1(_2429_),
    .X(_2630_));
 sky130_fd_sc_hd__nand2_1 _6642_ (.A(_2416_),
    .B(_2517_),
    .Y(_2631_));
 sky130_fd_sc_hd__or2_1 _6643_ (.A(_2425_),
    .B(_2505_),
    .X(_2632_));
 sky130_fd_sc_hd__a21o_1 _6644_ (.A1(_2338_),
    .A2(_2429_),
    .B1(_2487_),
    .X(_2633_));
 sky130_fd_sc_hd__a2111o_1 _6645_ (.A1(_2620_),
    .A2(_2630_),
    .B1(_2631_),
    .C1(_2632_),
    .D1(_2633_),
    .X(_2634_));
 sky130_fd_sc_hd__or4_1 _6646_ (.A(_2626_),
    .B(_2627_),
    .C(_2628_),
    .D(_2634_),
    .X(_2635_));
 sky130_fd_sc_hd__a21oi_1 _6647_ (.A1(_2134_),
    .A2(_2387_),
    .B1(_2409_),
    .Y(_2636_));
 sky130_fd_sc_hd__nand2_1 _6648_ (.A(_2443_),
    .B(_2518_),
    .Y(_2637_));
 sky130_fd_sc_hd__nand2_1 _6649_ (.A(_2360_),
    .B(_2361_),
    .Y(_2638_));
 sky130_fd_sc_hd__nor2_1 _6650_ (.A(_2108_),
    .B(_2638_),
    .Y(_2639_));
 sky130_fd_sc_hd__nor2_1 _6651_ (.A(_2396_),
    .B(_2412_),
    .Y(_2640_));
 sky130_fd_sc_hd__a31o_1 _6652_ (.A1(_2360_),
    .A2(_2364_),
    .A3(_2493_),
    .B1(_2496_),
    .X(_2641_));
 sky130_fd_sc_hd__or2_1 _6653_ (.A(_2640_),
    .B(_2641_),
    .X(_2642_));
 sky130_fd_sc_hd__or2b_1 _6654_ (.A(_2404_),
    .B_N(_2519_),
    .X(_2643_));
 sky130_fd_sc_hd__or3_1 _6655_ (.A(_2101_),
    .B(_2363_),
    .C(_2494_),
    .X(_2644_));
 sky130_fd_sc_hd__o21ai_1 _6656_ (.A1(_2389_),
    .A2(_2511_),
    .B1(_2644_),
    .Y(_2645_));
 sky130_fd_sc_hd__or4_1 _6657_ (.A(_2442_),
    .B(_2512_),
    .C(_2643_),
    .D(_2645_),
    .X(_2646_));
 sky130_fd_sc_hd__or2_1 _6658_ (.A(_2638_),
    .B(_2387_),
    .X(_2647_));
 sky130_fd_sc_hd__or4b_1 _6659_ (.A(_2639_),
    .B(_2642_),
    .C(_2646_),
    .D_N(_2647_),
    .X(_2648_));
 sky130_fd_sc_hd__nand2_1 _6660_ (.A(_2525_),
    .B(_2620_),
    .Y(_2649_));
 sky130_fd_sc_hd__or4b_1 _6661_ (.A(_2636_),
    .B(_2637_),
    .C(_2648_),
    .D_N(_2649_),
    .X(_2650_));
 sky130_fd_sc_hd__a211o_1 _6662_ (.A1(_2493_),
    .A2(_2623_),
    .B1(_2635_),
    .C1(_2650_),
    .X(_2651_));
 sky130_fd_sc_hd__o21a_1 _6663_ (.A1(_2619_),
    .A2(_2651_),
    .B1(_2476_),
    .X(_2652_));
 sky130_fd_sc_hd__or2_2 _6664_ (.A(_2124_),
    .B(_2358_),
    .X(_2653_));
 sky130_fd_sc_hd__nor2_1 _6665_ (.A(_2553_),
    .B(_2462_),
    .Y(_2654_));
 sky130_fd_sc_hd__xnor2_1 _6666_ (.A(_2149_),
    .B(_2315_),
    .Y(_2655_));
 sky130_fd_sc_hd__or2_1 _6667_ (.A(_2378_),
    .B(_2655_),
    .X(_2656_));
 sky130_fd_sc_hd__or3_1 _6668_ (.A(_2371_),
    .B(_2460_),
    .C(_2656_),
    .X(_2657_));
 sky130_fd_sc_hd__nor2_1 _6669_ (.A(_2097_),
    .B(_2657_),
    .Y(_2658_));
 sky130_fd_sc_hd__and3_1 _6670_ (.A(_2373_),
    .B(_2380_),
    .C(_2381_),
    .X(_2659_));
 sky130_fd_sc_hd__or2_1 _6671_ (.A(_2383_),
    .B(_2659_),
    .X(_2660_));
 sky130_fd_sc_hd__and3_1 _6672_ (.A(_2099_),
    .B(_2307_),
    .C(_2381_),
    .X(_2661_));
 sky130_fd_sc_hd__nand2_1 _6673_ (.A(_2270_),
    .B(_2373_),
    .Y(_2662_));
 sky130_fd_sc_hd__o21ai_1 _6674_ (.A1(_2357_),
    .A2(_2415_),
    .B1(_2662_),
    .Y(_2663_));
 sky130_fd_sc_hd__o21bai_1 _6675_ (.A1(_2428_),
    .A2(_2431_),
    .B1_N(_2312_),
    .Y(_2664_));
 sky130_fd_sc_hd__a22o_1 _6676_ (.A1(_2305_),
    .A2(_2373_),
    .B1(_2411_),
    .B2(_2429_),
    .X(_2665_));
 sky130_fd_sc_hd__a32o_1 _6677_ (.A1(_2411_),
    .A2(_2493_),
    .A3(_2402_),
    .B1(_2373_),
    .B2(_2318_),
    .X(_2666_));
 sky130_fd_sc_hd__a32o_1 _6678_ (.A1(_2411_),
    .A2(_2401_),
    .A3(_2449_),
    .B1(_2373_),
    .B2(_2206_),
    .X(_2667_));
 sky130_fd_sc_hd__a31o_1 _6679_ (.A1(_2401_),
    .A2(_2430_),
    .A3(_2449_),
    .B1(_2319_),
    .X(_2668_));
 sky130_fd_sc_hd__a31o_1 _6680_ (.A1(_2401_),
    .A2(_2430_),
    .A3(_2418_),
    .B1(_2323_),
    .X(_2669_));
 sky130_fd_sc_hd__nor2_1 _6681_ (.A(_2253_),
    .B(_2097_),
    .Y(_2670_));
 sky130_fd_sc_hd__a31o_1 _6682_ (.A1(_2411_),
    .A2(_2401_),
    .A3(_2418_),
    .B1(_2670_),
    .X(_2671_));
 sky130_fd_sc_hd__a31o_1 _6683_ (.A1(_2174_),
    .A2(_2411_),
    .A3(_2401_),
    .B1(_2326_),
    .X(_2672_));
 sky130_fd_sc_hd__a22o_1 _6684_ (.A1(_2330_),
    .A2(_2373_),
    .B1(_2411_),
    .B2(_2508_),
    .X(_2673_));
 sky130_fd_sc_hd__nor2_1 _6685_ (.A(_2391_),
    .B(_2431_),
    .Y(_2674_));
 sky130_fd_sc_hd__a21o_1 _6686_ (.A1(_2335_),
    .A2(_2220_),
    .B1(_2674_),
    .X(_2675_));
 sky130_fd_sc_hd__a21o_1 _6687_ (.A1(_2430_),
    .A2(_2435_),
    .B1(_2331_),
    .X(_2676_));
 sky130_fd_sc_hd__a22o_1 _6688_ (.A1(_2335_),
    .A2(_2373_),
    .B1(_2410_),
    .B2(_2435_),
    .X(_2677_));
 sky130_fd_sc_hd__o211a_1 _6689_ (.A1(_2410_),
    .A2(_2430_),
    .B1(_2470_),
    .C1(_2310_),
    .X(_2678_));
 sky130_fd_sc_hd__a31o_1 _6690_ (.A1(_2373_),
    .A2(_2310_),
    .A3(_2380_),
    .B1(_2468_),
    .X(_2679_));
 sky130_fd_sc_hd__or2b_1 _6691_ (.A(_2376_),
    .B_N(_2375_),
    .X(_2680_));
 sky130_fd_sc_hd__nand2_1 _6692_ (.A(_2086_),
    .B(_2655_),
    .Y(_2681_));
 sky130_fd_sc_hd__nor2_1 _6693_ (.A(_2680_),
    .B(_2681_),
    .Y(_2682_));
 sky130_fd_sc_hd__a21oi_1 _6694_ (.A1(_2217_),
    .A2(_2497_),
    .B1(_2382_),
    .Y(_2683_));
 sky130_fd_sc_hd__or2_1 _6695_ (.A(_2656_),
    .B(_2680_),
    .X(_2684_));
 sky130_fd_sc_hd__o22a_1 _6696_ (.A1(_2356_),
    .A2(_2391_),
    .B1(_2684_),
    .B2(_2097_),
    .X(_2685_));
 sky130_fd_sc_hd__nor2_1 _6697_ (.A(_2382_),
    .B(_2685_),
    .Y(_2686_));
 sky130_fd_sc_hd__a311o_1 _6698_ (.A1(_2373_),
    .A2(_2310_),
    .A3(_2682_),
    .B1(_2683_),
    .C1(_2686_),
    .X(_2687_));
 sky130_fd_sc_hd__a2111o_1 _6699_ (.A1(_2220_),
    .A2(_2545_),
    .B1(_2678_),
    .C1(_2679_),
    .D1(_2687_),
    .X(_2688_));
 sky130_fd_sc_hd__or4_1 _6700_ (.A(_2675_),
    .B(_2676_),
    .C(_2677_),
    .D(_2688_),
    .X(_2689_));
 sky130_fd_sc_hd__a2111o_1 _6701_ (.A1(_2508_),
    .A2(_2430_),
    .B1(_2673_),
    .C1(_2689_),
    .D1(_2327_),
    .X(_2690_));
 sky130_fd_sc_hd__a31o_1 _6702_ (.A1(_2174_),
    .A2(_2401_),
    .A3(_2430_),
    .B1(_2324_),
    .X(_2691_));
 sky130_fd_sc_hd__or4_1 _6703_ (.A(_2671_),
    .B(_2672_),
    .C(_2690_),
    .D(_2691_),
    .X(_2692_));
 sky130_fd_sc_hd__or4_1 _6704_ (.A(_2667_),
    .B(_2668_),
    .C(_2669_),
    .D(_2692_),
    .X(_2693_));
 sky130_fd_sc_hd__a31o_1 _6705_ (.A1(_2493_),
    .A2(_2402_),
    .A3(_2430_),
    .B1(_2313_),
    .X(_2694_));
 sky130_fd_sc_hd__or4_1 _6706_ (.A(_2665_),
    .B(_2666_),
    .C(_2693_),
    .D(_2694_),
    .X(_2695_));
 sky130_fd_sc_hd__or4_1 _6707_ (.A(_2661_),
    .B(_2663_),
    .C(_2664_),
    .D(_2695_),
    .X(_2696_));
 sky130_fd_sc_hd__or2_1 _6708_ (.A(_2154_),
    .B(_2298_),
    .X(_2697_));
 sky130_fd_sc_hd__or4_1 _6709_ (.A(_2658_),
    .B(_2660_),
    .C(_2696_),
    .D(_2697_),
    .X(_2698_));
 sky130_fd_sc_hd__or4_1 _6710_ (.A(_2278_),
    .B(_2296_),
    .C(_2654_),
    .D(_2698_),
    .X(_2699_));
 sky130_fd_sc_hd__o41a_1 _6711_ (.A1(_2098_),
    .A2(_2365_),
    .A3(_2653_),
    .A4(_2699_),
    .B1(_2372_),
    .X(_2700_));
 sky130_fd_sc_hd__a2111o_1 _6712_ (.A1(_2282_),
    .A2(_2618_),
    .B1(_2652_),
    .C1(_2533_),
    .D1(_2700_),
    .X(_2701_));
 sky130_fd_sc_hd__o22a_1 _6713_ (.A1(\wbbd_addr[1] ),
    .A2(_1949_),
    .B1(_2573_),
    .B2(_2701_),
    .X(_0378_));
 sky130_fd_sc_hd__or3b_2 _6714_ (.A(_2098_),
    .B(_2574_),
    .C_N(_2282_),
    .X(_2702_));
 sky130_fd_sc_hd__nor2_1 _6715_ (.A(_2215_),
    .B(_2301_),
    .Y(_2703_));
 sky130_fd_sc_hd__or3_2 _6716_ (.A(_2099_),
    .B(_2082_),
    .C(_2703_),
    .X(_2704_));
 sky130_fd_sc_hd__inv_2 _6717_ (.A(_2704_),
    .Y(_2705_));
 sky130_fd_sc_hd__a211o_1 _6718_ (.A1(_2612_),
    .A2(_2705_),
    .B1(_2482_),
    .C1(_2254_),
    .X(_2706_));
 sky130_fd_sc_hd__inv_2 _6719_ (.A(_2214_),
    .Y(_2707_));
 sky130_fd_sc_hd__a31o_1 _6720_ (.A1(_2707_),
    .A2(_2118_),
    .A3(_2705_),
    .B1(_2583_),
    .X(_2708_));
 sky130_fd_sc_hd__and2_2 _6721_ (.A(_2086_),
    .B(_2085_),
    .X(_2709_));
 sky130_fd_sc_hd__a311o_1 _6722_ (.A1(_2707_),
    .A2(_2709_),
    .A3(_2705_),
    .B1(_2505_),
    .C1(_2589_),
    .X(_2710_));
 sky130_fd_sc_hd__or3_1 _6723_ (.A(_2706_),
    .B(_2708_),
    .C(_2710_),
    .X(_2711_));
 sky130_fd_sc_hd__or3_2 _6724_ (.A(_2085_),
    .B(_2088_),
    .C(_2214_),
    .X(_2712_));
 sky130_fd_sc_hd__nor2_1 _6725_ (.A(_2712_),
    .B(_2704_),
    .Y(_2713_));
 sky130_fd_sc_hd__or3_1 _6726_ (.A(_2581_),
    .B(_2487_),
    .C(_2713_),
    .X(_2714_));
 sky130_fd_sc_hd__or2_1 _6727_ (.A(_2214_),
    .B(_2235_),
    .X(_2715_));
 sky130_fd_sc_hd__or3_1 _6728_ (.A(_2084_),
    .B(_2715_),
    .C(_2703_),
    .X(_2716_));
 sky130_fd_sc_hd__nand3b_1 _6729_ (.A_N(_2610_),
    .B(_2518_),
    .C(_2716_),
    .Y(_2717_));
 sky130_fd_sc_hd__or2_1 _6730_ (.A(_2233_),
    .B(_2703_),
    .X(_2718_));
 sky130_fd_sc_hd__o21bai_1 _6731_ (.A1(_2712_),
    .A2(_2718_),
    .B1_N(_2604_),
    .Y(_2719_));
 sky130_fd_sc_hd__nor2_1 _6732_ (.A(_2084_),
    .B(_2115_),
    .Y(_2720_));
 sky130_fd_sc_hd__a21o_1 _6733_ (.A1(_2612_),
    .A2(_2720_),
    .B1(_2613_),
    .X(_2721_));
 sky130_fd_sc_hd__a221o_1 _6734_ (.A1(_2301_),
    .A2(_2270_),
    .B1(_2184_),
    .B2(_2275_),
    .C1(_2721_),
    .X(_2722_));
 sky130_fd_sc_hd__or4_1 _6735_ (.A(_2714_),
    .B(_2717_),
    .C(_2719_),
    .D(_2722_),
    .X(_2723_));
 sky130_fd_sc_hd__nand2_1 _6736_ (.A(_2263_),
    .B(_2134_),
    .Y(_2724_));
 sky130_fd_sc_hd__a21o_1 _6737_ (.A1(_2218_),
    .A2(_2724_),
    .B1(_2597_),
    .X(_2725_));
 sky130_fd_sc_hd__or3_1 _6738_ (.A(_2639_),
    .B(_2285_),
    .C(_2653_),
    .X(_2726_));
 sky130_fd_sc_hd__nor2_1 _6739_ (.A(_2067_),
    .B(_2079_),
    .Y(_2727_));
 sky130_fd_sc_hd__a31o_1 _6740_ (.A1(_2727_),
    .A2(_2709_),
    .A3(_2720_),
    .B1(_2399_),
    .X(_2728_));
 sky130_fd_sc_hd__or4_1 _6741_ (.A(_2577_),
    .B(_2725_),
    .C(_2726_),
    .D(_2728_),
    .X(_2729_));
 sky130_fd_sc_hd__nor2_1 _6742_ (.A(_2233_),
    .B(_2703_),
    .Y(_2730_));
 sky130_fd_sc_hd__a311o_1 _6743_ (.A1(_2707_),
    .A2(_2118_),
    .A3(_2730_),
    .B1(_2512_),
    .C1(_2592_),
    .X(_2731_));
 sky130_fd_sc_hd__or3_1 _6744_ (.A(_2233_),
    .B(_2235_),
    .C(_2284_),
    .X(_2732_));
 sky130_fd_sc_hd__a21o_1 _6745_ (.A1(_2598_),
    .A2(_2732_),
    .B1(_2214_),
    .X(_2733_));
 sky130_fd_sc_hd__o21ai_1 _6746_ (.A1(_2715_),
    .A2(_2718_),
    .B1(_2733_),
    .Y(_2734_));
 sky130_fd_sc_hd__a21o_1 _6747_ (.A1(_2612_),
    .A2(_2730_),
    .B1(_2596_),
    .X(_2735_));
 sky130_fd_sc_hd__nor2_1 _6748_ (.A(_2132_),
    .B(_2108_),
    .Y(_2736_));
 sky130_fd_sc_hd__a21oi_1 _6749_ (.A1(_2225_),
    .A2(_2134_),
    .B1(_2120_),
    .Y(_2737_));
 sky130_fd_sc_hd__or4_1 _6750_ (.A(_2734_),
    .B(_2735_),
    .C(_2736_),
    .D(_2737_),
    .X(_2738_));
 sky130_fd_sc_hd__or4_1 _6751_ (.A(_2723_),
    .B(_2729_),
    .C(_2731_),
    .D(_2738_),
    .X(_2739_));
 sky130_fd_sc_hd__nor2_1 _6752_ (.A(_2711_),
    .B(_2739_),
    .Y(_2740_));
 sky130_fd_sc_hd__nor2_1 _6753_ (.A(_2702_),
    .B(_2740_),
    .Y(_2741_));
 sky130_fd_sc_hd__or4b_4 _6754_ (.A(_2098_),
    .B(_2111_),
    .C(_2365_),
    .D_N(_2372_),
    .X(_2742_));
 sky130_fd_sc_hd__a21oi_1 _6755_ (.A1(_2357_),
    .A2(_2387_),
    .B1(_2420_),
    .Y(_2743_));
 sky130_fd_sc_hd__o22a_1 _6756_ (.A1(_2198_),
    .A2(_2097_),
    .B1(_2357_),
    .B2(_2403_),
    .X(_2744_));
 sky130_fd_sc_hd__o221a_1 _6757_ (.A1(_2198_),
    .A2(_2316_),
    .B1(_2387_),
    .B2(_2403_),
    .C1(_2744_),
    .X(_2745_));
 sky130_fd_sc_hd__or4b_1 _6758_ (.A(_2322_),
    .B(_2670_),
    .C(_2743_),
    .D_N(_2745_),
    .X(_2746_));
 sky130_fd_sc_hd__or3_1 _6759_ (.A(_2329_),
    .B(_2439_),
    .C(_2673_),
    .X(_2747_));
 sky130_fd_sc_hd__a211o_1 _6760_ (.A1(_2364_),
    .A2(_2429_),
    .B1(_2665_),
    .C1(_2311_),
    .X(_2748_));
 sky130_fd_sc_hd__or3_1 _6761_ (.A(_2746_),
    .B(_2747_),
    .C(_2748_),
    .X(_2749_));
 sky130_fd_sc_hd__o211a_1 _6762_ (.A1(_2220_),
    .A2(_2338_),
    .B1(_2310_),
    .C1(_2360_),
    .X(_2750_));
 sky130_fd_sc_hd__or2_1 _6763_ (.A(_2679_),
    .B(_2750_),
    .X(_2751_));
 sky130_fd_sc_hd__nor2_1 _6764_ (.A(_2123_),
    .B(_2657_),
    .Y(_2752_));
 sky130_fd_sc_hd__or3_1 _6765_ (.A(_2397_),
    .B(_2535_),
    .C(_2752_),
    .X(_2753_));
 sky130_fd_sc_hd__nand2_1 _6766_ (.A(_2097_),
    .B(_2316_),
    .Y(_2754_));
 sky130_fd_sc_hd__a2bb2o_1 _6767_ (.A1_N(_2412_),
    .A2_N(_2509_),
    .B1(_2335_),
    .B2(_2754_),
    .X(_2755_));
 sky130_fd_sc_hd__inv_2 _6768_ (.A(_2754_),
    .Y(_2756_));
 sky130_fd_sc_hd__o21ba_1 _6769_ (.A1(_2249_),
    .A2(_2756_),
    .B1_N(_2413_),
    .X(_2757_));
 sky130_fd_sc_hd__or4b_1 _6770_ (.A(_2751_),
    .B(_2753_),
    .C(_2755_),
    .D_N(_2757_),
    .X(_2758_));
 sky130_fd_sc_hd__a311o_1 _6771_ (.A1(_2364_),
    .A2(_2493_),
    .A3(_2449_),
    .B1(_2667_),
    .C1(_2320_),
    .X(_2759_));
 sky130_fd_sc_hd__nor2_1 _6772_ (.A(_2412_),
    .B(_2471_),
    .Y(_2760_));
 sky130_fd_sc_hd__a31o_1 _6773_ (.A1(_2310_),
    .A2(_2754_),
    .A3(_2682_),
    .B1(_2760_),
    .X(_2761_));
 sky130_fd_sc_hd__a32o_1 _6774_ (.A1(_2220_),
    .A2(_2360_),
    .A3(_2381_),
    .B1(_2525_),
    .B2(_2364_),
    .X(_2762_));
 sky130_fd_sc_hd__or3_1 _6775_ (.A(_2097_),
    .B(_2460_),
    .C(_2681_),
    .X(_2763_));
 sky130_fd_sc_hd__a2bb2o_1 _6776_ (.A1_N(_2371_),
    .A2_N(_2763_),
    .B1(_2293_),
    .B2(_2624_),
    .X(_2764_));
 sky130_fd_sc_hd__or4_1 _6777_ (.A(_2663_),
    .B(_2761_),
    .C(_2762_),
    .D(_2764_),
    .X(_2765_));
 sky130_fd_sc_hd__or2_2 _6778_ (.A(_2124_),
    .B(_2619_),
    .X(_2766_));
 sky130_fd_sc_hd__or3_1 _6779_ (.A(_2097_),
    .B(_2382_),
    .C(_2684_),
    .X(_2767_));
 sky130_fd_sc_hd__o31a_1 _6780_ (.A1(_2357_),
    .A2(_2382_),
    .A3(_2391_),
    .B1(_2767_),
    .X(_2768_));
 sky130_fd_sc_hd__or4_1 _6781_ (.A(_2149_),
    .B(_2387_),
    .C(_2382_),
    .D(_2389_),
    .X(_2769_));
 sky130_fd_sc_hd__o211a_1 _6782_ (.A1(_2229_),
    .A2(_2316_),
    .B1(_2768_),
    .C1(_2769_),
    .X(_2770_));
 sky130_fd_sc_hd__or3b_1 _6783_ (.A(_2484_),
    .B(_2766_),
    .C_N(_2770_),
    .X(_2771_));
 sky130_fd_sc_hd__or4_1 _6784_ (.A(_2758_),
    .B(_2759_),
    .C(_2765_),
    .D(_2771_),
    .X(_2772_));
 sky130_fd_sc_hd__nor2_1 _6785_ (.A(_2749_),
    .B(_2772_),
    .Y(_2773_));
 sky130_fd_sc_hd__nor2_1 _6786_ (.A(_2742_),
    .B(_2773_),
    .Y(_2774_));
 sky130_fd_sc_hd__a21o_1 _6787_ (.A1(_2209_),
    .A2(_2123_),
    .B1(_2180_),
    .X(_2775_));
 sky130_fd_sc_hd__or3_2 _6788_ (.A(_2287_),
    .B(_2302_),
    .C(_2483_),
    .X(_2776_));
 sky130_fd_sc_hd__nand2_1 _6789_ (.A(_2775_),
    .B(_2776_),
    .Y(_2777_));
 sky130_fd_sc_hd__and3_1 _6790_ (.A(_2209_),
    .B(_2191_),
    .C(_2553_),
    .X(_2778_));
 sky130_fd_sc_hd__clkbuf_4 _6791_ (.A(_2778_),
    .X(_2779_));
 sky130_fd_sc_hd__nor2_1 _6792_ (.A(_2552_),
    .B(_2779_),
    .Y(_2780_));
 sky130_fd_sc_hd__nor2_1 _6793_ (.A(_2284_),
    .B(_2536_),
    .Y(_2781_));
 sky130_fd_sc_hd__nor2_1 _6794_ (.A(_2105_),
    .B(_2622_),
    .Y(_2782_));
 sky130_fd_sc_hd__and3_1 _6795_ (.A(net395),
    .B(_2126_),
    .C(_2360_),
    .X(_2783_));
 sky130_fd_sc_hd__a211o_1 _6796_ (.A1(_2782_),
    .A2(_2303_),
    .B1(_2548_),
    .C1(_2783_),
    .X(_2784_));
 sky130_fd_sc_hd__a32o_1 _6797_ (.A1(_2301_),
    .A2(_2186_),
    .A3(net394),
    .B1(_2624_),
    .B2(_2095_),
    .X(_2785_));
 sky130_fd_sc_hd__or4_1 _6798_ (.A(_2285_),
    .B(_2781_),
    .C(_2784_),
    .D(_2785_),
    .X(_2786_));
 sky130_fd_sc_hd__nor2_1 _6799_ (.A(_2198_),
    .B(_2779_),
    .Y(_2787_));
 sky130_fd_sc_hd__nor2_1 _6800_ (.A(_2189_),
    .B(_2779_),
    .Y(_2788_));
 sky130_fd_sc_hd__a21oi_2 _6801_ (.A1(_2225_),
    .A2(_2295_),
    .B1(_2120_),
    .Y(_2789_));
 sky130_fd_sc_hd__nor2_1 _6802_ (.A(_2253_),
    .B(_2779_),
    .Y(_2790_));
 sky130_fd_sc_hd__a41o_1 _6803_ (.A1(_2223_),
    .A2(_2212_),
    .A3(_2203_),
    .A4(_2249_),
    .B1(_2779_),
    .X(_2791_));
 sky130_fd_sc_hd__or3b_1 _6804_ (.A(_2789_),
    .B(_2790_),
    .C_N(_2791_),
    .X(_2792_));
 sky130_fd_sc_hd__or3_1 _6805_ (.A(_2787_),
    .B(_2788_),
    .C(_2792_),
    .X(_2793_));
 sky130_fd_sc_hd__or4_1 _6806_ (.A(_2766_),
    .B(_2780_),
    .C(_2786_),
    .D(_2793_),
    .X(_2794_));
 sky130_fd_sc_hd__or3b_1 _6807_ (.A(_2777_),
    .B(_2794_),
    .C_N(_2662_),
    .X(_2795_));
 sky130_fd_sc_hd__o31a_1 _6808_ (.A1(_2104_),
    .A2(_2091_),
    .A3(_2094_),
    .B1(_2367_),
    .X(_2796_));
 sky130_fd_sc_hd__and4bb_1 _6809_ (.A_N(_2111_),
    .B_N(_2285_),
    .C(_2647_),
    .D(_2476_),
    .X(_2797_));
 sky130_fd_sc_hd__or3_1 _6810_ (.A(_2397_),
    .B(_2481_),
    .C(_2296_),
    .X(_2798_));
 sky130_fd_sc_hd__and3_1 _6811_ (.A(_2126_),
    .B(_2360_),
    .C(_2361_),
    .X(_2799_));
 sky130_fd_sc_hd__nand2_2 _6812_ (.A(_2363_),
    .B(_2490_),
    .Y(_2800_));
 sky130_fd_sc_hd__a21o_1 _6813_ (.A1(_2276_),
    .A2(_2629_),
    .B1(_2508_),
    .X(_2801_));
 sky130_fd_sc_hd__o221a_1 _6814_ (.A1(_2151_),
    .A2(_2479_),
    .B1(_2494_),
    .B2(_2500_),
    .C1(_2649_),
    .X(_2802_));
 sky130_fd_sc_hd__nor3_1 _6815_ (.A(_2110_),
    .B(_2363_),
    .C(_2428_),
    .Y(_2803_));
 sky130_fd_sc_hd__a21oi_1 _6816_ (.A1(_2075_),
    .A2(_2624_),
    .B1(_2803_),
    .Y(_2804_));
 sky130_fd_sc_hd__nand2_1 _6817_ (.A(_2802_),
    .B(_2804_),
    .Y(_2805_));
 sky130_fd_sc_hd__or3b_1 _6818_ (.A(_2388_),
    .B(_2414_),
    .C_N(_2100_),
    .X(_2806_));
 sky130_fd_sc_hd__a21boi_1 _6819_ (.A1(_2450_),
    .A2(_2806_),
    .B1_N(_2800_),
    .Y(_2807_));
 sky130_fd_sc_hd__nor2_1 _6820_ (.A(_2153_),
    .B(_2357_),
    .Y(_2808_));
 sky130_fd_sc_hd__a211o_1 _6821_ (.A1(_2429_),
    .A2(_2800_),
    .B1(_2807_),
    .C1(_2808_),
    .X(_2809_));
 sky130_fd_sc_hd__or2_1 _6822_ (.A(_2546_),
    .B(_2641_),
    .X(_2810_));
 sky130_fd_sc_hd__a2111o_1 _6823_ (.A1(_2800_),
    .A2(_2801_),
    .B1(_2805_),
    .C1(_2809_),
    .D1(_2810_),
    .X(_2811_));
 sky130_fd_sc_hd__or4_1 _6824_ (.A(_2619_),
    .B(_2798_),
    .C(_2799_),
    .D(_2811_),
    .X(_2812_));
 sky130_fd_sc_hd__a21o_1 _6825_ (.A1(_2797_),
    .A2(_2812_),
    .B1(_2533_),
    .X(_2813_));
 sky130_fd_sc_hd__a31o_1 _6826_ (.A1(_2647_),
    .A2(_2795_),
    .A3(_2796_),
    .B1(_2813_),
    .X(_2814_));
 sky130_fd_sc_hd__o32a_1 _6827_ (.A1(_2741_),
    .A2(_2774_),
    .A3(_2814_),
    .B1(_1949_),
    .B2(net1557),
    .X(_0379_));
 sky130_fd_sc_hd__or3b_2 _6828_ (.A(_2095_),
    .B(_2113_),
    .C_N(_2138_),
    .X(_2815_));
 sky130_fd_sc_hd__o211a_1 _6829_ (.A1(_2189_),
    .A2(_2815_),
    .B1(_2447_),
    .C1(_2452_),
    .X(_2816_));
 sky130_fd_sc_hd__inv_2 _6830_ (.A(_2420_),
    .Y(_2817_));
 sky130_fd_sc_hd__a2111oi_1 _6831_ (.A1(_2411_),
    .A2(_2817_),
    .B1(_2456_),
    .C1(_2670_),
    .D1(_2322_),
    .Y(_2818_));
 sky130_fd_sc_hd__o221a_1 _6832_ (.A1(_2128_),
    .A2(_2203_),
    .B1(_2417_),
    .B2(_2420_),
    .C1(_2451_),
    .X(_2819_));
 sky130_fd_sc_hd__o211a_1 _6833_ (.A1(_2203_),
    .A2(_2123_),
    .B1(_2818_),
    .C1(_2819_),
    .X(_2820_));
 sky130_fd_sc_hd__and3_1 _6834_ (.A(_2745_),
    .B(_2816_),
    .C(_2820_),
    .X(_2821_));
 sky130_fd_sc_hd__or2_1 _6835_ (.A(_2661_),
    .B(_2663_),
    .X(_2822_));
 sky130_fd_sc_hd__or3_1 _6836_ (.A(_2659_),
    .B(_2822_),
    .C(_2762_),
    .X(_2823_));
 sky130_fd_sc_hd__a311o_1 _6837_ (.A1(_2554_),
    .A2(_2310_),
    .A3(_2682_),
    .B1(_2683_),
    .C1(_2436_),
    .X(_2824_));
 sky130_fd_sc_hd__nor2_1 _6838_ (.A(_2751_),
    .B(_2824_),
    .Y(_2825_));
 sky130_fd_sc_hd__nor2_1 _6839_ (.A(_2122_),
    .B(_2306_),
    .Y(_2826_));
 sky130_fd_sc_hd__o22a_1 _6840_ (.A1(_2128_),
    .A2(_2638_),
    .B1(_2826_),
    .B2(_2462_),
    .X(_2827_));
 sky130_fd_sc_hd__and4bb_1 _6841_ (.A_N(_2577_),
    .B_N(_2753_),
    .C(_2825_),
    .D(_2827_),
    .X(_2828_));
 sky130_fd_sc_hd__nor2_1 _6842_ (.A(_2327_),
    .B(_2432_),
    .Y(_2829_));
 sky130_fd_sc_hd__and4bb_1 _6843_ (.A_N(_2328_),
    .B_N(_2747_),
    .C(_2416_),
    .D(_2829_),
    .X(_2830_));
 sky130_fd_sc_hd__nor2_1 _6844_ (.A(_2441_),
    .B(_2674_),
    .Y(_2831_));
 sky130_fd_sc_hd__o211a_1 _6845_ (.A1(_2223_),
    .A2(_2815_),
    .B1(_2770_),
    .C1(_2831_),
    .X(_2832_));
 sky130_fd_sc_hd__and4b_1 _6846_ (.A_N(_2823_),
    .B(_2828_),
    .C(_2830_),
    .D(_2832_),
    .X(_2833_));
 sky130_fd_sc_hd__a21oi_1 _6847_ (.A1(_2821_),
    .A2(_2833_),
    .B1(_2742_),
    .Y(_2834_));
 sky130_fd_sc_hd__o21a_1 _6848_ (.A1(_2215_),
    .A2(_2181_),
    .B1(_2184_),
    .X(_2835_));
 sky130_fd_sc_hd__a221o_1 _6849_ (.A1(_2301_),
    .A2(_2270_),
    .B1(_2184_),
    .B2(_2275_),
    .C1(_2721_),
    .X(_2836_));
 sky130_fd_sc_hd__nor3_1 _6850_ (.A(_2171_),
    .B(_2173_),
    .C(_2479_),
    .Y(_2837_));
 sky130_fd_sc_hd__or4_1 _6851_ (.A(_2250_),
    .B(_2837_),
    .C(_2588_),
    .D(_2719_),
    .X(_2838_));
 sky130_fd_sc_hd__nor2_1 _6852_ (.A(_2585_),
    .B(_2479_),
    .Y(_2839_));
 sky130_fd_sc_hd__or4_1 _6853_ (.A(_2259_),
    .B(_2839_),
    .C(_2587_),
    .D(_2706_),
    .X(_2840_));
 sky130_fd_sc_hd__or4_1 _6854_ (.A(_2835_),
    .B(_2836_),
    .C(_2838_),
    .D(_2840_),
    .X(_2841_));
 sky130_fd_sc_hd__o32a_1 _6855_ (.A1(_2171_),
    .A2(_2388_),
    .A3(_2479_),
    .B1(_2147_),
    .B2(_2295_),
    .X(_2842_));
 sky130_fd_sc_hd__or3b_1 _6856_ (.A(_2221_),
    .B(_2725_),
    .C_N(_2842_),
    .X(_2843_));
 sky130_fd_sc_hd__or4_1 _6857_ (.A(_2228_),
    .B(_2230_),
    .C(_2510_),
    .D(_2735_),
    .X(_2844_));
 sky130_fd_sc_hd__nor2_1 _6858_ (.A(_2140_),
    .B(_2120_),
    .Y(_2845_));
 sky130_fd_sc_hd__or4b_2 _6859_ (.A(_2845_),
    .B(_2469_),
    .C(_2736_),
    .D_N(_2617_),
    .X(_2846_));
 sky130_fd_sc_hd__and2b_1 _6860_ (.A_N(_2132_),
    .B(_2724_),
    .X(_2847_));
 sky130_fd_sc_hd__or4_1 _6861_ (.A(_2737_),
    .B(_2844_),
    .C(_2846_),
    .D(_2847_),
    .X(_2848_));
 sky130_fd_sc_hd__nor2_1 _6862_ (.A(_2428_),
    .B(_2479_),
    .Y(_2849_));
 sky130_fd_sc_hd__or4_1 _6863_ (.A(_2266_),
    .B(_2849_),
    .C(_2582_),
    .D(_2714_),
    .X(_2850_));
 sky130_fd_sc_hd__or3_1 _6864_ (.A(_2843_),
    .B(_2848_),
    .C(_2850_),
    .X(_2851_));
 sky130_fd_sc_hd__or2_1 _6865_ (.A(_2575_),
    .B(_2702_),
    .X(_2852_));
 sky130_fd_sc_hd__o21ba_1 _6866_ (.A1(_2841_),
    .A2(_2851_),
    .B1_N(_2852_),
    .X(_2853_));
 sky130_fd_sc_hd__or4bb_2 _6867_ (.A(_2285_),
    .B(_2766_),
    .C_N(_2796_),
    .D_N(_2647_),
    .X(_2854_));
 sky130_fd_sc_hd__inv_2 _6868_ (.A(_2854_),
    .Y(_2855_));
 sky130_fd_sc_hd__or4_1 _6869_ (.A(_2266_),
    .B(_2610_),
    .C(_2313_),
    .D(_2317_),
    .X(_2856_));
 sky130_fd_sc_hd__or2_1 _6870_ (.A(_2787_),
    .B(_2856_),
    .X(_2857_));
 sky130_fd_sc_hd__nor2_1 _6871_ (.A(_2284_),
    .B(_2203_),
    .Y(_2858_));
 sky130_fd_sc_hd__or4_1 _6872_ (.A(_2858_),
    .B(_2323_),
    .C(_2544_),
    .D(_2790_),
    .X(_2859_));
 sky130_fd_sc_hd__nand2_1 _6873_ (.A(_2225_),
    .B(_2284_),
    .Y(_2860_));
 sky130_fd_sc_hd__nand2_1 _6874_ (.A(_2316_),
    .B(_2779_),
    .Y(_2861_));
 sky130_fd_sc_hd__a22o_1 _6875_ (.A1(_2335_),
    .A2(_2860_),
    .B1(_2861_),
    .B2(_2545_),
    .X(_2862_));
 sky130_fd_sc_hd__nor2_1 _6876_ (.A(_2225_),
    .B(_2132_),
    .Y(_2863_));
 sky130_fd_sc_hd__or4_1 _6877_ (.A(_2355_),
    .B(_2290_),
    .C(_2484_),
    .D(_2781_),
    .X(_2864_));
 sky130_fd_sc_hd__or3_1 _6878_ (.A(_2789_),
    .B(_2863_),
    .C(_2864_),
    .X(_2865_));
 sky130_fd_sc_hd__a41o_1 _6879_ (.A1(_2217_),
    .A2(_2500_),
    .A3(_2497_),
    .A4(_2599_),
    .B1(_2194_),
    .X(_2866_));
 sky130_fd_sc_hd__or4b_1 _6880_ (.A(_2784_),
    .B(_2862_),
    .C(_2865_),
    .D_N(_2866_),
    .X(_2867_));
 sky130_fd_sc_hd__nor2_1 _6881_ (.A(_2212_),
    .B(_2779_),
    .Y(_2868_));
 sky130_fd_sc_hd__or4_1 _6882_ (.A(_2589_),
    .B(_2327_),
    .C(_2559_),
    .D(_2868_),
    .X(_2869_));
 sky130_fd_sc_hd__o211ai_2 _6883_ (.A1(_2301_),
    .A2(_2205_),
    .B1(_2303_),
    .C1(_2299_),
    .Y(_2870_));
 sky130_fd_sc_hd__o211a_1 _6884_ (.A1(_2180_),
    .A2(_2555_),
    .B1(_2776_),
    .C1(_2662_),
    .X(_2871_));
 sky130_fd_sc_hd__nand3b_1 _6885_ (.A_N(_2869_),
    .B(_2870_),
    .C(_2871_),
    .Y(_2872_));
 sky130_fd_sc_hd__or4_1 _6886_ (.A(_2857_),
    .B(_2859_),
    .C(_2867_),
    .D(_2872_),
    .X(_2873_));
 sky130_fd_sc_hd__nor2_1 _6887_ (.A(_2389_),
    .B(_2414_),
    .Y(_2874_));
 sky130_fd_sc_hd__a31o_1 _6888_ (.A1(_2149_),
    .A2(_2411_),
    .A3(_2874_),
    .B1(_2436_),
    .X(_2875_));
 sky130_fd_sc_hd__a211o_1 _6889_ (.A1(_2493_),
    .A2(_2498_),
    .B1(_2810_),
    .C1(_2875_),
    .X(_2876_));
 sky130_fd_sc_hd__a21o_1 _6890_ (.A1(_2538_),
    .A2(_2357_),
    .B1(_2434_),
    .X(_2877_));
 sky130_fd_sc_hd__or2_1 _6891_ (.A(_2075_),
    .B(_2094_),
    .X(_2878_));
 sky130_fd_sc_hd__a31o_1 _6892_ (.A1(_2878_),
    .A2(_2387_),
    .A3(_2490_),
    .B1(_2391_),
    .X(_2879_));
 sky130_fd_sc_hd__a21oi_1 _6893_ (.A1(_2877_),
    .A2(_2879_),
    .B1(_2414_),
    .Y(_2880_));
 sky130_fd_sc_hd__nor2_1 _6894_ (.A(_2538_),
    .B(_2153_),
    .Y(_2881_));
 sky130_fd_sc_hd__nand2_2 _6895_ (.A(_2140_),
    .B(_2357_),
    .Y(_2882_));
 sky130_fd_sc_hd__a221o_1 _6896_ (.A1(_2504_),
    .A2(_2800_),
    .B1(_2882_),
    .B2(_2429_),
    .C1(_2633_),
    .X(_2883_));
 sky130_fd_sc_hd__nor2_1 _6897_ (.A(_2215_),
    .B(_2411_),
    .Y(_2884_));
 sky130_fd_sc_hd__nor2_1 _6898_ (.A(_2450_),
    .B(_2884_),
    .Y(_2885_));
 sky130_fd_sc_hd__a211o_1 _6899_ (.A1(_2817_),
    .A2(_2800_),
    .B1(_2885_),
    .C1(_2625_),
    .X(_2886_));
 sky130_fd_sc_hd__nor2_1 _6900_ (.A(_2409_),
    .B(_2884_),
    .Y(_2887_));
 sky130_fd_sc_hd__a211o_1 _6901_ (.A1(_2508_),
    .A2(_2800_),
    .B1(_2887_),
    .C1(_2631_),
    .X(_2888_));
 sky130_fd_sc_hd__or4_1 _6902_ (.A(_2881_),
    .B(_2883_),
    .C(_2886_),
    .D(_2888_),
    .X(_2889_));
 sky130_fd_sc_hd__a311o_1 _6903_ (.A1(_2360_),
    .A2(_2361_),
    .A3(_2338_),
    .B1(_2640_),
    .C1(_2808_),
    .X(_2890_));
 sky130_fd_sc_hd__and4b_1 _6904_ (.A_N(_2890_),
    .B(_2644_),
    .C(_2514_),
    .D(_2802_),
    .X(_2891_));
 sky130_fd_sc_hd__or3b_1 _6905_ (.A(_2880_),
    .B(_2889_),
    .C_N(_2891_),
    .X(_2892_));
 sky130_fd_sc_hd__or3_1 _6906_ (.A(_2225_),
    .B(_2101_),
    .C(_2110_),
    .X(_2893_));
 sky130_fd_sc_hd__and3b_1 _6907_ (.A_N(_2619_),
    .B(_2797_),
    .C(_2893_),
    .X(_2894_));
 sky130_fd_sc_hd__and2_1 _6908_ (.A(_1949_),
    .B(_2894_),
    .X(_2895_));
 sky130_fd_sc_hd__o31a_1 _6909_ (.A1(_2798_),
    .A2(_2876_),
    .A3(_2892_),
    .B1(_2895_),
    .X(_2896_));
 sky130_fd_sc_hd__a221o_1 _6910_ (.A1(\wbbd_addr[3] ),
    .A2(_2533_),
    .B1(_2855_),
    .B2(_2873_),
    .C1(_2896_),
    .X(_2897_));
 sky130_fd_sc_hd__or3_1 _6911_ (.A(_2834_),
    .B(_2853_),
    .C(_2897_),
    .X(_2898_));
 sky130_fd_sc_hd__clkbuf_1 _6912_ (.A(_2898_),
    .X(_0380_));
 sky130_fd_sc_hd__a2111o_1 _6913_ (.A1(_2385_),
    .A2(_2435_),
    .B1(_2513_),
    .C1(_2880_),
    .D1(_2408_),
    .X(_2899_));
 sky130_fd_sc_hd__a32o_1 _6914_ (.A1(_2493_),
    .A2(_2449_),
    .A3(_2800_),
    .B1(_2882_),
    .B2(_2504_),
    .X(_2900_));
 sky130_fd_sc_hd__or3_1 _6915_ (.A(_2643_),
    .B(_2886_),
    .C(_2900_),
    .X(_2901_));
 sky130_fd_sc_hd__a21o_1 _6916_ (.A1(_2538_),
    .A2(_2363_),
    .B1(_2153_),
    .X(_2902_));
 sky130_fd_sc_hd__and4b_1 _6917_ (.A_N(_2455_),
    .B(_2516_),
    .C(_2804_),
    .D(_2902_),
    .X(_2903_));
 sky130_fd_sc_hd__and3_1 _6918_ (.A(_2644_),
    .B(_2802_),
    .C(_2903_),
    .X(_2904_));
 sky130_fd_sc_hd__or3b_1 _6919_ (.A(_2899_),
    .B(_2901_),
    .C_N(_2904_),
    .X(_2905_));
 sky130_fd_sc_hd__a22o_1 _6920_ (.A1(\wbbd_addr[4] ),
    .A2(_2533_),
    .B1(_2895_),
    .B2(_2905_),
    .X(_2906_));
 sky130_fd_sc_hd__o22ai_1 _6921_ (.A1(_2198_),
    .A2(_2815_),
    .B1(_2431_),
    .B2(_2585_),
    .Y(_2907_));
 sky130_fd_sc_hd__nor3_1 _6922_ (.A(_2404_),
    .B(_2759_),
    .C(_2907_),
    .Y(_2908_));
 sky130_fd_sc_hd__nand2_1 _6923_ (.A(_2820_),
    .B(_2908_),
    .Y(_2909_));
 sky130_fd_sc_hd__or4_1 _6924_ (.A(_2455_),
    .B(_2658_),
    .C(_2577_),
    .D(_2764_),
    .X(_2910_));
 sky130_fd_sc_hd__or4_1 _6925_ (.A(_2481_),
    .B(_2383_),
    .C(_2823_),
    .D(_2910_),
    .X(_2911_));
 sky130_fd_sc_hd__or2_1 _6926_ (.A(_2431_),
    .B(_2434_),
    .X(_2912_));
 sky130_fd_sc_hd__o22a_1 _6927_ (.A1(_2212_),
    .A2(_2123_),
    .B1(_2295_),
    .B2(_2407_),
    .X(_2913_));
 sky130_fd_sc_hd__and3b_1 _6928_ (.A_N(_2331_),
    .B(_2912_),
    .C(_2913_),
    .X(_2914_));
 sky130_fd_sc_hd__nand3b_1 _6929_ (.A_N(_2755_),
    .B(_2832_),
    .C(_2914_),
    .Y(_2915_));
 sky130_fd_sc_hd__a211o_1 _6930_ (.A1(_2102_),
    .A2(_2463_),
    .B1(_2654_),
    .C1(_2766_),
    .X(_2916_));
 sky130_fd_sc_hd__or3b_1 _6931_ (.A(_2742_),
    .B(_2752_),
    .C_N(_2893_),
    .X(_2917_));
 sky130_fd_sc_hd__nor2_1 _6932_ (.A(_2916_),
    .B(_2917_),
    .Y(_2918_));
 sky130_fd_sc_hd__o31a_1 _6933_ (.A1(_2909_),
    .A2(_2911_),
    .A3(_2915_),
    .B1(_2918_),
    .X(_2919_));
 sky130_fd_sc_hd__o22a_1 _6934_ (.A1(_2284_),
    .A2(_2198_),
    .B1(_2203_),
    .B2(_2779_),
    .X(_2920_));
 sky130_fd_sc_hd__or4b_2 _6935_ (.A(_2319_),
    .B(_2543_),
    .C(_2859_),
    .D_N(_2920_),
    .X(_2921_));
 sky130_fd_sc_hd__o21ai_1 _6936_ (.A1(_2223_),
    .A2(_2779_),
    .B1(_2245_),
    .Y(_2922_));
 sky130_fd_sc_hd__or4_1 _6937_ (.A(_2331_),
    .B(_2560_),
    .C(_2862_),
    .D(_2922_),
    .X(_2923_));
 sky130_fd_sc_hd__or4_1 _6938_ (.A(_2537_),
    .B(_2627_),
    .C(_2863_),
    .D(_2923_),
    .X(_2924_));
 sky130_fd_sc_hd__nand4_1 _6939_ (.A(_2662_),
    .B(_2870_),
    .C(_2775_),
    .D(_2776_),
    .Y(_2925_));
 sky130_fd_sc_hd__a311o_1 _6940_ (.A1(net395),
    .A2(_2205_),
    .A3(_2299_),
    .B1(_2785_),
    .C1(_2925_),
    .X(_2926_));
 sky130_fd_sc_hd__or3_1 _6941_ (.A(_2921_),
    .B(_2924_),
    .C(_2926_),
    .X(_2927_));
 sky130_fd_sc_hd__and2_1 _6942_ (.A(_2855_),
    .B(_2927_),
    .X(_2928_));
 sky130_fd_sc_hd__o31a_1 _6943_ (.A1(_2173_),
    .A2(_2100_),
    .A3(_2479_),
    .B1(_2264_),
    .X(_2929_));
 sky130_fd_sc_hd__or4b_2 _6944_ (.A(_2584_),
    .B(_2708_),
    .C(_2840_),
    .D_N(_2929_),
    .X(_2930_));
 sky130_fd_sc_hd__o22a_1 _6945_ (.A1(_2212_),
    .A2(_2263_),
    .B1(_2108_),
    .B2(_2407_),
    .X(_2931_));
 sky130_fd_sc_hd__or4b_1 _6946_ (.A(_2591_),
    .B(_2731_),
    .C(_2844_),
    .D_N(_2931_),
    .X(_2932_));
 sky130_fd_sc_hd__a31o_1 _6947_ (.A1(_2263_),
    .A2(_2115_),
    .A3(_2134_),
    .B1(_2132_),
    .X(_2933_));
 sky130_fd_sc_hd__or3b_1 _6948_ (.A(_2397_),
    .B(_2296_),
    .C_N(_2933_),
    .X(_2934_));
 sky130_fd_sc_hd__a311o_1 _6949_ (.A1(_2727_),
    .A2(_2709_),
    .A3(_2720_),
    .B1(_2577_),
    .C1(_2399_),
    .X(_2935_));
 sky130_fd_sc_hd__or4_1 _6950_ (.A(_2148_),
    .B(_2835_),
    .C(_2836_),
    .D(_2935_),
    .X(_2936_));
 sky130_fd_sc_hd__or4_1 _6951_ (.A(_2930_),
    .B(_2932_),
    .C(_2934_),
    .D(_2936_),
    .X(_2937_));
 sky130_fd_sc_hd__or4b_1 _6952_ (.A(_2653_),
    .B(_2846_),
    .C(_2852_),
    .D_N(_2937_),
    .X(_2938_));
 sky130_fd_sc_hd__or4b_1 _6953_ (.A(_2906_),
    .B(_2919_),
    .C(_2928_),
    .D_N(_2938_),
    .X(_2939_));
 sky130_fd_sc_hd__clkbuf_1 _6954_ (.A(_2939_),
    .X(_0381_));
 sky130_fd_sc_hd__or4_1 _6955_ (.A(_2355_),
    .B(_2290_),
    .C(_2484_),
    .D(_2781_),
    .X(_2940_));
 sky130_fd_sc_hd__or3_1 _6956_ (.A(_2537_),
    .B(_2627_),
    .C(_2863_),
    .X(_2941_));
 sky130_fd_sc_hd__or3_1 _6957_ (.A(_2789_),
    .B(_2940_),
    .C(_2941_),
    .X(_2942_));
 sky130_fd_sc_hd__nor3_1 _6958_ (.A(_2854_),
    .B(_2926_),
    .C(_2942_),
    .Y(_2943_));
 sky130_fd_sc_hd__or4_1 _6959_ (.A(_2613_),
    .B(_2312_),
    .C(_2542_),
    .D(_2788_),
    .X(_2944_));
 sky130_fd_sc_hd__or3b_1 _6960_ (.A(_2549_),
    .B(_2783_),
    .C_N(_2866_),
    .X(_2945_));
 sky130_fd_sc_hd__a221o_1 _6961_ (.A1(_2545_),
    .A2(_2860_),
    .B1(_2861_),
    .B2(_2551_),
    .C1(_2945_),
    .X(_2946_));
 sky130_fd_sc_hd__or4_1 _6962_ (.A(_2857_),
    .B(_2921_),
    .C(_2944_),
    .D(_2946_),
    .X(_2947_));
 sky130_fd_sc_hd__a21oi_1 _6963_ (.A1(_2225_),
    .A2(_2134_),
    .B1(_2120_),
    .Y(_2948_));
 sky130_fd_sc_hd__or4_1 _6964_ (.A(_2653_),
    .B(_2948_),
    .C(_2846_),
    .D(_2934_),
    .X(_2949_));
 sky130_fd_sc_hd__nor3_1 _6965_ (.A(_2852_),
    .B(_2936_),
    .C(_2949_),
    .Y(_2950_));
 sky130_fd_sc_hd__or4_1 _6966_ (.A(_2541_),
    .B(_2480_),
    .C(_2580_),
    .D(_2717_),
    .X(_2951_));
 sky130_fd_sc_hd__nor3_1 _6967_ (.A(_2214_),
    .B(_2391_),
    .C(_2490_),
    .Y(_2952_));
 sky130_fd_sc_hd__o32a_1 _6968_ (.A1(_2233_),
    .A2(_2715_),
    .A3(_2191_),
    .B1(_2263_),
    .B2(_2229_),
    .X(_2953_));
 sky130_fd_sc_hd__or4b_1 _6969_ (.A(_2734_),
    .B(_2952_),
    .C(_2843_),
    .D_N(_2953_),
    .X(_2954_));
 sky130_fd_sc_hd__or4_1 _6970_ (.A(_2850_),
    .B(_2930_),
    .C(_2951_),
    .D(_2954_),
    .X(_2955_));
 sky130_fd_sc_hd__a221o_1 _6971_ (.A1(_2429_),
    .A2(_2800_),
    .B1(_2882_),
    .B2(_2525_),
    .C1(_2637_),
    .X(_2956_));
 sky130_fd_sc_hd__or3_1 _6972_ (.A(_2883_),
    .B(_2901_),
    .C(_2956_),
    .X(_2957_));
 sky130_fd_sc_hd__or3_1 _6973_ (.A(_2149_),
    .B(_2338_),
    .C(_2882_),
    .X(_2958_));
 sky130_fd_sc_hd__o211ai_1 _6974_ (.A1(_2075_),
    .A2(_2102_),
    .B1(_2149_),
    .C1(_2134_),
    .Y(_2959_));
 sky130_fd_sc_hd__a31o_1 _6975_ (.A1(_2874_),
    .A2(_2958_),
    .A3(_2959_),
    .B1(_2876_),
    .X(_2960_));
 sky130_fd_sc_hd__or4_1 _6976_ (.A(_2533_),
    .B(_2624_),
    .C(_2455_),
    .D(_2803_),
    .X(_2961_));
 sky130_fd_sc_hd__nor3_1 _6977_ (.A(_2627_),
    .B(_2628_),
    .C(_2961_),
    .Y(_2962_));
 sky130_fd_sc_hd__and4_1 _6978_ (.A(_2477_),
    .B(_2894_),
    .C(_2891_),
    .D(_2962_),
    .X(_2963_));
 sky130_fd_sc_hd__o21a_1 _6979_ (.A1(_2957_),
    .A2(_2960_),
    .B1(_2963_),
    .X(_2964_));
 sky130_fd_sc_hd__a221o_1 _6980_ (.A1(\wbbd_addr[5] ),
    .A2(_2533_),
    .B1(_2950_),
    .B2(_2955_),
    .C1(_2964_),
    .X(_2965_));
 sky130_fd_sc_hd__o221a_1 _6981_ (.A1(_2180_),
    .A2(_2815_),
    .B1(_2428_),
    .B2(_2431_),
    .C1(_2443_),
    .X(_2966_));
 sky130_fd_sc_hd__and4b_1 _6982_ (.A_N(_2748_),
    .B(_2821_),
    .C(_2908_),
    .D(_2966_),
    .X(_2967_));
 sky130_fd_sc_hd__inv_2 _6983_ (.A(_2761_),
    .Y(_2968_));
 sky130_fd_sc_hd__o32a_1 _6984_ (.A1(_2123_),
    .A2(_2382_),
    .A3(_2684_),
    .B1(_2440_),
    .B2(_2391_),
    .X(_2969_));
 sky130_fd_sc_hd__o211a_1 _6985_ (.A1(_2417_),
    .A2(_2471_),
    .B1(_2968_),
    .C1(_2969_),
    .X(_2970_));
 sky130_fd_sc_hd__o311a_1 _6986_ (.A1(_2125_),
    .A2(_2095_),
    .A3(_2229_),
    .B1(_2825_),
    .C1(_2970_),
    .X(_2971_));
 sky130_fd_sc_hd__or4_1 _6987_ (.A(_2384_),
    .B(_2535_),
    .C(_2627_),
    .D(_2762_),
    .X(_2972_));
 sky130_fd_sc_hd__or3_1 _6988_ (.A(_2822_),
    .B(_2910_),
    .C(_2972_),
    .X(_2973_));
 sky130_fd_sc_hd__or3_1 _6989_ (.A(_2916_),
    .B(_2917_),
    .C(_2973_),
    .X(_2974_));
 sky130_fd_sc_hd__a21oi_1 _6990_ (.A1(_2967_),
    .A2(_2971_),
    .B1(_2974_),
    .Y(_2975_));
 sky130_fd_sc_hd__a211o_1 _6991_ (.A1(_2943_),
    .A2(_2947_),
    .B1(_2965_),
    .C1(_2975_),
    .X(_0382_));
 sky130_fd_sc_hd__o21ai_1 _6992_ (.A1(_2420_),
    .A2(_2490_),
    .B1(_2256_),
    .Y(_2976_));
 sky130_fd_sc_hd__or4_1 _6993_ (.A(_2255_),
    .B(_2710_),
    .C(_2838_),
    .D(_2976_),
    .X(_2977_));
 sky130_fd_sc_hd__nor3_1 _6994_ (.A(_2850_),
    .B(_2930_),
    .C(_2951_),
    .Y(_2978_));
 sky130_fd_sc_hd__o311a_1 _6995_ (.A1(_2932_),
    .A2(_2954_),
    .A3(_2977_),
    .B1(_2950_),
    .C1(_2978_),
    .X(_2979_));
 sky130_fd_sc_hd__a32o_1 _6996_ (.A1(_2174_),
    .A2(_2493_),
    .A3(_2800_),
    .B1(_2882_),
    .B2(_2817_),
    .X(_2980_));
 sky130_fd_sc_hd__or4_1 _6997_ (.A(_2632_),
    .B(_2888_),
    .C(_2899_),
    .D(_2980_),
    .X(_2981_));
 sky130_fd_sc_hd__or2_1 _6998_ (.A(_2960_),
    .B(_2981_),
    .X(_2982_));
 sky130_fd_sc_hd__a22o_1 _6999_ (.A1(\wbbd_addr[6] ),
    .A2(_2533_),
    .B1(_2963_),
    .B2(_2982_),
    .X(_2983_));
 sky130_fd_sc_hd__nor3_1 _7000_ (.A(_2857_),
    .B(_2921_),
    .C(_2944_),
    .Y(_2984_));
 sky130_fd_sc_hd__nor2_1 _7001_ (.A(_2249_),
    .B(_2779_),
    .Y(_2985_));
 sky130_fd_sc_hd__or4_1 _7002_ (.A(_2254_),
    .B(_2324_),
    .C(_2562_),
    .D(_2985_),
    .X(_2986_));
 sky130_fd_sc_hd__or4_1 _7003_ (.A(_2869_),
    .B(_2923_),
    .C(_2946_),
    .D(_2986_),
    .X(_2987_));
 sky130_fd_sc_hd__and3_1 _7004_ (.A(_2943_),
    .B(_2984_),
    .C(_2987_),
    .X(_2988_));
 sky130_fd_sc_hd__a211oi_1 _7005_ (.A1(_2321_),
    .A2(_2554_),
    .B1(_2424_),
    .C1(_2425_),
    .Y(_2989_));
 sky130_fd_sc_hd__and4b_1 _7006_ (.A_N(_2324_),
    .B(_2757_),
    .C(_2830_),
    .D(_2989_),
    .X(_2990_));
 sky130_fd_sc_hd__and3b_1 _7007_ (.A_N(_2915_),
    .B(_2971_),
    .C(_2990_),
    .X(_2991_));
 sky130_fd_sc_hd__or3b_1 _7008_ (.A(_2974_),
    .B(_2991_),
    .C_N(_2967_),
    .X(_2992_));
 sky130_fd_sc_hd__or4b_1 _7009_ (.A(_2979_),
    .B(_2983_),
    .C(_2988_),
    .D_N(_2992_),
    .X(_2993_));
 sky130_fd_sc_hd__clkbuf_1 _7010_ (.A(_2993_),
    .X(_0383_));
 sky130_fd_sc_hd__and2_1 _7011_ (.A(_1652_),
    .B(_1654_),
    .X(_2994_));
 sky130_fd_sc_hd__clkbuf_1 _7012_ (.A(_2994_),
    .X(_0057_));
 sky130_fd_sc_hd__and2_1 _7013_ (.A(_1627_),
    .B(_1654_),
    .X(_2995_));
 sky130_fd_sc_hd__clkbuf_1 _7014_ (.A(_2995_),
    .X(_0058_));
 sky130_fd_sc_hd__and2_1 _7015_ (.A(_1627_),
    .B(_1508_),
    .X(_2996_));
 sky130_fd_sc_hd__clkbuf_1 _7016_ (.A(_2996_),
    .X(_0059_));
 sky130_fd_sc_hd__and2_1 _7017_ (.A(_1627_),
    .B(_1508_),
    .X(_2997_));
 sky130_fd_sc_hd__clkbuf_1 _7018_ (.A(_2997_),
    .X(_0060_));
 sky130_fd_sc_hd__and2_1 _7019_ (.A(_1627_),
    .B(_1508_),
    .X(_2998_));
 sky130_fd_sc_hd__clkbuf_1 _7020_ (.A(_2998_),
    .X(_0061_));
 sky130_fd_sc_hd__and2_1 _7021_ (.A(_1627_),
    .B(_1508_),
    .X(_2999_));
 sky130_fd_sc_hd__clkbuf_1 _7022_ (.A(_2999_),
    .X(_0062_));
 sky130_fd_sc_hd__and2_1 _7023_ (.A(_1627_),
    .B(_1508_),
    .X(_3000_));
 sky130_fd_sc_hd__clkbuf_1 _7024_ (.A(_3000_),
    .X(_0063_));
 sky130_fd_sc_hd__and2_1 _7025_ (.A(_1627_),
    .B(_1508_),
    .X(_3001_));
 sky130_fd_sc_hd__clkbuf_1 _7026_ (.A(_3001_),
    .X(_0064_));
 sky130_fd_sc_hd__nand2_1 _7027_ (.A(_1345_),
    .B(_1602_),
    .Y(_3002_));
 sky130_fd_sc_hd__mux2_1 _7028_ (.A0(_1993_),
    .A1(net270),
    .S(_3002_),
    .X(_3003_));
 sky130_fd_sc_hd__clkbuf_1 _7029_ (.A(net1360),
    .X(_0392_));
 sky130_fd_sc_hd__mux2_1 _7030_ (.A0(_1996_),
    .A1(net264),
    .S(_3002_),
    .X(_3004_));
 sky130_fd_sc_hd__clkbuf_1 _7031_ (.A(net1316),
    .X(_0393_));
 sky130_fd_sc_hd__nand2_2 _7032_ (.A(_1140_),
    .B(_1858_),
    .Y(_3005_));
 sky130_fd_sc_hd__mux2_1 _7033_ (.A0(_1993_),
    .A1(net265),
    .S(_3005_),
    .X(_3006_));
 sky130_fd_sc_hd__clkbuf_1 _7034_ (.A(net1369),
    .X(_0394_));
 sky130_fd_sc_hd__mux2_1 _7035_ (.A0(_1996_),
    .A1(net266),
    .S(_3005_),
    .X(_3007_));
 sky130_fd_sc_hd__clkbuf_1 _7036_ (.A(net1298),
    .X(_0395_));
 sky130_fd_sc_hd__mux2_1 _7037_ (.A0(_2030_),
    .A1(net267),
    .S(_3005_),
    .X(_3008_));
 sky130_fd_sc_hd__clkbuf_1 _7038_ (.A(net1282),
    .X(_0396_));
 sky130_fd_sc_hd__mux2_1 _7039_ (.A0(_2032_),
    .A1(net268),
    .S(_3005_),
    .X(_3009_));
 sky130_fd_sc_hd__clkbuf_1 _7040_ (.A(net1202),
    .X(_0397_));
 sky130_fd_sc_hd__mux2_1 _7041_ (.A0(_2034_),
    .A1(net269),
    .S(_3005_),
    .X(_3010_));
 sky130_fd_sc_hd__clkbuf_1 _7042_ (.A(net847),
    .X(_0398_));
 sky130_fd_sc_hd__nand2_2 _7043_ (.A(_1028_),
    .B(_1858_),
    .Y(_3011_));
 sky130_fd_sc_hd__mux2_1 _7044_ (.A0(_1993_),
    .A1(net271),
    .S(_3011_),
    .X(_3012_));
 sky130_fd_sc_hd__clkbuf_1 _7045_ (.A(net1391),
    .X(_0399_));
 sky130_fd_sc_hd__mux2_1 _7046_ (.A0(_1996_),
    .A1(net272),
    .S(_3011_),
    .X(_3013_));
 sky130_fd_sc_hd__clkbuf_1 _7047_ (.A(net1289),
    .X(_0400_));
 sky130_fd_sc_hd__mux2_1 _7048_ (.A0(_2030_),
    .A1(net273),
    .S(_3011_),
    .X(_3014_));
 sky130_fd_sc_hd__clkbuf_1 _7049_ (.A(net1251),
    .X(_0401_));
 sky130_fd_sc_hd__mux2_1 _7050_ (.A0(_2032_),
    .A1(net260),
    .S(_3011_),
    .X(_3015_));
 sky130_fd_sc_hd__clkbuf_1 _7051_ (.A(net1215),
    .X(_0402_));
 sky130_fd_sc_hd__mux2_1 _7052_ (.A0(_2034_),
    .A1(net261),
    .S(_3011_),
    .X(_3016_));
 sky130_fd_sc_hd__clkbuf_1 _7053_ (.A(net850),
    .X(_0403_));
 sky130_fd_sc_hd__mux2_1 _7054_ (.A0(_1708_),
    .A1(net262),
    .S(_3011_),
    .X(_3017_));
 sky130_fd_sc_hd__clkbuf_1 _7055_ (.A(net1264),
    .X(_0404_));
 sky130_fd_sc_hd__and2_1 _7056_ (.A(_0946_),
    .B(net525),
    .X(_3018_));
 sky130_fd_sc_hd__clkbuf_4 _7057_ (.A(_3018_),
    .X(_3019_));
 sky130_fd_sc_hd__mux2_1 _7058_ (.A0(net281),
    .A1(_1878_),
    .S(_3019_),
    .X(_3020_));
 sky130_fd_sc_hd__clkbuf_1 _7059_ (.A(net1367),
    .X(_0405_));
 sky130_fd_sc_hd__mux2_1 _7060_ (.A0(net282),
    .A1(_1905_),
    .S(_3019_),
    .X(_3021_));
 sky130_fd_sc_hd__clkbuf_1 _7061_ (.A(net999),
    .X(_0406_));
 sky130_fd_sc_hd__mux2_1 _7062_ (.A0(net283),
    .A1(_2051_),
    .S(_3019_),
    .X(_3022_));
 sky130_fd_sc_hd__clkbuf_1 _7063_ (.A(net1055),
    .X(_0407_));
 sky130_fd_sc_hd__mux2_1 _7064_ (.A0(net284),
    .A1(net552),
    .S(_3019_),
    .X(_3023_));
 sky130_fd_sc_hd__clkbuf_1 _7065_ (.A(net585),
    .X(_0408_));
 sky130_fd_sc_hd__mux2_1 _7066_ (.A0(net286),
    .A1(_1668_),
    .S(_3019_),
    .X(_3024_));
 sky130_fd_sc_hd__clkbuf_1 _7067_ (.A(net670),
    .X(_0409_));
 sky130_fd_sc_hd__mux2_1 _7068_ (.A0(net287),
    .A1(_1672_),
    .S(_3019_),
    .X(_3025_));
 sky130_fd_sc_hd__clkbuf_1 _7069_ (.A(net845),
    .X(_0410_));
 sky130_fd_sc_hd__mux2_1 _7070_ (.A0(net288),
    .A1(_1689_),
    .S(_3019_),
    .X(_3026_));
 sky130_fd_sc_hd__clkbuf_1 _7071_ (.A(net891),
    .X(_0411_));
 sky130_fd_sc_hd__mux2_1 _7072_ (.A0(net289),
    .A1(_1678_),
    .S(_3019_),
    .X(_3027_));
 sky130_fd_sc_hd__clkbuf_1 _7073_ (.A(net734),
    .X(_0412_));
 sky130_fd_sc_hd__nand2_1 _7074_ (.A(_1421_),
    .B(_1602_),
    .Y(_3028_));
 sky130_fd_sc_hd__mux2_1 _7075_ (.A0(_1993_),
    .A1(net263),
    .S(_3028_),
    .X(_3029_));
 sky130_fd_sc_hd__clkbuf_1 _7076_ (.A(net1314),
    .X(_0413_));
 sky130_fd_sc_hd__and2_1 _7077_ (.A(_1217_),
    .B(net526),
    .X(_3030_));
 sky130_fd_sc_hd__mux2_1 _7078_ (.A0(net300),
    .A1(_1878_),
    .S(net571),
    .X(_3031_));
 sky130_fd_sc_hd__clkbuf_1 _7079_ (.A(net1381),
    .X(_0414_));
 sky130_fd_sc_hd__mux2_1 _7080_ (.A0(net301),
    .A1(_1905_),
    .S(net571),
    .X(_3032_));
 sky130_fd_sc_hd__clkbuf_1 _7081_ (.A(net1579),
    .X(_0415_));
 sky130_fd_sc_hd__mux2_1 _7082_ (.A0(net302),
    .A1(_2051_),
    .S(net571),
    .X(_3033_));
 sky130_fd_sc_hd__clkbuf_1 _7083_ (.A(net971),
    .X(_0416_));
 sky130_fd_sc_hd__mux2_1 _7084_ (.A0(net303),
    .A1(net552),
    .S(net571),
    .X(_3034_));
 sky130_fd_sc_hd__clkbuf_1 _7085_ (.A(net572),
    .X(_0417_));
 sky130_fd_sc_hd__nand2_1 _7086_ (.A(_1325_),
    .B(_1602_),
    .Y(_3035_));
 sky130_fd_sc_hd__mux2_1 _7087_ (.A0(_1996_),
    .A1(net324),
    .S(_3035_),
    .X(_3036_));
 sky130_fd_sc_hd__clkbuf_1 _7088_ (.A(net1308),
    .X(_0418_));
 sky130_fd_sc_hd__mux2_1 _7089_ (.A0(_1993_),
    .A1(net325),
    .S(_3035_),
    .X(_3037_));
 sky130_fd_sc_hd__clkbuf_1 _7090_ (.A(net1370),
    .X(_0419_));
 sky130_fd_sc_hd__nand2_4 _7091_ (.A(_0851_),
    .B(_1967_),
    .Y(_3038_));
 sky130_fd_sc_hd__mux2_1 _7092_ (.A0(_1993_),
    .A1(net316),
    .S(_3038_),
    .X(_3039_));
 sky130_fd_sc_hd__clkbuf_1 _7093_ (.A(net1413),
    .X(_0420_));
 sky130_fd_sc_hd__mux2_1 _7094_ (.A0(_1996_),
    .A1(net317),
    .S(_3038_),
    .X(_3040_));
 sky130_fd_sc_hd__clkbuf_1 _7095_ (.A(net1313),
    .X(_0421_));
 sky130_fd_sc_hd__mux2_1 _7096_ (.A0(_2030_),
    .A1(net318),
    .S(_3038_),
    .X(_3041_));
 sky130_fd_sc_hd__clkbuf_1 _7097_ (.A(net1254),
    .X(_0422_));
 sky130_fd_sc_hd__mux2_1 _7098_ (.A0(_2032_),
    .A1(net319),
    .S(_3038_),
    .X(_3042_));
 sky130_fd_sc_hd__clkbuf_1 _7099_ (.A(net1208),
    .X(_0423_));
 sky130_fd_sc_hd__mux2_1 _7100_ (.A0(_2034_),
    .A1(net320),
    .S(_3038_),
    .X(_3043_));
 sky130_fd_sc_hd__clkbuf_1 _7101_ (.A(net833),
    .X(_0424_));
 sky130_fd_sc_hd__mux2_1 _7102_ (.A0(_1708_),
    .A1(net321),
    .S(_3038_),
    .X(_3044_));
 sky130_fd_sc_hd__clkbuf_1 _7103_ (.A(net1273),
    .X(_0425_));
 sky130_fd_sc_hd__mux2_1 _7104_ (.A0(_1710_),
    .A1(net322),
    .S(_3038_),
    .X(_3045_));
 sky130_fd_sc_hd__clkbuf_1 _7105_ (.A(net1258),
    .X(_0426_));
 sky130_fd_sc_hd__mux2_1 _7106_ (.A0(_1712_),
    .A1(net323),
    .S(_3038_),
    .X(_3046_));
 sky130_fd_sc_hd__clkbuf_1 _7107_ (.A(net1204),
    .X(_0427_));
 sky130_fd_sc_hd__nand2_1 _7108_ (.A(_1381_),
    .B(_1602_),
    .Y(_3047_));
 sky130_fd_sc_hd__mux2_1 _7109_ (.A0(_1993_),
    .A1(reset_reg),
    .S(_3047_),
    .X(_3048_));
 sky130_fd_sc_hd__clkbuf_1 _7110_ (.A(net1415),
    .X(_0428_));
 sky130_fd_sc_hd__or3_1 _7111_ (.A(_0893_),
    .B(_0974_),
    .C(net939),
    .X(_3049_));
 sky130_fd_sc_hd__o211a_1 _7112_ (.A1(net204),
    .A2(_1409_),
    .B1(_1602_),
    .C1(_3049_),
    .X(_0429_));
 sky130_fd_sc_hd__nand2_2 _7113_ (.A(_1011_),
    .B(_1967_),
    .Y(_3050_));
 sky130_fd_sc_hd__mux2_1 _7114_ (.A0(_2034_),
    .A1(net657),
    .S(_3050_),
    .X(_3051_));
 sky130_fd_sc_hd__clkbuf_1 _7115_ (.A(net658),
    .X(_0430_));
 sky130_fd_sc_hd__mux2_1 _7116_ (.A0(_2032_),
    .A1(serial_bb_load),
    .S(_3050_),
    .X(_3052_));
 sky130_fd_sc_hd__clkbuf_1 _7117_ (.A(net931),
    .X(_0431_));
 sky130_fd_sc_hd__mux2_1 _7118_ (.A0(_2030_),
    .A1(serial_bb_resetn),
    .S(_3050_),
    .X(_3053_));
 sky130_fd_sc_hd__clkbuf_1 _7119_ (.A(net1097),
    .X(_0432_));
 sky130_fd_sc_hd__mux2_1 _7120_ (.A0(_1708_),
    .A1(serial_bb_data_1),
    .S(_3050_),
    .X(_3054_));
 sky130_fd_sc_hd__clkbuf_1 _7121_ (.A(net1095),
    .X(_0433_));
 sky130_fd_sc_hd__mux2_1 _7122_ (.A0(_1710_),
    .A1(serial_bb_data_2),
    .S(_3050_),
    .X(_3055_));
 sky130_fd_sc_hd__clkbuf_1 _7123_ (.A(net1134),
    .X(_0434_));
 sky130_fd_sc_hd__mux2_1 _7124_ (.A0(_1996_),
    .A1(serial_bb_enable),
    .S(_3050_),
    .X(_3056_));
 sky130_fd_sc_hd__clkbuf_1 _7125_ (.A(net1056),
    .X(_0435_));
 sky130_fd_sc_hd__or3_1 _7126_ (.A(_0917_),
    .B(_1010_),
    .C(net939),
    .X(_3057_));
 sky130_fd_sc_hd__o211a_1 _7127_ (.A1(net1195),
    .A2(_1011_),
    .B1(_1602_),
    .C1(_3057_),
    .X(_0436_));
 sky130_fd_sc_hd__clkbuf_4 _7128_ (.A(_1597_),
    .X(_3058_));
 sky130_fd_sc_hd__nand2_1 _7129_ (.A(_1357_),
    .B(_1602_),
    .Y(_3059_));
 sky130_fd_sc_hd__mux2_1 _7130_ (.A0(_3058_),
    .A1(net1422),
    .S(_3059_),
    .X(_3060_));
 sky130_fd_sc_hd__clkbuf_1 _7131_ (.A(_3060_),
    .X(_0437_));
 sky130_fd_sc_hd__and2_1 _7132_ (.A(_1226_),
    .B(_1871_),
    .X(_3061_));
 sky130_fd_sc_hd__mux2_1 _7133_ (.A0(clk1_output_dest),
    .A1(_2051_),
    .S(_3061_),
    .X(_3062_));
 sky130_fd_sc_hd__clkbuf_1 _7134_ (.A(net1211),
    .X(_0438_));
 sky130_fd_sc_hd__mux2_1 _7135_ (.A0(clk2_output_dest),
    .A1(_1905_),
    .S(_3061_),
    .X(_3063_));
 sky130_fd_sc_hd__clkbuf_1 _7136_ (.A(net1299),
    .X(_0439_));
 sky130_fd_sc_hd__mux2_1 _7137_ (.A0(trap_output_dest),
    .A1(net939),
    .S(_3061_),
    .X(_3064_));
 sky130_fd_sc_hd__clkbuf_1 _7138_ (.A(net1374),
    .X(_0440_));
 sky130_fd_sc_hd__nand2_1 _7139_ (.A(_1297_),
    .B(_1602_),
    .Y(_3065_));
 sky130_fd_sc_hd__mux2_1 _7140_ (.A0(_3058_),
    .A1(irq_1_inputsrc),
    .S(_3065_),
    .X(_3066_));
 sky130_fd_sc_hd__clkbuf_1 _7141_ (.A(net1373),
    .X(_0441_));
 sky130_fd_sc_hd__mux2_1 _7142_ (.A0(_1996_),
    .A1(irq_2_inputsrc),
    .S(_3065_),
    .X(_3067_));
 sky130_fd_sc_hd__clkbuf_1 _7143_ (.A(net1309),
    .X(_0442_));
 sky130_fd_sc_hd__nand2_8 _7144_ (.A(net370),
    .B(_1967_),
    .Y(_3068_));
 sky130_fd_sc_hd__mux2_1 _7145_ (.A0(_3058_),
    .A1(\mgmt_gpio_data[32] ),
    .S(_3068_),
    .X(_3069_));
 sky130_fd_sc_hd__clkbuf_1 _7146_ (.A(net1439),
    .X(_0443_));
 sky130_fd_sc_hd__clkbuf_8 _7147_ (.A(net543),
    .X(_3070_));
 sky130_fd_sc_hd__mux2_1 _7148_ (.A0(_3070_),
    .A1(\mgmt_gpio_data[33] ),
    .S(_3068_),
    .X(_3071_));
 sky130_fd_sc_hd__clkbuf_1 _7149_ (.A(net652),
    .X(_0444_));
 sky130_fd_sc_hd__mux2_1 _7150_ (.A0(_2030_),
    .A1(\mgmt_gpio_data[34] ),
    .S(_3068_),
    .X(_3072_));
 sky130_fd_sc_hd__clkbuf_1 _7151_ (.A(net922),
    .X(_0445_));
 sky130_fd_sc_hd__mux2_1 _7152_ (.A0(_2032_),
    .A1(\mgmt_gpio_data[35] ),
    .S(_3068_),
    .X(_3073_));
 sky130_fd_sc_hd__clkbuf_1 _7153_ (.A(net966),
    .X(_0446_));
 sky130_fd_sc_hd__mux2_1 _7154_ (.A0(_2034_),
    .A1(\mgmt_gpio_data[36] ),
    .S(_3068_),
    .X(_3074_));
 sky130_fd_sc_hd__clkbuf_1 _7155_ (.A(net787),
    .X(_0447_));
 sky130_fd_sc_hd__mux2_1 _7156_ (.A0(_1708_),
    .A1(\mgmt_gpio_data[37] ),
    .S(_3068_),
    .X(_3075_));
 sky130_fd_sc_hd__clkbuf_1 _7157_ (.A(net1324),
    .X(_0448_));
 sky130_fd_sc_hd__or4_1 _7158_ (.A(_0909_),
    .B(_0940_),
    .C(_1506_),
    .D(net611),
    .X(_3076_));
 sky130_fd_sc_hd__buf_6 _7159_ (.A(_3076_),
    .X(_3077_));
 sky130_fd_sc_hd__mux2_1 _7160_ (.A0(_3058_),
    .A1(net1320),
    .S(_3077_),
    .X(_3078_));
 sky130_fd_sc_hd__clkbuf_1 _7161_ (.A(net1321),
    .X(_0449_));
 sky130_fd_sc_hd__mux2_1 _7162_ (.A0(_3070_),
    .A1(net688),
    .S(_3077_),
    .X(_3079_));
 sky130_fd_sc_hd__clkbuf_1 _7163_ (.A(net689),
    .X(_0450_));
 sky130_fd_sc_hd__mux2_1 _7164_ (.A0(_2030_),
    .A1(net992),
    .S(_3077_),
    .X(_3080_));
 sky130_fd_sc_hd__clkbuf_1 _7165_ (.A(net993),
    .X(_0451_));
 sky130_fd_sc_hd__mux2_1 _7166_ (.A0(_2032_),
    .A1(net880),
    .S(_3077_),
    .X(_3081_));
 sky130_fd_sc_hd__clkbuf_1 _7167_ (.A(net881),
    .X(_0452_));
 sky130_fd_sc_hd__mux2_1 _7168_ (.A0(_2034_),
    .A1(\mgmt_gpio_data_buf[4] ),
    .S(_3077_),
    .X(_3082_));
 sky130_fd_sc_hd__clkbuf_1 _7169_ (.A(net612),
    .X(_0453_));
 sky130_fd_sc_hd__mux2_1 _7170_ (.A0(_1708_),
    .A1(net1145),
    .S(_3077_),
    .X(_3083_));
 sky130_fd_sc_hd__clkbuf_1 _7171_ (.A(net1146),
    .X(_0454_));
 sky130_fd_sc_hd__mux2_1 _7172_ (.A0(_1710_),
    .A1(net1187),
    .S(_3077_),
    .X(_3084_));
 sky130_fd_sc_hd__clkbuf_1 _7173_ (.A(net1188),
    .X(_0455_));
 sky130_fd_sc_hd__mux2_1 _7174_ (.A0(_1712_),
    .A1(net1073),
    .S(_3077_),
    .X(_3085_));
 sky130_fd_sc_hd__clkbuf_1 _7175_ (.A(net1074),
    .X(_0456_));
 sky130_fd_sc_hd__and2_1 _7176_ (.A(_0971_),
    .B(net525),
    .X(_3086_));
 sky130_fd_sc_hd__buf_4 _7177_ (.A(_3086_),
    .X(_3087_));
 sky130_fd_sc_hd__mux2_1 _7178_ (.A0(net1333),
    .A1(net939),
    .S(_3087_),
    .X(_3088_));
 sky130_fd_sc_hd__clkbuf_1 _7179_ (.A(_3088_),
    .X(_0457_));
 sky130_fd_sc_hd__mux2_1 _7180_ (.A0(net1080),
    .A1(_1905_),
    .S(_3087_),
    .X(_3089_));
 sky130_fd_sc_hd__clkbuf_1 _7181_ (.A(_3089_),
    .X(_0458_));
 sky130_fd_sc_hd__mux2_1 _7182_ (.A0(net1249),
    .A1(_2051_),
    .S(_3087_),
    .X(_3090_));
 sky130_fd_sc_hd__clkbuf_1 _7183_ (.A(net1250),
    .X(_0459_));
 sky130_fd_sc_hd__mux2_1 _7184_ (.A0(\gpio_configure[0][3] ),
    .A1(net552),
    .S(_3087_),
    .X(_3091_));
 sky130_fd_sc_hd__clkbuf_1 _7185_ (.A(net709),
    .X(_0460_));
 sky130_fd_sc_hd__mux2_1 _7186_ (.A0(net851),
    .A1(_1668_),
    .S(_3087_),
    .X(_3092_));
 sky130_fd_sc_hd__clkbuf_1 _7187_ (.A(_3092_),
    .X(_0461_));
 sky130_fd_sc_hd__mux2_1 _7188_ (.A0(net836),
    .A1(_1672_),
    .S(_3087_),
    .X(_3093_));
 sky130_fd_sc_hd__clkbuf_1 _7189_ (.A(net837),
    .X(_0462_));
 sky130_fd_sc_hd__mux2_1 _7190_ (.A0(net828),
    .A1(_1689_),
    .S(_3087_),
    .X(_3094_));
 sky130_fd_sc_hd__clkbuf_1 _7191_ (.A(net829),
    .X(_0463_));
 sky130_fd_sc_hd__mux2_1 _7192_ (.A0(net711),
    .A1(_1678_),
    .S(_3087_),
    .X(_3095_));
 sky130_fd_sc_hd__clkbuf_1 _7193_ (.A(net712),
    .X(_0464_));
 sky130_fd_sc_hd__nand2_8 _7194_ (.A(net383),
    .B(_1967_),
    .Y(_3096_));
 sky130_fd_sc_hd__mux2_1 _7195_ (.A0(_3058_),
    .A1(net1414),
    .S(_3096_),
    .X(_3097_));
 sky130_fd_sc_hd__clkbuf_1 _7196_ (.A(_3097_),
    .X(_0465_));
 sky130_fd_sc_hd__mux2_1 _7197_ (.A0(_3070_),
    .A1(net822),
    .S(_3096_),
    .X(_3098_));
 sky130_fd_sc_hd__clkbuf_1 _7198_ (.A(net823),
    .X(_0466_));
 sky130_fd_sc_hd__mux2_1 _7199_ (.A0(_2030_),
    .A1(net1306),
    .S(_3096_),
    .X(_3099_));
 sky130_fd_sc_hd__clkbuf_1 _7200_ (.A(net1307),
    .X(_0467_));
 sky130_fd_sc_hd__mux2_1 _7201_ (.A0(_2032_),
    .A1(net1206),
    .S(_3096_),
    .X(_3100_));
 sky130_fd_sc_hd__clkbuf_1 _7202_ (.A(net1207),
    .X(_0468_));
 sky130_fd_sc_hd__mux2_1 _7203_ (.A0(_2034_),
    .A1(net858),
    .S(_3096_),
    .X(_3101_));
 sky130_fd_sc_hd__clkbuf_1 _7204_ (.A(net859),
    .X(_0469_));
 sky130_fd_sc_hd__mux2_1 _7205_ (.A0(_1708_),
    .A1(net1311),
    .S(_3096_),
    .X(_3102_));
 sky130_fd_sc_hd__clkbuf_1 _7206_ (.A(net1312),
    .X(_0470_));
 sky130_fd_sc_hd__mux2_1 _7207_ (.A0(_1710_),
    .A1(net1182),
    .S(_3096_),
    .X(_3103_));
 sky130_fd_sc_hd__clkbuf_1 _7208_ (.A(net1183),
    .X(_0471_));
 sky130_fd_sc_hd__mux2_1 _7209_ (.A0(_1712_),
    .A1(net1137),
    .S(_3096_),
    .X(_3104_));
 sky130_fd_sc_hd__clkbuf_1 _7210_ (.A(net1138),
    .X(_0472_));
 sky130_fd_sc_hd__nand2_8 _7211_ (.A(net385),
    .B(_1967_),
    .Y(_3105_));
 sky130_fd_sc_hd__mux2_1 _7212_ (.A0(_3058_),
    .A1(net1417),
    .S(_3105_),
    .X(_3106_));
 sky130_fd_sc_hd__clkbuf_1 _7213_ (.A(_3106_),
    .X(_0473_));
 sky130_fd_sc_hd__mux2_1 _7214_ (.A0(_3070_),
    .A1(net641),
    .S(_3105_),
    .X(_3107_));
 sky130_fd_sc_hd__clkbuf_1 _7215_ (.A(net642),
    .X(_0474_));
 sky130_fd_sc_hd__mux2_1 _7216_ (.A0(_2030_),
    .A1(net1285),
    .S(_3105_),
    .X(_3108_));
 sky130_fd_sc_hd__clkbuf_1 _7217_ (.A(net1286),
    .X(_0475_));
 sky130_fd_sc_hd__mux2_1 _7218_ (.A0(_2032_),
    .A1(\gpio_configure[2][3] ),
    .S(_3105_),
    .X(_3109_));
 sky130_fd_sc_hd__clkbuf_1 _7219_ (.A(net1232),
    .X(_0476_));
 sky130_fd_sc_hd__mux2_1 _7220_ (.A0(_2034_),
    .A1(net720),
    .S(_3105_),
    .X(_3110_));
 sky130_fd_sc_hd__clkbuf_1 _7221_ (.A(net721),
    .X(_0477_));
 sky130_fd_sc_hd__mux2_1 _7222_ (.A0(_1708_),
    .A1(net1185),
    .S(_3105_),
    .X(_3111_));
 sky130_fd_sc_hd__clkbuf_1 _7223_ (.A(net1186),
    .X(_0478_));
 sky130_fd_sc_hd__mux2_1 _7224_ (.A0(_1710_),
    .A1(net1189),
    .S(_3105_),
    .X(_3112_));
 sky130_fd_sc_hd__clkbuf_1 _7225_ (.A(net1190),
    .X(_0479_));
 sky130_fd_sc_hd__mux2_1 _7226_ (.A0(_1712_),
    .A1(net1132),
    .S(_3105_),
    .X(_3113_));
 sky130_fd_sc_hd__clkbuf_1 _7227_ (.A(net1133),
    .X(_0480_));
 sky130_fd_sc_hd__nand2_8 _7228_ (.A(_0857_),
    .B(_1967_),
    .Y(_3114_));
 sky130_fd_sc_hd__mux2_1 _7229_ (.A0(_3058_),
    .A1(\gpio_configure[3][0] ),
    .S(_3114_),
    .X(_3115_));
 sky130_fd_sc_hd__clkbuf_1 _7230_ (.A(net1364),
    .X(_0481_));
 sky130_fd_sc_hd__mux2_1 _7231_ (.A0(_3070_),
    .A1(net801),
    .S(_3114_),
    .X(_3116_));
 sky130_fd_sc_hd__clkbuf_1 _7232_ (.A(net802),
    .X(_0482_));
 sky130_fd_sc_hd__buf_4 _7233_ (.A(_1610_),
    .X(_3117_));
 sky130_fd_sc_hd__mux2_1 _7234_ (.A0(_3117_),
    .A1(net1371),
    .S(_3114_),
    .X(_3118_));
 sky130_fd_sc_hd__clkbuf_1 _7235_ (.A(_3118_),
    .X(_0483_));
 sky130_fd_sc_hd__clkbuf_4 _7236_ (.A(_1614_),
    .X(_3119_));
 sky130_fd_sc_hd__mux2_1 _7237_ (.A0(_3119_),
    .A1(\gpio_configure[3][3] ),
    .S(_3114_),
    .X(_3120_));
 sky130_fd_sc_hd__clkbuf_1 _7238_ (.A(net1194),
    .X(_0484_));
 sky130_fd_sc_hd__buf_6 _7239_ (.A(net530),
    .X(_3121_));
 sky130_fd_sc_hd__mux2_1 _7240_ (.A0(_3121_),
    .A1(net792),
    .S(_3114_),
    .X(_3122_));
 sky130_fd_sc_hd__clkbuf_1 _7241_ (.A(net793),
    .X(_0485_));
 sky130_fd_sc_hd__buf_4 _7242_ (.A(net521),
    .X(_3123_));
 sky130_fd_sc_hd__mux2_1 _7243_ (.A0(_3123_),
    .A1(net686),
    .S(_3114_),
    .X(_3124_));
 sky130_fd_sc_hd__clkbuf_1 _7244_ (.A(net687),
    .X(_0486_));
 sky130_fd_sc_hd__mux2_1 _7245_ (.A0(_1710_),
    .A1(net1291),
    .S(_3114_),
    .X(_3125_));
 sky130_fd_sc_hd__clkbuf_1 _7246_ (.A(net1292),
    .X(_0487_));
 sky130_fd_sc_hd__mux2_1 _7247_ (.A0(_1712_),
    .A1(net1222),
    .S(_3114_),
    .X(_3126_));
 sky130_fd_sc_hd__clkbuf_1 _7248_ (.A(net1223),
    .X(_0488_));
 sky130_fd_sc_hd__nand2_8 _7249_ (.A(_0967_),
    .B(_1967_),
    .Y(_3127_));
 sky130_fd_sc_hd__mux2_1 _7250_ (.A0(_3058_),
    .A1(net1377),
    .S(_3127_),
    .X(_3128_));
 sky130_fd_sc_hd__clkbuf_1 _7251_ (.A(_3128_),
    .X(_0489_));
 sky130_fd_sc_hd__mux2_1 _7252_ (.A0(_3070_),
    .A1(net748),
    .S(_3127_),
    .X(_3129_));
 sky130_fd_sc_hd__clkbuf_1 _7253_ (.A(net749),
    .X(_0490_));
 sky130_fd_sc_hd__mux2_1 _7254_ (.A0(_3117_),
    .A1(net1076),
    .S(_3127_),
    .X(_3130_));
 sky130_fd_sc_hd__clkbuf_1 _7255_ (.A(net1077),
    .X(_0491_));
 sky130_fd_sc_hd__mux2_1 _7256_ (.A0(_3119_),
    .A1(\gpio_configure[4][3] ),
    .S(_3127_),
    .X(_3131_));
 sky130_fd_sc_hd__clkbuf_1 _7257_ (.A(net1199),
    .X(_0492_));
 sky130_fd_sc_hd__mux2_1 _7258_ (.A0(_3121_),
    .A1(net671),
    .S(_3127_),
    .X(_3132_));
 sky130_fd_sc_hd__clkbuf_1 _7259_ (.A(net672),
    .X(_0493_));
 sky130_fd_sc_hd__mux2_1 _7260_ (.A0(_3123_),
    .A1(net766),
    .S(_3127_),
    .X(_3133_));
 sky130_fd_sc_hd__clkbuf_1 _7261_ (.A(net767),
    .X(_0494_));
 sky130_fd_sc_hd__mux2_1 _7262_ (.A0(_1710_),
    .A1(net1300),
    .S(_3127_),
    .X(_3134_));
 sky130_fd_sc_hd__clkbuf_1 _7263_ (.A(net1301),
    .X(_0495_));
 sky130_fd_sc_hd__mux2_1 _7264_ (.A0(_1712_),
    .A1(net1176),
    .S(_3127_),
    .X(_3135_));
 sky130_fd_sc_hd__clkbuf_1 _7265_ (.A(net1177),
    .X(_0496_));
 sky130_fd_sc_hd__nand2_8 _7266_ (.A(net363),
    .B(_1967_),
    .Y(_3136_));
 sky130_fd_sc_hd__mux2_1 _7267_ (.A0(_3058_),
    .A1(net1418),
    .S(_3136_),
    .X(_3137_));
 sky130_fd_sc_hd__clkbuf_1 _7268_ (.A(_3137_),
    .X(_0497_));
 sky130_fd_sc_hd__mux2_1 _7269_ (.A0(_3070_),
    .A1(net640),
    .S(_3136_),
    .X(_3138_));
 sky130_fd_sc_hd__clkbuf_1 _7270_ (.A(_3138_),
    .X(_0498_));
 sky130_fd_sc_hd__mux2_1 _7271_ (.A0(_3117_),
    .A1(net1270),
    .S(_3136_),
    .X(_3139_));
 sky130_fd_sc_hd__clkbuf_1 _7272_ (.A(_3139_),
    .X(_0499_));
 sky130_fd_sc_hd__mux2_1 _7273_ (.A0(_3119_),
    .A1(\gpio_configure[5][3] ),
    .S(_3136_),
    .X(_3140_));
 sky130_fd_sc_hd__clkbuf_1 _7274_ (.A(net1193),
    .X(_0500_));
 sky130_fd_sc_hd__mux2_1 _7275_ (.A0(_3121_),
    .A1(net673),
    .S(_3136_),
    .X(_3141_));
 sky130_fd_sc_hd__clkbuf_1 _7276_ (.A(net674),
    .X(_0501_));
 sky130_fd_sc_hd__mux2_1 _7277_ (.A0(_3123_),
    .A1(net728),
    .S(_3136_),
    .X(_3142_));
 sky130_fd_sc_hd__clkbuf_1 _7278_ (.A(net729),
    .X(_0502_));
 sky130_fd_sc_hd__clkbuf_4 _7279_ (.A(_1689_),
    .X(_3143_));
 sky130_fd_sc_hd__mux2_1 _7280_ (.A0(_3143_),
    .A1(net1271),
    .S(_3136_),
    .X(_3144_));
 sky130_fd_sc_hd__clkbuf_1 _7281_ (.A(net1272),
    .X(_0503_));
 sky130_fd_sc_hd__mux2_1 _7282_ (.A0(_1712_),
    .A1(net1130),
    .S(_3136_),
    .X(_3145_));
 sky130_fd_sc_hd__clkbuf_1 _7283_ (.A(net1131),
    .X(_0504_));
 sky130_fd_sc_hd__nand2_8 _7284_ (.A(net382),
    .B(_1967_),
    .Y(_3146_));
 sky130_fd_sc_hd__mux2_1 _7285_ (.A0(_3058_),
    .A1(net1399),
    .S(_3146_),
    .X(_3147_));
 sky130_fd_sc_hd__clkbuf_1 _7286_ (.A(_3147_),
    .X(_0505_));
 sky130_fd_sc_hd__mux2_1 _7287_ (.A0(_3070_),
    .A1(net621),
    .S(_3146_),
    .X(_3148_));
 sky130_fd_sc_hd__clkbuf_1 _7288_ (.A(net622),
    .X(_0506_));
 sky130_fd_sc_hd__mux2_1 _7289_ (.A0(_3117_),
    .A1(net1275),
    .S(_3146_),
    .X(_3149_));
 sky130_fd_sc_hd__clkbuf_1 _7290_ (.A(net1276),
    .X(_0507_));
 sky130_fd_sc_hd__mux2_1 _7291_ (.A0(_3119_),
    .A1(\gpio_configure[6][3] ),
    .S(_3146_),
    .X(_3150_));
 sky130_fd_sc_hd__clkbuf_1 _7292_ (.A(net946),
    .X(_0508_));
 sky130_fd_sc_hd__mux2_1 _7293_ (.A0(_3121_),
    .A1(net795),
    .S(_3146_),
    .X(_3151_));
 sky130_fd_sc_hd__clkbuf_1 _7294_ (.A(net796),
    .X(_0509_));
 sky130_fd_sc_hd__mux2_1 _7295_ (.A0(_3123_),
    .A1(net724),
    .S(_3146_),
    .X(_3152_));
 sky130_fd_sc_hd__clkbuf_1 _7296_ (.A(net725),
    .X(_0510_));
 sky130_fd_sc_hd__mux2_1 _7297_ (.A0(_3143_),
    .A1(net1304),
    .S(_3146_),
    .X(_3153_));
 sky130_fd_sc_hd__clkbuf_1 _7298_ (.A(net1305),
    .X(_0511_));
 sky130_fd_sc_hd__buf_4 _7299_ (.A(_1678_),
    .X(_3154_));
 sky130_fd_sc_hd__mux2_1 _7300_ (.A0(_3154_),
    .A1(net1068),
    .S(_3146_),
    .X(_3155_));
 sky130_fd_sc_hd__clkbuf_1 _7301_ (.A(net1069),
    .X(_0512_));
 sky130_fd_sc_hd__buf_4 _7302_ (.A(_1597_),
    .X(_3156_));
 sky130_fd_sc_hd__buf_12 _7303_ (.A(net526),
    .X(_3157_));
 sky130_fd_sc_hd__nand2_8 _7304_ (.A(net377),
    .B(_3157_),
    .Y(_3158_));
 sky130_fd_sc_hd__mux2_1 _7305_ (.A0(_3156_),
    .A1(net1426),
    .S(_3158_),
    .X(_3159_));
 sky130_fd_sc_hd__clkbuf_1 _7306_ (.A(_3159_),
    .X(_0513_));
 sky130_fd_sc_hd__mux2_1 _7307_ (.A0(_3070_),
    .A1(net774),
    .S(_3158_),
    .X(_3160_));
 sky130_fd_sc_hd__clkbuf_1 _7308_ (.A(net775),
    .X(_0514_));
 sky130_fd_sc_hd__mux2_1 _7309_ (.A0(_3117_),
    .A1(net1066),
    .S(_3158_),
    .X(_3161_));
 sky130_fd_sc_hd__clkbuf_1 _7310_ (.A(net1067),
    .X(_0515_));
 sky130_fd_sc_hd__mux2_1 _7311_ (.A0(_3119_),
    .A1(\gpio_configure[7][3] ),
    .S(_3158_),
    .X(_3162_));
 sky130_fd_sc_hd__clkbuf_1 _7312_ (.A(net1295),
    .X(_0516_));
 sky130_fd_sc_hd__mux2_1 _7313_ (.A0(_3121_),
    .A1(net813),
    .S(_3158_),
    .X(_3163_));
 sky130_fd_sc_hd__clkbuf_1 _7314_ (.A(net814),
    .X(_0517_));
 sky130_fd_sc_hd__mux2_1 _7315_ (.A0(_3123_),
    .A1(net771),
    .S(_3158_),
    .X(_3164_));
 sky130_fd_sc_hd__clkbuf_1 _7316_ (.A(net772),
    .X(_0518_));
 sky130_fd_sc_hd__mux2_1 _7317_ (.A0(_3143_),
    .A1(net1268),
    .S(_3158_),
    .X(_3165_));
 sky130_fd_sc_hd__clkbuf_1 _7318_ (.A(net1269),
    .X(_0519_));
 sky130_fd_sc_hd__mux2_1 _7319_ (.A0(_3154_),
    .A1(net1033),
    .S(_3158_),
    .X(_3166_));
 sky130_fd_sc_hd__clkbuf_1 _7320_ (.A(net1034),
    .X(_0520_));
 sky130_fd_sc_hd__and2_1 _7321_ (.A(_0973_),
    .B(net525),
    .X(_3167_));
 sky130_fd_sc_hd__buf_8 _7322_ (.A(_3167_),
    .X(_3168_));
 sky130_fd_sc_hd__mux2_1 _7323_ (.A0(net1346),
    .A1(net939),
    .S(_3168_),
    .X(_3169_));
 sky130_fd_sc_hd__clkbuf_1 _7324_ (.A(_3169_),
    .X(_0521_));
 sky130_fd_sc_hd__mux2_1 _7325_ (.A0(net614),
    .A1(_1606_),
    .S(_3168_),
    .X(_3170_));
 sky130_fd_sc_hd__clkbuf_1 _7326_ (.A(_3170_),
    .X(_0522_));
 sky130_fd_sc_hd__mux2_1 _7327_ (.A0(net1226),
    .A1(_2051_),
    .S(_3168_),
    .X(_3171_));
 sky130_fd_sc_hd__clkbuf_1 _7328_ (.A(net1227),
    .X(_0523_));
 sky130_fd_sc_hd__mux2_1 _7329_ (.A0(\gpio_configure[8][3] ),
    .A1(net552),
    .S(_3168_),
    .X(_3172_));
 sky130_fd_sc_hd__clkbuf_1 _7330_ (.A(net573),
    .X(_0524_));
 sky130_fd_sc_hd__mux2_1 _7331_ (.A0(net815),
    .A1(_1668_),
    .S(_3168_),
    .X(_3173_));
 sky130_fd_sc_hd__clkbuf_1 _7332_ (.A(net1625),
    .X(_0525_));
 sky130_fd_sc_hd__mux2_1 _7333_ (.A0(net799),
    .A1(_1672_),
    .S(_3168_),
    .X(_3174_));
 sky130_fd_sc_hd__clkbuf_1 _7334_ (.A(net800),
    .X(_0526_));
 sky130_fd_sc_hd__mux2_1 _7335_ (.A0(net864),
    .A1(_1689_),
    .S(_3168_),
    .X(_3175_));
 sky130_fd_sc_hd__clkbuf_1 _7336_ (.A(net865),
    .X(_0527_));
 sky130_fd_sc_hd__mux2_1 _7337_ (.A0(net713),
    .A1(_1678_),
    .S(_3168_),
    .X(_3176_));
 sky130_fd_sc_hd__clkbuf_1 _7338_ (.A(net714),
    .X(_0528_));
 sky130_fd_sc_hd__nand2_4 _7339_ (.A(net366),
    .B(_3157_),
    .Y(_3177_));
 sky130_fd_sc_hd__mux2_1 _7340_ (.A0(_3156_),
    .A1(net1432),
    .S(_3177_),
    .X(_3178_));
 sky130_fd_sc_hd__clkbuf_1 _7341_ (.A(_3178_),
    .X(_0529_));
 sky130_fd_sc_hd__mux2_1 _7342_ (.A0(_3070_),
    .A1(net625),
    .S(_3177_),
    .X(_3179_));
 sky130_fd_sc_hd__clkbuf_1 _7343_ (.A(net626),
    .X(_0530_));
 sky130_fd_sc_hd__mux2_1 _7344_ (.A0(_3117_),
    .A1(net1287),
    .S(_3177_),
    .X(_3180_));
 sky130_fd_sc_hd__clkbuf_1 _7345_ (.A(_3180_),
    .X(_0531_));
 sky130_fd_sc_hd__mux2_1 _7346_ (.A0(_3119_),
    .A1(\gpio_configure[9][3] ),
    .S(_3177_),
    .X(_3181_));
 sky130_fd_sc_hd__clkbuf_1 _7347_ (.A(net930),
    .X(_0532_));
 sky130_fd_sc_hd__mux2_1 _7348_ (.A0(_3121_),
    .A1(net820),
    .S(_3177_),
    .X(_3182_));
 sky130_fd_sc_hd__clkbuf_1 _7349_ (.A(net821),
    .X(_0533_));
 sky130_fd_sc_hd__mux2_1 _7350_ (.A0(_3123_),
    .A1(net803),
    .S(_3177_),
    .X(_3183_));
 sky130_fd_sc_hd__clkbuf_1 _7351_ (.A(net804),
    .X(_0534_));
 sky130_fd_sc_hd__mux2_1 _7352_ (.A0(_3143_),
    .A1(net1338),
    .S(_3177_),
    .X(_3184_));
 sky130_fd_sc_hd__clkbuf_1 _7353_ (.A(net1339),
    .X(_0535_));
 sky130_fd_sc_hd__mux2_1 _7354_ (.A0(_3154_),
    .A1(net1197),
    .S(_3177_),
    .X(_3185_));
 sky130_fd_sc_hd__clkbuf_1 _7355_ (.A(net1198),
    .X(_0536_));
 sky130_fd_sc_hd__nand2_8 _7356_ (.A(net362),
    .B(_3157_),
    .Y(_3186_));
 sky130_fd_sc_hd__mux2_1 _7357_ (.A0(_3156_),
    .A1(net1428),
    .S(_3186_),
    .X(_3187_));
 sky130_fd_sc_hd__clkbuf_1 _7358_ (.A(_3187_),
    .X(_0537_));
 sky130_fd_sc_hd__buf_2 _7359_ (.A(net543),
    .X(_3188_));
 sky130_fd_sc_hd__mux2_1 _7360_ (.A0(_3188_),
    .A1(net650),
    .S(_3186_),
    .X(_3189_));
 sky130_fd_sc_hd__clkbuf_1 _7361_ (.A(net651),
    .X(_0538_));
 sky130_fd_sc_hd__mux2_1 _7362_ (.A0(_3117_),
    .A1(net1284),
    .S(_3186_),
    .X(_3190_));
 sky130_fd_sc_hd__clkbuf_1 _7363_ (.A(_3190_),
    .X(_0539_));
 sky130_fd_sc_hd__mux2_1 _7364_ (.A0(_3119_),
    .A1(\gpio_configure[10][3] ),
    .S(_3186_),
    .X(_3191_));
 sky130_fd_sc_hd__clkbuf_1 _7365_ (.A(net935),
    .X(_0540_));
 sky130_fd_sc_hd__mux2_1 _7366_ (.A0(_3121_),
    .A1(net783),
    .S(_3186_),
    .X(_3192_));
 sky130_fd_sc_hd__clkbuf_1 _7367_ (.A(net784),
    .X(_0541_));
 sky130_fd_sc_hd__mux2_1 _7368_ (.A0(_3123_),
    .A1(net722),
    .S(_3186_),
    .X(_3193_));
 sky130_fd_sc_hd__clkbuf_1 _7369_ (.A(net723),
    .X(_0542_));
 sky130_fd_sc_hd__mux2_1 _7370_ (.A0(_3143_),
    .A1(net1330),
    .S(_3186_),
    .X(_3194_));
 sky130_fd_sc_hd__clkbuf_1 _7371_ (.A(net1331),
    .X(_0543_));
 sky130_fd_sc_hd__mux2_1 _7372_ (.A0(_3154_),
    .A1(net1174),
    .S(_3186_),
    .X(_3195_));
 sky130_fd_sc_hd__clkbuf_1 _7373_ (.A(net1175),
    .X(_0544_));
 sky130_fd_sc_hd__nand2_8 _7374_ (.A(_0923_),
    .B(_3157_),
    .Y(_3196_));
 sky130_fd_sc_hd__mux2_1 _7375_ (.A0(_3156_),
    .A1(net1359),
    .S(_3196_),
    .X(_3197_));
 sky130_fd_sc_hd__clkbuf_1 _7376_ (.A(_3197_),
    .X(_0545_));
 sky130_fd_sc_hd__mux2_1 _7377_ (.A0(_3188_),
    .A1(net899),
    .S(_3196_),
    .X(_3198_));
 sky130_fd_sc_hd__clkbuf_1 _7378_ (.A(_3198_),
    .X(_0546_));
 sky130_fd_sc_hd__mux2_1 _7379_ (.A0(_3117_),
    .A1(net1288),
    .S(_3196_),
    .X(_3199_));
 sky130_fd_sc_hd__clkbuf_1 _7380_ (.A(_3199_),
    .X(_0547_));
 sky130_fd_sc_hd__mux2_1 _7381_ (.A0(_3119_),
    .A1(\gpio_configure[11][3] ),
    .S(_3196_),
    .X(_3200_));
 sky130_fd_sc_hd__clkbuf_1 _7382_ (.A(net1203),
    .X(_0548_));
 sky130_fd_sc_hd__mux2_1 _7383_ (.A0(_3121_),
    .A1(net824),
    .S(_3196_),
    .X(_3201_));
 sky130_fd_sc_hd__clkbuf_1 _7384_ (.A(net825),
    .X(_0549_));
 sky130_fd_sc_hd__mux2_1 _7385_ (.A0(_3123_),
    .A1(net779),
    .S(_3196_),
    .X(_3202_));
 sky130_fd_sc_hd__clkbuf_1 _7386_ (.A(net780),
    .X(_0550_));
 sky130_fd_sc_hd__mux2_1 _7387_ (.A0(_3143_),
    .A1(net1256),
    .S(_3196_),
    .X(_3203_));
 sky130_fd_sc_hd__clkbuf_1 _7388_ (.A(net1257),
    .X(_0551_));
 sky130_fd_sc_hd__mux2_1 _7389_ (.A0(_3154_),
    .A1(net1039),
    .S(_3196_),
    .X(_3204_));
 sky130_fd_sc_hd__clkbuf_1 _7390_ (.A(net1040),
    .X(_0552_));
 sky130_fd_sc_hd__nand2_4 _7391_ (.A(net387),
    .B(_3157_),
    .Y(_3205_));
 sky130_fd_sc_hd__mux2_1 _7392_ (.A0(_3156_),
    .A1(net1444),
    .S(_3205_),
    .X(_3206_));
 sky130_fd_sc_hd__clkbuf_1 _7393_ (.A(_3206_),
    .X(_0553_));
 sky130_fd_sc_hd__mux2_1 _7394_ (.A0(_3188_),
    .A1(net649),
    .S(_3205_),
    .X(_3207_));
 sky130_fd_sc_hd__clkbuf_1 _7395_ (.A(_3207_),
    .X(_0554_));
 sky130_fd_sc_hd__mux2_1 _7396_ (.A0(_3117_),
    .A1(net1277),
    .S(_3205_),
    .X(_3208_));
 sky130_fd_sc_hd__clkbuf_1 _7397_ (.A(_3208_),
    .X(_0555_));
 sky130_fd_sc_hd__mux2_1 _7398_ (.A0(_3119_),
    .A1(\gpio_configure[12][3] ),
    .S(_3205_),
    .X(_3209_));
 sky130_fd_sc_hd__clkbuf_1 _7399_ (.A(net936),
    .X(_0556_));
 sky130_fd_sc_hd__mux2_1 _7400_ (.A0(_3121_),
    .A1(net791),
    .S(_3205_),
    .X(_3210_));
 sky130_fd_sc_hd__clkbuf_1 _7401_ (.A(net1648),
    .X(_0557_));
 sky130_fd_sc_hd__mux2_1 _7402_ (.A0(_3123_),
    .A1(net785),
    .S(_3205_),
    .X(_3211_));
 sky130_fd_sc_hd__clkbuf_1 _7403_ (.A(net786),
    .X(_0558_));
 sky130_fd_sc_hd__mux2_1 _7404_ (.A0(_3143_),
    .A1(net1340),
    .S(_3205_),
    .X(_3212_));
 sky130_fd_sc_hd__clkbuf_1 _7405_ (.A(net1341),
    .X(_0559_));
 sky130_fd_sc_hd__mux2_1 _7406_ (.A0(_3154_),
    .A1(net1200),
    .S(_3205_),
    .X(_3213_));
 sky130_fd_sc_hd__clkbuf_1 _7407_ (.A(net1201),
    .X(_0560_));
 sky130_fd_sc_hd__nand2_8 _7408_ (.A(net371),
    .B(_3157_),
    .Y(_3214_));
 sky130_fd_sc_hd__mux2_1 _7409_ (.A0(_3156_),
    .A1(net1411),
    .S(_3214_),
    .X(_3215_));
 sky130_fd_sc_hd__clkbuf_1 _7410_ (.A(_3215_),
    .X(_0561_));
 sky130_fd_sc_hd__mux2_1 _7411_ (.A0(_3188_),
    .A1(net895),
    .S(_3214_),
    .X(_3216_));
 sky130_fd_sc_hd__clkbuf_1 _7412_ (.A(_3216_),
    .X(_0562_));
 sky130_fd_sc_hd__mux2_1 _7413_ (.A0(_3117_),
    .A1(net1293),
    .S(_3214_),
    .X(_3217_));
 sky130_fd_sc_hd__clkbuf_1 _7414_ (.A(_3217_),
    .X(_0563_));
 sky130_fd_sc_hd__mux2_1 _7415_ (.A0(_3119_),
    .A1(\gpio_configure[13][3] ),
    .S(_3214_),
    .X(_3218_));
 sky130_fd_sc_hd__clkbuf_1 _7416_ (.A(net1205),
    .X(_0564_));
 sky130_fd_sc_hd__mux2_1 _7417_ (.A0(_3121_),
    .A1(net765),
    .S(_3214_),
    .X(_3219_));
 sky130_fd_sc_hd__clkbuf_1 _7418_ (.A(net1600),
    .X(_0565_));
 sky130_fd_sc_hd__mux2_1 _7419_ (.A0(_3123_),
    .A1(net777),
    .S(_3214_),
    .X(_3220_));
 sky130_fd_sc_hd__clkbuf_1 _7420_ (.A(net778),
    .X(_0566_));
 sky130_fd_sc_hd__mux2_1 _7421_ (.A0(_3143_),
    .A1(net1239),
    .S(_3214_),
    .X(_3221_));
 sky130_fd_sc_hd__clkbuf_1 _7422_ (.A(net1240),
    .X(_0567_));
 sky130_fd_sc_hd__mux2_1 _7423_ (.A0(_3154_),
    .A1(net1036),
    .S(_3214_),
    .X(_3222_));
 sky130_fd_sc_hd__clkbuf_1 _7424_ (.A(net1037),
    .X(_0568_));
 sky130_fd_sc_hd__nand2_8 _7425_ (.A(net375),
    .B(_3157_),
    .Y(_3223_));
 sky130_fd_sc_hd__mux2_1 _7426_ (.A0(_3156_),
    .A1(net1420),
    .S(_3223_),
    .X(_3224_));
 sky130_fd_sc_hd__clkbuf_1 _7427_ (.A(_3224_),
    .X(_0569_));
 sky130_fd_sc_hd__mux2_1 _7428_ (.A0(_3188_),
    .A1(net639),
    .S(_3223_),
    .X(_3225_));
 sky130_fd_sc_hd__clkbuf_1 _7429_ (.A(_3225_),
    .X(_0570_));
 sky130_fd_sc_hd__clkbuf_2 _7430_ (.A(_1610_),
    .X(_3226_));
 sky130_fd_sc_hd__mux2_1 _7431_ (.A0(_3226_),
    .A1(net908),
    .S(_3223_),
    .X(_3227_));
 sky130_fd_sc_hd__clkbuf_1 _7432_ (.A(net909),
    .X(_0571_));
 sky130_fd_sc_hd__clkbuf_2 _7433_ (.A(_1614_),
    .X(_3228_));
 sky130_fd_sc_hd__mux2_1 _7434_ (.A0(_3228_),
    .A1(\gpio_configure[14][3] ),
    .S(_3223_),
    .X(_3229_));
 sky130_fd_sc_hd__clkbuf_1 _7435_ (.A(net861),
    .X(_0572_));
 sky130_fd_sc_hd__clkbuf_2 _7436_ (.A(net530),
    .X(_3230_));
 sky130_fd_sc_hd__mux2_1 _7437_ (.A0(_3230_),
    .A1(net794),
    .S(_3223_),
    .X(_3231_));
 sky130_fd_sc_hd__clkbuf_1 _7438_ (.A(_3231_),
    .X(_0573_));
 sky130_fd_sc_hd__buf_2 _7439_ (.A(net521),
    .X(_3232_));
 sky130_fd_sc_hd__mux2_1 _7440_ (.A0(_3232_),
    .A1(net817),
    .S(_3223_),
    .X(_3233_));
 sky130_fd_sc_hd__clkbuf_1 _7441_ (.A(net818),
    .X(_0574_));
 sky130_fd_sc_hd__mux2_1 _7442_ (.A0(_3143_),
    .A1(net1342),
    .S(_3223_),
    .X(_3234_));
 sky130_fd_sc_hd__clkbuf_1 _7443_ (.A(net1343),
    .X(_0575_));
 sky130_fd_sc_hd__mux2_1 _7444_ (.A0(_3154_),
    .A1(net1354),
    .S(_3223_),
    .X(_3235_));
 sky130_fd_sc_hd__clkbuf_1 _7445_ (.A(_3235_),
    .X(_0576_));
 sky130_fd_sc_hd__nand2_8 _7446_ (.A(_0876_),
    .B(_3157_),
    .Y(_3236_));
 sky130_fd_sc_hd__mux2_1 _7447_ (.A0(_3156_),
    .A1(net1382),
    .S(_3236_),
    .X(_3237_));
 sky130_fd_sc_hd__clkbuf_1 _7448_ (.A(_3237_),
    .X(_0577_));
 sky130_fd_sc_hd__mux2_1 _7449_ (.A0(_3188_),
    .A1(net900),
    .S(_3236_),
    .X(_3238_));
 sky130_fd_sc_hd__clkbuf_1 _7450_ (.A(_3238_),
    .X(_0578_));
 sky130_fd_sc_hd__mux2_1 _7451_ (.A0(_3226_),
    .A1(net1212),
    .S(_3236_),
    .X(_3239_));
 sky130_fd_sc_hd__clkbuf_1 _7452_ (.A(_3239_),
    .X(_0579_));
 sky130_fd_sc_hd__mux2_1 _7453_ (.A0(_3228_),
    .A1(\gpio_configure[15][3] ),
    .S(_3236_),
    .X(_3240_));
 sky130_fd_sc_hd__clkbuf_1 _7454_ (.A(net854),
    .X(_0580_));
 sky130_fd_sc_hd__mux2_1 _7455_ (.A0(_3230_),
    .A1(net832),
    .S(_3236_),
    .X(_3241_));
 sky130_fd_sc_hd__clkbuf_1 _7456_ (.A(_3241_),
    .X(_0581_));
 sky130_fd_sc_hd__mux2_1 _7457_ (.A0(_3232_),
    .A1(net737),
    .S(_3236_),
    .X(_3242_));
 sky130_fd_sc_hd__clkbuf_1 _7458_ (.A(net738),
    .X(_0582_));
 sky130_fd_sc_hd__mux2_1 _7459_ (.A0(_3143_),
    .A1(net1265),
    .S(_3236_),
    .X(_3243_));
 sky130_fd_sc_hd__clkbuf_1 _7460_ (.A(net1266),
    .X(_0583_));
 sky130_fd_sc_hd__mux2_1 _7461_ (.A0(_3154_),
    .A1(net1026),
    .S(_3236_),
    .X(_3244_));
 sky130_fd_sc_hd__clkbuf_1 _7462_ (.A(net1027),
    .X(_0584_));
 sky130_fd_sc_hd__and2_1 _7463_ (.A(_0872_),
    .B(net525),
    .X(_3245_));
 sky130_fd_sc_hd__buf_6 _7464_ (.A(net567),
    .X(_3246_));
 sky130_fd_sc_hd__mux2_1 _7465_ (.A0(net1358),
    .A1(net939),
    .S(_3246_),
    .X(_3247_));
 sky130_fd_sc_hd__clkbuf_1 _7466_ (.A(_3247_),
    .X(_0585_));
 sky130_fd_sc_hd__mux2_1 _7467_ (.A0(net615),
    .A1(_1606_),
    .S(_3246_),
    .X(_3248_));
 sky130_fd_sc_hd__clkbuf_1 _7468_ (.A(_3248_),
    .X(_0586_));
 sky130_fd_sc_hd__mux2_1 _7469_ (.A0(net1072),
    .A1(_2051_),
    .S(_3246_),
    .X(_3249_));
 sky130_fd_sc_hd__clkbuf_1 _7470_ (.A(_3249_),
    .X(_0587_));
 sky130_fd_sc_hd__mux2_1 _7471_ (.A0(\gpio_configure[16][3] ),
    .A1(net552),
    .S(_3246_),
    .X(_3250_));
 sky130_fd_sc_hd__clkbuf_1 _7472_ (.A(net1592),
    .X(_0588_));
 sky130_fd_sc_hd__mux2_1 _7473_ (.A0(net840),
    .A1(_1668_),
    .S(_3246_),
    .X(_3251_));
 sky130_fd_sc_hd__clkbuf_1 _7474_ (.A(net1613),
    .X(_0589_));
 sky130_fd_sc_hd__mux2_1 _7475_ (.A0(net838),
    .A1(_1672_),
    .S(_3246_),
    .X(_3252_));
 sky130_fd_sc_hd__clkbuf_1 _7476_ (.A(net839),
    .X(_0590_));
 sky130_fd_sc_hd__mux2_1 _7477_ (.A0(net904),
    .A1(_1689_),
    .S(_3246_),
    .X(_3253_));
 sky130_fd_sc_hd__clkbuf_1 _7478_ (.A(_3253_),
    .X(_0591_));
 sky130_fd_sc_hd__mux2_1 _7479_ (.A0(net741),
    .A1(_1678_),
    .S(_3246_),
    .X(_3254_));
 sky130_fd_sc_hd__clkbuf_1 _7480_ (.A(_3254_),
    .X(_0592_));
 sky130_fd_sc_hd__nand2_8 _7481_ (.A(net376),
    .B(_3157_),
    .Y(_3255_));
 sky130_fd_sc_hd__mux2_1 _7482_ (.A0(_3156_),
    .A1(net1433),
    .S(_3255_),
    .X(_3256_));
 sky130_fd_sc_hd__clkbuf_1 _7483_ (.A(_3256_),
    .X(_0593_));
 sky130_fd_sc_hd__mux2_1 _7484_ (.A0(_3188_),
    .A1(net631),
    .S(_3255_),
    .X(_3257_));
 sky130_fd_sc_hd__clkbuf_1 _7485_ (.A(net632),
    .X(_0594_));
 sky130_fd_sc_hd__mux2_1 _7486_ (.A0(_3226_),
    .A1(net1228),
    .S(_3255_),
    .X(_3258_));
 sky130_fd_sc_hd__clkbuf_1 _7487_ (.A(_3258_),
    .X(_0595_));
 sky130_fd_sc_hd__mux2_1 _7488_ (.A0(_3228_),
    .A1(\gpio_configure[17][3] ),
    .S(_3255_),
    .X(_3259_));
 sky130_fd_sc_hd__clkbuf_1 _7489_ (.A(net853),
    .X(_0596_));
 sky130_fd_sc_hd__mux2_1 _7490_ (.A0(_3230_),
    .A1(net809),
    .S(_3255_),
    .X(_3260_));
 sky130_fd_sc_hd__clkbuf_1 _7491_ (.A(net810),
    .X(_0597_));
 sky130_fd_sc_hd__mux2_1 _7492_ (.A0(_3232_),
    .A1(net807),
    .S(_3255_),
    .X(_3261_));
 sky130_fd_sc_hd__clkbuf_1 _7493_ (.A(net808),
    .X(_0598_));
 sky130_fd_sc_hd__buf_2 _7494_ (.A(_1689_),
    .X(_3262_));
 sky130_fd_sc_hd__mux2_1 _7495_ (.A0(_3262_),
    .A1(net1260),
    .S(_3255_),
    .X(_3263_));
 sky130_fd_sc_hd__clkbuf_1 _7496_ (.A(net1261),
    .X(_0599_));
 sky130_fd_sc_hd__mux2_1 _7497_ (.A0(_3154_),
    .A1(net1070),
    .S(_3255_),
    .X(_3264_));
 sky130_fd_sc_hd__clkbuf_1 _7498_ (.A(net1071),
    .X(_0600_));
 sky130_fd_sc_hd__nand2_8 _7499_ (.A(net361),
    .B(_3157_),
    .Y(_3265_));
 sky130_fd_sc_hd__mux2_1 _7500_ (.A0(_3156_),
    .A1(net1434),
    .S(_3265_),
    .X(_3266_));
 sky130_fd_sc_hd__clkbuf_1 _7501_ (.A(_3266_),
    .X(_0601_));
 sky130_fd_sc_hd__mux2_1 _7502_ (.A0(_3188_),
    .A1(net633),
    .S(_3265_),
    .X(_3267_));
 sky130_fd_sc_hd__clkbuf_1 _7503_ (.A(net634),
    .X(_0602_));
 sky130_fd_sc_hd__mux2_1 _7504_ (.A0(_3226_),
    .A1(net1225),
    .S(_3265_),
    .X(_3268_));
 sky130_fd_sc_hd__clkbuf_1 _7505_ (.A(_3268_),
    .X(_0603_));
 sky130_fd_sc_hd__mux2_1 _7506_ (.A0(_3228_),
    .A1(\gpio_configure[18][3] ),
    .S(_3265_),
    .X(_3269_));
 sky130_fd_sc_hd__clkbuf_1 _7507_ (.A(net871),
    .X(_0604_));
 sky130_fd_sc_hd__mux2_1 _7508_ (.A0(_3230_),
    .A1(net789),
    .S(_3265_),
    .X(_3270_));
 sky130_fd_sc_hd__clkbuf_1 _7509_ (.A(net790),
    .X(_0605_));
 sky130_fd_sc_hd__mux2_1 _7510_ (.A0(_3232_),
    .A1(net768),
    .S(_3265_),
    .X(_3271_));
 sky130_fd_sc_hd__clkbuf_1 _7511_ (.A(net769),
    .X(_0606_));
 sky130_fd_sc_hd__mux2_1 _7512_ (.A0(_3262_),
    .A1(net1278),
    .S(_3265_),
    .X(_3272_));
 sky130_fd_sc_hd__clkbuf_1 _7513_ (.A(net1279),
    .X(_0607_));
 sky130_fd_sc_hd__clkbuf_4 _7514_ (.A(_1678_),
    .X(_3273_));
 sky130_fd_sc_hd__mux2_1 _7515_ (.A0(_3273_),
    .A1(net1142),
    .S(_3265_),
    .X(_3274_));
 sky130_fd_sc_hd__clkbuf_1 _7516_ (.A(net1143),
    .X(_0608_));
 sky130_fd_sc_hd__clkbuf_4 _7517_ (.A(_1597_),
    .X(_3275_));
 sky130_fd_sc_hd__buf_12 _7518_ (.A(_1601_),
    .X(_3276_));
 sky130_fd_sc_hd__nand2_8 _7519_ (.A(net386),
    .B(_3276_),
    .Y(_3277_));
 sky130_fd_sc_hd__mux2_1 _7520_ (.A0(_3275_),
    .A1(net1431),
    .S(_3277_),
    .X(_3278_));
 sky130_fd_sc_hd__clkbuf_1 _7521_ (.A(_3278_),
    .X(_0609_));
 sky130_fd_sc_hd__mux2_1 _7522_ (.A0(_3188_),
    .A1(net654),
    .S(_3277_),
    .X(_3279_));
 sky130_fd_sc_hd__clkbuf_1 _7523_ (.A(_3279_),
    .X(_0610_));
 sky130_fd_sc_hd__mux2_1 _7524_ (.A0(_3226_),
    .A1(net1219),
    .S(_3277_),
    .X(_3280_));
 sky130_fd_sc_hd__clkbuf_1 _7525_ (.A(_3280_),
    .X(_0611_));
 sky130_fd_sc_hd__mux2_1 _7526_ (.A0(_3228_),
    .A1(\gpio_configure[19][3] ),
    .S(_3277_),
    .X(_3281_));
 sky130_fd_sc_hd__clkbuf_1 _7527_ (.A(net848),
    .X(_0612_));
 sky130_fd_sc_hd__mux2_1 _7528_ (.A0(_3230_),
    .A1(net746),
    .S(_3277_),
    .X(_3282_));
 sky130_fd_sc_hd__clkbuf_1 _7529_ (.A(_3282_),
    .X(_0613_));
 sky130_fd_sc_hd__mux2_1 _7530_ (.A0(_3232_),
    .A1(net744),
    .S(_3277_),
    .X(_3283_));
 sky130_fd_sc_hd__clkbuf_1 _7531_ (.A(net745),
    .X(_0614_));
 sky130_fd_sc_hd__mux2_1 _7532_ (.A0(_3262_),
    .A1(net1236),
    .S(_3277_),
    .X(_3284_));
 sky130_fd_sc_hd__clkbuf_1 _7533_ (.A(net1237),
    .X(_0615_));
 sky130_fd_sc_hd__mux2_1 _7534_ (.A0(_3273_),
    .A1(net1104),
    .S(_3277_),
    .X(_3285_));
 sky130_fd_sc_hd__clkbuf_1 _7535_ (.A(net1105),
    .X(_0616_));
 sky130_fd_sc_hd__nand2_8 _7536_ (.A(net360),
    .B(_3276_),
    .Y(_3286_));
 sky130_fd_sc_hd__mux2_1 _7537_ (.A0(_3275_),
    .A1(net1435),
    .S(_3286_),
    .X(_3287_));
 sky130_fd_sc_hd__clkbuf_1 _7538_ (.A(_3287_),
    .X(_0617_));
 sky130_fd_sc_hd__mux2_1 _7539_ (.A0(_3188_),
    .A1(net667),
    .S(_3286_),
    .X(_3288_));
 sky130_fd_sc_hd__clkbuf_1 _7540_ (.A(_3288_),
    .X(_0618_));
 sky130_fd_sc_hd__mux2_1 _7541_ (.A0(_3226_),
    .A1(net1224),
    .S(_3286_),
    .X(_3289_));
 sky130_fd_sc_hd__clkbuf_1 _7542_ (.A(_3289_),
    .X(_0619_));
 sky130_fd_sc_hd__mux2_1 _7543_ (.A0(_3228_),
    .A1(\gpio_configure[20][3] ),
    .S(_3286_),
    .X(_3290_));
 sky130_fd_sc_hd__clkbuf_1 _7544_ (.A(net855),
    .X(_0620_));
 sky130_fd_sc_hd__mux2_1 _7545_ (.A0(_3230_),
    .A1(net773),
    .S(_3286_),
    .X(_3291_));
 sky130_fd_sc_hd__clkbuf_1 _7546_ (.A(_3291_),
    .X(_0621_));
 sky130_fd_sc_hd__mux2_1 _7547_ (.A0(_3232_),
    .A1(net742),
    .S(_3286_),
    .X(_3292_));
 sky130_fd_sc_hd__clkbuf_1 _7548_ (.A(net743),
    .X(_0622_));
 sky130_fd_sc_hd__mux2_1 _7549_ (.A0(_3262_),
    .A1(net1252),
    .S(_3286_),
    .X(_3293_));
 sky130_fd_sc_hd__clkbuf_1 _7550_ (.A(net1253),
    .X(_0623_));
 sky130_fd_sc_hd__mux2_1 _7551_ (.A0(_3273_),
    .A1(net1101),
    .S(_3286_),
    .X(_3294_));
 sky130_fd_sc_hd__clkbuf_1 _7552_ (.A(net1102),
    .X(_0624_));
 sky130_fd_sc_hd__nand2_8 _7553_ (.A(net365),
    .B(_3276_),
    .Y(_3295_));
 sky130_fd_sc_hd__mux2_1 _7554_ (.A0(_3275_),
    .A1(net1395),
    .S(_3295_),
    .X(_3296_));
 sky130_fd_sc_hd__clkbuf_1 _7555_ (.A(_3296_),
    .X(_0625_));
 sky130_fd_sc_hd__clkbuf_2 _7556_ (.A(net543),
    .X(_3297_));
 sky130_fd_sc_hd__mux2_1 _7557_ (.A0(_3297_),
    .A1(\gpio_configure[21][1] ),
    .S(net605),
    .X(_3298_));
 sky130_fd_sc_hd__clkbuf_1 _7558_ (.A(net606),
    .X(_0626_));
 sky130_fd_sc_hd__mux2_1 _7559_ (.A0(_3226_),
    .A1(net1229),
    .S(_3295_),
    .X(_3299_));
 sky130_fd_sc_hd__clkbuf_1 _7560_ (.A(_3299_),
    .X(_0627_));
 sky130_fd_sc_hd__mux2_1 _7561_ (.A0(_3228_),
    .A1(\gpio_configure[21][3] ),
    .S(net605),
    .X(_3300_));
 sky130_fd_sc_hd__clkbuf_1 _7562_ (.A(net849),
    .X(_0628_));
 sky130_fd_sc_hd__mux2_1 _7563_ (.A0(_3230_),
    .A1(net764),
    .S(_3295_),
    .X(_3301_));
 sky130_fd_sc_hd__clkbuf_1 _7564_ (.A(net1669),
    .X(_0629_));
 sky130_fd_sc_hd__mux2_1 _7565_ (.A0(_3232_),
    .A1(net739),
    .S(_3295_),
    .X(_3302_));
 sky130_fd_sc_hd__clkbuf_1 _7566_ (.A(net740),
    .X(_0630_));
 sky130_fd_sc_hd__mux2_1 _7567_ (.A0(_3262_),
    .A1(net1262),
    .S(_3295_),
    .X(_3303_));
 sky130_fd_sc_hd__clkbuf_1 _7568_ (.A(net1263),
    .X(_0631_));
 sky130_fd_sc_hd__mux2_1 _7569_ (.A0(_3273_),
    .A1(net1347),
    .S(_3295_),
    .X(_3304_));
 sky130_fd_sc_hd__clkbuf_1 _7570_ (.A(_3304_),
    .X(_0632_));
 sky130_fd_sc_hd__nand2_8 _7571_ (.A(net384),
    .B(_3276_),
    .Y(_3305_));
 sky130_fd_sc_hd__mux2_1 _7572_ (.A0(_3275_),
    .A1(net1410),
    .S(net584),
    .X(_3306_));
 sky130_fd_sc_hd__clkbuf_1 _7573_ (.A(_3306_),
    .X(_0633_));
 sky130_fd_sc_hd__mux2_1 _7574_ (.A0(_3297_),
    .A1(net1549),
    .S(net584),
    .X(_3307_));
 sky130_fd_sc_hd__clkbuf_1 _7575_ (.A(_3307_),
    .X(_0634_));
 sky130_fd_sc_hd__mux2_1 _7576_ (.A0(_3226_),
    .A1(net1220),
    .S(net584),
    .X(_3308_));
 sky130_fd_sc_hd__clkbuf_1 _7577_ (.A(_3308_),
    .X(_0635_));
 sky130_fd_sc_hd__mux2_1 _7578_ (.A0(_3228_),
    .A1(\gpio_configure[22][3] ),
    .S(net584),
    .X(_3309_));
 sky130_fd_sc_hd__clkbuf_1 _7579_ (.A(net1593),
    .X(_0636_));
 sky130_fd_sc_hd__mux2_1 _7580_ (.A0(_3230_),
    .A1(net770),
    .S(net584),
    .X(_3310_));
 sky130_fd_sc_hd__clkbuf_1 _7581_ (.A(_3310_),
    .X(_0637_));
 sky130_fd_sc_hd__mux2_1 _7582_ (.A0(_3232_),
    .A1(net754),
    .S(net584),
    .X(_3311_));
 sky130_fd_sc_hd__clkbuf_1 _7583_ (.A(net755),
    .X(_0638_));
 sky130_fd_sc_hd__mux2_1 _7584_ (.A0(_3262_),
    .A1(net1283),
    .S(net584),
    .X(_3312_));
 sky130_fd_sc_hd__clkbuf_1 _7585_ (.A(_3312_),
    .X(_0639_));
 sky130_fd_sc_hd__mux2_1 _7586_ (.A0(_3273_),
    .A1(net1152),
    .S(net584),
    .X(_3313_));
 sky130_fd_sc_hd__clkbuf_1 _7587_ (.A(net1153),
    .X(_0640_));
 sky130_fd_sc_hd__nand2_8 _7588_ (.A(net373),
    .B(_3276_),
    .Y(_3314_));
 sky130_fd_sc_hd__mux2_1 _7589_ (.A0(_3275_),
    .A1(net1437),
    .S(net581),
    .X(_3315_));
 sky130_fd_sc_hd__clkbuf_1 _7590_ (.A(_3315_),
    .X(_0641_));
 sky130_fd_sc_hd__mux2_1 _7591_ (.A0(_3297_),
    .A1(net1551),
    .S(net581),
    .X(_3316_));
 sky130_fd_sc_hd__clkbuf_1 _7592_ (.A(_3316_),
    .X(_0642_));
 sky130_fd_sc_hd__mux2_1 _7593_ (.A0(_3226_),
    .A1(net1217),
    .S(net581),
    .X(_3317_));
 sky130_fd_sc_hd__clkbuf_1 _7594_ (.A(_3317_),
    .X(_0643_));
 sky130_fd_sc_hd__mux2_1 _7595_ (.A0(_3228_),
    .A1(\gpio_configure[23][3] ),
    .S(net581),
    .X(_3318_));
 sky130_fd_sc_hd__clkbuf_1 _7596_ (.A(net1595),
    .X(_0644_));
 sky130_fd_sc_hd__mux2_1 _7597_ (.A0(_3230_),
    .A1(net776),
    .S(net581),
    .X(_3319_));
 sky130_fd_sc_hd__clkbuf_1 _7598_ (.A(_3319_),
    .X(_0645_));
 sky130_fd_sc_hd__mux2_1 _7599_ (.A0(_3232_),
    .A1(net733),
    .S(net581),
    .X(_3320_));
 sky130_fd_sc_hd__clkbuf_1 _7600_ (.A(_3320_),
    .X(_0646_));
 sky130_fd_sc_hd__mux2_1 _7601_ (.A0(_3262_),
    .A1(net1233),
    .S(net581),
    .X(_3321_));
 sky130_fd_sc_hd__clkbuf_1 _7602_ (.A(_3321_),
    .X(_0647_));
 sky130_fd_sc_hd__mux2_1 _7603_ (.A0(_3273_),
    .A1(net1090),
    .S(net581),
    .X(_3322_));
 sky130_fd_sc_hd__clkbuf_1 _7604_ (.A(net1091),
    .X(_0648_));
 sky130_fd_sc_hd__and2_1 _7605_ (.A(_0890_),
    .B(net525),
    .X(_3323_));
 sky130_fd_sc_hd__buf_6 _7606_ (.A(net560),
    .X(_3324_));
 sky130_fd_sc_hd__mux2_1 _7607_ (.A0(net1384),
    .A1(_1731_),
    .S(_3324_),
    .X(_3325_));
 sky130_fd_sc_hd__clkbuf_1 _7608_ (.A(net1385),
    .X(_0649_));
 sky130_fd_sc_hd__mux2_1 _7609_ (.A0(net620),
    .A1(_1606_),
    .S(_3324_),
    .X(_3326_));
 sky130_fd_sc_hd__clkbuf_1 _7610_ (.A(_3326_),
    .X(_0650_));
 sky130_fd_sc_hd__mux2_1 _7611_ (.A0(net1221),
    .A1(_2051_),
    .S(_3324_),
    .X(_3327_));
 sky130_fd_sc_hd__clkbuf_1 _7612_ (.A(_3327_),
    .X(_0651_));
 sky130_fd_sc_hd__mux2_1 _7613_ (.A0(\gpio_configure[24][3] ),
    .A1(net552),
    .S(_3324_),
    .X(_3328_));
 sky130_fd_sc_hd__clkbuf_1 _7614_ (.A(net1591),
    .X(_0652_));
 sky130_fd_sc_hd__mux2_1 _7615_ (.A0(net816),
    .A1(_1668_),
    .S(_3324_),
    .X(_3329_));
 sky130_fd_sc_hd__clkbuf_1 _7616_ (.A(net1604),
    .X(_0653_));
 sky130_fd_sc_hd__mux2_1 _7617_ (.A0(net811),
    .A1(_1672_),
    .S(_3324_),
    .X(_3330_));
 sky130_fd_sc_hd__clkbuf_1 _7618_ (.A(net812),
    .X(_0654_));
 sky130_fd_sc_hd__mux2_1 _7619_ (.A0(net892),
    .A1(_1689_),
    .S(_3324_),
    .X(_3331_));
 sky130_fd_sc_hd__clkbuf_1 _7620_ (.A(_3331_),
    .X(_0655_));
 sky130_fd_sc_hd__mux2_1 _7621_ (.A0(net730),
    .A1(_1678_),
    .S(_3324_),
    .X(_3332_));
 sky130_fd_sc_hd__clkbuf_1 _7622_ (.A(_3332_),
    .X(_0656_));
 sky130_fd_sc_hd__nand2_8 _7623_ (.A(net380),
    .B(_3276_),
    .Y(_3333_));
 sky130_fd_sc_hd__mux2_1 _7624_ (.A0(_3275_),
    .A1(net1393),
    .S(_3333_),
    .X(_3334_));
 sky130_fd_sc_hd__clkbuf_1 _7625_ (.A(_3334_),
    .X(_0657_));
 sky130_fd_sc_hd__mux2_1 _7626_ (.A0(_3297_),
    .A1(net596),
    .S(_3333_),
    .X(_3335_));
 sky130_fd_sc_hd__clkbuf_1 _7627_ (.A(net597),
    .X(_0658_));
 sky130_fd_sc_hd__mux2_1 _7628_ (.A0(_3226_),
    .A1(net914),
    .S(_3333_),
    .X(_3336_));
 sky130_fd_sc_hd__clkbuf_1 _7629_ (.A(net915),
    .X(_0659_));
 sky130_fd_sc_hd__mux2_1 _7630_ (.A0(_3228_),
    .A1(\gpio_configure[25][3] ),
    .S(_3333_),
    .X(_3337_));
 sky130_fd_sc_hd__clkbuf_1 _7631_ (.A(net846),
    .X(_0660_));
 sky130_fd_sc_hd__mux2_1 _7632_ (.A0(_3230_),
    .A1(net760),
    .S(_3333_),
    .X(_3338_));
 sky130_fd_sc_hd__clkbuf_1 _7633_ (.A(net761),
    .X(_0661_));
 sky130_fd_sc_hd__mux2_1 _7634_ (.A0(_3232_),
    .A1(net735),
    .S(_3333_),
    .X(_3339_));
 sky130_fd_sc_hd__clkbuf_1 _7635_ (.A(net736),
    .X(_0662_));
 sky130_fd_sc_hd__mux2_1 _7636_ (.A0(_3262_),
    .A1(net1241),
    .S(_3333_),
    .X(_3340_));
 sky130_fd_sc_hd__clkbuf_1 _7637_ (.A(net1242),
    .X(_0663_));
 sky130_fd_sc_hd__mux2_1 _7638_ (.A0(_3273_),
    .A1(net1171),
    .S(_3333_),
    .X(_3341_));
 sky130_fd_sc_hd__clkbuf_1 _7639_ (.A(net1172),
    .X(_0664_));
 sky130_fd_sc_hd__nand2_8 _7640_ (.A(net392),
    .B(_3276_),
    .Y(_3342_));
 sky130_fd_sc_hd__mux2_1 _7641_ (.A0(_3275_),
    .A1(net1430),
    .S(net590),
    .X(_3343_));
 sky130_fd_sc_hd__clkbuf_1 _7642_ (.A(_3343_),
    .X(_0665_));
 sky130_fd_sc_hd__mux2_1 _7643_ (.A0(_3297_),
    .A1(net1550),
    .S(net590),
    .X(_3344_));
 sky130_fd_sc_hd__clkbuf_1 _7644_ (.A(_3344_),
    .X(_0666_));
 sky130_fd_sc_hd__buf_6 _7645_ (.A(_1610_),
    .X(_3345_));
 sky130_fd_sc_hd__mux2_1 _7646_ (.A0(_3345_),
    .A1(net1127),
    .S(net590),
    .X(_3346_));
 sky130_fd_sc_hd__clkbuf_1 _7647_ (.A(_3346_),
    .X(_0667_));
 sky130_fd_sc_hd__buf_2 _7648_ (.A(_1614_),
    .X(_3347_));
 sky130_fd_sc_hd__mux2_1 _7649_ (.A0(_3347_),
    .A1(\gpio_configure[26][3] ),
    .S(net590),
    .X(_3348_));
 sky130_fd_sc_hd__clkbuf_1 _7650_ (.A(net1594),
    .X(_0668_));
 sky130_fd_sc_hd__buf_4 _7651_ (.A(net530),
    .X(_3349_));
 sky130_fd_sc_hd__mux2_1 _7652_ (.A0(_3349_),
    .A1(net872),
    .S(net590),
    .X(_3350_));
 sky130_fd_sc_hd__clkbuf_1 _7653_ (.A(_3350_),
    .X(_0669_));
 sky130_fd_sc_hd__buf_4 _7654_ (.A(net521),
    .X(_3351_));
 sky130_fd_sc_hd__mux2_1 _7655_ (.A0(_3351_),
    .A1(net747),
    .S(net590),
    .X(_3352_));
 sky130_fd_sc_hd__clkbuf_1 _7656_ (.A(_3352_),
    .X(_0670_));
 sky130_fd_sc_hd__mux2_1 _7657_ (.A0(_3262_),
    .A1(net1238),
    .S(net590),
    .X(_3353_));
 sky130_fd_sc_hd__clkbuf_1 _7658_ (.A(_3353_),
    .X(_0671_));
 sky130_fd_sc_hd__mux2_1 _7659_ (.A0(_3273_),
    .A1(net1163),
    .S(net590),
    .X(_3354_));
 sky130_fd_sc_hd__clkbuf_1 _7660_ (.A(_3354_),
    .X(_0672_));
 sky130_fd_sc_hd__nand2_8 _7661_ (.A(net388),
    .B(_3276_),
    .Y(_3355_));
 sky130_fd_sc_hd__mux2_1 _7662_ (.A0(_3275_),
    .A1(net1441),
    .S(_3355_),
    .X(_3356_));
 sky130_fd_sc_hd__clkbuf_1 _7663_ (.A(_3356_),
    .X(_0673_));
 sky130_fd_sc_hd__mux2_1 _7664_ (.A0(_3297_),
    .A1(net598),
    .S(_3355_),
    .X(_3357_));
 sky130_fd_sc_hd__clkbuf_1 _7665_ (.A(net599),
    .X(_0674_));
 sky130_fd_sc_hd__mux2_1 _7666_ (.A0(_3345_),
    .A1(net920),
    .S(_3355_),
    .X(_3358_));
 sky130_fd_sc_hd__clkbuf_1 _7667_ (.A(net921),
    .X(_0675_));
 sky130_fd_sc_hd__mux2_1 _7668_ (.A0(_3347_),
    .A1(\gpio_configure[27][3] ),
    .S(_3355_),
    .X(_3359_));
 sky130_fd_sc_hd__clkbuf_1 _7669_ (.A(net888),
    .X(_0676_));
 sky130_fd_sc_hd__mux2_1 _7670_ (.A0(_3349_),
    .A1(net879),
    .S(_3355_),
    .X(_3360_));
 sky130_fd_sc_hd__clkbuf_1 _7671_ (.A(_3360_),
    .X(_0677_));
 sky130_fd_sc_hd__mux2_1 _7672_ (.A0(_3351_),
    .A1(net731),
    .S(_3355_),
    .X(_3361_));
 sky130_fd_sc_hd__clkbuf_1 _7673_ (.A(net732),
    .X(_0678_));
 sky130_fd_sc_hd__mux2_1 _7674_ (.A0(_3262_),
    .A1(net1246),
    .S(_3355_),
    .X(_3362_));
 sky130_fd_sc_hd__clkbuf_1 _7675_ (.A(net1247),
    .X(_0679_));
 sky130_fd_sc_hd__mux2_1 _7676_ (.A0(_3273_),
    .A1(net1109),
    .S(_3355_),
    .X(_3363_));
 sky130_fd_sc_hd__clkbuf_1 _7677_ (.A(net1110),
    .X(_0680_));
 sky130_fd_sc_hd__nand2_8 _7678_ (.A(net381),
    .B(_3276_),
    .Y(_3364_));
 sky130_fd_sc_hd__mux2_1 _7679_ (.A0(_3275_),
    .A1(net1425),
    .S(_3364_),
    .X(_3365_));
 sky130_fd_sc_hd__clkbuf_1 _7680_ (.A(_3365_),
    .X(_0681_));
 sky130_fd_sc_hd__mux2_1 _7681_ (.A0(_3297_),
    .A1(net602),
    .S(_3364_),
    .X(_3366_));
 sky130_fd_sc_hd__clkbuf_1 _7682_ (.A(net603),
    .X(_0682_));
 sky130_fd_sc_hd__mux2_1 _7683_ (.A0(_3345_),
    .A1(net932),
    .S(_3364_),
    .X(_3367_));
 sky130_fd_sc_hd__clkbuf_1 _7684_ (.A(net933),
    .X(_0683_));
 sky130_fd_sc_hd__mux2_1 _7685_ (.A0(_3347_),
    .A1(\gpio_configure[28][3] ),
    .S(_3364_),
    .X(_3368_));
 sky130_fd_sc_hd__clkbuf_1 _7686_ (.A(net877),
    .X(_0684_));
 sky130_fd_sc_hd__mux2_1 _7687_ (.A0(_3349_),
    .A1(net878),
    .S(_3364_),
    .X(_3369_));
 sky130_fd_sc_hd__clkbuf_1 _7688_ (.A(_3369_),
    .X(_0685_));
 sky130_fd_sc_hd__mux2_1 _7689_ (.A0(_3351_),
    .A1(net756),
    .S(_3364_),
    .X(_3370_));
 sky130_fd_sc_hd__clkbuf_1 _7690_ (.A(net757),
    .X(_0686_));
 sky130_fd_sc_hd__mux2_1 _7691_ (.A0(_1675_),
    .A1(net707),
    .S(_3364_),
    .X(_3371_));
 sky130_fd_sc_hd__clkbuf_1 _7692_ (.A(net708),
    .X(_0687_));
 sky130_fd_sc_hd__mux2_1 _7693_ (.A0(_3273_),
    .A1(net1092),
    .S(_3364_),
    .X(_3372_));
 sky130_fd_sc_hd__clkbuf_1 _7694_ (.A(net1093),
    .X(_0688_));
 sky130_fd_sc_hd__nand2_8 _7695_ (.A(net390),
    .B(_3276_),
    .Y(_3373_));
 sky130_fd_sc_hd__mux2_1 _7696_ (.A0(_3275_),
    .A1(net1408),
    .S(_3373_),
    .X(_3374_));
 sky130_fd_sc_hd__clkbuf_1 _7697_ (.A(_3374_),
    .X(_0689_));
 sky130_fd_sc_hd__mux2_1 _7698_ (.A0(_3297_),
    .A1(net594),
    .S(_3373_),
    .X(_3375_));
 sky130_fd_sc_hd__clkbuf_1 _7699_ (.A(net595),
    .X(_0690_));
 sky130_fd_sc_hd__mux2_1 _7700_ (.A0(_3345_),
    .A1(net1230),
    .S(_3373_),
    .X(_3376_));
 sky130_fd_sc_hd__clkbuf_1 _7701_ (.A(_3376_),
    .X(_0691_));
 sky130_fd_sc_hd__mux2_1 _7702_ (.A0(_3347_),
    .A1(\gpio_configure[29][3] ),
    .S(_3373_),
    .X(_3377_));
 sky130_fd_sc_hd__clkbuf_1 _7703_ (.A(net882),
    .X(_0692_));
 sky130_fd_sc_hd__mux2_1 _7704_ (.A0(_3349_),
    .A1(net876),
    .S(_3373_),
    .X(_3378_));
 sky130_fd_sc_hd__clkbuf_1 _7705_ (.A(_3378_),
    .X(_0693_));
 sky130_fd_sc_hd__mux2_1 _7706_ (.A0(_3351_),
    .A1(net718),
    .S(_3373_),
    .X(_3379_));
 sky130_fd_sc_hd__clkbuf_1 _7707_ (.A(net719),
    .X(_0694_));
 sky130_fd_sc_hd__mux2_1 _7708_ (.A0(_1675_),
    .A1(net694),
    .S(_3373_),
    .X(_3380_));
 sky130_fd_sc_hd__clkbuf_1 _7709_ (.A(net695),
    .X(_0695_));
 sky130_fd_sc_hd__mux2_1 _7710_ (.A0(_1679_),
    .A1(net1149),
    .S(_3373_),
    .X(_3381_));
 sky130_fd_sc_hd__clkbuf_1 _7711_ (.A(net1150),
    .X(_0696_));
 sky130_fd_sc_hd__nand2_8 _7712_ (.A(net391),
    .B(_1912_),
    .Y(_3382_));
 sky130_fd_sc_hd__mux2_1 _7713_ (.A0(_1658_),
    .A1(net1394),
    .S(net601),
    .X(_3383_));
 sky130_fd_sc_hd__clkbuf_1 _7714_ (.A(_3383_),
    .X(_0697_));
 sky130_fd_sc_hd__mux2_1 _7715_ (.A0(_3297_),
    .A1(net1552),
    .S(net601),
    .X(_3384_));
 sky130_fd_sc_hd__clkbuf_1 _7716_ (.A(_3384_),
    .X(_0698_));
 sky130_fd_sc_hd__mux2_1 _7717_ (.A0(_3345_),
    .A1(net924),
    .S(net601),
    .X(_3385_));
 sky130_fd_sc_hd__clkbuf_1 _7718_ (.A(_3385_),
    .X(_0699_));
 sky130_fd_sc_hd__mux2_1 _7719_ (.A0(_3347_),
    .A1(\gpio_configure[30][3] ),
    .S(net601),
    .X(_3386_));
 sky130_fd_sc_hd__clkbuf_1 _7720_ (.A(net1597),
    .X(_0700_));
 sky130_fd_sc_hd__mux2_1 _7721_ (.A0(_3349_),
    .A1(net860),
    .S(_3382_),
    .X(_3387_));
 sky130_fd_sc_hd__clkbuf_1 _7722_ (.A(_3387_),
    .X(_0701_));
 sky130_fd_sc_hd__mux2_1 _7723_ (.A0(_3351_),
    .A1(net758),
    .S(_3382_),
    .X(_3388_));
 sky130_fd_sc_hd__clkbuf_1 _7724_ (.A(net759),
    .X(_0702_));
 sky130_fd_sc_hd__mux2_1 _7725_ (.A0(_1675_),
    .A1(net702),
    .S(net601),
    .X(_3389_));
 sky130_fd_sc_hd__clkbuf_1 _7726_ (.A(_3389_),
    .X(_0703_));
 sky130_fd_sc_hd__mux2_1 _7727_ (.A0(_1679_),
    .A1(net1161),
    .S(net601),
    .X(_3390_));
 sky130_fd_sc_hd__clkbuf_1 _7728_ (.A(net1162),
    .X(_0704_));
 sky130_fd_sc_hd__nand2_8 _7729_ (.A(_0949_),
    .B(_1912_),
    .Y(_3391_));
 sky130_fd_sc_hd__mux2_1 _7730_ (.A0(_1658_),
    .A1(net1406),
    .S(net592),
    .X(_3392_));
 sky130_fd_sc_hd__clkbuf_1 _7731_ (.A(_3392_),
    .X(_0705_));
 sky130_fd_sc_hd__mux2_1 _7732_ (.A0(_3297_),
    .A1(\gpio_configure[31][1] ),
    .S(net592),
    .X(_3393_));
 sky130_fd_sc_hd__clkbuf_1 _7733_ (.A(net593),
    .X(_0706_));
 sky130_fd_sc_hd__mux2_1 _7734_ (.A0(_3345_),
    .A1(net1243),
    .S(net592),
    .X(_3394_));
 sky130_fd_sc_hd__clkbuf_1 _7735_ (.A(_3394_),
    .X(_0707_));
 sky130_fd_sc_hd__mux2_1 _7736_ (.A0(_3347_),
    .A1(\gpio_configure[31][3] ),
    .S(net592),
    .X(_3395_));
 sky130_fd_sc_hd__clkbuf_1 _7737_ (.A(net1596),
    .X(_0708_));
 sky130_fd_sc_hd__mux2_1 _7738_ (.A0(_3349_),
    .A1(net887),
    .S(net592),
    .X(_3396_));
 sky130_fd_sc_hd__clkbuf_1 _7739_ (.A(_3396_),
    .X(_0709_));
 sky130_fd_sc_hd__mux2_1 _7740_ (.A0(_3351_),
    .A1(net684),
    .S(net592),
    .X(_3397_));
 sky130_fd_sc_hd__clkbuf_1 _7741_ (.A(net685),
    .X(_0710_));
 sky130_fd_sc_hd__mux2_1 _7742_ (.A0(_1675_),
    .A1(net841),
    .S(net592),
    .X(_3398_));
 sky130_fd_sc_hd__clkbuf_1 _7743_ (.A(_3398_),
    .X(_0711_));
 sky130_fd_sc_hd__mux2_1 _7744_ (.A0(_1679_),
    .A1(net1296),
    .S(net592),
    .X(_3399_));
 sky130_fd_sc_hd__clkbuf_1 _7745_ (.A(net1297),
    .X(_0712_));
 sky130_fd_sc_hd__and2_1 _7746_ (.A(_0898_),
    .B(net525),
    .X(_3400_));
 sky130_fd_sc_hd__buf_6 _7747_ (.A(_3400_),
    .X(_3401_));
 sky130_fd_sc_hd__mux2_1 _7748_ (.A0(net1379),
    .A1(_1731_),
    .S(_3401_),
    .X(_3402_));
 sky130_fd_sc_hd__clkbuf_1 _7749_ (.A(net1380),
    .X(_0713_));
 sky130_fd_sc_hd__mux2_1 _7750_ (.A0(net681),
    .A1(_1606_),
    .S(_3401_),
    .X(_3403_));
 sky130_fd_sc_hd__clkbuf_1 _7751_ (.A(_3403_),
    .X(_0714_));
 sky130_fd_sc_hd__mux2_1 _7752_ (.A0(net1009),
    .A1(_2051_),
    .S(_3401_),
    .X(_3404_));
 sky130_fd_sc_hd__clkbuf_1 _7753_ (.A(net1010),
    .X(_0715_));
 sky130_fd_sc_hd__mux2_1 _7754_ (.A0(\gpio_configure[32][3] ),
    .A1(net552),
    .S(_3401_),
    .X(_3405_));
 sky130_fd_sc_hd__clkbuf_1 _7755_ (.A(net553),
    .X(_0716_));
 sky130_fd_sc_hd__mux2_1 _7756_ (.A0(net623),
    .A1(_1668_),
    .S(_3401_),
    .X(_3406_));
 sky130_fd_sc_hd__clkbuf_1 _7757_ (.A(net624),
    .X(_0717_));
 sky130_fd_sc_hd__mux2_1 _7758_ (.A0(net797),
    .A1(_1672_),
    .S(_3401_),
    .X(_3407_));
 sky130_fd_sc_hd__clkbuf_1 _7759_ (.A(net798),
    .X(_0718_));
 sky130_fd_sc_hd__mux2_1 _7760_ (.A0(net885),
    .A1(_1689_),
    .S(_3401_),
    .X(_3408_));
 sky130_fd_sc_hd__clkbuf_1 _7761_ (.A(net886),
    .X(_0719_));
 sky130_fd_sc_hd__mux2_1 _7762_ (.A0(net715),
    .A1(_1678_),
    .S(_3401_),
    .X(_3409_));
 sky130_fd_sc_hd__clkbuf_1 _7763_ (.A(net716),
    .X(_0720_));
 sky130_fd_sc_hd__nand2_8 _7764_ (.A(_0957_),
    .B(_1912_),
    .Y(_3410_));
 sky130_fd_sc_hd__mux2_1 _7765_ (.A0(_1658_),
    .A1(net1332),
    .S(_3410_),
    .X(_3411_));
 sky130_fd_sc_hd__clkbuf_1 _7766_ (.A(_3411_),
    .X(_0721_));
 sky130_fd_sc_hd__mux2_1 _7767_ (.A0(_1662_),
    .A1(net1005),
    .S(_3410_),
    .X(_3412_));
 sky130_fd_sc_hd__clkbuf_1 _7768_ (.A(_3412_),
    .X(_0722_));
 sky130_fd_sc_hd__mux2_1 _7769_ (.A0(_3345_),
    .A1(net994),
    .S(_3410_),
    .X(_3413_));
 sky130_fd_sc_hd__clkbuf_1 _7770_ (.A(net995),
    .X(_0723_));
 sky130_fd_sc_hd__mux2_1 _7771_ (.A0(_3347_),
    .A1(\gpio_configure[33][3] ),
    .S(_3410_),
    .X(_3414_));
 sky130_fd_sc_hd__clkbuf_1 _7772_ (.A(net870),
    .X(_0724_));
 sky130_fd_sc_hd__mux2_1 _7773_ (.A0(_3349_),
    .A1(net698),
    .S(_3410_),
    .X(_3415_));
 sky130_fd_sc_hd__clkbuf_1 _7774_ (.A(net699),
    .X(_0725_));
 sky130_fd_sc_hd__mux2_1 _7775_ (.A0(_3351_),
    .A1(net750),
    .S(_3410_),
    .X(_3416_));
 sky130_fd_sc_hd__clkbuf_1 _7776_ (.A(net751),
    .X(_0726_));
 sky130_fd_sc_hd__mux2_1 _7777_ (.A0(_1675_),
    .A1(net805),
    .S(_3410_),
    .X(_3417_));
 sky130_fd_sc_hd__clkbuf_1 _7778_ (.A(net806),
    .X(_0727_));
 sky130_fd_sc_hd__mux2_1 _7779_ (.A0(_1679_),
    .A1(net1159),
    .S(_3410_),
    .X(_3418_));
 sky130_fd_sc_hd__clkbuf_1 _7780_ (.A(net1160),
    .X(_0728_));
 sky130_fd_sc_hd__nand2_8 _7781_ (.A(net364),
    .B(_1912_),
    .Y(_3419_));
 sky130_fd_sc_hd__mux2_1 _7782_ (.A0(_1658_),
    .A1(net1442),
    .S(_3419_),
    .X(_3420_));
 sky130_fd_sc_hd__clkbuf_1 _7783_ (.A(_3420_),
    .X(_0729_));
 sky130_fd_sc_hd__mux2_1 _7784_ (.A0(_1662_),
    .A1(net982),
    .S(_3419_),
    .X(_3421_));
 sky130_fd_sc_hd__clkbuf_1 _7785_ (.A(_3421_),
    .X(_0730_));
 sky130_fd_sc_hd__mux2_1 _7786_ (.A0(_3345_),
    .A1(net1016),
    .S(_3419_),
    .X(_3422_));
 sky130_fd_sc_hd__clkbuf_1 _7787_ (.A(net1017),
    .X(_0731_));
 sky130_fd_sc_hd__mux2_1 _7788_ (.A0(_3347_),
    .A1(\gpio_configure[34][3] ),
    .S(_3419_),
    .X(_3423_));
 sky130_fd_sc_hd__clkbuf_1 _7789_ (.A(net868),
    .X(_0732_));
 sky130_fd_sc_hd__mux2_1 _7790_ (.A0(_3349_),
    .A1(net690),
    .S(_3419_),
    .X(_3424_));
 sky130_fd_sc_hd__clkbuf_1 _7791_ (.A(net691),
    .X(_0733_));
 sky130_fd_sc_hd__mux2_1 _7792_ (.A0(_3351_),
    .A1(net682),
    .S(_3419_),
    .X(_3425_));
 sky130_fd_sc_hd__clkbuf_1 _7793_ (.A(net683),
    .X(_0734_));
 sky130_fd_sc_hd__mux2_1 _7794_ (.A0(_1675_),
    .A1(net830),
    .S(_3419_),
    .X(_3426_));
 sky130_fd_sc_hd__clkbuf_1 _7795_ (.A(net831),
    .X(_0735_));
 sky130_fd_sc_hd__mux2_1 _7796_ (.A0(_1679_),
    .A1(net1191),
    .S(_3419_),
    .X(_3427_));
 sky130_fd_sc_hd__clkbuf_1 _7797_ (.A(net1192),
    .X(_0736_));
 sky130_fd_sc_hd__nand2_8 _7798_ (.A(net379),
    .B(net527),
    .Y(_3428_));
 sky130_fd_sc_hd__mux2_1 _7799_ (.A0(_1658_),
    .A1(net1427),
    .S(_3428_),
    .X(_3429_));
 sky130_fd_sc_hd__clkbuf_1 _7800_ (.A(_3429_),
    .X(_0737_));
 sky130_fd_sc_hd__mux2_1 _7801_ (.A0(_1662_),
    .A1(net1023),
    .S(_3428_),
    .X(_3430_));
 sky130_fd_sc_hd__clkbuf_1 _7802_ (.A(_3430_),
    .X(_0738_));
 sky130_fd_sc_hd__mux2_1 _7803_ (.A0(_3345_),
    .A1(net1231),
    .S(_3428_),
    .X(_3431_));
 sky130_fd_sc_hd__clkbuf_1 _7804_ (.A(_3431_),
    .X(_0739_));
 sky130_fd_sc_hd__mux2_1 _7805_ (.A0(_3347_),
    .A1(\gpio_configure[35][3] ),
    .S(_3428_),
    .X(_3432_));
 sky130_fd_sc_hd__clkbuf_1 _7806_ (.A(net857),
    .X(_0740_));
 sky130_fd_sc_hd__mux2_1 _7807_ (.A0(_3349_),
    .A1(net856),
    .S(_3428_),
    .X(_3433_));
 sky130_fd_sc_hd__clkbuf_1 _7808_ (.A(_3433_),
    .X(_0741_));
 sky130_fd_sc_hd__mux2_1 _7809_ (.A0(_3351_),
    .A1(net726),
    .S(_3428_),
    .X(_3434_));
 sky130_fd_sc_hd__clkbuf_1 _7810_ (.A(net727),
    .X(_0742_));
 sky130_fd_sc_hd__mux2_1 _7811_ (.A0(_1675_),
    .A1(net700),
    .S(_3428_),
    .X(_3435_));
 sky130_fd_sc_hd__clkbuf_1 _7812_ (.A(net701),
    .X(_0743_));
 sky130_fd_sc_hd__mux2_1 _7813_ (.A0(_1679_),
    .A1(net1155),
    .S(_3428_),
    .X(_3436_));
 sky130_fd_sc_hd__clkbuf_1 _7814_ (.A(net1156),
    .X(_0744_));
 sky130_fd_sc_hd__nand2_8 _7815_ (.A(_0942_),
    .B(_1912_),
    .Y(_3437_));
 sky130_fd_sc_hd__mux2_1 _7816_ (.A0(_1658_),
    .A1(net1348),
    .S(_3437_),
    .X(_3438_));
 sky130_fd_sc_hd__clkbuf_1 _7817_ (.A(_3438_),
    .X(_0745_));
 sky130_fd_sc_hd__mux2_1 _7818_ (.A0(_1662_),
    .A1(net981),
    .S(_3437_),
    .X(_3439_));
 sky130_fd_sc_hd__clkbuf_1 _7819_ (.A(_3439_),
    .X(_0746_));
 sky130_fd_sc_hd__mux2_1 _7820_ (.A0(_3345_),
    .A1(net1002),
    .S(_3437_),
    .X(_3440_));
 sky130_fd_sc_hd__clkbuf_1 _7821_ (.A(net1003),
    .X(_0747_));
 sky130_fd_sc_hd__mux2_1 _7822_ (.A0(_3347_),
    .A1(\gpio_configure[36][3] ),
    .S(_3437_),
    .X(_3441_));
 sky130_fd_sc_hd__clkbuf_1 _7823_ (.A(net852),
    .X(_0748_));
 sky130_fd_sc_hd__mux2_1 _7824_ (.A0(_3349_),
    .A1(net696),
    .S(_3437_),
    .X(_3442_));
 sky130_fd_sc_hd__clkbuf_1 _7825_ (.A(net697),
    .X(_0749_));
 sky130_fd_sc_hd__mux2_1 _7826_ (.A0(_3351_),
    .A1(net762),
    .S(_3437_),
    .X(_3443_));
 sky130_fd_sc_hd__clkbuf_1 _7827_ (.A(net763),
    .X(_0750_));
 sky130_fd_sc_hd__mux2_1 _7828_ (.A0(_1675_),
    .A1(net752),
    .S(_3437_),
    .X(_3444_));
 sky130_fd_sc_hd__clkbuf_1 _7829_ (.A(net753),
    .X(_0751_));
 sky130_fd_sc_hd__mux2_1 _7830_ (.A0(_1679_),
    .A1(net1209),
    .S(_3437_),
    .X(_3445_));
 sky130_fd_sc_hd__clkbuf_1 _7831_ (.A(net1210),
    .X(_0752_));
 sky130_fd_sc_hd__nand2_8 _7832_ (.A(_0939_),
    .B(_1912_),
    .Y(_3446_));
 sky130_fd_sc_hd__mux2_1 _7833_ (.A0(_1658_),
    .A1(net1365),
    .S(_3446_),
    .X(_3447_));
 sky130_fd_sc_hd__clkbuf_1 _7834_ (.A(_3447_),
    .X(_0753_));
 sky130_fd_sc_hd__mux2_1 _7835_ (.A0(_1662_),
    .A1(net1043),
    .S(_3446_),
    .X(_3448_));
 sky130_fd_sc_hd__clkbuf_1 _7836_ (.A(_3448_),
    .X(_0754_));
 sky130_fd_sc_hd__mux2_1 _7837_ (.A0(_1664_),
    .A1(net1139),
    .S(_3446_),
    .X(_3449_));
 sky130_fd_sc_hd__clkbuf_1 _7838_ (.A(net1140),
    .X(_0755_));
 sky130_fd_sc_hd__mux2_1 _7839_ (.A0(_1666_),
    .A1(\gpio_configure[37][3] ),
    .S(_3446_),
    .X(_3450_));
 sky130_fd_sc_hd__clkbuf_1 _7840_ (.A(net884),
    .X(_0756_));
 sky130_fd_sc_hd__mux2_1 _7841_ (.A0(_1669_),
    .A1(net1079),
    .S(_3446_),
    .X(_3451_));
 sky130_fd_sc_hd__clkbuf_1 _7842_ (.A(_3451_),
    .X(_0757_));
 sky130_fd_sc_hd__mux2_1 _7843_ (.A0(_1672_),
    .A1(net781),
    .S(_3446_),
    .X(_3452_));
 sky130_fd_sc_hd__clkbuf_1 _7844_ (.A(net782),
    .X(_0758_));
 sky130_fd_sc_hd__mux2_1 _7845_ (.A0(_1675_),
    .A1(net826),
    .S(_3446_),
    .X(_3453_));
 sky130_fd_sc_hd__clkbuf_1 _7846_ (.A(net827),
    .X(_0759_));
 sky130_fd_sc_hd__mux2_1 _7847_ (.A0(_1679_),
    .A1(net1244),
    .S(_3446_),
    .X(_3454_));
 sky130_fd_sc_hd__clkbuf_1 _7848_ (.A(net1245),
    .X(_0760_));
 sky130_fd_sc_hd__nor2_1 _7849_ (.A(\xfer_state[1] ),
    .B(\xfer_state[2] ),
    .Y(_3455_));
 sky130_fd_sc_hd__or3_1 _7850_ (.A(\xfer_state[3] ),
    .B(_1547_),
    .C(_3455_),
    .X(_3456_));
 sky130_fd_sc_hd__nand2_1 _7851_ (.A(\xfer_state[1] ),
    .B(net306),
    .Y(_3457_));
 sky130_fd_sc_hd__o31a_1 _7852_ (.A1(\xfer_state[1] ),
    .A2(\xfer_state[3] ),
    .A3(\xfer_state[2] ),
    .B1(_3457_),
    .X(_3458_));
 sky130_fd_sc_hd__nand2_1 _7853_ (.A(\xfer_count[0] ),
    .B(_3458_),
    .Y(_3459_));
 sky130_fd_sc_hd__or2_1 _7854_ (.A(\xfer_count[0] ),
    .B(_3458_),
    .X(_3460_));
 sky130_fd_sc_hd__and3_1 _7855_ (.A(_3456_),
    .B(_3459_),
    .C(_3460_),
    .X(_3461_));
 sky130_fd_sc_hd__clkbuf_1 _7856_ (.A(_3461_),
    .X(_0761_));
 sky130_fd_sc_hd__inv_2 _7857_ (.A(_3458_),
    .Y(_3462_));
 sky130_fd_sc_hd__nor2_1 _7858_ (.A(\xfer_state[1] ),
    .B(\xfer_state[3] ),
    .Y(_3463_));
 sky130_fd_sc_hd__a21o_1 _7859_ (.A1(\xfer_count[0] ),
    .A2(\xfer_count[1] ),
    .B1(_3463_),
    .X(_3464_));
 sky130_fd_sc_hd__nor2_1 _7860_ (.A(_1532_),
    .B(_3464_),
    .Y(_3465_));
 sky130_fd_sc_hd__a22o_1 _7861_ (.A1(net1531),
    .A2(_3462_),
    .B1(_3465_),
    .B2(_3457_),
    .X(_0762_));
 sky130_fd_sc_hd__a31o_1 _7862_ (.A1(\xfer_count[0] ),
    .A2(\xfer_count[1] ),
    .A3(_3458_),
    .B1(\xfer_count[2] ),
    .X(_3466_));
 sky130_fd_sc_hd__and4_1 _7863_ (.A(\xfer_count[0] ),
    .B(\xfer_count[1] ),
    .C(\xfer_count[2] ),
    .D(_3458_),
    .X(_3467_));
 sky130_fd_sc_hd__clkinv_2 _7864_ (.A(_3467_),
    .Y(_3468_));
 sky130_fd_sc_hd__and3_1 _7865_ (.A(_3456_),
    .B(_3466_),
    .C(_3468_),
    .X(_3469_));
 sky130_fd_sc_hd__clkbuf_1 _7866_ (.A(_3469_),
    .X(_0763_));
 sky130_fd_sc_hd__a21boi_1 _7867_ (.A1(net1517),
    .A2(_3467_),
    .B1_N(_3456_),
    .Y(_3470_));
 sky130_fd_sc_hd__o21a_1 _7868_ (.A1(net1517),
    .A2(_3467_),
    .B1(_3470_),
    .X(_0764_));
 sky130_fd_sc_hd__nor2_2 _7869_ (.A(\xfer_state[0] ),
    .B(_1545_),
    .Y(_3471_));
 sky130_fd_sc_hd__mux2_1 _7870_ (.A0(_1545_),
    .A1(_3471_),
    .S(\pad_count_1[0] ),
    .X(_3472_));
 sky130_fd_sc_hd__clkbuf_1 _7871_ (.A(_3472_),
    .X(_0765_));
 sky130_fd_sc_hd__inv_2 _7872_ (.A(_1545_),
    .Y(_3473_));
 sky130_fd_sc_hd__nor2_8 _7873_ (.A(\pad_count_1[1] ),
    .B(\pad_count_1[0] ),
    .Y(_3474_));
 sky130_fd_sc_hd__and2_4 _7874_ (.A(\pad_count_1[1] ),
    .B(\pad_count_1[0] ),
    .X(_3475_));
 sky130_fd_sc_hd__or2_1 _7875_ (.A(\xfer_state[0] ),
    .B(_1545_),
    .X(_3476_));
 sky130_fd_sc_hd__o32a_1 _7876_ (.A1(_3473_),
    .A2(_3474_),
    .A3(_3475_),
    .B1(net1516),
    .B2(_3476_),
    .X(_0766_));
 sky130_fd_sc_hd__inv_2 _7877_ (.A(\pad_count_1[2] ),
    .Y(_3477_));
 sky130_fd_sc_hd__nand2_1 _7878_ (.A(_1545_),
    .B(_3474_),
    .Y(_3478_));
 sky130_fd_sc_hd__nand2_2 _7879_ (.A(\xfer_state[0] ),
    .B(_3473_),
    .Y(_3479_));
 sky130_fd_sc_hd__nand2_1 _7880_ (.A(_3478_),
    .B(_3479_),
    .Y(_3480_));
 sky130_fd_sc_hd__or2_1 _7881_ (.A(\pad_count_1[2] ),
    .B(_3478_),
    .X(_3481_));
 sky130_fd_sc_hd__o21ai_1 _7882_ (.A1(_3477_),
    .A2(_3480_),
    .B1(_3481_),
    .Y(_0767_));
 sky130_fd_sc_hd__nor2_1 _7883_ (.A(\pad_count_1[3] ),
    .B(_3481_),
    .Y(_3482_));
 sky130_fd_sc_hd__a31o_1 _7884_ (.A1(\pad_count_1[3] ),
    .A2(_3479_),
    .A3(_3481_),
    .B1(_3482_),
    .X(_0768_));
 sky130_fd_sc_hd__clkinv_4 _7885_ (.A(\pad_count_1[4] ),
    .Y(_3483_));
 sky130_fd_sc_hd__buf_6 _7886_ (.A(_3483_),
    .X(_3484_));
 sky130_fd_sc_hd__nand2_1 _7887_ (.A(_3484_),
    .B(_3479_),
    .Y(_3485_));
 sky130_fd_sc_hd__mux2_1 _7888_ (.A0(_3485_),
    .A1(_3484_),
    .S(_3482_),
    .X(_3486_));
 sky130_fd_sc_hd__clkbuf_1 _7889_ (.A(_3486_),
    .X(_0769_));
 sky130_fd_sc_hd__mux2_1 _7890_ (.A0(_3476_),
    .A1(_3473_),
    .S(\pad_count_2[0] ),
    .X(_3487_));
 sky130_fd_sc_hd__clkbuf_1 _7891_ (.A(_3487_),
    .X(_0770_));
 sky130_fd_sc_hd__nor2b_2 _7892_ (.A(\pad_count_2[1] ),
    .B_N(\pad_count_2[0] ),
    .Y(_3488_));
 sky130_fd_sc_hd__o32a_1 _7893_ (.A1(_3473_),
    .A2(_1528_),
    .A3(_3488_),
    .B1(_3476_),
    .B2(net1519),
    .X(_0771_));
 sky130_fd_sc_hd__and3_1 _7894_ (.A(\pad_count_2[1] ),
    .B(\pad_count_2[0] ),
    .C(_1545_),
    .X(_3489_));
 sky130_fd_sc_hd__a21oi_1 _7895_ (.A1(\pad_count_2[2] ),
    .A2(_3479_),
    .B1(_3489_),
    .Y(_3490_));
 sky130_fd_sc_hd__a21oi_1 _7896_ (.A1(net1499),
    .A2(_3489_),
    .B1(_3490_),
    .Y(_0772_));
 sky130_fd_sc_hd__and2_2 _7897_ (.A(\pad_count_2[3] ),
    .B(\pad_count_2[2] ),
    .X(_3491_));
 sky130_fd_sc_hd__nand2_1 _7898_ (.A(_3489_),
    .B(_3491_),
    .Y(_3492_));
 sky130_fd_sc_hd__and2_2 _7899_ (.A(\pad_count_2[1] ),
    .B(\pad_count_2[0] ),
    .X(_3493_));
 sky130_fd_sc_hd__and3_1 _7900_ (.A(_1545_),
    .B(_1529_),
    .C(_3493_),
    .X(_3494_));
 sky130_fd_sc_hd__a31o_1 _7901_ (.A1(net1529),
    .A2(_3479_),
    .A3(_3492_),
    .B1(_3494_),
    .X(_0773_));
 sky130_fd_sc_hd__nor2_1 _7902_ (.A(_1542_),
    .B(_1545_),
    .Y(_3495_));
 sky130_fd_sc_hd__nor2_1 _7903_ (.A(net1524),
    .B(_3495_),
    .Y(_3496_));
 sky130_fd_sc_hd__and3_1 _7904_ (.A(\pad_count_2[4] ),
    .B(_3489_),
    .C(_3491_),
    .X(_3497_));
 sky130_fd_sc_hd__a21oi_1 _7905_ (.A1(_3492_),
    .A2(_3496_),
    .B1(_3497_),
    .Y(_0774_));
 sky130_fd_sc_hd__and2b_1 _7906_ (.A_N(\pad_count_2[5] ),
    .B(\pad_count_2[4] ),
    .X(_3498_));
 sky130_fd_sc_hd__and3_2 _7907_ (.A(_3493_),
    .B(_3491_),
    .C(_3498_),
    .X(_3499_));
 sky130_fd_sc_hd__clkbuf_16 _7908_ (.A(_3499_),
    .X(_3500_));
 sky130_fd_sc_hd__nor2_1 _7909_ (.A(_3495_),
    .B(_3497_),
    .Y(_3501_));
 sky130_fd_sc_hd__a22o_1 _7910_ (.A1(_1545_),
    .A2(_3500_),
    .B1(_3501_),
    .B2(net1527),
    .X(_0775_));
 sky130_fd_sc_hd__nor2_1 _7911_ (.A(_1546_),
    .B(net306),
    .Y(_3502_));
 sky130_fd_sc_hd__a211o_1 _7912_ (.A1(\xfer_count[0] ),
    .A2(\xfer_count[1] ),
    .B1(\xfer_count[2] ),
    .C1(\xfer_count[3] ),
    .X(_3503_));
 sky130_fd_sc_hd__a22o_1 _7913_ (.A1(_3463_),
    .A2(_3471_),
    .B1(_3503_),
    .B2(\xfer_state[3] ),
    .X(_3504_));
 sky130_fd_sc_hd__mux2_1 _7914_ (.A0(_3502_),
    .A1(net1510),
    .S(_3504_),
    .X(_3505_));
 sky130_fd_sc_hd__clkbuf_1 _7915_ (.A(_3505_),
    .X(_0776_));
 sky130_fd_sc_hd__or4b_1 _7916_ (.A(\xfer_count[2] ),
    .B(\xfer_count[3] ),
    .C(_1543_),
    .D_N(\xfer_count[0] ),
    .X(_3506_));
 sky130_fd_sc_hd__a2bb2o_1 _7917_ (.A1_N(\xfer_count[1] ),
    .A2_N(_3506_),
    .B1(_3504_),
    .B2(serial_load_pre),
    .X(_0777_));
 sky130_fd_sc_hd__a21o_1 _7918_ (.A1(\xfer_state[0] ),
    .A2(_1543_),
    .B1(serial_busy),
    .X(_3507_));
 sky130_fd_sc_hd__o311a_1 _7919_ (.A1(serial_xfer),
    .A2(_1542_),
    .A3(net1525),
    .B1(_1544_),
    .C1(_3507_),
    .X(_0778_));
 sky130_fd_sc_hd__nor2_1 _7920_ (.A(\xfer_state[1] ),
    .B(_3473_),
    .Y(_3508_));
 sky130_fd_sc_hd__nor2_4 _7921_ (.A(\pad_count_1[3] ),
    .B(\pad_count_1[2] ),
    .Y(_3509_));
 sky130_fd_sc_hd__and3_2 _7922_ (.A(_3483_),
    .B(_3475_),
    .C(_3509_),
    .X(_3510_));
 sky130_fd_sc_hd__buf_8 _7923_ (.A(_3510_),
    .X(_3511_));
 sky130_fd_sc_hd__clkbuf_4 _7924_ (.A(_3483_),
    .X(_3512_));
 sky130_fd_sc_hd__nor2_4 _7925_ (.A(\pad_count_1[3] ),
    .B(_3477_),
    .Y(_3513_));
 sky130_fd_sc_hd__and3_2 _7926_ (.A(_3512_),
    .B(_3474_),
    .C(_3513_),
    .X(_3514_));
 sky130_fd_sc_hd__buf_8 _7927_ (.A(_3514_),
    .X(_3515_));
 sky130_fd_sc_hd__clkbuf_2 _7928_ (.A(\pad_count_1[4] ),
    .X(_3516_));
 sky130_fd_sc_hd__and2_2 _7929_ (.A(\pad_count_1[3] ),
    .B(_3477_),
    .X(_3517_));
 sky130_fd_sc_hd__and3_1 _7930_ (.A(_3516_),
    .B(_3475_),
    .C(_3517_),
    .X(_3518_));
 sky130_fd_sc_hd__buf_8 _7931_ (.A(_3518_),
    .X(_3519_));
 sky130_fd_sc_hd__and3_1 _7932_ (.A(_3516_),
    .B(_3475_),
    .C(_3509_),
    .X(_3520_));
 sky130_fd_sc_hd__buf_6 _7933_ (.A(_3520_),
    .X(_3521_));
 sky130_fd_sc_hd__a22o_1 _7934_ (.A1(\gpio_configure[27][0] ),
    .A2(_3519_),
    .B1(_3521_),
    .B2(\gpio_configure[19][0] ),
    .X(_3522_));
 sky130_fd_sc_hd__a221o_1 _7935_ (.A1(\gpio_configure[3][0] ),
    .A2(_3511_),
    .B1(_3515_),
    .B2(\gpio_configure[4][0] ),
    .C1(_3522_),
    .X(_3523_));
 sky130_fd_sc_hd__and2b_4 _7936_ (.A_N(\pad_count_1[0] ),
    .B(\pad_count_1[1] ),
    .X(_3524_));
 sky130_fd_sc_hd__and3_2 _7937_ (.A(_3512_),
    .B(_3509_),
    .C(_3524_),
    .X(_3525_));
 sky130_fd_sc_hd__buf_6 _7938_ (.A(_3525_),
    .X(_3526_));
 sky130_fd_sc_hd__and3_2 _7939_ (.A(_3512_),
    .B(_3474_),
    .C(_3517_),
    .X(_3527_));
 sky130_fd_sc_hd__buf_8 _7940_ (.A(_3527_),
    .X(_3528_));
 sky130_fd_sc_hd__and2b_4 _7941_ (.A_N(\pad_count_1[1] ),
    .B(\pad_count_1[0] ),
    .X(_3529_));
 sky130_fd_sc_hd__and3_2 _7942_ (.A(_3516_),
    .B(_3513_),
    .C(_3529_),
    .X(_3530_));
 sky130_fd_sc_hd__and3_4 _7943_ (.A(_3484_),
    .B(_3513_),
    .C(_3524_),
    .X(_3531_));
 sky130_fd_sc_hd__a22o_1 _7944_ (.A1(\gpio_configure[21][0] ),
    .A2(_3530_),
    .B1(_3531_),
    .B2(\gpio_configure[6][0] ),
    .X(_3532_));
 sky130_fd_sc_hd__a221o_1 _7945_ (.A1(\gpio_configure[2][0] ),
    .A2(_3526_),
    .B1(_3528_),
    .B2(\gpio_configure[8][0] ),
    .C1(_3532_),
    .X(_3533_));
 sky130_fd_sc_hd__and3_2 _7946_ (.A(\pad_count_1[4] ),
    .B(_3474_),
    .C(_3517_),
    .X(_3534_));
 sky130_fd_sc_hd__buf_6 _7947_ (.A(_3534_),
    .X(_3535_));
 sky130_fd_sc_hd__and3_2 _7948_ (.A(_3512_),
    .B(_3475_),
    .C(_3513_),
    .X(_3536_));
 sky130_fd_sc_hd__buf_6 _7949_ (.A(_3536_),
    .X(_3537_));
 sky130_fd_sc_hd__and2_2 _7950_ (.A(\pad_count_1[3] ),
    .B(\pad_count_1[2] ),
    .X(_3538_));
 sky130_fd_sc_hd__and3_1 _7951_ (.A(_3483_),
    .B(_3474_),
    .C(_3538_),
    .X(_3539_));
 sky130_fd_sc_hd__buf_6 _7952_ (.A(_3539_),
    .X(_3540_));
 sky130_fd_sc_hd__and2_1 _7953_ (.A(\gpio_configure[12][0] ),
    .B(_3540_),
    .X(_3541_));
 sky130_fd_sc_hd__a221o_1 _7954_ (.A1(\gpio_configure[24][0] ),
    .A2(_3535_),
    .B1(_3537_),
    .B2(\gpio_configure[7][0] ),
    .C1(_3541_),
    .X(_3542_));
 sky130_fd_sc_hd__and3_4 _7955_ (.A(_3483_),
    .B(_3475_),
    .C(_3538_),
    .X(_3543_));
 sky130_fd_sc_hd__buf_8 _7956_ (.A(_3543_),
    .X(_3544_));
 sky130_fd_sc_hd__and3_4 _7957_ (.A(_3483_),
    .B(_3517_),
    .C(_3529_),
    .X(_3545_));
 sky130_fd_sc_hd__buf_6 _7958_ (.A(_3545_),
    .X(_3546_));
 sky130_fd_sc_hd__and3_4 _7959_ (.A(_3516_),
    .B(_3475_),
    .C(_3513_),
    .X(_3547_));
 sky130_fd_sc_hd__buf_8 _7960_ (.A(_3547_),
    .X(_3548_));
 sky130_fd_sc_hd__and3_2 _7961_ (.A(\pad_count_1[4] ),
    .B(_3509_),
    .C(_3529_),
    .X(_3549_));
 sky130_fd_sc_hd__buf_6 _7962_ (.A(_3549_),
    .X(_3550_));
 sky130_fd_sc_hd__a22o_1 _7963_ (.A1(\gpio_configure[23][0] ),
    .A2(_3548_),
    .B1(_3550_),
    .B2(\gpio_configure[17][0] ),
    .X(_3551_));
 sky130_fd_sc_hd__a221o_1 _7964_ (.A1(\gpio_configure[15][0] ),
    .A2(_3544_),
    .B1(_3546_),
    .B2(\gpio_configure[9][0] ),
    .C1(_3551_),
    .X(_3552_));
 sky130_fd_sc_hd__or4_1 _7965_ (.A(_3523_),
    .B(_3533_),
    .C(_3542_),
    .D(_3552_),
    .X(_3553_));
 sky130_fd_sc_hd__and3_2 _7966_ (.A(_3516_),
    .B(_3474_),
    .C(_3538_),
    .X(_3554_));
 sky130_fd_sc_hd__buf_6 _7967_ (.A(_3554_),
    .X(_3555_));
 sky130_fd_sc_hd__and3_2 _7968_ (.A(_3512_),
    .B(_3529_),
    .C(_3538_),
    .X(_3556_));
 sky130_fd_sc_hd__buf_6 _7969_ (.A(_3556_),
    .X(_3557_));
 sky130_fd_sc_hd__and3_4 _7970_ (.A(\pad_count_1[4] ),
    .B(_3529_),
    .C(_3538_),
    .X(_3558_));
 sky130_fd_sc_hd__buf_6 _7971_ (.A(_3558_),
    .X(_3559_));
 sky130_fd_sc_hd__and3_4 _7972_ (.A(_3512_),
    .B(_3509_),
    .C(_3529_),
    .X(_3560_));
 sky130_fd_sc_hd__buf_6 _7973_ (.A(_3560_),
    .X(_3561_));
 sky130_fd_sc_hd__a22o_1 _7974_ (.A1(\gpio_configure[29][0] ),
    .A2(_3559_),
    .B1(_3561_),
    .B2(\gpio_configure[1][0] ),
    .X(_3562_));
 sky130_fd_sc_hd__a221o_1 _7975_ (.A1(\gpio_configure[28][0] ),
    .A2(_3555_),
    .B1(_3557_),
    .B2(\gpio_configure[13][0] ),
    .C1(_3562_),
    .X(_3563_));
 sky130_fd_sc_hd__and3_2 _7976_ (.A(\pad_count_1[4] ),
    .B(_3517_),
    .C(_3524_),
    .X(_3564_));
 sky130_fd_sc_hd__buf_6 _7977_ (.A(_3564_),
    .X(_3565_));
 sky130_fd_sc_hd__and3_2 _7978_ (.A(_3483_),
    .B(_3513_),
    .C(_3529_),
    .X(_3566_));
 sky130_fd_sc_hd__buf_6 _7979_ (.A(_3566_),
    .X(_3567_));
 sky130_fd_sc_hd__and3_2 _7980_ (.A(_3516_),
    .B(_3509_),
    .C(_3524_),
    .X(_3568_));
 sky130_fd_sc_hd__buf_6 _7981_ (.A(_3568_),
    .X(_3569_));
 sky130_fd_sc_hd__and2_4 _7982_ (.A(_3474_),
    .B(_3509_),
    .X(_3570_));
 sky130_fd_sc_hd__buf_8 _7983_ (.A(_3570_),
    .X(_3571_));
 sky130_fd_sc_hd__and3_2 _7984_ (.A(_3512_),
    .B(_3474_),
    .C(_3509_),
    .X(_3572_));
 sky130_fd_sc_hd__a221o_1 _7985_ (.A1(\gpio_configure[18][0] ),
    .A2(_3569_),
    .B1(_3571_),
    .B2(\gpio_configure[16][0] ),
    .C1(_3572_),
    .X(_3573_));
 sky130_fd_sc_hd__a221o_1 _7986_ (.A1(\gpio_configure[26][0] ),
    .A2(_3565_),
    .B1(_3567_),
    .B2(\gpio_configure[5][0] ),
    .C1(_3573_),
    .X(_3574_));
 sky130_fd_sc_hd__and3_2 _7987_ (.A(\pad_count_1[4] ),
    .B(_3475_),
    .C(_3538_),
    .X(_3575_));
 sky130_fd_sc_hd__buf_8 _7988_ (.A(_3575_),
    .X(_3576_));
 sky130_fd_sc_hd__and3_2 _7989_ (.A(_3484_),
    .B(_3475_),
    .C(_3517_),
    .X(_3577_));
 sky130_fd_sc_hd__buf_8 _7990_ (.A(_3577_),
    .X(_3578_));
 sky130_fd_sc_hd__and3_2 _7991_ (.A(_3516_),
    .B(_3474_),
    .C(_3513_),
    .X(_3579_));
 sky130_fd_sc_hd__and3_4 _7992_ (.A(_3516_),
    .B(_3517_),
    .C(_3529_),
    .X(_3580_));
 sky130_fd_sc_hd__buf_8 _7993_ (.A(_3580_),
    .X(_3581_));
 sky130_fd_sc_hd__a22o_1 _7994_ (.A1(\gpio_configure[20][0] ),
    .A2(_3579_),
    .B1(_3581_),
    .B2(\gpio_configure[25][0] ),
    .X(_3582_));
 sky130_fd_sc_hd__a221o_1 _7995_ (.A1(\gpio_configure[31][0] ),
    .A2(_3576_),
    .B1(_3578_),
    .B2(\gpio_configure[11][0] ),
    .C1(_3582_),
    .X(_3583_));
 sky130_fd_sc_hd__and3_2 _7996_ (.A(_3516_),
    .B(_3513_),
    .C(_3524_),
    .X(_3584_));
 sky130_fd_sc_hd__buf_8 _7997_ (.A(_3584_),
    .X(_3585_));
 sky130_fd_sc_hd__and3_1 _7998_ (.A(_3516_),
    .B(_3524_),
    .C(_3538_),
    .X(_3586_));
 sky130_fd_sc_hd__buf_6 _7999_ (.A(_3586_),
    .X(_3587_));
 sky130_fd_sc_hd__and3_2 _8000_ (.A(_3512_),
    .B(_3517_),
    .C(_3524_),
    .X(_3588_));
 sky130_fd_sc_hd__buf_8 _8001_ (.A(_3588_),
    .X(_3589_));
 sky130_fd_sc_hd__and3_1 _8002_ (.A(_3483_),
    .B(_3524_),
    .C(_3538_),
    .X(_3590_));
 sky130_fd_sc_hd__buf_6 _8003_ (.A(_3590_),
    .X(_3591_));
 sky130_fd_sc_hd__a22o_1 _8004_ (.A1(\gpio_configure[10][0] ),
    .A2(_3589_),
    .B1(_3591_),
    .B2(\gpio_configure[14][0] ),
    .X(_3592_));
 sky130_fd_sc_hd__a221o_1 _8005_ (.A1(\gpio_configure[22][0] ),
    .A2(_3585_),
    .B1(_3587_),
    .B2(\gpio_configure[30][0] ),
    .C1(_3592_),
    .X(_3593_));
 sky130_fd_sc_hd__or4_1 _8006_ (.A(_3563_),
    .B(_3574_),
    .C(_3583_),
    .D(_3593_),
    .X(_3594_));
 sky130_fd_sc_hd__or2_1 _8007_ (.A(_3553_),
    .B(_3594_),
    .X(_3595_));
 sky130_fd_sc_hd__nand2_2 _8008_ (.A(_3484_),
    .B(_3571_),
    .Y(_3596_));
 sky130_fd_sc_hd__buf_4 _8009_ (.A(_3596_),
    .X(_3597_));
 sky130_fd_sc_hd__or2_1 _8010_ (.A(\gpio_configure[0][0] ),
    .B(_3597_),
    .X(_3598_));
 sky130_fd_sc_hd__or2_1 _8011_ (.A(_3502_),
    .B(_3455_),
    .X(_3599_));
 sky130_fd_sc_hd__clkbuf_4 _8012_ (.A(_3599_),
    .X(_3600_));
 sky130_fd_sc_hd__buf_2 _8013_ (.A(_3600_),
    .X(_3601_));
 sky130_fd_sc_hd__a32o_1 _8014_ (.A1(_3508_),
    .A2(_3595_),
    .A3(_3598_),
    .B1(_3601_),
    .B2(net1459),
    .X(_0779_));
 sky130_fd_sc_hd__nor2_2 _8015_ (.A(_3502_),
    .B(_3455_),
    .Y(_3602_));
 sky130_fd_sc_hd__clkbuf_4 _8016_ (.A(_3602_),
    .X(_3603_));
 sky130_fd_sc_hd__clkbuf_4 _8017_ (.A(_3603_),
    .X(_3604_));
 sky130_fd_sc_hd__a22o_1 _8018_ (.A1(\gpio_configure[27][1] ),
    .A2(_3518_),
    .B1(_3587_),
    .B2(\gpio_configure[30][1] ),
    .X(_3605_));
 sky130_fd_sc_hd__a221o_1 _8019_ (.A1(\gpio_configure[18][1] ),
    .A2(_3569_),
    .B1(_3585_),
    .B2(\gpio_configure[22][1] ),
    .C1(_3605_),
    .X(_3606_));
 sky130_fd_sc_hd__buf_6 _8020_ (.A(_3530_),
    .X(_3607_));
 sky130_fd_sc_hd__a22o_1 _8021_ (.A1(\gpio_configure[19][1] ),
    .A2(_3520_),
    .B1(_3577_),
    .B2(\gpio_configure[11][1] ),
    .X(_3608_));
 sky130_fd_sc_hd__a221o_1 _8022_ (.A1(\gpio_configure[21][1] ),
    .A2(_3607_),
    .B1(_3546_),
    .B2(\gpio_configure[9][1] ),
    .C1(_3608_),
    .X(_3609_));
 sky130_fd_sc_hd__and2_1 _8023_ (.A(\gpio_configure[15][1] ),
    .B(_3544_),
    .X(_3610_));
 sky130_fd_sc_hd__a221o_1 _8024_ (.A1(\gpio_configure[23][1] ),
    .A2(_3548_),
    .B1(_3561_),
    .B2(\gpio_configure[1][1] ),
    .C1(_3610_),
    .X(_3611_));
 sky130_fd_sc_hd__a22o_1 _8025_ (.A1(\gpio_configure[24][1] ),
    .A2(_3535_),
    .B1(_3565_),
    .B2(\gpio_configure[26][1] ),
    .X(_3612_));
 sky130_fd_sc_hd__a221o_1 _8026_ (.A1(\gpio_configure[4][1] ),
    .A2(_3515_),
    .B1(_3550_),
    .B2(\gpio_configure[17][1] ),
    .C1(_3612_),
    .X(_3613_));
 sky130_fd_sc_hd__or4_2 _8027_ (.A(_3606_),
    .B(_3609_),
    .C(_3611_),
    .D(_3613_),
    .X(_3614_));
 sky130_fd_sc_hd__a22o_1 _8028_ (.A1(\gpio_configure[29][1] ),
    .A2(_3559_),
    .B1(_3555_),
    .B2(\gpio_configure[28][1] ),
    .X(_3615_));
 sky130_fd_sc_hd__a221o_1 _8029_ (.A1(\gpio_configure[8][1] ),
    .A2(_3528_),
    .B1(_3589_),
    .B2(\gpio_configure[10][1] ),
    .C1(_3615_),
    .X(_3616_));
 sky130_fd_sc_hd__a221o_1 _8030_ (.A1(\gpio_configure[16][1] ),
    .A2(_3571_),
    .B1(_3579_),
    .B2(\gpio_configure[20][1] ),
    .C1(_3572_),
    .X(_3617_));
 sky130_fd_sc_hd__a221o_1 _8031_ (.A1(\gpio_configure[12][1] ),
    .A2(_3540_),
    .B1(_3557_),
    .B2(\gpio_configure[13][1] ),
    .C1(_3617_),
    .X(_3618_));
 sky130_fd_sc_hd__a22o_1 _8032_ (.A1(\gpio_configure[3][1] ),
    .A2(_3511_),
    .B1(_3576_),
    .B2(\gpio_configure[31][1] ),
    .X(_3619_));
 sky130_fd_sc_hd__a221o_1 _8033_ (.A1(\gpio_configure[2][1] ),
    .A2(_3526_),
    .B1(_3537_),
    .B2(\gpio_configure[7][1] ),
    .C1(_3619_),
    .X(_3620_));
 sky130_fd_sc_hd__buf_6 _8034_ (.A(_3531_),
    .X(_3621_));
 sky130_fd_sc_hd__a22o_1 _8035_ (.A1(\gpio_configure[5][1] ),
    .A2(_3567_),
    .B1(_3591_),
    .B2(\gpio_configure[14][1] ),
    .X(_3622_));
 sky130_fd_sc_hd__a221o_1 _8036_ (.A1(\gpio_configure[6][1] ),
    .A2(_3621_),
    .B1(_3581_),
    .B2(\gpio_configure[25][1] ),
    .C1(_3622_),
    .X(_3623_));
 sky130_fd_sc_hd__or4_2 _8037_ (.A(_3616_),
    .B(_3618_),
    .C(_3620_),
    .D(_3623_),
    .X(_3624_));
 sky130_fd_sc_hd__buf_6 _8038_ (.A(_1546_),
    .X(_3625_));
 sky130_fd_sc_hd__o221a_1 _8039_ (.A1(\gpio_configure[0][1] ),
    .A2(_3597_),
    .B1(_3614_),
    .B2(_3624_),
    .C1(_3625_),
    .X(_3626_));
 sky130_fd_sc_hd__a211o_1 _8040_ (.A1(_1525_),
    .A2(\serial_data_staging_1[0] ),
    .B1(_3600_),
    .C1(_3626_),
    .X(_3627_));
 sky130_fd_sc_hd__o21a_1 _8041_ (.A1(net1453),
    .A2(_3604_),
    .B1(_3627_),
    .X(_0780_));
 sky130_fd_sc_hd__a22o_1 _8042_ (.A1(\gpio_configure[24][2] ),
    .A2(_3534_),
    .B1(_3568_),
    .B2(\gpio_configure[18][2] ),
    .X(_3628_));
 sky130_fd_sc_hd__a221o_1 _8043_ (.A1(\gpio_configure[23][2] ),
    .A2(_3547_),
    .B1(_3588_),
    .B2(\gpio_configure[10][2] ),
    .C1(_3628_),
    .X(_3629_));
 sky130_fd_sc_hd__a22o_1 _8044_ (.A1(\gpio_configure[12][2] ),
    .A2(_3539_),
    .B1(_3590_),
    .B2(\gpio_configure[14][2] ),
    .X(_3630_));
 sky130_fd_sc_hd__a221o_1 _8045_ (.A1(\gpio_configure[8][2] ),
    .A2(_3527_),
    .B1(_3556_),
    .B2(\gpio_configure[13][2] ),
    .C1(_3630_),
    .X(_3631_));
 sky130_fd_sc_hd__a22o_1 _8046_ (.A1(\gpio_configure[17][2] ),
    .A2(_3549_),
    .B1(_3575_),
    .B2(\gpio_configure[31][2] ),
    .X(_3632_));
 sky130_fd_sc_hd__a221o_1 _8047_ (.A1(\gpio_configure[3][2] ),
    .A2(_3510_),
    .B1(_3584_),
    .B2(\gpio_configure[22][2] ),
    .C1(_3632_),
    .X(_3633_));
 sky130_fd_sc_hd__a221o_1 _8048_ (.A1(\gpio_configure[16][2] ),
    .A2(_3570_),
    .B1(_3564_),
    .B2(\gpio_configure[26][2] ),
    .C1(_3572_),
    .X(_3634_));
 sky130_fd_sc_hd__a221o_1 _8049_ (.A1(\gpio_configure[4][2] ),
    .A2(_3514_),
    .B1(_3543_),
    .B2(\gpio_configure[15][2] ),
    .C1(_3634_),
    .X(_3635_));
 sky130_fd_sc_hd__or4_1 _8050_ (.A(_3629_),
    .B(_3631_),
    .C(_3633_),
    .D(_3635_),
    .X(_3636_));
 sky130_fd_sc_hd__a22o_1 _8051_ (.A1(\gpio_configure[5][2] ),
    .A2(_3567_),
    .B1(_3581_),
    .B2(\gpio_configure[25][2] ),
    .X(_3637_));
 sky130_fd_sc_hd__a22o_1 _8052_ (.A1(\gpio_configure[7][2] ),
    .A2(_3536_),
    .B1(_3560_),
    .B2(\gpio_configure[1][2] ),
    .X(_3638_));
 sky130_fd_sc_hd__a22o_1 _8053_ (.A1(\gpio_configure[9][2] ),
    .A2(_3545_),
    .B1(_3558_),
    .B2(\gpio_configure[29][2] ),
    .X(_3639_));
 sky130_fd_sc_hd__a211o_1 _8054_ (.A1(\gpio_configure[6][2] ),
    .A2(_3531_),
    .B1(_3638_),
    .C1(_3639_),
    .X(_3640_));
 sky130_fd_sc_hd__a22o_1 _8055_ (.A1(\gpio_configure[28][2] ),
    .A2(_3554_),
    .B1(_3586_),
    .B2(\gpio_configure[30][2] ),
    .X(_3641_));
 sky130_fd_sc_hd__a221o_1 _8056_ (.A1(\gpio_configure[2][2] ),
    .A2(_3525_),
    .B1(_3579_),
    .B2(\gpio_configure[20][2] ),
    .C1(_3641_),
    .X(_3642_));
 sky130_fd_sc_hd__a22o_1 _8057_ (.A1(\gpio_configure[27][2] ),
    .A2(_3518_),
    .B1(_3520_),
    .B2(\gpio_configure[19][2] ),
    .X(_3643_));
 sky130_fd_sc_hd__a221o_1 _8058_ (.A1(\gpio_configure[21][2] ),
    .A2(_3530_),
    .B1(_3577_),
    .B2(\gpio_configure[11][2] ),
    .C1(_3643_),
    .X(_3644_));
 sky130_fd_sc_hd__or4_2 _8059_ (.A(_3637_),
    .B(_3640_),
    .C(_3642_),
    .D(_3644_),
    .X(_3645_));
 sky130_fd_sc_hd__o22a_1 _8060_ (.A1(\gpio_configure[0][2] ),
    .A2(_3596_),
    .B1(_3636_),
    .B2(_3645_),
    .X(_3646_));
 sky130_fd_sc_hd__o22a_1 _8061_ (.A1(\serial_data_staging_1[1] ),
    .A2(_3508_),
    .B1(_3646_),
    .B2(\xfer_state[1] ),
    .X(_3647_));
 sky130_fd_sc_hd__mux2_1 _8062_ (.A0(net1513),
    .A1(_3647_),
    .S(_3603_),
    .X(_3648_));
 sky130_fd_sc_hd__clkbuf_1 _8063_ (.A(_3648_),
    .X(_0781_));
 sky130_fd_sc_hd__a22o_1 _8064_ (.A1(\gpio_configure[17][3] ),
    .A2(_3550_),
    .B1(_3544_),
    .B2(\gpio_configure[15][3] ),
    .X(_3649_));
 sky130_fd_sc_hd__a221o_1 _8065_ (.A1(\gpio_configure[4][3] ),
    .A2(_3515_),
    .B1(_3565_),
    .B2(\gpio_configure[26][3] ),
    .C1(_3649_),
    .X(_3650_));
 sky130_fd_sc_hd__a22o_1 _8066_ (.A1(\gpio_configure[2][3] ),
    .A2(_3525_),
    .B1(_3557_),
    .B2(\gpio_configure[13][3] ),
    .X(_3651_));
 sky130_fd_sc_hd__a221o_1 _8067_ (.A1(\gpio_configure[6][3] ),
    .A2(_3621_),
    .B1(_3576_),
    .B2(\gpio_configure[31][3] ),
    .C1(_3651_),
    .X(_3652_));
 sky130_fd_sc_hd__and2_1 _8068_ (.A(\gpio_configure[30][3] ),
    .B(_3586_),
    .X(_3653_));
 sky130_fd_sc_hd__a221o_1 _8069_ (.A1(\gpio_configure[27][3] ),
    .A2(_3519_),
    .B1(_3521_),
    .B2(\gpio_configure[19][3] ),
    .C1(_3653_),
    .X(_3654_));
 sky130_fd_sc_hd__a22o_1 _8070_ (.A1(\gpio_configure[24][3] ),
    .A2(_3535_),
    .B1(_3577_),
    .B2(\gpio_configure[11][3] ),
    .X(_3655_));
 sky130_fd_sc_hd__a221o_1 _8071_ (.A1(\gpio_configure[18][3] ),
    .A2(_3569_),
    .B1(_3581_),
    .B2(\gpio_configure[25][3] ),
    .C1(_3655_),
    .X(_3656_));
 sky130_fd_sc_hd__or4_2 _8072_ (.A(_3650_),
    .B(_3652_),
    .C(_3654_),
    .D(_3656_),
    .X(_3657_));
 sky130_fd_sc_hd__a22o_1 _8073_ (.A1(\gpio_configure[12][3] ),
    .A2(_3540_),
    .B1(_3591_),
    .B2(\gpio_configure[14][3] ),
    .X(_3658_));
 sky130_fd_sc_hd__a221o_1 _8074_ (.A1(\gpio_configure[8][3] ),
    .A2(_3528_),
    .B1(_3589_),
    .B2(\gpio_configure[10][3] ),
    .C1(_3658_),
    .X(_3659_));
 sky130_fd_sc_hd__a221o_1 _8075_ (.A1(\gpio_configure[16][3] ),
    .A2(_3571_),
    .B1(_3566_),
    .B2(\gpio_configure[5][3] ),
    .C1(_3572_),
    .X(_3660_));
 sky130_fd_sc_hd__a221o_1 _8076_ (.A1(\gpio_configure[7][3] ),
    .A2(_3537_),
    .B1(_3559_),
    .B2(\gpio_configure[29][3] ),
    .C1(_3660_),
    .X(_3661_));
 sky130_fd_sc_hd__buf_6 _8077_ (.A(_3579_),
    .X(_3662_));
 sky130_fd_sc_hd__a22o_1 _8078_ (.A1(\gpio_configure[21][3] ),
    .A2(_3530_),
    .B1(_3561_),
    .B2(\gpio_configure[1][3] ),
    .X(_3663_));
 sky130_fd_sc_hd__a221o_1 _8079_ (.A1(\gpio_configure[9][3] ),
    .A2(_3546_),
    .B1(_3662_),
    .B2(\gpio_configure[20][3] ),
    .C1(_3663_),
    .X(_3664_));
 sky130_fd_sc_hd__a22o_1 _8080_ (.A1(\gpio_configure[3][3] ),
    .A2(_3511_),
    .B1(_3585_),
    .B2(\gpio_configure[22][3] ),
    .X(_3665_));
 sky130_fd_sc_hd__a221o_1 _8081_ (.A1(\gpio_configure[23][3] ),
    .A2(_3548_),
    .B1(_3555_),
    .B2(\gpio_configure[28][3] ),
    .C1(_3665_),
    .X(_3666_));
 sky130_fd_sc_hd__or4_2 _8082_ (.A(_3659_),
    .B(_3661_),
    .C(_3664_),
    .D(_3666_),
    .X(_3667_));
 sky130_fd_sc_hd__o221a_1 _8083_ (.A1(\gpio_configure[0][3] ),
    .A2(_3597_),
    .B1(_3657_),
    .B2(_3667_),
    .C1(_3625_),
    .X(_3668_));
 sky130_fd_sc_hd__a211o_1 _8084_ (.A1(_1525_),
    .A2(\serial_data_staging_1[2] ),
    .B1(_3600_),
    .C1(_3668_),
    .X(_3669_));
 sky130_fd_sc_hd__o21a_1 _8085_ (.A1(net1480),
    .A2(_3604_),
    .B1(_3669_),
    .X(_0782_));
 sky130_fd_sc_hd__a22o_1 _8086_ (.A1(\gpio_configure[27][4] ),
    .A2(_3519_),
    .B1(_3521_),
    .B2(\gpio_configure[19][4] ),
    .X(_3670_));
 sky130_fd_sc_hd__a221o_1 _8087_ (.A1(\gpio_configure[21][4] ),
    .A2(_3607_),
    .B1(_3578_),
    .B2(\gpio_configure[11][4] ),
    .C1(_3670_),
    .X(_3671_));
 sky130_fd_sc_hd__a22o_1 _8088_ (.A1(\gpio_configure[24][4] ),
    .A2(_3535_),
    .B1(_3569_),
    .B2(\gpio_configure[18][4] ),
    .X(_3672_));
 sky130_fd_sc_hd__a221o_1 _8089_ (.A1(\gpio_configure[23][4] ),
    .A2(_3548_),
    .B1(_3589_),
    .B2(\gpio_configure[10][4] ),
    .C1(_3672_),
    .X(_3673_));
 sky130_fd_sc_hd__a22o_1 _8090_ (.A1(\gpio_configure[12][4] ),
    .A2(_3540_),
    .B1(_3591_),
    .B2(\gpio_configure[14][4] ),
    .X(_3674_));
 sky130_fd_sc_hd__a221o_1 _8091_ (.A1(\gpio_configure[8][4] ),
    .A2(_3528_),
    .B1(_3557_),
    .B2(\gpio_configure[13][4] ),
    .C1(_3674_),
    .X(_3675_));
 sky130_fd_sc_hd__a22o_1 _8092_ (.A1(\gpio_configure[17][4] ),
    .A2(_3550_),
    .B1(_3576_),
    .B2(\gpio_configure[31][4] ),
    .X(_3676_));
 sky130_fd_sc_hd__a221o_1 _8093_ (.A1(\gpio_configure[3][4] ),
    .A2(_3511_),
    .B1(_3585_),
    .B2(\gpio_configure[22][4] ),
    .C1(_3676_),
    .X(_3677_));
 sky130_fd_sc_hd__or2_1 _8094_ (.A(\gpio_configure[16][4] ),
    .B(_3512_),
    .X(_3678_));
 sky130_fd_sc_hd__a22o_1 _8095_ (.A1(\gpio_configure[26][4] ),
    .A2(_3565_),
    .B1(_3678_),
    .B2(_3571_),
    .X(_3679_));
 sky130_fd_sc_hd__a221o_1 _8096_ (.A1(\gpio_configure[4][4] ),
    .A2(_3515_),
    .B1(_3544_),
    .B2(\gpio_configure[15][4] ),
    .C1(_3679_),
    .X(_3680_));
 sky130_fd_sc_hd__or4_1 _8097_ (.A(_3673_),
    .B(_3675_),
    .C(_3677_),
    .D(_3680_),
    .X(_3681_));
 sky130_fd_sc_hd__a22o_1 _8098_ (.A1(\gpio_configure[5][4] ),
    .A2(_3567_),
    .B1(_3581_),
    .B2(\gpio_configure[25][4] ),
    .X(_3682_));
 sky130_fd_sc_hd__a22o_1 _8099_ (.A1(\gpio_configure[9][4] ),
    .A2(_3546_),
    .B1(_3559_),
    .B2(\gpio_configure[29][4] ),
    .X(_3683_));
 sky130_fd_sc_hd__a221o_1 _8100_ (.A1(\gpio_configure[7][4] ),
    .A2(_3537_),
    .B1(_3561_),
    .B2(\gpio_configure[1][4] ),
    .C1(_3683_),
    .X(_3684_));
 sky130_fd_sc_hd__a211o_1 _8101_ (.A1(\gpio_configure[6][4] ),
    .A2(_3621_),
    .B1(_3682_),
    .C1(_3684_),
    .X(_3685_));
 sky130_fd_sc_hd__a22o_1 _8102_ (.A1(\gpio_configure[28][4] ),
    .A2(_3555_),
    .B1(_3587_),
    .B2(\gpio_configure[30][4] ),
    .X(_3686_));
 sky130_fd_sc_hd__a221o_1 _8103_ (.A1(\gpio_configure[2][4] ),
    .A2(_3526_),
    .B1(_3662_),
    .B2(\gpio_configure[20][4] ),
    .C1(_3686_),
    .X(_3687_));
 sky130_fd_sc_hd__or4_4 _8104_ (.A(_3671_),
    .B(_3681_),
    .C(_3685_),
    .D(_3687_),
    .X(_3688_));
 sky130_fd_sc_hd__buf_4 _8105_ (.A(_1546_),
    .X(_3689_));
 sky130_fd_sc_hd__o211a_1 _8106_ (.A1(\gpio_configure[0][4] ),
    .A2(_3597_),
    .B1(_3688_),
    .C1(_3689_),
    .X(_3690_));
 sky130_fd_sc_hd__a21o_1 _8107_ (.A1(_1526_),
    .A2(net1480),
    .B1(_3601_),
    .X(_3691_));
 sky130_fd_sc_hd__o22a_1 _8108_ (.A1(net1495),
    .A2(_3604_),
    .B1(_3690_),
    .B2(_3691_),
    .X(_0783_));
 sky130_fd_sc_hd__a22o_1 _8109_ (.A1(\gpio_configure[2][5] ),
    .A2(_3526_),
    .B1(_3548_),
    .B2(\gpio_configure[23][5] ),
    .X(_3692_));
 sky130_fd_sc_hd__a221o_1 _8110_ (.A1(\gpio_configure[28][5] ),
    .A2(_3555_),
    .B1(_3581_),
    .B2(\gpio_configure[25][5] ),
    .C1(_3692_),
    .X(_3693_));
 sky130_fd_sc_hd__a22o_1 _8111_ (.A1(\gpio_configure[12][5] ),
    .A2(_3540_),
    .B1(_3569_),
    .B2(\gpio_configure[18][5] ),
    .X(_3694_));
 sky130_fd_sc_hd__a221o_1 _8112_ (.A1(\gpio_configure[27][5] ),
    .A2(_3519_),
    .B1(_3578_),
    .B2(\gpio_configure[11][5] ),
    .C1(_3694_),
    .X(_3695_));
 sky130_fd_sc_hd__a22o_1 _8113_ (.A1(\gpio_configure[20][5] ),
    .A2(_3662_),
    .B1(_3585_),
    .B2(\gpio_configure[22][5] ),
    .X(_3696_));
 sky130_fd_sc_hd__a21o_1 _8114_ (.A1(\gpio_configure[8][5] ),
    .A2(_3528_),
    .B1(_3696_),
    .X(_3697_));
 sky130_fd_sc_hd__a22o_1 _8115_ (.A1(\gpio_configure[7][5] ),
    .A2(_3537_),
    .B1(_3587_),
    .B2(\gpio_configure[30][5] ),
    .X(_3698_));
 sky130_fd_sc_hd__a221o_1 _8116_ (.A1(\gpio_configure[4][5] ),
    .A2(_3515_),
    .B1(_3535_),
    .B2(\gpio_configure[24][5] ),
    .C1(_3698_),
    .X(_3699_));
 sky130_fd_sc_hd__or4_1 _8117_ (.A(_3693_),
    .B(_3695_),
    .C(_3697_),
    .D(_3699_),
    .X(_3700_));
 sky130_fd_sc_hd__a22o_1 _8118_ (.A1(\gpio_configure[19][5] ),
    .A2(_3521_),
    .B1(_3576_),
    .B2(\gpio_configure[31][5] ),
    .X(_3701_));
 sky130_fd_sc_hd__a221o_1 _8119_ (.A1(\gpio_configure[5][5] ),
    .A2(_3567_),
    .B1(_3589_),
    .B2(\gpio_configure[10][5] ),
    .C1(_3701_),
    .X(_3702_));
 sky130_fd_sc_hd__or2_1 _8120_ (.A(\gpio_configure[16][5] ),
    .B(_3484_),
    .X(_3703_));
 sky130_fd_sc_hd__a22o_1 _8121_ (.A1(\gpio_configure[21][5] ),
    .A2(_3607_),
    .B1(_3571_),
    .B2(_3703_),
    .X(_3704_));
 sky130_fd_sc_hd__a221o_1 _8122_ (.A1(\gpio_configure[9][5] ),
    .A2(_3546_),
    .B1(_3557_),
    .B2(\gpio_configure[13][5] ),
    .C1(_3704_),
    .X(_3705_));
 sky130_fd_sc_hd__a22o_1 _8123_ (.A1(\gpio_configure[17][5] ),
    .A2(_3550_),
    .B1(_3591_),
    .B2(\gpio_configure[14][5] ),
    .X(_3706_));
 sky130_fd_sc_hd__a221o_1 _8124_ (.A1(\gpio_configure[6][5] ),
    .A2(_3621_),
    .B1(_3559_),
    .B2(\gpio_configure[29][5] ),
    .C1(_3706_),
    .X(_3707_));
 sky130_fd_sc_hd__a22o_1 _8125_ (.A1(\gpio_configure[3][5] ),
    .A2(_3511_),
    .B1(_3561_),
    .B2(\gpio_configure[1][5] ),
    .X(_3708_));
 sky130_fd_sc_hd__a221o_1 _8126_ (.A1(\gpio_configure[15][5] ),
    .A2(_3544_),
    .B1(_3565_),
    .B2(\gpio_configure[26][5] ),
    .C1(_3708_),
    .X(_3709_));
 sky130_fd_sc_hd__or4_1 _8127_ (.A(_3702_),
    .B(_3705_),
    .C(_3707_),
    .D(_3709_),
    .X(_3710_));
 sky130_fd_sc_hd__o221a_2 _8128_ (.A1(\gpio_configure[0][5] ),
    .A2(_3597_),
    .B1(_3700_),
    .B2(_3710_),
    .C1(_3689_),
    .X(_3711_));
 sky130_fd_sc_hd__a21o_1 _8129_ (.A1(_1526_),
    .A2(net1495),
    .B1(_3601_),
    .X(_3712_));
 sky130_fd_sc_hd__o22a_1 _8130_ (.A1(net1503),
    .A2(_3604_),
    .B1(_3711_),
    .B2(_3712_),
    .X(_0784_));
 sky130_fd_sc_hd__a22o_1 _8131_ (.A1(\gpio_configure[24][6] ),
    .A2(_3534_),
    .B1(_3568_),
    .B2(\gpio_configure[18][6] ),
    .X(_3713_));
 sky130_fd_sc_hd__a221o_1 _8132_ (.A1(\gpio_configure[23][6] ),
    .A2(_3547_),
    .B1(_3588_),
    .B2(\gpio_configure[10][6] ),
    .C1(_3713_),
    .X(_3714_));
 sky130_fd_sc_hd__a22o_1 _8133_ (.A1(\gpio_configure[12][6] ),
    .A2(_3539_),
    .B1(_3590_),
    .B2(\gpio_configure[14][6] ),
    .X(_3715_));
 sky130_fd_sc_hd__a221o_1 _8134_ (.A1(\gpio_configure[8][6] ),
    .A2(_3527_),
    .B1(_3556_),
    .B2(\gpio_configure[13][6] ),
    .C1(_3715_),
    .X(_3716_));
 sky130_fd_sc_hd__a22o_1 _8135_ (.A1(\gpio_configure[17][6] ),
    .A2(_3549_),
    .B1(_3575_),
    .B2(\gpio_configure[31][6] ),
    .X(_3717_));
 sky130_fd_sc_hd__a221o_1 _8136_ (.A1(\gpio_configure[3][6] ),
    .A2(_3510_),
    .B1(_3584_),
    .B2(\gpio_configure[22][6] ),
    .C1(_3717_),
    .X(_3718_));
 sky130_fd_sc_hd__or2_1 _8137_ (.A(\gpio_configure[16][6] ),
    .B(_3483_),
    .X(_3719_));
 sky130_fd_sc_hd__a22o_1 _8138_ (.A1(\gpio_configure[26][6] ),
    .A2(_3564_),
    .B1(_3719_),
    .B2(_3570_),
    .X(_3720_));
 sky130_fd_sc_hd__a221o_1 _8139_ (.A1(\gpio_configure[4][6] ),
    .A2(_3514_),
    .B1(_3543_),
    .B2(\gpio_configure[15][6] ),
    .C1(_3720_),
    .X(_3721_));
 sky130_fd_sc_hd__or4_1 _8140_ (.A(_3714_),
    .B(_3716_),
    .C(_3718_),
    .D(_3721_),
    .X(_3722_));
 sky130_fd_sc_hd__a22o_1 _8141_ (.A1(\gpio_configure[5][6] ),
    .A2(_3567_),
    .B1(_3581_),
    .B2(\gpio_configure[25][6] ),
    .X(_3723_));
 sky130_fd_sc_hd__a22o_1 _8142_ (.A1(\gpio_configure[9][6] ),
    .A2(_3546_),
    .B1(_3559_),
    .B2(\gpio_configure[29][6] ),
    .X(_3724_));
 sky130_fd_sc_hd__a221o_1 _8143_ (.A1(\gpio_configure[7][6] ),
    .A2(_3537_),
    .B1(_3561_),
    .B2(\gpio_configure[1][6] ),
    .C1(_3724_),
    .X(_3725_));
 sky130_fd_sc_hd__a211o_1 _8144_ (.A1(\gpio_configure[6][6] ),
    .A2(_3621_),
    .B1(_3723_),
    .C1(_3725_),
    .X(_3726_));
 sky130_fd_sc_hd__a22o_1 _8145_ (.A1(\gpio_configure[28][6] ),
    .A2(_3555_),
    .B1(_3587_),
    .B2(\gpio_configure[30][6] ),
    .X(_3727_));
 sky130_fd_sc_hd__a221o_1 _8146_ (.A1(\gpio_configure[2][6] ),
    .A2(_3526_),
    .B1(_3662_),
    .B2(\gpio_configure[20][6] ),
    .C1(_3727_),
    .X(_3728_));
 sky130_fd_sc_hd__a22o_1 _8147_ (.A1(\gpio_configure[27][6] ),
    .A2(_3519_),
    .B1(_3521_),
    .B2(\gpio_configure[19][6] ),
    .X(_3729_));
 sky130_fd_sc_hd__a221o_1 _8148_ (.A1(\gpio_configure[21][6] ),
    .A2(_3607_),
    .B1(_3578_),
    .B2(\gpio_configure[11][6] ),
    .C1(_3729_),
    .X(_3730_));
 sky130_fd_sc_hd__or4_4 _8149_ (.A(_3722_),
    .B(_3726_),
    .C(_3728_),
    .D(_3730_),
    .X(_3731_));
 sky130_fd_sc_hd__o211a_1 _8150_ (.A1(\gpio_configure[0][6] ),
    .A2(_3597_),
    .B1(_3731_),
    .C1(_3689_),
    .X(_3732_));
 sky130_fd_sc_hd__a211o_1 _8151_ (.A1(_1525_),
    .A2(\serial_data_staging_1[5] ),
    .B1(_3600_),
    .C1(_3732_),
    .X(_3733_));
 sky130_fd_sc_hd__o21a_1 _8152_ (.A1(net1482),
    .A2(_3604_),
    .B1(_3733_),
    .X(_0785_));
 sky130_fd_sc_hd__a22o_1 _8153_ (.A1(\gpio_configure[24][7] ),
    .A2(_3535_),
    .B1(_3569_),
    .B2(\gpio_configure[18][7] ),
    .X(_3734_));
 sky130_fd_sc_hd__a221o_1 _8154_ (.A1(\gpio_configure[23][7] ),
    .A2(_3548_),
    .B1(_3589_),
    .B2(\gpio_configure[10][7] ),
    .C1(_3734_),
    .X(_3735_));
 sky130_fd_sc_hd__a22o_2 _8155_ (.A1(\gpio_configure[12][7] ),
    .A2(_3540_),
    .B1(_3591_),
    .B2(\gpio_configure[14][7] ),
    .X(_3736_));
 sky130_fd_sc_hd__a221o_1 _8156_ (.A1(\gpio_configure[8][7] ),
    .A2(_3528_),
    .B1(_3557_),
    .B2(\gpio_configure[13][7] ),
    .C1(_3736_),
    .X(_3737_));
 sky130_fd_sc_hd__a22o_1 _8157_ (.A1(\gpio_configure[17][7] ),
    .A2(_3550_),
    .B1(_3576_),
    .B2(\gpio_configure[31][7] ),
    .X(_3738_));
 sky130_fd_sc_hd__a221o_1 _8158_ (.A1(\gpio_configure[3][7] ),
    .A2(_3511_),
    .B1(_3585_),
    .B2(\gpio_configure[22][7] ),
    .C1(_3738_),
    .X(_3739_));
 sky130_fd_sc_hd__or2_1 _8159_ (.A(\gpio_configure[16][7] ),
    .B(_3484_),
    .X(_3740_));
 sky130_fd_sc_hd__a22o_1 _8160_ (.A1(\gpio_configure[26][7] ),
    .A2(_3565_),
    .B1(_3740_),
    .B2(_3571_),
    .X(_3741_));
 sky130_fd_sc_hd__a221o_1 _8161_ (.A1(\gpio_configure[4][7] ),
    .A2(_3515_),
    .B1(_3544_),
    .B2(\gpio_configure[15][7] ),
    .C1(_3741_),
    .X(_3742_));
 sky130_fd_sc_hd__or4_1 _8162_ (.A(_3735_),
    .B(_3737_),
    .C(_3739_),
    .D(_3742_),
    .X(_3743_));
 sky130_fd_sc_hd__a22o_1 _8163_ (.A1(\gpio_configure[27][7] ),
    .A2(_3519_),
    .B1(_3521_),
    .B2(\gpio_configure[19][7] ),
    .X(_3744_));
 sky130_fd_sc_hd__a22o_1 _8164_ (.A1(\gpio_configure[21][7] ),
    .A2(_3607_),
    .B1(_3578_),
    .B2(\gpio_configure[11][7] ),
    .X(_3745_));
 sky130_fd_sc_hd__a22o_1 _8165_ (.A1(\gpio_configure[5][7] ),
    .A2(_3567_),
    .B1(_3580_),
    .B2(\gpio_configure[25][7] ),
    .X(_3746_));
 sky130_fd_sc_hd__a22o_1 _8166_ (.A1(\gpio_configure[9][7] ),
    .A2(_3545_),
    .B1(_3558_),
    .B2(\gpio_configure[29][7] ),
    .X(_3747_));
 sky130_fd_sc_hd__a221o_1 _8167_ (.A1(\gpio_configure[7][7] ),
    .A2(_3536_),
    .B1(_3560_),
    .B2(\gpio_configure[1][7] ),
    .C1(_3747_),
    .X(_3748_));
 sky130_fd_sc_hd__a211o_1 _8168_ (.A1(\gpio_configure[6][7] ),
    .A2(_3621_),
    .B1(_3746_),
    .C1(_3748_),
    .X(_3749_));
 sky130_fd_sc_hd__a22o_1 _8169_ (.A1(\gpio_configure[28][7] ),
    .A2(_3554_),
    .B1(_3587_),
    .B2(\gpio_configure[30][7] ),
    .X(_3750_));
 sky130_fd_sc_hd__a221o_1 _8170_ (.A1(\gpio_configure[2][7] ),
    .A2(_3526_),
    .B1(_3662_),
    .B2(\gpio_configure[20][7] ),
    .C1(_3750_),
    .X(_3751_));
 sky130_fd_sc_hd__or4_1 _8171_ (.A(_3744_),
    .B(_3745_),
    .C(_3749_),
    .D(_3751_),
    .X(_3752_));
 sky130_fd_sc_hd__o221a_2 _8172_ (.A1(\gpio_configure[0][7] ),
    .A2(_3597_),
    .B1(_3743_),
    .B2(_3752_),
    .C1(_3625_),
    .X(_3753_));
 sky130_fd_sc_hd__a211o_1 _8173_ (.A1(_1525_),
    .A2(net1482),
    .B1(_3600_),
    .C1(_3753_),
    .X(_3754_));
 sky130_fd_sc_hd__o21a_1 _8174_ (.A1(net1488),
    .A2(_3604_),
    .B1(_3754_),
    .X(_0786_));
 sky130_fd_sc_hd__a22o_1 _8175_ (.A1(\gpio_configure[24][8] ),
    .A2(_3534_),
    .B1(_3568_),
    .B2(\gpio_configure[18][8] ),
    .X(_3755_));
 sky130_fd_sc_hd__a221o_1 _8176_ (.A1(\gpio_configure[23][8] ),
    .A2(_3547_),
    .B1(_3588_),
    .B2(\gpio_configure[10][8] ),
    .C1(_3755_),
    .X(_3756_));
 sky130_fd_sc_hd__a22o_1 _8177_ (.A1(\gpio_configure[12][8] ),
    .A2(_3539_),
    .B1(_3590_),
    .B2(\gpio_configure[14][8] ),
    .X(_3757_));
 sky130_fd_sc_hd__a221o_1 _8178_ (.A1(\gpio_configure[8][8] ),
    .A2(_3527_),
    .B1(_3556_),
    .B2(\gpio_configure[13][8] ),
    .C1(_3757_),
    .X(_3758_));
 sky130_fd_sc_hd__a22o_1 _8179_ (.A1(\gpio_configure[17][8] ),
    .A2(_3549_),
    .B1(_3575_),
    .B2(\gpio_configure[31][8] ),
    .X(_3759_));
 sky130_fd_sc_hd__a221o_1 _8180_ (.A1(\gpio_configure[3][8] ),
    .A2(_3510_),
    .B1(_3584_),
    .B2(\gpio_configure[22][8] ),
    .C1(_3759_),
    .X(_3760_));
 sky130_fd_sc_hd__or2_1 _8181_ (.A(\gpio_configure[16][8] ),
    .B(_3483_),
    .X(_3761_));
 sky130_fd_sc_hd__a22o_1 _8182_ (.A1(\gpio_configure[26][8] ),
    .A2(_3564_),
    .B1(_3761_),
    .B2(_3570_),
    .X(_3762_));
 sky130_fd_sc_hd__a221o_1 _8183_ (.A1(\gpio_configure[4][8] ),
    .A2(_3514_),
    .B1(_3543_),
    .B2(\gpio_configure[15][8] ),
    .C1(_3762_),
    .X(_3763_));
 sky130_fd_sc_hd__or4_1 _8184_ (.A(_3756_),
    .B(_3758_),
    .C(_3760_),
    .D(_3763_),
    .X(_3764_));
 sky130_fd_sc_hd__a22o_1 _8185_ (.A1(\gpio_configure[5][8] ),
    .A2(_3566_),
    .B1(_3580_),
    .B2(\gpio_configure[25][8] ),
    .X(_3765_));
 sky130_fd_sc_hd__a22o_1 _8186_ (.A1(\gpio_configure[9][8] ),
    .A2(_3545_),
    .B1(_3558_),
    .B2(\gpio_configure[29][8] ),
    .X(_3766_));
 sky130_fd_sc_hd__a221o_1 _8187_ (.A1(\gpio_configure[7][8] ),
    .A2(_3536_),
    .B1(_3560_),
    .B2(\gpio_configure[1][8] ),
    .C1(_3766_),
    .X(_3767_));
 sky130_fd_sc_hd__a211o_1 _8188_ (.A1(\gpio_configure[6][8] ),
    .A2(_3621_),
    .B1(_3765_),
    .C1(_3767_),
    .X(_3768_));
 sky130_fd_sc_hd__a22o_1 _8189_ (.A1(\gpio_configure[28][8] ),
    .A2(_3554_),
    .B1(_3586_),
    .B2(\gpio_configure[30][8] ),
    .X(_3769_));
 sky130_fd_sc_hd__a221o_1 _8190_ (.A1(\gpio_configure[2][8] ),
    .A2(_3526_),
    .B1(_3662_),
    .B2(\gpio_configure[20][8] ),
    .C1(_3769_),
    .X(_3770_));
 sky130_fd_sc_hd__a22o_1 _8191_ (.A1(\gpio_configure[27][8] ),
    .A2(_3518_),
    .B1(_3521_),
    .B2(\gpio_configure[19][8] ),
    .X(_3771_));
 sky130_fd_sc_hd__a221o_1 _8192_ (.A1(\gpio_configure[21][8] ),
    .A2(_3607_),
    .B1(_3578_),
    .B2(\gpio_configure[11][8] ),
    .C1(_3771_),
    .X(_3772_));
 sky130_fd_sc_hd__or4_2 _8193_ (.A(_3764_),
    .B(_3768_),
    .C(_3770_),
    .D(_3772_),
    .X(_3773_));
 sky130_fd_sc_hd__o21a_1 _8194_ (.A1(\gpio_configure[0][8] ),
    .A2(_3596_),
    .B1(_1546_),
    .X(_3774_));
 sky130_fd_sc_hd__a22o_1 _8195_ (.A1(\xfer_state[1] ),
    .A2(\serial_data_staging_1[7] ),
    .B1(_3773_),
    .B2(_3774_),
    .X(_3775_));
 sky130_fd_sc_hd__mux2_1 _8196_ (.A0(net1511),
    .A1(_3775_),
    .S(_3603_),
    .X(_3776_));
 sky130_fd_sc_hd__clkbuf_1 _8197_ (.A(_3776_),
    .X(_0787_));
 sky130_fd_sc_hd__a22o_1 _8198_ (.A1(\gpio_configure[27][9] ),
    .A2(_3519_),
    .B1(_3578_),
    .B2(\gpio_configure[11][9] ),
    .X(_3777_));
 sky130_fd_sc_hd__a221o_1 _8199_ (.A1(\gpio_configure[19][9] ),
    .A2(_3521_),
    .B1(_3607_),
    .B2(\gpio_configure[21][9] ),
    .C1(_3777_),
    .X(_3778_));
 sky130_fd_sc_hd__a22o_1 _8200_ (.A1(\gpio_configure[24][9] ),
    .A2(_3535_),
    .B1(_3569_),
    .B2(\gpio_configure[18][9] ),
    .X(_3779_));
 sky130_fd_sc_hd__a221o_1 _8201_ (.A1(\gpio_configure[23][9] ),
    .A2(_3548_),
    .B1(_3589_),
    .B2(\gpio_configure[10][9] ),
    .C1(_3779_),
    .X(_3780_));
 sky130_fd_sc_hd__a22o_1 _8202_ (.A1(\gpio_configure[12][9] ),
    .A2(_3540_),
    .B1(_3591_),
    .B2(\gpio_configure[14][9] ),
    .X(_3781_));
 sky130_fd_sc_hd__a221o_1 _8203_ (.A1(\gpio_configure[8][9] ),
    .A2(_3528_),
    .B1(_3557_),
    .B2(\gpio_configure[13][9] ),
    .C1(_3781_),
    .X(_3782_));
 sky130_fd_sc_hd__a22o_1 _8204_ (.A1(\gpio_configure[17][9] ),
    .A2(_3550_),
    .B1(_3576_),
    .B2(\gpio_configure[31][9] ),
    .X(_3783_));
 sky130_fd_sc_hd__a221o_1 _8205_ (.A1(\gpio_configure[3][9] ),
    .A2(_3511_),
    .B1(_3585_),
    .B2(\gpio_configure[22][9] ),
    .C1(_3783_),
    .X(_3784_));
 sky130_fd_sc_hd__or2_1 _8206_ (.A(\gpio_configure[16][9] ),
    .B(_3512_),
    .X(_3785_));
 sky130_fd_sc_hd__a22o_1 _8207_ (.A1(\gpio_configure[26][9] ),
    .A2(_3565_),
    .B1(_3785_),
    .B2(_3570_),
    .X(_3786_));
 sky130_fd_sc_hd__a221o_1 _8208_ (.A1(\gpio_configure[4][9] ),
    .A2(_3515_),
    .B1(_3544_),
    .B2(\gpio_configure[15][9] ),
    .C1(_3786_),
    .X(_3787_));
 sky130_fd_sc_hd__or4_1 _8209_ (.A(_3780_),
    .B(_3782_),
    .C(_3784_),
    .D(_3787_),
    .X(_3788_));
 sky130_fd_sc_hd__a22o_1 _8210_ (.A1(\gpio_configure[5][9] ),
    .A2(_3567_),
    .B1(_3581_),
    .B2(\gpio_configure[25][9] ),
    .X(_3789_));
 sky130_fd_sc_hd__a22o_1 _8211_ (.A1(\gpio_configure[9][9] ),
    .A2(_3546_),
    .B1(_3559_),
    .B2(\gpio_configure[29][9] ),
    .X(_3790_));
 sky130_fd_sc_hd__a221o_1 _8212_ (.A1(\gpio_configure[7][9] ),
    .A2(_3537_),
    .B1(_3561_),
    .B2(\gpio_configure[1][9] ),
    .C1(_3790_),
    .X(_3791_));
 sky130_fd_sc_hd__a211o_1 _8213_ (.A1(\gpio_configure[6][9] ),
    .A2(_3621_),
    .B1(_3789_),
    .C1(_3791_),
    .X(_3792_));
 sky130_fd_sc_hd__a22o_1 _8214_ (.A1(\gpio_configure[28][9] ),
    .A2(_3555_),
    .B1(_3587_),
    .B2(\gpio_configure[30][9] ),
    .X(_3793_));
 sky130_fd_sc_hd__a221o_1 _8215_ (.A1(\gpio_configure[2][9] ),
    .A2(_3526_),
    .B1(_3662_),
    .B2(\gpio_configure[20][9] ),
    .C1(_3793_),
    .X(_3794_));
 sky130_fd_sc_hd__or4_1 _8216_ (.A(_3778_),
    .B(_3788_),
    .C(_3792_),
    .D(_3794_),
    .X(_3795_));
 sky130_fd_sc_hd__o211a_1 _8217_ (.A1(\gpio_configure[0][9] ),
    .A2(_3597_),
    .B1(_3795_),
    .C1(_3689_),
    .X(_3796_));
 sky130_fd_sc_hd__a21o_1 _8218_ (.A1(_1526_),
    .A2(\serial_data_staging_1[8] ),
    .B1(_3601_),
    .X(_3797_));
 sky130_fd_sc_hd__o22a_1 _8219_ (.A1(net1484),
    .A2(_3603_),
    .B1(_3796_),
    .B2(_3797_),
    .X(_0788_));
 sky130_fd_sc_hd__a22o_1 _8220_ (.A1(\gpio_configure[7][10] ),
    .A2(_3537_),
    .B1(_3576_),
    .B2(\gpio_configure[31][10] ),
    .X(_3798_));
 sky130_fd_sc_hd__a221o_1 _8221_ (.A1(\gpio_configure[4][10] ),
    .A2(_3515_),
    .B1(_3589_),
    .B2(\gpio_configure[10][10] ),
    .C1(_3798_),
    .X(_3799_));
 sky130_fd_sc_hd__a22o_1 _8222_ (.A1(\gpio_configure[23][10] ),
    .A2(_3548_),
    .B1(_3569_),
    .B2(\gpio_configure[18][10] ),
    .X(_3800_));
 sky130_fd_sc_hd__a221o_1 _8223_ (.A1(\gpio_configure[15][10] ),
    .A2(_3544_),
    .B1(_3546_),
    .B2(\gpio_configure[9][10] ),
    .C1(_3800_),
    .X(_3801_));
 sky130_fd_sc_hd__and2_1 _8224_ (.A(\gpio_configure[29][10] ),
    .B(_3559_),
    .X(_3802_));
 sky130_fd_sc_hd__a221o_1 _8225_ (.A1(\gpio_configure[27][10] ),
    .A2(_3519_),
    .B1(_3567_),
    .B2(\gpio_configure[5][10] ),
    .C1(_3802_),
    .X(_3803_));
 sky130_fd_sc_hd__a22o_1 _8226_ (.A1(\gpio_configure[13][10] ),
    .A2(_3557_),
    .B1(_3565_),
    .B2(\gpio_configure[26][10] ),
    .X(_3804_));
 sky130_fd_sc_hd__a221o_1 _8227_ (.A1(\gpio_configure[2][10] ),
    .A2(_3526_),
    .B1(_3585_),
    .B2(\gpio_configure[22][10] ),
    .C1(_3804_),
    .X(_3805_));
 sky130_fd_sc_hd__or4_1 _8228_ (.A(_3799_),
    .B(_3801_),
    .C(_3803_),
    .D(_3805_),
    .X(_3806_));
 sky130_fd_sc_hd__a22o_1 _8229_ (.A1(\gpio_configure[3][10] ),
    .A2(_3511_),
    .B1(_3607_),
    .B2(\gpio_configure[21][10] ),
    .X(_3807_));
 sky130_fd_sc_hd__a221o_1 _8230_ (.A1(\gpio_configure[28][10] ),
    .A2(_3555_),
    .B1(_3578_),
    .B2(\gpio_configure[11][10] ),
    .C1(_3807_),
    .X(_3808_));
 sky130_fd_sc_hd__or2_1 _8231_ (.A(\gpio_configure[16][10] ),
    .B(_3484_),
    .X(_3809_));
 sky130_fd_sc_hd__a22o_1 _8232_ (.A1(\gpio_configure[24][10] ),
    .A2(_3535_),
    .B1(_3571_),
    .B2(_3809_),
    .X(_3810_));
 sky130_fd_sc_hd__a221o_1 _8233_ (.A1(\gpio_configure[8][10] ),
    .A2(_3528_),
    .B1(_3581_),
    .B2(\gpio_configure[25][10] ),
    .C1(_3810_),
    .X(_3811_));
 sky130_fd_sc_hd__a22o_1 _8234_ (.A1(\gpio_configure[12][10] ),
    .A2(_3540_),
    .B1(_3591_),
    .B2(\gpio_configure[14][10] ),
    .X(_3812_));
 sky130_fd_sc_hd__a221o_1 _8235_ (.A1(\gpio_configure[17][10] ),
    .A2(_3550_),
    .B1(_3662_),
    .B2(\gpio_configure[20][10] ),
    .C1(_3812_),
    .X(_3813_));
 sky130_fd_sc_hd__a22o_1 _8236_ (.A1(\gpio_configure[19][10] ),
    .A2(_3521_),
    .B1(_3561_),
    .B2(\gpio_configure[1][10] ),
    .X(_3814_));
 sky130_fd_sc_hd__a221o_1 _8237_ (.A1(\gpio_configure[6][10] ),
    .A2(_3621_),
    .B1(_3587_),
    .B2(\gpio_configure[30][10] ),
    .C1(_3814_),
    .X(_3815_));
 sky130_fd_sc_hd__or4_2 _8238_ (.A(_3808_),
    .B(_3811_),
    .C(_3813_),
    .D(_3815_),
    .X(_3816_));
 sky130_fd_sc_hd__o221a_1 _8239_ (.A1(\gpio_configure[0][10] ),
    .A2(_3597_),
    .B1(_3806_),
    .B2(_3816_),
    .C1(_3689_),
    .X(_3817_));
 sky130_fd_sc_hd__a21o_1 _8240_ (.A1(_1526_),
    .A2(net1484),
    .B1(_3601_),
    .X(_3818_));
 sky130_fd_sc_hd__o22a_1 _8241_ (.A1(net1493),
    .A2(_3603_),
    .B1(_3817_),
    .B2(_3818_),
    .X(_0789_));
 sky130_fd_sc_hd__a22o_1 _8242_ (.A1(\gpio_configure[3][11] ),
    .A2(_3511_),
    .B1(_3526_),
    .B2(\gpio_configure[2][11] ),
    .X(_3819_));
 sky130_fd_sc_hd__a221o_1 _8243_ (.A1(\gpio_configure[25][11] ),
    .A2(_3581_),
    .B1(_3587_),
    .B2(\gpio_configure[30][11] ),
    .C1(_3819_),
    .X(_3820_));
 sky130_fd_sc_hd__a22o_1 _8244_ (.A1(\gpio_configure[7][11] ),
    .A2(_3537_),
    .B1(_3589_),
    .B2(\gpio_configure[10][11] ),
    .X(_3821_));
 sky130_fd_sc_hd__a221o_1 _8245_ (.A1(\gpio_configure[5][11] ),
    .A2(_3567_),
    .B1(_3662_),
    .B2(\gpio_configure[20][11] ),
    .C1(_3821_),
    .X(_3822_));
 sky130_fd_sc_hd__a22o_1 _8246_ (.A1(\gpio_configure[24][11] ),
    .A2(_3535_),
    .B1(_3585_),
    .B2(\gpio_configure[22][11] ),
    .X(_3823_));
 sky130_fd_sc_hd__a22o_1 _8247_ (.A1(\gpio_configure[13][11] ),
    .A2(_3557_),
    .B1(_3569_),
    .B2(\gpio_configure[18][11] ),
    .X(_3824_));
 sky130_fd_sc_hd__a221o_1 _8248_ (.A1(\gpio_configure[23][11] ),
    .A2(_3548_),
    .B1(_3576_),
    .B2(\gpio_configure[31][11] ),
    .C1(_3824_),
    .X(_3825_));
 sky130_fd_sc_hd__a211o_1 _8249_ (.A1(\gpio_configure[15][11] ),
    .A2(_3544_),
    .B1(_3823_),
    .C1(_3825_),
    .X(_3826_));
 sky130_fd_sc_hd__or3_1 _8250_ (.A(_3820_),
    .B(_3822_),
    .C(_3826_),
    .X(_3827_));
 sky130_fd_sc_hd__a22o_1 _8251_ (.A1(\gpio_configure[12][11] ),
    .A2(_3540_),
    .B1(_3561_),
    .B2(\gpio_configure[1][11] ),
    .X(_3828_));
 sky130_fd_sc_hd__a221o_1 _8252_ (.A1(\gpio_configure[19][11] ),
    .A2(_3521_),
    .B1(_3607_),
    .B2(\gpio_configure[21][11] ),
    .C1(_3828_),
    .X(_3829_));
 sky130_fd_sc_hd__or2_1 _8253_ (.A(\gpio_configure[16][11] ),
    .B(_3484_),
    .X(_3830_));
 sky130_fd_sc_hd__a22o_1 _8254_ (.A1(\gpio_configure[28][11] ),
    .A2(_3555_),
    .B1(_3571_),
    .B2(_3830_),
    .X(_3831_));
 sky130_fd_sc_hd__a221o_1 _8255_ (.A1(\gpio_configure[27][11] ),
    .A2(_3519_),
    .B1(_3621_),
    .B2(\gpio_configure[6][11] ),
    .C1(_3831_),
    .X(_3832_));
 sky130_fd_sc_hd__a22o_1 _8256_ (.A1(\gpio_configure[9][11] ),
    .A2(_3546_),
    .B1(_3559_),
    .B2(\gpio_configure[29][11] ),
    .X(_3833_));
 sky130_fd_sc_hd__a221o_1 _8257_ (.A1(\gpio_configure[4][11] ),
    .A2(_3515_),
    .B1(_3578_),
    .B2(\gpio_configure[11][11] ),
    .C1(_3833_),
    .X(_3834_));
 sky130_fd_sc_hd__a22o_1 _8258_ (.A1(\gpio_configure[17][11] ),
    .A2(_3550_),
    .B1(_3565_),
    .B2(\gpio_configure[26][11] ),
    .X(_3835_));
 sky130_fd_sc_hd__a221o_1 _8259_ (.A1(\gpio_configure[8][11] ),
    .A2(_3528_),
    .B1(_3591_),
    .B2(\gpio_configure[14][11] ),
    .C1(_3835_),
    .X(_3836_));
 sky130_fd_sc_hd__or4_1 _8260_ (.A(_3829_),
    .B(_3832_),
    .C(_3834_),
    .D(_3836_),
    .X(_3837_));
 sky130_fd_sc_hd__o221a_1 _8261_ (.A1(\gpio_configure[0][11] ),
    .A2(_3597_),
    .B1(_3827_),
    .B2(_3837_),
    .C1(_3689_),
    .X(_3838_));
 sky130_fd_sc_hd__a21o_1 _8262_ (.A1(_1526_),
    .A2(\serial_data_staging_1[10] ),
    .B1(_3601_),
    .X(_3839_));
 sky130_fd_sc_hd__o22a_1 _8263_ (.A1(net1491),
    .A2(_3603_),
    .B1(_3838_),
    .B2(_3839_),
    .X(_0790_));
 sky130_fd_sc_hd__a22o_1 _8264_ (.A1(\gpio_configure[5][12] ),
    .A2(_3566_),
    .B1(_3580_),
    .B2(\gpio_configure[25][12] ),
    .X(_3840_));
 sky130_fd_sc_hd__a221o_1 _8265_ (.A1(\gpio_configure[31][12] ),
    .A2(_3576_),
    .B1(_3578_),
    .B2(\gpio_configure[11][12] ),
    .C1(_3840_),
    .X(_3841_));
 sky130_fd_sc_hd__a22o_1 _8266_ (.A1(\gpio_configure[19][12] ),
    .A2(_3520_),
    .B1(_3587_),
    .B2(\gpio_configure[30][12] ),
    .X(_3842_));
 sky130_fd_sc_hd__a221o_1 _8267_ (.A1(\gpio_configure[4][12] ),
    .A2(_3515_),
    .B1(_3544_),
    .B2(\gpio_configure[15][12] ),
    .C1(_3842_),
    .X(_3843_));
 sky130_fd_sc_hd__a22o_1 _8268_ (.A1(\gpio_configure[9][12] ),
    .A2(_3546_),
    .B1(_3589_),
    .B2(\gpio_configure[10][12] ),
    .X(_3844_));
 sky130_fd_sc_hd__a21o_1 _8269_ (.A1(\gpio_configure[27][12] ),
    .A2(_3519_),
    .B1(_3844_),
    .X(_3845_));
 sky130_fd_sc_hd__a22o_1 _8270_ (.A1(\gpio_configure[7][12] ),
    .A2(_3537_),
    .B1(_3550_),
    .B2(\gpio_configure[17][12] ),
    .X(_3846_));
 sky130_fd_sc_hd__a221o_1 _8271_ (.A1(\gpio_configure[23][12] ),
    .A2(_3548_),
    .B1(_3555_),
    .B2(\gpio_configure[28][12] ),
    .C1(_3846_),
    .X(_3847_));
 sky130_fd_sc_hd__or4_1 _8272_ (.A(_3841_),
    .B(_3843_),
    .C(_3845_),
    .D(_3847_),
    .X(_3848_));
 sky130_fd_sc_hd__a22o_1 _8273_ (.A1(\gpio_configure[29][12] ),
    .A2(_3559_),
    .B1(_3569_),
    .B2(\gpio_configure[18][12] ),
    .X(_3849_));
 sky130_fd_sc_hd__a221o_1 _8274_ (.A1(\gpio_configure[8][12] ),
    .A2(_3528_),
    .B1(_3585_),
    .B2(\gpio_configure[22][12] ),
    .C1(_3849_),
    .X(_3850_));
 sky130_fd_sc_hd__or2_1 _8275_ (.A(\gpio_configure[16][12] ),
    .B(_3484_),
    .X(_3851_));
 sky130_fd_sc_hd__a22o_1 _8276_ (.A1(\gpio_configure[6][12] ),
    .A2(_3531_),
    .B1(_3571_),
    .B2(_3851_),
    .X(_3852_));
 sky130_fd_sc_hd__a221o_1 _8277_ (.A1(\gpio_configure[24][12] ),
    .A2(_3535_),
    .B1(_3561_),
    .B2(\gpio_configure[1][12] ),
    .C1(_3852_),
    .X(_3853_));
 sky130_fd_sc_hd__a22o_1 _8278_ (.A1(\gpio_configure[2][12] ),
    .A2(_3525_),
    .B1(_3565_),
    .B2(\gpio_configure[26][12] ),
    .X(_3854_));
 sky130_fd_sc_hd__a221o_1 _8279_ (.A1(\gpio_configure[21][12] ),
    .A2(_3607_),
    .B1(_3591_),
    .B2(\gpio_configure[14][12] ),
    .C1(_3854_),
    .X(_3855_));
 sky130_fd_sc_hd__a22o_1 _8280_ (.A1(\gpio_configure[3][12] ),
    .A2(_3511_),
    .B1(_3540_),
    .B2(\gpio_configure[12][12] ),
    .X(_3856_));
 sky130_fd_sc_hd__a221o_1 _8281_ (.A1(\gpio_configure[13][12] ),
    .A2(_3557_),
    .B1(_3662_),
    .B2(\gpio_configure[20][12] ),
    .C1(_3856_),
    .X(_3857_));
 sky130_fd_sc_hd__or4_1 _8282_ (.A(_3850_),
    .B(_3853_),
    .C(_3855_),
    .D(_3857_),
    .X(_3858_));
 sky130_fd_sc_hd__o221a_1 _8283_ (.A1(\gpio_configure[0][12] ),
    .A2(_3596_),
    .B1(_3848_),
    .B2(_3858_),
    .C1(_3625_),
    .X(_3859_));
 sky130_fd_sc_hd__a211o_1 _8284_ (.A1(_1525_),
    .A2(\serial_data_staging_1[11] ),
    .B1(_3600_),
    .C1(_3859_),
    .X(_3860_));
 sky130_fd_sc_hd__o21a_1 _8285_ (.A1(\serial_data_staging_1[12] ),
    .A2(_3604_),
    .B1(_3860_),
    .X(_0791_));
 sky130_fd_sc_hd__nor2_2 _8286_ (.A(\pad_count_2[4] ),
    .B(\pad_count_2[5] ),
    .Y(_3861_));
 sky130_fd_sc_hd__nor2_4 _8287_ (.A(\pad_count_2[3] ),
    .B(\pad_count_2[2] ),
    .Y(_3862_));
 sky130_fd_sc_hd__and3_2 _8288_ (.A(_3493_),
    .B(_3861_),
    .C(_3862_),
    .X(_3863_));
 sky130_fd_sc_hd__buf_6 _8289_ (.A(_3863_),
    .X(_3864_));
 sky130_fd_sc_hd__and2b_1 _8290_ (.A_N(\pad_count_2[2] ),
    .B(\pad_count_2[3] ),
    .X(_3865_));
 sky130_fd_sc_hd__and3_2 _8291_ (.A(_3488_),
    .B(_3498_),
    .C(_3865_),
    .X(_3866_));
 sky130_fd_sc_hd__buf_6 _8292_ (.A(_3866_),
    .X(_3867_));
 sky130_fd_sc_hd__and3_2 _8293_ (.A(_3488_),
    .B(_3491_),
    .C(_3861_),
    .X(_3868_));
 sky130_fd_sc_hd__buf_6 _8294_ (.A(_3868_),
    .X(_3869_));
 sky130_fd_sc_hd__nand2b_4 _8295_ (.A_N(\pad_count_2[5] ),
    .B(\pad_count_2[4] ),
    .Y(_3870_));
 sky130_fd_sc_hd__nand2_2 _8296_ (.A(_1528_),
    .B(_3862_),
    .Y(_3871_));
 sky130_fd_sc_hd__nor2_2 _8297_ (.A(_3870_),
    .B(_3871_),
    .Y(_3872_));
 sky130_fd_sc_hd__buf_8 _8298_ (.A(_3872_),
    .X(_3873_));
 sky130_fd_sc_hd__nor2_2 _8299_ (.A(\pad_count_2[1] ),
    .B(\pad_count_2[0] ),
    .Y(_3874_));
 sky130_fd_sc_hd__and3b_4 _8300_ (.A_N(_1527_),
    .B(_3862_),
    .C(_3874_),
    .X(_3875_));
 sky130_fd_sc_hd__buf_6 _8301_ (.A(_3875_),
    .X(_3876_));
 sky130_fd_sc_hd__buf_2 _8302_ (.A(_3498_),
    .X(_3877_));
 sky130_fd_sc_hd__and3_2 _8303_ (.A(_1528_),
    .B(_3877_),
    .C(_3865_),
    .X(_3878_));
 sky130_fd_sc_hd__buf_6 _8304_ (.A(_3878_),
    .X(_3879_));
 sky130_fd_sc_hd__a22o_1 _8305_ (.A1(\gpio_configure[32][0] ),
    .A2(_3876_),
    .B1(_3879_),
    .B2(\gpio_configure[26][0] ),
    .X(_3880_));
 sky130_fd_sc_hd__a221o_1 _8306_ (.A1(\gpio_configure[13][0] ),
    .A2(_3869_),
    .B1(_3873_),
    .B2(\gpio_configure[18][0] ),
    .C1(_3880_),
    .X(_3881_));
 sky130_fd_sc_hd__a221o_1 _8307_ (.A1(\gpio_configure[3][0] ),
    .A2(_3864_),
    .B1(_3867_),
    .B2(\gpio_configure[25][0] ),
    .C1(_3881_),
    .X(_3882_));
 sky130_fd_sc_hd__nand2_4 _8308_ (.A(_3488_),
    .B(_3862_),
    .Y(_3883_));
 sky130_fd_sc_hd__nor2_8 _8309_ (.A(_1527_),
    .B(_3883_),
    .Y(_3884_));
 sky130_fd_sc_hd__buf_6 _8310_ (.A(_3884_),
    .X(_3885_));
 sky130_fd_sc_hd__and3b_4 _8311_ (.A_N(_1527_),
    .B(_3493_),
    .C(_3862_),
    .X(_3886_));
 sky130_fd_sc_hd__buf_6 _8312_ (.A(_3886_),
    .X(_3887_));
 sky130_fd_sc_hd__and3_4 _8313_ (.A(_1528_),
    .B(_3491_),
    .C(_3861_),
    .X(_3888_));
 sky130_fd_sc_hd__buf_6 _8314_ (.A(_3888_),
    .X(_3889_));
 sky130_fd_sc_hd__and3_2 _8315_ (.A(_3491_),
    .B(_3861_),
    .C(_3874_),
    .X(_3890_));
 sky130_fd_sc_hd__buf_6 _8316_ (.A(_3890_),
    .X(_3891_));
 sky130_fd_sc_hd__a22o_1 _8317_ (.A1(\gpio_configure[14][0] ),
    .A2(_3889_),
    .B1(_3891_),
    .B2(\gpio_configure[12][0] ),
    .X(_3892_));
 sky130_fd_sc_hd__a221o_1 _8318_ (.A1(\gpio_configure[33][0] ),
    .A2(_3885_),
    .B1(_3887_),
    .B2(\gpio_configure[35][0] ),
    .C1(_3892_),
    .X(_3893_));
 sky130_fd_sc_hd__or2_1 _8319_ (.A(\pad_count_2[4] ),
    .B(\pad_count_2[5] ),
    .X(_3894_));
 sky130_fd_sc_hd__buf_2 _8320_ (.A(_3894_),
    .X(_3895_));
 sky130_fd_sc_hd__nor2_2 _8321_ (.A(_1530_),
    .B(_3895_),
    .Y(_3896_));
 sky130_fd_sc_hd__buf_8 _8322_ (.A(_3896_),
    .X(_3897_));
 sky130_fd_sc_hd__and3_2 _8323_ (.A(_1529_),
    .B(_3493_),
    .C(_3861_),
    .X(_3898_));
 sky130_fd_sc_hd__buf_6 _8324_ (.A(_3898_),
    .X(_3899_));
 sky130_fd_sc_hd__and3_4 _8325_ (.A(_3488_),
    .B(_3491_),
    .C(_3877_),
    .X(_3900_));
 sky130_fd_sc_hd__and3_2 _8326_ (.A(_3488_),
    .B(_3861_),
    .C(_3865_),
    .X(_3901_));
 sky130_fd_sc_hd__buf_8 _8327_ (.A(_3901_),
    .X(_3902_));
 sky130_fd_sc_hd__a22o_1 _8328_ (.A1(\gpio_configure[29][0] ),
    .A2(_3900_),
    .B1(_3902_),
    .B2(\gpio_configure[9][0] ),
    .X(_3903_));
 sky130_fd_sc_hd__a221o_1 _8329_ (.A1(\gpio_configure[6][0] ),
    .A2(_3897_),
    .B1(_3899_),
    .B2(\gpio_configure[7][0] ),
    .C1(_3903_),
    .X(_3904_));
 sky130_fd_sc_hd__and3_2 _8330_ (.A(_3493_),
    .B(_3877_),
    .C(_3865_),
    .X(_3905_));
 sky130_fd_sc_hd__buf_6 _8331_ (.A(_3905_),
    .X(_3906_));
 sky130_fd_sc_hd__and3_2 _8332_ (.A(_1528_),
    .B(_3861_),
    .C(_3865_),
    .X(_3907_));
 sky130_fd_sc_hd__buf_8 _8333_ (.A(_3907_),
    .X(_3908_));
 sky130_fd_sc_hd__and3_2 _8334_ (.A(_3493_),
    .B(_3861_),
    .C(_3865_),
    .X(_3909_));
 sky130_fd_sc_hd__buf_8 _8335_ (.A(_3909_),
    .X(_3910_));
 sky130_fd_sc_hd__and3_2 _8336_ (.A(_3498_),
    .B(_3865_),
    .C(_3874_),
    .X(_3911_));
 sky130_fd_sc_hd__buf_8 _8337_ (.A(_3911_),
    .X(_3912_));
 sky130_fd_sc_hd__a22o_1 _8338_ (.A1(\gpio_configure[11][0] ),
    .A2(_3910_),
    .B1(_3912_),
    .B2(\gpio_configure[24][0] ),
    .X(_3913_));
 sky130_fd_sc_hd__a221o_1 _8339_ (.A1(\gpio_configure[27][0] ),
    .A2(_3906_),
    .B1(_3908_),
    .B2(\gpio_configure[10][0] ),
    .C1(_3913_),
    .X(_3914_));
 sky130_fd_sc_hd__and3_2 _8340_ (.A(_3493_),
    .B(_3491_),
    .C(_3861_),
    .X(_3915_));
 sky130_fd_sc_hd__buf_6 _8341_ (.A(_3915_),
    .X(_3916_));
 sky130_fd_sc_hd__nand2_2 _8342_ (.A(_1529_),
    .B(_3488_),
    .Y(_3917_));
 sky130_fd_sc_hd__nor2_4 _8343_ (.A(_1527_),
    .B(_3917_),
    .Y(_3918_));
 sky130_fd_sc_hd__buf_4 _8344_ (.A(_3918_),
    .X(_3919_));
 sky130_fd_sc_hd__and3_4 _8345_ (.A(_1529_),
    .B(_3493_),
    .C(_3877_),
    .X(_3920_));
 sky130_fd_sc_hd__buf_8 _8346_ (.A(_3920_),
    .X(_3921_));
 sky130_fd_sc_hd__nor2_4 _8347_ (.A(_1527_),
    .B(_3871_),
    .Y(_3922_));
 sky130_fd_sc_hd__buf_6 _8348_ (.A(_3922_),
    .X(_3923_));
 sky130_fd_sc_hd__a22o_1 _8349_ (.A1(\gpio_configure[23][0] ),
    .A2(_3921_),
    .B1(_3923_),
    .B2(\gpio_configure[34][0] ),
    .X(_3924_));
 sky130_fd_sc_hd__a221o_1 _8350_ (.A1(\gpio_configure[15][0] ),
    .A2(_3916_),
    .B1(_3919_),
    .B2(\gpio_configure[37][0] ),
    .C1(_3924_),
    .X(_3925_));
 sky130_fd_sc_hd__or4_1 _8351_ (.A(_3893_),
    .B(_3904_),
    .C(_3914_),
    .D(_3925_),
    .X(_3926_));
 sky130_fd_sc_hd__nand2_2 _8352_ (.A(_1529_),
    .B(_3874_),
    .Y(_3927_));
 sky130_fd_sc_hd__nor2_4 _8353_ (.A(_3895_),
    .B(_3927_),
    .Y(_3928_));
 sky130_fd_sc_hd__or4_1 _8354_ (.A(_3886_),
    .B(_3888_),
    .C(_3898_),
    .D(_3928_),
    .X(_3929_));
 sky130_fd_sc_hd__nor2_4 _8355_ (.A(_1527_),
    .B(_3927_),
    .Y(_3930_));
 sky130_fd_sc_hd__or4_1 _8356_ (.A(_3863_),
    .B(_3896_),
    .C(_3918_),
    .D(_3930_),
    .X(_3931_));
 sky130_fd_sc_hd__and3_2 _8357_ (.A(_3861_),
    .B(_3865_),
    .C(_3874_),
    .X(_3932_));
 sky130_fd_sc_hd__or4_1 _8358_ (.A(_3868_),
    .B(_3890_),
    .C(_3909_),
    .D(_3932_),
    .X(_3933_));
 sky130_fd_sc_hd__nor2_2 _8359_ (.A(_3895_),
    .B(_3871_),
    .Y(_3934_));
 sky130_fd_sc_hd__or4_1 _8360_ (.A(_3884_),
    .B(_3915_),
    .C(_3922_),
    .D(_3934_),
    .X(_3935_));
 sky130_fd_sc_hd__or4_1 _8361_ (.A(_3929_),
    .B(_3931_),
    .C(_3933_),
    .D(_3935_),
    .X(_3936_));
 sky130_fd_sc_hd__nor2_2 _8362_ (.A(_3895_),
    .B(_3917_),
    .Y(_3937_));
 sky130_fd_sc_hd__nor2_2 _8363_ (.A(_3895_),
    .B(_3883_),
    .Y(_3938_));
 sky130_fd_sc_hd__or4_1 _8364_ (.A(_3901_),
    .B(_3907_),
    .C(_3937_),
    .D(_3938_),
    .X(_3939_));
 sky130_fd_sc_hd__nor4_1 _8365_ (.A(_3877_),
    .B(_3876_),
    .C(_3936_),
    .D(_3939_),
    .Y(_3940_));
 sky130_fd_sc_hd__clkbuf_8 _8366_ (.A(net393),
    .X(_3941_));
 sky130_fd_sc_hd__clkbuf_8 _8367_ (.A(_3930_),
    .X(_3942_));
 sky130_fd_sc_hd__nor2_4 _8368_ (.A(_3870_),
    .B(_3883_),
    .Y(_3943_));
 sky130_fd_sc_hd__buf_6 _8369_ (.A(_3943_),
    .X(_3944_));
 sky130_fd_sc_hd__buf_6 _8370_ (.A(_3932_),
    .X(_3945_));
 sky130_fd_sc_hd__and3_4 _8371_ (.A(_3877_),
    .B(_3862_),
    .C(_3874_),
    .X(_3946_));
 sky130_fd_sc_hd__buf_6 _8372_ (.A(_3946_),
    .X(_3947_));
 sky130_fd_sc_hd__a22o_1 _8373_ (.A1(\gpio_configure[8][0] ),
    .A2(_3945_),
    .B1(_3947_),
    .B2(\gpio_configure[16][0] ),
    .X(_3948_));
 sky130_fd_sc_hd__a221o_1 _8374_ (.A1(\gpio_configure[36][0] ),
    .A2(_3942_),
    .B1(_3944_),
    .B2(\gpio_configure[17][0] ),
    .C1(_3948_),
    .X(_3949_));
 sky130_fd_sc_hd__and3_4 _8375_ (.A(_1528_),
    .B(_3491_),
    .C(_3877_),
    .X(_3950_));
 sky130_fd_sc_hd__buf_6 _8376_ (.A(_3950_),
    .X(_3951_));
 sky130_fd_sc_hd__nor2_4 _8377_ (.A(_3870_),
    .B(_3917_),
    .Y(_3952_));
 sky130_fd_sc_hd__buf_6 _8378_ (.A(_3952_),
    .X(_3953_));
 sky130_fd_sc_hd__buf_8 _8379_ (.A(_3934_),
    .X(_3954_));
 sky130_fd_sc_hd__nor2_8 _8380_ (.A(_1530_),
    .B(_3870_),
    .Y(_3955_));
 sky130_fd_sc_hd__buf_8 _8381_ (.A(_3955_),
    .X(_3956_));
 sky130_fd_sc_hd__a22o_1 _8382_ (.A1(\gpio_configure[2][0] ),
    .A2(_3954_),
    .B1(_3956_),
    .B2(\gpio_configure[22][0] ),
    .X(_3957_));
 sky130_fd_sc_hd__a221o_1 _8383_ (.A1(\gpio_configure[30][0] ),
    .A2(_3951_),
    .B1(_3953_),
    .B2(\gpio_configure[21][0] ),
    .C1(_3957_),
    .X(_3958_));
 sky130_fd_sc_hd__buf_8 _8384_ (.A(_3938_),
    .X(_3959_));
 sky130_fd_sc_hd__nor2_4 _8385_ (.A(_3870_),
    .B(_3927_),
    .Y(_3960_));
 sky130_fd_sc_hd__buf_6 _8386_ (.A(_3960_),
    .X(_3961_));
 sky130_fd_sc_hd__a22o_1 _8387_ (.A1(\gpio_configure[1][0] ),
    .A2(_3959_),
    .B1(_3961_),
    .B2(\gpio_configure[20][0] ),
    .X(_3962_));
 sky130_fd_sc_hd__buf_8 _8388_ (.A(_3937_),
    .X(_3963_));
 sky130_fd_sc_hd__and3_4 _8389_ (.A(_3491_),
    .B(_3877_),
    .C(_3874_),
    .X(_3964_));
 sky130_fd_sc_hd__buf_6 _8390_ (.A(_3964_),
    .X(_3965_));
 sky130_fd_sc_hd__buf_4 _8391_ (.A(_3928_),
    .X(_3966_));
 sky130_fd_sc_hd__and3_4 _8392_ (.A(_3493_),
    .B(_3877_),
    .C(_3862_),
    .X(_3967_));
 sky130_fd_sc_hd__a22o_1 _8393_ (.A1(\gpio_configure[4][0] ),
    .A2(_3966_),
    .B1(_3967_),
    .B2(\gpio_configure[19][0] ),
    .X(_3968_));
 sky130_fd_sc_hd__a221o_1 _8394_ (.A1(\gpio_configure[5][0] ),
    .A2(_3963_),
    .B1(_3965_),
    .B2(\gpio_configure[28][0] ),
    .C1(_3968_),
    .X(_3969_));
 sky130_fd_sc_hd__a211o_1 _8395_ (.A1(\gpio_configure[31][0] ),
    .A2(_3500_),
    .B1(_3962_),
    .C1(_3969_),
    .X(_3970_));
 sky130_fd_sc_hd__or4_1 _8396_ (.A(_3941_),
    .B(_3949_),
    .C(_3958_),
    .D(_3970_),
    .X(_3971_));
 sky130_fd_sc_hd__or3_2 _8397_ (.A(_3882_),
    .B(_3926_),
    .C(_3971_),
    .X(_3972_));
 sky130_fd_sc_hd__or4_4 _8398_ (.A(_3877_),
    .B(_3876_),
    .C(_3936_),
    .D(_3939_),
    .X(_3973_));
 sky130_fd_sc_hd__buf_6 _8399_ (.A(_3973_),
    .X(_3974_));
 sky130_fd_sc_hd__or2_1 _8400_ (.A(\gpio_configure[0][0] ),
    .B(_3974_),
    .X(_3975_));
 sky130_fd_sc_hd__a32o_1 _8401_ (.A1(_3508_),
    .A2(_3972_),
    .A3(_3975_),
    .B1(_3601_),
    .B2(net1452),
    .X(_0792_));
 sky130_fd_sc_hd__buf_8 _8402_ (.A(_3900_),
    .X(_3976_));
 sky130_fd_sc_hd__a22o_1 _8403_ (.A1(\gpio_configure[35][1] ),
    .A2(_3887_),
    .B1(_3951_),
    .B2(\gpio_configure[30][1] ),
    .X(_3977_));
 sky130_fd_sc_hd__a221o_2 _8404_ (.A1(\gpio_configure[29][1] ),
    .A2(_3976_),
    .B1(_3953_),
    .B2(\gpio_configure[21][1] ),
    .C1(_3977_),
    .X(_3978_));
 sky130_fd_sc_hd__a22o_1 _8405_ (.A1(\gpio_configure[23][1] ),
    .A2(_3921_),
    .B1(_3961_),
    .B2(\gpio_configure[20][1] ),
    .X(_3979_));
 sky130_fd_sc_hd__a22o_1 _8406_ (.A1(\gpio_configure[18][1] ),
    .A2(_3873_),
    .B1(_3945_),
    .B2(\gpio_configure[8][1] ),
    .X(_3980_));
 sky130_fd_sc_hd__a221o_1 _8407_ (.A1(\gpio_configure[33][1] ),
    .A2(_3885_),
    .B1(_3956_),
    .B2(\gpio_configure[22][1] ),
    .C1(_3980_),
    .X(_3981_));
 sky130_fd_sc_hd__a22o_1 _8408_ (.A1(\gpio_configure[14][1] ),
    .A2(_3889_),
    .B1(_3906_),
    .B2(\gpio_configure[27][1] ),
    .X(_3982_));
 sky130_fd_sc_hd__a221o_1 _8409_ (.A1(\gpio_configure[16][1] ),
    .A2(_3947_),
    .B1(_3944_),
    .B2(\gpio_configure[17][1] ),
    .C1(_3982_),
    .X(_3983_));
 sky130_fd_sc_hd__a2111o_2 _8410_ (.A1(\gpio_configure[28][1] ),
    .A2(_3965_),
    .B1(_3979_),
    .C1(_3981_),
    .D1(_3983_),
    .X(_3984_));
 sky130_fd_sc_hd__buf_6 _8411_ (.A(_3967_),
    .X(_3985_));
 sky130_fd_sc_hd__a22o_1 _8412_ (.A1(\gpio_configure[4][1] ),
    .A2(_3928_),
    .B1(_3930_),
    .B2(\gpio_configure[36][1] ),
    .X(_3986_));
 sky130_fd_sc_hd__a221o_1 _8413_ (.A1(\gpio_configure[32][1] ),
    .A2(_3875_),
    .B1(_3919_),
    .B2(\gpio_configure[37][1] ),
    .C1(_3986_),
    .X(_3987_));
 sky130_fd_sc_hd__a221o_1 _8414_ (.A1(\gpio_configure[34][1] ),
    .A2(_3923_),
    .B1(_3985_),
    .B2(\gpio_configure[19][1] ),
    .C1(_3987_),
    .X(_3988_));
 sky130_fd_sc_hd__a22o_1 _8415_ (.A1(\gpio_configure[12][1] ),
    .A2(_3890_),
    .B1(_3901_),
    .B2(\gpio_configure[9][1] ),
    .X(_3989_));
 sky130_fd_sc_hd__a221o_1 _8416_ (.A1(\gpio_configure[6][1] ),
    .A2(_3896_),
    .B1(_3907_),
    .B2(\gpio_configure[10][1] ),
    .C1(_3989_),
    .X(_3990_));
 sky130_fd_sc_hd__a22o_1 _8417_ (.A1(\gpio_configure[25][1] ),
    .A2(_3867_),
    .B1(_3869_),
    .B2(\gpio_configure[13][1] ),
    .X(_3991_));
 sky130_fd_sc_hd__a221o_1 _8418_ (.A1(\gpio_configure[5][1] ),
    .A2(_3963_),
    .B1(_3954_),
    .B2(\gpio_configure[2][1] ),
    .C1(_3991_),
    .X(_3992_));
 sky130_fd_sc_hd__a22o_1 _8419_ (.A1(\gpio_configure[31][1] ),
    .A2(_3499_),
    .B1(_3910_),
    .B2(\gpio_configure[11][1] ),
    .X(_3993_));
 sky130_fd_sc_hd__a221o_1 _8420_ (.A1(\gpio_configure[24][1] ),
    .A2(_3912_),
    .B1(_3959_),
    .B2(\gpio_configure[1][1] ),
    .C1(_3993_),
    .X(_3994_));
 sky130_fd_sc_hd__a22o_1 _8421_ (.A1(\gpio_configure[26][1] ),
    .A2(_3878_),
    .B1(_3898_),
    .B2(\gpio_configure[7][1] ),
    .X(_3995_));
 sky130_fd_sc_hd__a221o_1 _8422_ (.A1(\gpio_configure[3][1] ),
    .A2(_3864_),
    .B1(_3916_),
    .B2(\gpio_configure[15][1] ),
    .C1(_3995_),
    .X(_3996_));
 sky130_fd_sc_hd__or4_1 _8423_ (.A(_3990_),
    .B(_3992_),
    .C(_3994_),
    .D(_3996_),
    .X(_3997_));
 sky130_fd_sc_hd__or3_1 _8424_ (.A(_3941_),
    .B(_3988_),
    .C(_3997_),
    .X(_3998_));
 sky130_fd_sc_hd__o32a_1 _8425_ (.A1(_3978_),
    .A2(_3984_),
    .A3(_3998_),
    .B1(_3974_),
    .B2(\gpio_configure[0][1] ),
    .X(_3999_));
 sky130_fd_sc_hd__mux2_1 _8426_ (.A0(\serial_data_staging_2[0] ),
    .A1(_3999_),
    .S(_3625_),
    .X(_4000_));
 sky130_fd_sc_hd__mux2_1 _8427_ (.A0(net1508),
    .A1(_4000_),
    .S(_3602_),
    .X(_4001_));
 sky130_fd_sc_hd__clkbuf_1 _8428_ (.A(_4001_),
    .X(_0793_));
 sky130_fd_sc_hd__a22o_1 _8429_ (.A1(\gpio_configure[35][2] ),
    .A2(_3887_),
    .B1(_3951_),
    .B2(\gpio_configure[30][2] ),
    .X(_4002_));
 sky130_fd_sc_hd__a221o_1 _8430_ (.A1(\gpio_configure[29][2] ),
    .A2(_3976_),
    .B1(_3953_),
    .B2(\gpio_configure[21][2] ),
    .C1(_4002_),
    .X(_4003_));
 sky130_fd_sc_hd__and2_1 _8431_ (.A(\gpio_configure[28][2] ),
    .B(_3965_),
    .X(_4004_));
 sky130_fd_sc_hd__a221o_1 _8432_ (.A1(\gpio_configure[23][2] ),
    .A2(_3921_),
    .B1(_3961_),
    .B2(\gpio_configure[20][2] ),
    .C1(_4004_),
    .X(_4005_));
 sky130_fd_sc_hd__a22o_1 _8433_ (.A1(\gpio_configure[18][2] ),
    .A2(_3873_),
    .B1(_3945_),
    .B2(\gpio_configure[8][2] ),
    .X(_4006_));
 sky130_fd_sc_hd__a221o_1 _8434_ (.A1(\gpio_configure[33][2] ),
    .A2(_3885_),
    .B1(_3956_),
    .B2(\gpio_configure[22][2] ),
    .C1(_4006_),
    .X(_4007_));
 sky130_fd_sc_hd__a22o_1 _8435_ (.A1(\gpio_configure[14][2] ),
    .A2(_3889_),
    .B1(_3906_),
    .B2(\gpio_configure[27][2] ),
    .X(_4008_));
 sky130_fd_sc_hd__a221o_1 _8436_ (.A1(\gpio_configure[16][2] ),
    .A2(_3947_),
    .B1(_3944_),
    .B2(\gpio_configure[17][2] ),
    .C1(_4008_),
    .X(_4009_));
 sky130_fd_sc_hd__or4_4 _8437_ (.A(_4003_),
    .B(_4005_),
    .C(_4007_),
    .D(_4009_),
    .X(_4010_));
 sky130_fd_sc_hd__a22o_1 _8438_ (.A1(\gpio_configure[32][2] ),
    .A2(_3876_),
    .B1(_3919_),
    .B2(\gpio_configure[37][2] ),
    .X(_4011_));
 sky130_fd_sc_hd__a221o_1 _8439_ (.A1(\gpio_configure[4][2] ),
    .A2(_3966_),
    .B1(_3942_),
    .B2(\gpio_configure[36][2] ),
    .C1(_4011_),
    .X(_4012_));
 sky130_fd_sc_hd__a221o_1 _8440_ (.A1(\gpio_configure[34][2] ),
    .A2(_3923_),
    .B1(_3985_),
    .B2(\gpio_configure[19][2] ),
    .C1(_4012_),
    .X(_4013_));
 sky130_fd_sc_hd__a22o_1 _8441_ (.A1(\gpio_configure[12][2] ),
    .A2(_3891_),
    .B1(_3902_),
    .B2(\gpio_configure[9][2] ),
    .X(_4014_));
 sky130_fd_sc_hd__a221o_1 _8442_ (.A1(\gpio_configure[6][2] ),
    .A2(_3897_),
    .B1(_3908_),
    .B2(\gpio_configure[10][2] ),
    .C1(_4014_),
    .X(_4015_));
 sky130_fd_sc_hd__a22o_1 _8443_ (.A1(\gpio_configure[25][2] ),
    .A2(_3867_),
    .B1(_3869_),
    .B2(\gpio_configure[13][2] ),
    .X(_4016_));
 sky130_fd_sc_hd__a221o_1 _8444_ (.A1(\gpio_configure[5][2] ),
    .A2(_3963_),
    .B1(_3954_),
    .B2(\gpio_configure[2][2] ),
    .C1(_4016_),
    .X(_4017_));
 sky130_fd_sc_hd__a22o_1 _8445_ (.A1(\gpio_configure[31][2] ),
    .A2(_3500_),
    .B1(_3910_),
    .B2(\gpio_configure[11][2] ),
    .X(_4018_));
 sky130_fd_sc_hd__a221o_1 _8446_ (.A1(\gpio_configure[24][2] ),
    .A2(_3912_),
    .B1(_3959_),
    .B2(\gpio_configure[1][2] ),
    .C1(_4018_),
    .X(_4019_));
 sky130_fd_sc_hd__a22o_1 _8447_ (.A1(\gpio_configure[26][2] ),
    .A2(_3879_),
    .B1(_3899_),
    .B2(\gpio_configure[7][2] ),
    .X(_4020_));
 sky130_fd_sc_hd__a221o_1 _8448_ (.A1(\gpio_configure[3][2] ),
    .A2(_3864_),
    .B1(_3916_),
    .B2(\gpio_configure[15][2] ),
    .C1(_4020_),
    .X(_4021_));
 sky130_fd_sc_hd__or4_1 _8449_ (.A(_4015_),
    .B(_4017_),
    .C(_4019_),
    .D(_4021_),
    .X(_4022_));
 sky130_fd_sc_hd__or3_1 _8450_ (.A(_3941_),
    .B(_4013_),
    .C(_4022_),
    .X(_4023_));
 sky130_fd_sc_hd__o221a_1 _8451_ (.A1(\gpio_configure[0][2] ),
    .A2(_3974_),
    .B1(_4010_),
    .B2(_4023_),
    .C1(_3689_),
    .X(_4024_));
 sky130_fd_sc_hd__a21o_1 _8452_ (.A1(_1526_),
    .A2(\serial_data_staging_2[1] ),
    .B1(_3601_),
    .X(_4025_));
 sky130_fd_sc_hd__o22a_1 _8453_ (.A1(net1474),
    .A2(_3603_),
    .B1(_4024_),
    .B2(_4025_),
    .X(_0794_));
 sky130_fd_sc_hd__a22o_1 _8454_ (.A1(\gpio_configure[35][3] ),
    .A2(_3887_),
    .B1(_3951_),
    .B2(\gpio_configure[30][3] ),
    .X(_4026_));
 sky130_fd_sc_hd__a221o_1 _8455_ (.A1(\gpio_configure[29][3] ),
    .A2(_3976_),
    .B1(_3953_),
    .B2(\gpio_configure[21][3] ),
    .C1(_4026_),
    .X(_4027_));
 sky130_fd_sc_hd__a22o_1 _8456_ (.A1(\gpio_configure[23][3] ),
    .A2(_3921_),
    .B1(_3961_),
    .B2(\gpio_configure[20][3] ),
    .X(_4028_));
 sky130_fd_sc_hd__a22o_1 _8457_ (.A1(\gpio_configure[18][3] ),
    .A2(_3872_),
    .B1(_3932_),
    .B2(\gpio_configure[8][3] ),
    .X(_4029_));
 sky130_fd_sc_hd__a221o_1 _8458_ (.A1(\gpio_configure[33][3] ),
    .A2(_3885_),
    .B1(_3956_),
    .B2(\gpio_configure[22][3] ),
    .C1(_4029_),
    .X(_4030_));
 sky130_fd_sc_hd__a22o_1 _8459_ (.A1(\gpio_configure[14][3] ),
    .A2(_3889_),
    .B1(_3906_),
    .B2(\gpio_configure[27][3] ),
    .X(_4031_));
 sky130_fd_sc_hd__a221o_1 _8460_ (.A1(\gpio_configure[16][3] ),
    .A2(_3947_),
    .B1(_3944_),
    .B2(\gpio_configure[17][3] ),
    .C1(_4031_),
    .X(_4032_));
 sky130_fd_sc_hd__a2111o_1 _8461_ (.A1(\gpio_configure[28][3] ),
    .A2(_3965_),
    .B1(_4028_),
    .C1(_4030_),
    .D1(_4032_),
    .X(_4033_));
 sky130_fd_sc_hd__a22o_1 _8462_ (.A1(\gpio_configure[32][3] ),
    .A2(_3875_),
    .B1(_3918_),
    .B2(\gpio_configure[37][3] ),
    .X(_4034_));
 sky130_fd_sc_hd__a221o_1 _8463_ (.A1(\gpio_configure[4][3] ),
    .A2(_3928_),
    .B1(_3930_),
    .B2(\gpio_configure[36][3] ),
    .C1(_4034_),
    .X(_4035_));
 sky130_fd_sc_hd__a221o_1 _8464_ (.A1(\gpio_configure[34][3] ),
    .A2(_3922_),
    .B1(_3967_),
    .B2(\gpio_configure[19][3] ),
    .C1(_4035_),
    .X(_4036_));
 sky130_fd_sc_hd__a22o_1 _8465_ (.A1(\gpio_configure[12][3] ),
    .A2(_3891_),
    .B1(_3902_),
    .B2(\gpio_configure[9][3] ),
    .X(_4037_));
 sky130_fd_sc_hd__a221o_1 _8466_ (.A1(\gpio_configure[6][3] ),
    .A2(_3897_),
    .B1(_3908_),
    .B2(\gpio_configure[10][3] ),
    .C1(_4037_),
    .X(_4038_));
 sky130_fd_sc_hd__a22o_1 _8467_ (.A1(\gpio_configure[3][3] ),
    .A2(_3863_),
    .B1(_3879_),
    .B2(\gpio_configure[26][3] ),
    .X(_4039_));
 sky130_fd_sc_hd__a22o_1 _8468_ (.A1(\gpio_configure[7][3] ),
    .A2(_3899_),
    .B1(_3915_),
    .B2(\gpio_configure[15][3] ),
    .X(_4040_));
 sky130_fd_sc_hd__a22o_1 _8469_ (.A1(\gpio_configure[25][3] ),
    .A2(_3866_),
    .B1(_3868_),
    .B2(\gpio_configure[13][3] ),
    .X(_4041_));
 sky130_fd_sc_hd__a221o_1 _8470_ (.A1(\gpio_configure[5][3] ),
    .A2(_3937_),
    .B1(_3934_),
    .B2(\gpio_configure[2][3] ),
    .C1(_4041_),
    .X(_4042_));
 sky130_fd_sc_hd__a22o_1 _8471_ (.A1(\gpio_configure[31][3] ),
    .A2(_3499_),
    .B1(_3909_),
    .B2(\gpio_configure[11][3] ),
    .X(_4043_));
 sky130_fd_sc_hd__a221o_1 _8472_ (.A1(\gpio_configure[24][3] ),
    .A2(_3911_),
    .B1(_3938_),
    .B2(\gpio_configure[1][3] ),
    .C1(_4043_),
    .X(_4044_));
 sky130_fd_sc_hd__or4_1 _8473_ (.A(_4039_),
    .B(_4040_),
    .C(_4042_),
    .D(_4044_),
    .X(_4045_));
 sky130_fd_sc_hd__or4_1 _8474_ (.A(_3940_),
    .B(_4036_),
    .C(_4038_),
    .D(_4045_),
    .X(_4046_));
 sky130_fd_sc_hd__o32a_2 _8475_ (.A1(_4027_),
    .A2(_4033_),
    .A3(_4046_),
    .B1(_3973_),
    .B2(\gpio_configure[0][3] ),
    .X(_4047_));
 sky130_fd_sc_hd__mux2_1 _8476_ (.A0(\serial_data_staging_2[2] ),
    .A1(_4047_),
    .S(_3625_),
    .X(_4048_));
 sky130_fd_sc_hd__mux2_1 _8477_ (.A0(net1512),
    .A1(_4048_),
    .S(_3602_),
    .X(_4049_));
 sky130_fd_sc_hd__clkbuf_1 _8478_ (.A(_4049_),
    .X(_0795_));
 sky130_fd_sc_hd__a22o_1 _8479_ (.A1(\gpio_configure[35][4] ),
    .A2(_3887_),
    .B1(_3951_),
    .B2(\gpio_configure[30][4] ),
    .X(_4050_));
 sky130_fd_sc_hd__a221o_1 _8480_ (.A1(\gpio_configure[29][4] ),
    .A2(_3976_),
    .B1(_3953_),
    .B2(\gpio_configure[21][4] ),
    .C1(_4050_),
    .X(_4051_));
 sky130_fd_sc_hd__and2_1 _8481_ (.A(\gpio_configure[28][4] ),
    .B(_3965_),
    .X(_4052_));
 sky130_fd_sc_hd__a221o_1 _8482_ (.A1(\gpio_configure[23][4] ),
    .A2(_3921_),
    .B1(_3961_),
    .B2(\gpio_configure[20][4] ),
    .C1(_4052_),
    .X(_4053_));
 sky130_fd_sc_hd__a22o_1 _8483_ (.A1(\gpio_configure[33][4] ),
    .A2(_3885_),
    .B1(_3956_),
    .B2(\gpio_configure[22][4] ),
    .X(_4054_));
 sky130_fd_sc_hd__a221o_1 _8484_ (.A1(\gpio_configure[18][4] ),
    .A2(_3873_),
    .B1(_3945_),
    .B2(\gpio_configure[8][4] ),
    .C1(_4054_),
    .X(_4055_));
 sky130_fd_sc_hd__a22o_1 _8485_ (.A1(\gpio_configure[14][4] ),
    .A2(_3889_),
    .B1(_3906_),
    .B2(\gpio_configure[27][4] ),
    .X(_4056_));
 sky130_fd_sc_hd__a221o_1 _8486_ (.A1(\gpio_configure[16][4] ),
    .A2(_3947_),
    .B1(_3944_),
    .B2(\gpio_configure[17][4] ),
    .C1(_4056_),
    .X(_4057_));
 sky130_fd_sc_hd__or4_4 _8487_ (.A(_4051_),
    .B(_4053_),
    .C(_4055_),
    .D(_4057_),
    .X(_4058_));
 sky130_fd_sc_hd__a22o_1 _8488_ (.A1(\gpio_configure[32][4] ),
    .A2(_3876_),
    .B1(_3919_),
    .B2(\gpio_configure[37][4] ),
    .X(_4059_));
 sky130_fd_sc_hd__a221o_1 _8489_ (.A1(\gpio_configure[4][4] ),
    .A2(_3966_),
    .B1(_3942_),
    .B2(\gpio_configure[36][4] ),
    .C1(_4059_),
    .X(_4060_));
 sky130_fd_sc_hd__a221o_1 _8490_ (.A1(\gpio_configure[34][4] ),
    .A2(_3923_),
    .B1(_3985_),
    .B2(\gpio_configure[19][4] ),
    .C1(_4060_),
    .X(_4061_));
 sky130_fd_sc_hd__a22o_1 _8491_ (.A1(\gpio_configure[12][4] ),
    .A2(_3891_),
    .B1(_3902_),
    .B2(\gpio_configure[9][4] ),
    .X(_4062_));
 sky130_fd_sc_hd__a221o_1 _8492_ (.A1(\gpio_configure[6][4] ),
    .A2(_3897_),
    .B1(_3908_),
    .B2(\gpio_configure[10][4] ),
    .C1(_4062_),
    .X(_4063_));
 sky130_fd_sc_hd__a22o_1 _8493_ (.A1(\gpio_configure[25][4] ),
    .A2(_3867_),
    .B1(_3869_),
    .B2(\gpio_configure[13][4] ),
    .X(_4064_));
 sky130_fd_sc_hd__a221o_1 _8494_ (.A1(\gpio_configure[5][4] ),
    .A2(_3963_),
    .B1(_3954_),
    .B2(\gpio_configure[2][4] ),
    .C1(_4064_),
    .X(_4065_));
 sky130_fd_sc_hd__a22o_1 _8495_ (.A1(\gpio_configure[31][4] ),
    .A2(_3500_),
    .B1(_3910_),
    .B2(\gpio_configure[11][4] ),
    .X(_4066_));
 sky130_fd_sc_hd__a221o_1 _8496_ (.A1(\gpio_configure[24][4] ),
    .A2(_3912_),
    .B1(_3959_),
    .B2(\gpio_configure[1][4] ),
    .C1(_4066_),
    .X(_4067_));
 sky130_fd_sc_hd__a22o_1 _8497_ (.A1(\gpio_configure[26][4] ),
    .A2(_3879_),
    .B1(_3899_),
    .B2(\gpio_configure[7][4] ),
    .X(_4068_));
 sky130_fd_sc_hd__a221o_1 _8498_ (.A1(\gpio_configure[3][4] ),
    .A2(_3864_),
    .B1(_3916_),
    .B2(\gpio_configure[15][4] ),
    .C1(_4068_),
    .X(_4069_));
 sky130_fd_sc_hd__or4_2 _8499_ (.A(_4063_),
    .B(_4065_),
    .C(_4067_),
    .D(_4069_),
    .X(_4070_));
 sky130_fd_sc_hd__or3_1 _8500_ (.A(_3941_),
    .B(_4061_),
    .C(_4070_),
    .X(_4071_));
 sky130_fd_sc_hd__o221a_1 _8501_ (.A1(\gpio_configure[0][4] ),
    .A2(_3974_),
    .B1(_4058_),
    .B2(_4071_),
    .C1(_3625_),
    .X(_4072_));
 sky130_fd_sc_hd__a211o_1 _8502_ (.A1(_1525_),
    .A2(\serial_data_staging_2[3] ),
    .B1(_3600_),
    .C1(_4072_),
    .X(_4073_));
 sky130_fd_sc_hd__o21a_1 _8503_ (.A1(net1460),
    .A2(_3604_),
    .B1(_4073_),
    .X(_0796_));
 sky130_fd_sc_hd__a22o_1 _8504_ (.A1(\gpio_configure[35][5] ),
    .A2(_3887_),
    .B1(_3951_),
    .B2(\gpio_configure[30][5] ),
    .X(_4074_));
 sky130_fd_sc_hd__a221o_1 _8505_ (.A1(\gpio_configure[29][5] ),
    .A2(_3976_),
    .B1(_3953_),
    .B2(\gpio_configure[21][5] ),
    .C1(_4074_),
    .X(_4075_));
 sky130_fd_sc_hd__and2_1 _8506_ (.A(\gpio_configure[28][5] ),
    .B(_3965_),
    .X(_4076_));
 sky130_fd_sc_hd__a221o_1 _8507_ (.A1(\gpio_configure[23][5] ),
    .A2(_3921_),
    .B1(_3961_),
    .B2(\gpio_configure[20][5] ),
    .C1(_4076_),
    .X(_4077_));
 sky130_fd_sc_hd__a22o_1 _8508_ (.A1(\gpio_configure[18][5] ),
    .A2(_3873_),
    .B1(_3945_),
    .B2(\gpio_configure[8][5] ),
    .X(_4078_));
 sky130_fd_sc_hd__a221o_1 _8509_ (.A1(\gpio_configure[33][5] ),
    .A2(_3885_),
    .B1(_3956_),
    .B2(\gpio_configure[22][5] ),
    .C1(_4078_),
    .X(_4079_));
 sky130_fd_sc_hd__a22o_1 _8510_ (.A1(\gpio_configure[14][5] ),
    .A2(_3889_),
    .B1(_3906_),
    .B2(\gpio_configure[27][5] ),
    .X(_4080_));
 sky130_fd_sc_hd__a221o_1 _8511_ (.A1(\gpio_configure[16][5] ),
    .A2(_3947_),
    .B1(_3944_),
    .B2(\gpio_configure[17][5] ),
    .C1(_4080_),
    .X(_4081_));
 sky130_fd_sc_hd__or4_1 _8512_ (.A(_4075_),
    .B(_4077_),
    .C(_4079_),
    .D(_4081_),
    .X(_4082_));
 sky130_fd_sc_hd__a22o_1 _8513_ (.A1(\gpio_configure[32][5] ),
    .A2(_3876_),
    .B1(_3919_),
    .B2(\gpio_configure[37][5] ),
    .X(_4083_));
 sky130_fd_sc_hd__a221o_2 _8514_ (.A1(\gpio_configure[4][5] ),
    .A2(_3966_),
    .B1(_3942_),
    .B2(\gpio_configure[36][5] ),
    .C1(_4083_),
    .X(_4084_));
 sky130_fd_sc_hd__a221o_1 _8515_ (.A1(\gpio_configure[34][5] ),
    .A2(_3923_),
    .B1(_3985_),
    .B2(\gpio_configure[19][5] ),
    .C1(_4084_),
    .X(_4085_));
 sky130_fd_sc_hd__a22o_1 _8516_ (.A1(\gpio_configure[31][5] ),
    .A2(_3500_),
    .B1(_3910_),
    .B2(\gpio_configure[11][5] ),
    .X(_4086_));
 sky130_fd_sc_hd__a221o_1 _8517_ (.A1(\gpio_configure[24][5] ),
    .A2(_3912_),
    .B1(_3959_),
    .B2(\gpio_configure[1][5] ),
    .C1(_4086_),
    .X(_4087_));
 sky130_fd_sc_hd__a22o_1 _8518_ (.A1(\gpio_configure[26][5] ),
    .A2(_3879_),
    .B1(_3899_),
    .B2(\gpio_configure[7][5] ),
    .X(_4088_));
 sky130_fd_sc_hd__a221o_1 _8519_ (.A1(\gpio_configure[3][5] ),
    .A2(_3864_),
    .B1(_3916_),
    .B2(\gpio_configure[15][5] ),
    .C1(_4088_),
    .X(_4089_));
 sky130_fd_sc_hd__a22o_1 _8520_ (.A1(\gpio_configure[12][5] ),
    .A2(_3891_),
    .B1(_3902_),
    .B2(\gpio_configure[9][5] ),
    .X(_4090_));
 sky130_fd_sc_hd__a221o_1 _8521_ (.A1(\gpio_configure[6][5] ),
    .A2(_3897_),
    .B1(_3908_),
    .B2(\gpio_configure[10][5] ),
    .C1(_4090_),
    .X(_4091_));
 sky130_fd_sc_hd__a22o_1 _8522_ (.A1(\gpio_configure[25][5] ),
    .A2(_3867_),
    .B1(_3869_),
    .B2(\gpio_configure[13][5] ),
    .X(_4092_));
 sky130_fd_sc_hd__a221o_1 _8523_ (.A1(\gpio_configure[5][5] ),
    .A2(_3963_),
    .B1(_3954_),
    .B2(\gpio_configure[2][5] ),
    .C1(_4092_),
    .X(_4093_));
 sky130_fd_sc_hd__or4_1 _8524_ (.A(_4087_),
    .B(_4089_),
    .C(_4091_),
    .D(_4093_),
    .X(_4094_));
 sky130_fd_sc_hd__or3_1 _8525_ (.A(_3941_),
    .B(_4085_),
    .C(_4094_),
    .X(_4095_));
 sky130_fd_sc_hd__o221a_2 _8526_ (.A1(\gpio_configure[0][5] ),
    .A2(_3974_),
    .B1(_4082_),
    .B2(_4095_),
    .C1(_3689_),
    .X(_4096_));
 sky130_fd_sc_hd__a21o_1 _8527_ (.A1(_1526_),
    .A2(net1460),
    .B1(_3601_),
    .X(_4097_));
 sky130_fd_sc_hd__o22a_1 _8528_ (.A1(net1489),
    .A2(_3603_),
    .B1(_4096_),
    .B2(_4097_),
    .X(_0797_));
 sky130_fd_sc_hd__a22o_1 _8529_ (.A1(\gpio_configure[35][6] ),
    .A2(_3886_),
    .B1(_3950_),
    .B2(\gpio_configure[30][6] ),
    .X(_4098_));
 sky130_fd_sc_hd__a221o_1 _8530_ (.A1(\gpio_configure[29][6] ),
    .A2(_3900_),
    .B1(_3952_),
    .B2(\gpio_configure[21][6] ),
    .C1(_4098_),
    .X(_4099_));
 sky130_fd_sc_hd__and2_1 _8531_ (.A(\gpio_configure[23][6] ),
    .B(_3920_),
    .X(_4100_));
 sky130_fd_sc_hd__a221o_1 _8532_ (.A1(\gpio_configure[20][6] ),
    .A2(_3960_),
    .B1(_3964_),
    .B2(\gpio_configure[28][6] ),
    .C1(_4100_),
    .X(_4101_));
 sky130_fd_sc_hd__a22o_1 _8533_ (.A1(\gpio_configure[33][6] ),
    .A2(_3884_),
    .B1(_3955_),
    .B2(\gpio_configure[22][6] ),
    .X(_4102_));
 sky130_fd_sc_hd__a221o_1 _8534_ (.A1(\gpio_configure[18][6] ),
    .A2(_3873_),
    .B1(_3945_),
    .B2(\gpio_configure[8][6] ),
    .C1(_4102_),
    .X(_4103_));
 sky130_fd_sc_hd__a22o_1 _8535_ (.A1(\gpio_configure[14][6] ),
    .A2(_3888_),
    .B1(_3905_),
    .B2(\gpio_configure[27][6] ),
    .X(_4104_));
 sky130_fd_sc_hd__a221o_1 _8536_ (.A1(\gpio_configure[16][6] ),
    .A2(_3946_),
    .B1(_3943_),
    .B2(\gpio_configure[17][6] ),
    .C1(_4104_),
    .X(_4105_));
 sky130_fd_sc_hd__or4_1 _8537_ (.A(_4099_),
    .B(_4101_),
    .C(_4103_),
    .D(_4105_),
    .X(_4106_));
 sky130_fd_sc_hd__a22o_1 _8538_ (.A1(\gpio_configure[32][6] ),
    .A2(_3875_),
    .B1(_3919_),
    .B2(\gpio_configure[37][6] ),
    .X(_4107_));
 sky130_fd_sc_hd__a221o_1 _8539_ (.A1(\gpio_configure[4][6] ),
    .A2(_3966_),
    .B1(_3942_),
    .B2(\gpio_configure[36][6] ),
    .C1(_4107_),
    .X(_4108_));
 sky130_fd_sc_hd__a221o_1 _8540_ (.A1(\gpio_configure[34][6] ),
    .A2(_3923_),
    .B1(_3985_),
    .B2(\gpio_configure[19][6] ),
    .C1(_4108_),
    .X(_4109_));
 sky130_fd_sc_hd__a22o_1 _8541_ (.A1(\gpio_configure[12][6] ),
    .A2(_3891_),
    .B1(_3902_),
    .B2(\gpio_configure[9][6] ),
    .X(_4110_));
 sky130_fd_sc_hd__a221o_1 _8542_ (.A1(\gpio_configure[6][6] ),
    .A2(_3897_),
    .B1(_3908_),
    .B2(\gpio_configure[10][6] ),
    .C1(_4110_),
    .X(_4111_));
 sky130_fd_sc_hd__a22o_1 _8543_ (.A1(\gpio_configure[25][6] ),
    .A2(_3867_),
    .B1(_3869_),
    .B2(\gpio_configure[13][6] ),
    .X(_4112_));
 sky130_fd_sc_hd__a221o_1 _8544_ (.A1(\gpio_configure[5][6] ),
    .A2(_3963_),
    .B1(_3954_),
    .B2(\gpio_configure[2][6] ),
    .C1(_4112_),
    .X(_4113_));
 sky130_fd_sc_hd__a22o_1 _8545_ (.A1(\gpio_configure[31][6] ),
    .A2(_3500_),
    .B1(_3910_),
    .B2(\gpio_configure[11][6] ),
    .X(_4114_));
 sky130_fd_sc_hd__a221o_1 _8546_ (.A1(\gpio_configure[24][6] ),
    .A2(_3912_),
    .B1(_3959_),
    .B2(\gpio_configure[1][6] ),
    .C1(_4114_),
    .X(_4115_));
 sky130_fd_sc_hd__a22o_1 _8547_ (.A1(\gpio_configure[26][6] ),
    .A2(_3879_),
    .B1(_3899_),
    .B2(\gpio_configure[7][6] ),
    .X(_4116_));
 sky130_fd_sc_hd__a221o_1 _8548_ (.A1(\gpio_configure[3][6] ),
    .A2(_3864_),
    .B1(_3916_),
    .B2(\gpio_configure[15][6] ),
    .C1(_4116_),
    .X(_4117_));
 sky130_fd_sc_hd__or4_1 _8549_ (.A(_4111_),
    .B(_4113_),
    .C(_4115_),
    .D(_4117_),
    .X(_4118_));
 sky130_fd_sc_hd__or4_4 _8550_ (.A(_3941_),
    .B(_4106_),
    .C(_4109_),
    .D(_4118_),
    .X(_4119_));
 sky130_fd_sc_hd__o21a_1 _8551_ (.A1(\gpio_configure[0][6] ),
    .A2(_3974_),
    .B1(_1546_),
    .X(_4120_));
 sky130_fd_sc_hd__a22o_1 _8552_ (.A1(\xfer_state[1] ),
    .A2(\serial_data_staging_2[5] ),
    .B1(_4119_),
    .B2(_4120_),
    .X(_4121_));
 sky130_fd_sc_hd__mux2_1 _8553_ (.A0(net1520),
    .A1(_4121_),
    .S(_3602_),
    .X(_4122_));
 sky130_fd_sc_hd__clkbuf_1 _8554_ (.A(_4122_),
    .X(_0798_));
 sky130_fd_sc_hd__a22o_1 _8555_ (.A1(\gpio_configure[35][7] ),
    .A2(_3886_),
    .B1(_3950_),
    .B2(\gpio_configure[30][7] ),
    .X(_4123_));
 sky130_fd_sc_hd__a221o_1 _8556_ (.A1(\gpio_configure[29][7] ),
    .A2(_3976_),
    .B1(_3952_),
    .B2(\gpio_configure[21][7] ),
    .C1(_4123_),
    .X(_4124_));
 sky130_fd_sc_hd__and2_1 _8557_ (.A(\gpio_configure[23][7] ),
    .B(_3920_),
    .X(_4125_));
 sky130_fd_sc_hd__a221o_1 _8558_ (.A1(\gpio_configure[20][7] ),
    .A2(_3961_),
    .B1(_3965_),
    .B2(\gpio_configure[28][7] ),
    .C1(_4125_),
    .X(_4126_));
 sky130_fd_sc_hd__a22o_1 _8559_ (.A1(\gpio_configure[33][7] ),
    .A2(_3884_),
    .B1(_3955_),
    .B2(\gpio_configure[22][7] ),
    .X(_4127_));
 sky130_fd_sc_hd__a221o_1 _8560_ (.A1(\gpio_configure[18][7] ),
    .A2(_3873_),
    .B1(_3945_),
    .B2(\gpio_configure[8][7] ),
    .C1(_4127_),
    .X(_4128_));
 sky130_fd_sc_hd__a22o_1 _8561_ (.A1(\gpio_configure[14][7] ),
    .A2(_3889_),
    .B1(_3906_),
    .B2(\gpio_configure[27][7] ),
    .X(_4129_));
 sky130_fd_sc_hd__a221o_1 _8562_ (.A1(\gpio_configure[16][7] ),
    .A2(_3947_),
    .B1(_3944_),
    .B2(\gpio_configure[17][7] ),
    .C1(_4129_),
    .X(_4130_));
 sky130_fd_sc_hd__or4_1 _8563_ (.A(_4124_),
    .B(_4126_),
    .C(_4128_),
    .D(_4130_),
    .X(_4131_));
 sky130_fd_sc_hd__a22o_1 _8564_ (.A1(\gpio_configure[4][7] ),
    .A2(_3966_),
    .B1(_3942_),
    .B2(\gpio_configure[36][7] ),
    .X(_4132_));
 sky130_fd_sc_hd__a221o_1 _8565_ (.A1(\gpio_configure[32][7] ),
    .A2(_3876_),
    .B1(_3919_),
    .B2(\gpio_configure[37][7] ),
    .C1(_4132_),
    .X(_4133_));
 sky130_fd_sc_hd__a221o_1 _8566_ (.A1(\gpio_configure[34][7] ),
    .A2(_3923_),
    .B1(_3985_),
    .B2(\gpio_configure[19][7] ),
    .C1(_4133_),
    .X(_4134_));
 sky130_fd_sc_hd__a22o_2 _8567_ (.A1(\gpio_configure[12][7] ),
    .A2(_3891_),
    .B1(_3902_),
    .B2(\gpio_configure[9][7] ),
    .X(_4135_));
 sky130_fd_sc_hd__a221o_1 _8568_ (.A1(\gpio_configure[6][7] ),
    .A2(_3897_),
    .B1(_3908_),
    .B2(\gpio_configure[10][7] ),
    .C1(_4135_),
    .X(_4136_));
 sky130_fd_sc_hd__a22o_1 _8569_ (.A1(\gpio_configure[25][7] ),
    .A2(_3867_),
    .B1(_3869_),
    .B2(\gpio_configure[13][7] ),
    .X(_4137_));
 sky130_fd_sc_hd__a221o_1 _8570_ (.A1(\gpio_configure[5][7] ),
    .A2(_3963_),
    .B1(_3954_),
    .B2(\gpio_configure[2][7] ),
    .C1(_4137_),
    .X(_4138_));
 sky130_fd_sc_hd__a22o_1 _8571_ (.A1(\gpio_configure[31][7] ),
    .A2(_3500_),
    .B1(_3910_),
    .B2(\gpio_configure[11][7] ),
    .X(_4139_));
 sky130_fd_sc_hd__a221o_1 _8572_ (.A1(\gpio_configure[24][7] ),
    .A2(_3912_),
    .B1(_3959_),
    .B2(\gpio_configure[1][7] ),
    .C1(_4139_),
    .X(_4140_));
 sky130_fd_sc_hd__a22o_1 _8573_ (.A1(\gpio_configure[26][7] ),
    .A2(_3879_),
    .B1(_3899_),
    .B2(\gpio_configure[7][7] ),
    .X(_4141_));
 sky130_fd_sc_hd__a221o_1 _8574_ (.A1(\gpio_configure[3][7] ),
    .A2(_3864_),
    .B1(_3916_),
    .B2(\gpio_configure[15][7] ),
    .C1(_4141_),
    .X(_4142_));
 sky130_fd_sc_hd__or4_1 _8575_ (.A(_4136_),
    .B(_4138_),
    .C(_4140_),
    .D(_4142_),
    .X(_4143_));
 sky130_fd_sc_hd__or4_1 _8576_ (.A(_3941_),
    .B(_4131_),
    .C(_4134_),
    .D(_4143_),
    .X(_4144_));
 sky130_fd_sc_hd__o211a_2 _8577_ (.A1(\gpio_configure[0][7] ),
    .A2(_3974_),
    .B1(_4144_),
    .C1(_3689_),
    .X(_4145_));
 sky130_fd_sc_hd__a21o_1 _8578_ (.A1(_1526_),
    .A2(\serial_data_staging_2[6] ),
    .B1(_3601_),
    .X(_4146_));
 sky130_fd_sc_hd__o22a_1 _8579_ (.A1(net1496),
    .A2(_3603_),
    .B1(_4145_),
    .B2(_4146_),
    .X(_0799_));
 sky130_fd_sc_hd__a22o_1 _8580_ (.A1(\gpio_configure[35][8] ),
    .A2(_3887_),
    .B1(_3951_),
    .B2(\gpio_configure[30][8] ),
    .X(_4147_));
 sky130_fd_sc_hd__a221o_1 _8581_ (.A1(\gpio_configure[29][8] ),
    .A2(_3976_),
    .B1(_3953_),
    .B2(\gpio_configure[21][8] ),
    .C1(_4147_),
    .X(_4148_));
 sky130_fd_sc_hd__and2_1 _8582_ (.A(\gpio_configure[28][8] ),
    .B(_3964_),
    .X(_4149_));
 sky130_fd_sc_hd__a221o_1 _8583_ (.A1(\gpio_configure[23][8] ),
    .A2(_3921_),
    .B1(_3961_),
    .B2(\gpio_configure[20][8] ),
    .C1(_4149_),
    .X(_4150_));
 sky130_fd_sc_hd__a22o_1 _8584_ (.A1(\gpio_configure[18][8] ),
    .A2(_3873_),
    .B1(_3945_),
    .B2(\gpio_configure[8][8] ),
    .X(_4151_));
 sky130_fd_sc_hd__a221o_1 _8585_ (.A1(\gpio_configure[33][8] ),
    .A2(_3885_),
    .B1(_3956_),
    .B2(\gpio_configure[22][8] ),
    .C1(_4151_),
    .X(_4152_));
 sky130_fd_sc_hd__a22o_1 _8586_ (.A1(\gpio_configure[14][8] ),
    .A2(_3889_),
    .B1(_3906_),
    .B2(\gpio_configure[27][8] ),
    .X(_4153_));
 sky130_fd_sc_hd__a221o_1 _8587_ (.A1(\gpio_configure[16][8] ),
    .A2(_3947_),
    .B1(_3944_),
    .B2(\gpio_configure[17][8] ),
    .C1(_4153_),
    .X(_4154_));
 sky130_fd_sc_hd__or4_1 _8588_ (.A(_4148_),
    .B(_4150_),
    .C(_4152_),
    .D(_4154_),
    .X(_4155_));
 sky130_fd_sc_hd__a22o_1 _8589_ (.A1(\gpio_configure[32][8] ),
    .A2(_3876_),
    .B1(_3919_),
    .B2(\gpio_configure[37][8] ),
    .X(_4156_));
 sky130_fd_sc_hd__a221o_1 _8590_ (.A1(\gpio_configure[4][8] ),
    .A2(_3966_),
    .B1(_3942_),
    .B2(\gpio_configure[36][8] ),
    .C1(_4156_),
    .X(_4157_));
 sky130_fd_sc_hd__a221o_1 _8591_ (.A1(\gpio_configure[34][8] ),
    .A2(_3923_),
    .B1(_3985_),
    .B2(\gpio_configure[19][8] ),
    .C1(_4157_),
    .X(_4158_));
 sky130_fd_sc_hd__a22o_1 _8592_ (.A1(\gpio_configure[12][8] ),
    .A2(_3891_),
    .B1(_3902_),
    .B2(\gpio_configure[9][8] ),
    .X(_4159_));
 sky130_fd_sc_hd__a221o_1 _8593_ (.A1(\gpio_configure[6][8] ),
    .A2(_3897_),
    .B1(_3908_),
    .B2(\gpio_configure[10][8] ),
    .C1(_4159_),
    .X(_4160_));
 sky130_fd_sc_hd__a22o_1 _8594_ (.A1(\gpio_configure[3][8] ),
    .A2(_3864_),
    .B1(_3879_),
    .B2(\gpio_configure[26][8] ),
    .X(_4161_));
 sky130_fd_sc_hd__a22o_1 _8595_ (.A1(\gpio_configure[7][8] ),
    .A2(_3899_),
    .B1(_3916_),
    .B2(\gpio_configure[15][8] ),
    .X(_4162_));
 sky130_fd_sc_hd__a22o_1 _8596_ (.A1(\gpio_configure[25][8] ),
    .A2(_3867_),
    .B1(_3869_),
    .B2(\gpio_configure[13][8] ),
    .X(_4163_));
 sky130_fd_sc_hd__a221o_1 _8597_ (.A1(\gpio_configure[5][8] ),
    .A2(_3963_),
    .B1(_3954_),
    .B2(\gpio_configure[2][8] ),
    .C1(_4163_),
    .X(_4164_));
 sky130_fd_sc_hd__a22o_1 _8598_ (.A1(\gpio_configure[31][8] ),
    .A2(_3500_),
    .B1(_3910_),
    .B2(\gpio_configure[11][8] ),
    .X(_4165_));
 sky130_fd_sc_hd__a221o_1 _8599_ (.A1(\gpio_configure[24][8] ),
    .A2(_3912_),
    .B1(_3959_),
    .B2(\gpio_configure[1][8] ),
    .C1(_4165_),
    .X(_4166_));
 sky130_fd_sc_hd__or4_1 _8600_ (.A(_4161_),
    .B(_4162_),
    .C(_4164_),
    .D(_4166_),
    .X(_4167_));
 sky130_fd_sc_hd__or4_1 _8601_ (.A(_3941_),
    .B(_4158_),
    .C(_4160_),
    .D(_4167_),
    .X(_4168_));
 sky130_fd_sc_hd__o221a_1 _8602_ (.A1(\gpio_configure[0][8] ),
    .A2(_3974_),
    .B1(_4155_),
    .B2(_4168_),
    .C1(_3625_),
    .X(_4169_));
 sky130_fd_sc_hd__a211o_1 _8603_ (.A1(_1525_),
    .A2(\serial_data_staging_2[7] ),
    .B1(_3600_),
    .C1(_4169_),
    .X(_4170_));
 sky130_fd_sc_hd__o21a_1 _8604_ (.A1(net1465),
    .A2(_3604_),
    .B1(_4170_),
    .X(_0800_));
 sky130_fd_sc_hd__a22o_1 _8605_ (.A1(\gpio_configure[35][9] ),
    .A2(_3887_),
    .B1(_3951_),
    .B2(\gpio_configure[30][9] ),
    .X(_4171_));
 sky130_fd_sc_hd__a221o_1 _8606_ (.A1(\gpio_configure[29][9] ),
    .A2(_3976_),
    .B1(_3953_),
    .B2(\gpio_configure[21][9] ),
    .C1(_4171_),
    .X(_4172_));
 sky130_fd_sc_hd__a22o_1 _8607_ (.A1(\gpio_configure[23][9] ),
    .A2(_3921_),
    .B1(_3960_),
    .B2(\gpio_configure[20][9] ),
    .X(_4173_));
 sky130_fd_sc_hd__a22o_1 _8608_ (.A1(\gpio_configure[18][9] ),
    .A2(_3872_),
    .B1(_3932_),
    .B2(\gpio_configure[8][9] ),
    .X(_4174_));
 sky130_fd_sc_hd__a221o_1 _8609_ (.A1(\gpio_configure[33][9] ),
    .A2(_3885_),
    .B1(_3956_),
    .B2(\gpio_configure[22][9] ),
    .C1(_4174_),
    .X(_4175_));
 sky130_fd_sc_hd__a22o_1 _8610_ (.A1(\gpio_configure[14][9] ),
    .A2(_3888_),
    .B1(_3905_),
    .B2(\gpio_configure[27][9] ),
    .X(_4176_));
 sky130_fd_sc_hd__a221o_1 _8611_ (.A1(\gpio_configure[16][9] ),
    .A2(_3946_),
    .B1(_3943_),
    .B2(\gpio_configure[17][9] ),
    .C1(_4176_),
    .X(_4177_));
 sky130_fd_sc_hd__a2111o_1 _8612_ (.A1(\gpio_configure[28][9] ),
    .A2(_3965_),
    .B1(_4173_),
    .C1(_4175_),
    .D1(_4177_),
    .X(_4178_));
 sky130_fd_sc_hd__a22o_1 _8613_ (.A1(\gpio_configure[4][9] ),
    .A2(_3928_),
    .B1(_3930_),
    .B2(\gpio_configure[36][9] ),
    .X(_4179_));
 sky130_fd_sc_hd__a221o_1 _8614_ (.A1(\gpio_configure[32][9] ),
    .A2(_3875_),
    .B1(_3918_),
    .B2(\gpio_configure[37][9] ),
    .C1(_4179_),
    .X(_4180_));
 sky130_fd_sc_hd__a221o_1 _8615_ (.A1(\gpio_configure[34][9] ),
    .A2(_3922_),
    .B1(_3985_),
    .B2(\gpio_configure[19][9] ),
    .C1(_4180_),
    .X(_4181_));
 sky130_fd_sc_hd__a22o_1 _8616_ (.A1(\gpio_configure[12][9] ),
    .A2(_3890_),
    .B1(_3901_),
    .B2(\gpio_configure[9][9] ),
    .X(_4182_));
 sky130_fd_sc_hd__a221o_1 _8617_ (.A1(\gpio_configure[6][9] ),
    .A2(_3896_),
    .B1(_3907_),
    .B2(\gpio_configure[10][9] ),
    .C1(_4182_),
    .X(_4183_));
 sky130_fd_sc_hd__a22o_1 _8618_ (.A1(\gpio_configure[25][9] ),
    .A2(_3866_),
    .B1(_3868_),
    .B2(\gpio_configure[13][9] ),
    .X(_4184_));
 sky130_fd_sc_hd__a221o_1 _8619_ (.A1(\gpio_configure[5][9] ),
    .A2(_3937_),
    .B1(_3934_),
    .B2(\gpio_configure[2][9] ),
    .C1(_4184_),
    .X(_4185_));
 sky130_fd_sc_hd__a22o_1 _8620_ (.A1(\gpio_configure[31][9] ),
    .A2(_3499_),
    .B1(_3909_),
    .B2(\gpio_configure[11][9] ),
    .X(_4186_));
 sky130_fd_sc_hd__a221o_1 _8621_ (.A1(\gpio_configure[24][9] ),
    .A2(_3911_),
    .B1(_3938_),
    .B2(\gpio_configure[1][9] ),
    .C1(_4186_),
    .X(_4187_));
 sky130_fd_sc_hd__a22o_1 _8622_ (.A1(\gpio_configure[26][9] ),
    .A2(_3878_),
    .B1(_3898_),
    .B2(\gpio_configure[7][9] ),
    .X(_4188_));
 sky130_fd_sc_hd__a221o_1 _8623_ (.A1(\gpio_configure[3][9] ),
    .A2(_3863_),
    .B1(_3915_),
    .B2(\gpio_configure[15][9] ),
    .C1(_4188_),
    .X(_4189_));
 sky130_fd_sc_hd__or4_1 _8624_ (.A(_4183_),
    .B(_4185_),
    .C(_4187_),
    .D(_4189_),
    .X(_4190_));
 sky130_fd_sc_hd__or3_1 _8625_ (.A(net393),
    .B(_4181_),
    .C(_4190_),
    .X(_4191_));
 sky130_fd_sc_hd__o32a_1 _8626_ (.A1(_4172_),
    .A2(_4178_),
    .A3(_4191_),
    .B1(_3973_),
    .B2(\gpio_configure[0][9] ),
    .X(_4192_));
 sky130_fd_sc_hd__mux2_1 _8627_ (.A0(\serial_data_staging_2[8] ),
    .A1(_4192_),
    .S(_3625_),
    .X(_4193_));
 sky130_fd_sc_hd__mux2_1 _8628_ (.A0(net1507),
    .A1(_4193_),
    .S(_3602_),
    .X(_4194_));
 sky130_fd_sc_hd__clkbuf_1 _8629_ (.A(_4194_),
    .X(_0801_));
 sky130_fd_sc_hd__a22o_1 _8630_ (.A1(\gpio_configure[35][10] ),
    .A2(_3887_),
    .B1(_3951_),
    .B2(\gpio_configure[30][10] ),
    .X(_4195_));
 sky130_fd_sc_hd__a221o_1 _8631_ (.A1(\gpio_configure[29][10] ),
    .A2(_3976_),
    .B1(_3953_),
    .B2(\gpio_configure[21][10] ),
    .C1(_4195_),
    .X(_4196_));
 sky130_fd_sc_hd__a22o_1 _8632_ (.A1(\gpio_configure[23][10] ),
    .A2(_3921_),
    .B1(_3960_),
    .B2(\gpio_configure[20][10] ),
    .X(_4197_));
 sky130_fd_sc_hd__a22o_1 _8633_ (.A1(\gpio_configure[18][10] ),
    .A2(_3872_),
    .B1(_3932_),
    .B2(\gpio_configure[8][10] ),
    .X(_4198_));
 sky130_fd_sc_hd__a221o_1 _8634_ (.A1(\gpio_configure[33][10] ),
    .A2(_3885_),
    .B1(_3956_),
    .B2(\gpio_configure[22][10] ),
    .C1(_4198_),
    .X(_4199_));
 sky130_fd_sc_hd__a22o_1 _8635_ (.A1(\gpio_configure[14][10] ),
    .A2(_3888_),
    .B1(_3905_),
    .B2(\gpio_configure[27][10] ),
    .X(_4200_));
 sky130_fd_sc_hd__a221o_1 _8636_ (.A1(\gpio_configure[16][10] ),
    .A2(_3946_),
    .B1(_3943_),
    .B2(\gpio_configure[17][10] ),
    .C1(_4200_),
    .X(_4201_));
 sky130_fd_sc_hd__a2111o_2 _8637_ (.A1(\gpio_configure[28][10] ),
    .A2(_3965_),
    .B1(_4197_),
    .C1(_4199_),
    .D1(_4201_),
    .X(_4202_));
 sky130_fd_sc_hd__a22o_1 _8638_ (.A1(\gpio_configure[32][10] ),
    .A2(_3875_),
    .B1(_3918_),
    .B2(\gpio_configure[37][10] ),
    .X(_4203_));
 sky130_fd_sc_hd__a221o_1 _8639_ (.A1(\gpio_configure[4][10] ),
    .A2(_3966_),
    .B1(_3942_),
    .B2(\gpio_configure[36][10] ),
    .C1(_4203_),
    .X(_4204_));
 sky130_fd_sc_hd__a221o_1 _8640_ (.A1(\gpio_configure[34][10] ),
    .A2(_3922_),
    .B1(_3967_),
    .B2(\gpio_configure[19][10] ),
    .C1(_4204_),
    .X(_4205_));
 sky130_fd_sc_hd__a22o_1 _8641_ (.A1(\gpio_configure[12][10] ),
    .A2(_3890_),
    .B1(_3901_),
    .B2(\gpio_configure[9][10] ),
    .X(_4206_));
 sky130_fd_sc_hd__a221o_1 _8642_ (.A1(\gpio_configure[6][10] ),
    .A2(_3896_),
    .B1(_3907_),
    .B2(\gpio_configure[10][10] ),
    .C1(_4206_),
    .X(_4207_));
 sky130_fd_sc_hd__a22o_1 _8643_ (.A1(\gpio_configure[25][10] ),
    .A2(_3866_),
    .B1(_3868_),
    .B2(\gpio_configure[13][10] ),
    .X(_4208_));
 sky130_fd_sc_hd__a221o_1 _8644_ (.A1(\gpio_configure[5][10] ),
    .A2(_3937_),
    .B1(_3934_),
    .B2(\gpio_configure[2][10] ),
    .C1(_4208_),
    .X(_4209_));
 sky130_fd_sc_hd__a22o_1 _8645_ (.A1(\gpio_configure[31][10] ),
    .A2(_3499_),
    .B1(_3909_),
    .B2(\gpio_configure[11][10] ),
    .X(_4210_));
 sky130_fd_sc_hd__a221o_1 _8646_ (.A1(\gpio_configure[24][10] ),
    .A2(_3911_),
    .B1(_3938_),
    .B2(\gpio_configure[1][10] ),
    .C1(_4210_),
    .X(_4211_));
 sky130_fd_sc_hd__a22o_1 _8647_ (.A1(\gpio_configure[26][10] ),
    .A2(_3878_),
    .B1(_3898_),
    .B2(\gpio_configure[7][10] ),
    .X(_4212_));
 sky130_fd_sc_hd__a221o_1 _8648_ (.A1(\gpio_configure[3][10] ),
    .A2(_3863_),
    .B1(_3915_),
    .B2(\gpio_configure[15][10] ),
    .C1(_4212_),
    .X(_4213_));
 sky130_fd_sc_hd__or4_1 _8649_ (.A(_4207_),
    .B(_4209_),
    .C(_4211_),
    .D(_4213_),
    .X(_4214_));
 sky130_fd_sc_hd__or3_1 _8650_ (.A(net393),
    .B(_4205_),
    .C(_4214_),
    .X(_4215_));
 sky130_fd_sc_hd__o32a_1 _8651_ (.A1(_4196_),
    .A2(_4202_),
    .A3(_4215_),
    .B1(_3973_),
    .B2(\gpio_configure[0][10] ),
    .X(_4216_));
 sky130_fd_sc_hd__mux2_1 _8652_ (.A0(\serial_data_staging_2[9] ),
    .A1(_4216_),
    .S(_1546_),
    .X(_4217_));
 sky130_fd_sc_hd__mux2_1 _8653_ (.A0(net1526),
    .A1(_4217_),
    .S(_3602_),
    .X(_4218_));
 sky130_fd_sc_hd__clkbuf_1 _8654_ (.A(_4218_),
    .X(_0802_));
 sky130_fd_sc_hd__a22o_1 _8655_ (.A1(\gpio_configure[35][11] ),
    .A2(_3887_),
    .B1(_3951_),
    .B2(\gpio_configure[30][11] ),
    .X(_4219_));
 sky130_fd_sc_hd__a221o_1 _8656_ (.A1(\gpio_configure[29][11] ),
    .A2(_3976_),
    .B1(_3953_),
    .B2(\gpio_configure[21][11] ),
    .C1(_4219_),
    .X(_4220_));
 sky130_fd_sc_hd__and2_1 _8657_ (.A(\gpio_configure[28][11] ),
    .B(_3964_),
    .X(_4221_));
 sky130_fd_sc_hd__a221o_2 _8658_ (.A1(\gpio_configure[23][11] ),
    .A2(_3921_),
    .B1(_3961_),
    .B2(\gpio_configure[20][11] ),
    .C1(_4221_),
    .X(_4222_));
 sky130_fd_sc_hd__a22o_1 _8659_ (.A1(\gpio_configure[18][11] ),
    .A2(_3873_),
    .B1(_3945_),
    .B2(\gpio_configure[8][11] ),
    .X(_4223_));
 sky130_fd_sc_hd__a221o_1 _8660_ (.A1(\gpio_configure[33][11] ),
    .A2(_3885_),
    .B1(_3956_),
    .B2(\gpio_configure[22][11] ),
    .C1(_4223_),
    .X(_4224_));
 sky130_fd_sc_hd__a22o_1 _8661_ (.A1(\gpio_configure[14][11] ),
    .A2(_3889_),
    .B1(_3906_),
    .B2(\gpio_configure[27][11] ),
    .X(_4225_));
 sky130_fd_sc_hd__a221o_1 _8662_ (.A1(\gpio_configure[16][11] ),
    .A2(_3947_),
    .B1(_3944_),
    .B2(\gpio_configure[17][11] ),
    .C1(_4225_),
    .X(_4226_));
 sky130_fd_sc_hd__or4_1 _8663_ (.A(_4220_),
    .B(_4222_),
    .C(_4224_),
    .D(_4226_),
    .X(_4227_));
 sky130_fd_sc_hd__a22o_1 _8664_ (.A1(\gpio_configure[32][11] ),
    .A2(_3876_),
    .B1(_3919_),
    .B2(\gpio_configure[37][11] ),
    .X(_4228_));
 sky130_fd_sc_hd__a221o_1 _8665_ (.A1(\gpio_configure[4][11] ),
    .A2(_3966_),
    .B1(_3942_),
    .B2(\gpio_configure[36][11] ),
    .C1(_4228_),
    .X(_4229_));
 sky130_fd_sc_hd__a221o_1 _8666_ (.A1(\gpio_configure[34][11] ),
    .A2(_3923_),
    .B1(_3985_),
    .B2(\gpio_configure[19][11] ),
    .C1(_4229_),
    .X(_4230_));
 sky130_fd_sc_hd__a22o_1 _8667_ (.A1(\gpio_configure[12][11] ),
    .A2(_3891_),
    .B1(_3902_),
    .B2(\gpio_configure[9][11] ),
    .X(_4231_));
 sky130_fd_sc_hd__a221o_1 _8668_ (.A1(\gpio_configure[6][11] ),
    .A2(_3897_),
    .B1(_3908_),
    .B2(\gpio_configure[10][11] ),
    .C1(_4231_),
    .X(_4232_));
 sky130_fd_sc_hd__a22o_1 _8669_ (.A1(\gpio_configure[25][11] ),
    .A2(_3867_),
    .B1(_3869_),
    .B2(\gpio_configure[13][11] ),
    .X(_4233_));
 sky130_fd_sc_hd__a221o_1 _8670_ (.A1(\gpio_configure[5][11] ),
    .A2(_3963_),
    .B1(_3954_),
    .B2(\gpio_configure[2][11] ),
    .C1(_4233_),
    .X(_4234_));
 sky130_fd_sc_hd__a22o_1 _8671_ (.A1(\gpio_configure[31][11] ),
    .A2(_3500_),
    .B1(_3910_),
    .B2(\gpio_configure[11][11] ),
    .X(_4235_));
 sky130_fd_sc_hd__a221o_1 _8672_ (.A1(\gpio_configure[24][11] ),
    .A2(_3912_),
    .B1(_3959_),
    .B2(\gpio_configure[1][11] ),
    .C1(_4235_),
    .X(_4236_));
 sky130_fd_sc_hd__a22o_1 _8673_ (.A1(\gpio_configure[3][11] ),
    .A2(_3864_),
    .B1(_3916_),
    .B2(\gpio_configure[15][11] ),
    .X(_4237_));
 sky130_fd_sc_hd__a221o_1 _8674_ (.A1(\gpio_configure[26][11] ),
    .A2(_3879_),
    .B1(_3899_),
    .B2(\gpio_configure[7][11] ),
    .C1(_4237_),
    .X(_4238_));
 sky130_fd_sc_hd__or4_1 _8675_ (.A(_4232_),
    .B(_4234_),
    .C(_4236_),
    .D(_4238_),
    .X(_4239_));
 sky130_fd_sc_hd__or3_1 _8676_ (.A(_3941_),
    .B(_4230_),
    .C(_4239_),
    .X(_4240_));
 sky130_fd_sc_hd__o221a_1 _8677_ (.A1(\gpio_configure[0][11] ),
    .A2(_3974_),
    .B1(_4227_),
    .B2(_4240_),
    .C1(_3625_),
    .X(_4241_));
 sky130_fd_sc_hd__a211o_1 _8678_ (.A1(_1525_),
    .A2(\serial_data_staging_2[10] ),
    .B1(_3600_),
    .C1(_4241_),
    .X(_4242_));
 sky130_fd_sc_hd__o21a_1 _8679_ (.A1(net1476),
    .A2(_3604_),
    .B1(_4242_),
    .X(_0803_));
 sky130_fd_sc_hd__a22o_1 _8680_ (.A1(\gpio_configure[35][12] ),
    .A2(_3886_),
    .B1(_3950_),
    .B2(\gpio_configure[30][12] ),
    .X(_4243_));
 sky130_fd_sc_hd__a221o_1 _8681_ (.A1(\gpio_configure[29][12] ),
    .A2(_3900_),
    .B1(_3952_),
    .B2(\gpio_configure[21][12] ),
    .C1(_4243_),
    .X(_4244_));
 sky130_fd_sc_hd__and2_1 _8682_ (.A(\gpio_configure[23][12] ),
    .B(_3920_),
    .X(_4245_));
 sky130_fd_sc_hd__a221o_1 _8683_ (.A1(\gpio_configure[20][12] ),
    .A2(_3961_),
    .B1(_3965_),
    .B2(\gpio_configure[28][12] ),
    .C1(_4245_),
    .X(_4246_));
 sky130_fd_sc_hd__a22o_1 _8684_ (.A1(\gpio_configure[33][12] ),
    .A2(_3884_),
    .B1(_3955_),
    .B2(\gpio_configure[22][12] ),
    .X(_4247_));
 sky130_fd_sc_hd__a221o_1 _8685_ (.A1(\gpio_configure[18][12] ),
    .A2(_3873_),
    .B1(_3945_),
    .B2(\gpio_configure[8][12] ),
    .C1(_4247_),
    .X(_4248_));
 sky130_fd_sc_hd__a22o_1 _8686_ (.A1(\gpio_configure[14][12] ),
    .A2(_3889_),
    .B1(_3906_),
    .B2(\gpio_configure[27][12] ),
    .X(_4249_));
 sky130_fd_sc_hd__a221o_1 _8687_ (.A1(\gpio_configure[16][12] ),
    .A2(_3947_),
    .B1(_3944_),
    .B2(\gpio_configure[17][12] ),
    .C1(_4249_),
    .X(_4250_));
 sky130_fd_sc_hd__or4_1 _8688_ (.A(_4244_),
    .B(_4246_),
    .C(_4248_),
    .D(_4250_),
    .X(_4251_));
 sky130_fd_sc_hd__a22o_1 _8689_ (.A1(\gpio_configure[4][12] ),
    .A2(_3966_),
    .B1(_3942_),
    .B2(\gpio_configure[36][12] ),
    .X(_4252_));
 sky130_fd_sc_hd__a221o_1 _8690_ (.A1(\gpio_configure[32][12] ),
    .A2(_3876_),
    .B1(_3919_),
    .B2(\gpio_configure[37][12] ),
    .C1(_4252_),
    .X(_4253_));
 sky130_fd_sc_hd__a221o_1 _8691_ (.A1(\gpio_configure[34][12] ),
    .A2(_3923_),
    .B1(_3985_),
    .B2(\gpio_configure[19][12] ),
    .C1(_4253_),
    .X(_4254_));
 sky130_fd_sc_hd__a22o_1 _8692_ (.A1(\gpio_configure[12][12] ),
    .A2(_3891_),
    .B1(_3902_),
    .B2(\gpio_configure[9][12] ),
    .X(_4255_));
 sky130_fd_sc_hd__a221o_1 _8693_ (.A1(\gpio_configure[6][12] ),
    .A2(_3897_),
    .B1(_3908_),
    .B2(\gpio_configure[10][12] ),
    .C1(_4255_),
    .X(_4256_));
 sky130_fd_sc_hd__a22o_1 _8694_ (.A1(\gpio_configure[25][12] ),
    .A2(_3867_),
    .B1(_3869_),
    .B2(\gpio_configure[13][12] ),
    .X(_4257_));
 sky130_fd_sc_hd__a221o_1 _8695_ (.A1(\gpio_configure[5][12] ),
    .A2(_3963_),
    .B1(_3954_),
    .B2(\gpio_configure[2][12] ),
    .C1(_4257_),
    .X(_4258_));
 sky130_fd_sc_hd__a22o_1 _8696_ (.A1(\gpio_configure[31][12] ),
    .A2(_3500_),
    .B1(_3910_),
    .B2(\gpio_configure[11][12] ),
    .X(_4259_));
 sky130_fd_sc_hd__a221o_1 _8697_ (.A1(\gpio_configure[24][12] ),
    .A2(_3912_),
    .B1(_3959_),
    .B2(\gpio_configure[1][12] ),
    .C1(_4259_),
    .X(_4260_));
 sky130_fd_sc_hd__a22o_1 _8698_ (.A1(\gpio_configure[26][12] ),
    .A2(_3879_),
    .B1(_3899_),
    .B2(\gpio_configure[7][12] ),
    .X(_4261_));
 sky130_fd_sc_hd__a221o_1 _8699_ (.A1(\gpio_configure[3][12] ),
    .A2(_3864_),
    .B1(_3916_),
    .B2(\gpio_configure[15][12] ),
    .C1(_4261_),
    .X(_4262_));
 sky130_fd_sc_hd__or4_1 _8700_ (.A(_4256_),
    .B(_4258_),
    .C(_4260_),
    .D(_4262_),
    .X(_4263_));
 sky130_fd_sc_hd__or4_1 _8701_ (.A(_3941_),
    .B(_4251_),
    .C(_4254_),
    .D(_4263_),
    .X(_4264_));
 sky130_fd_sc_hd__o211a_1 _8702_ (.A1(\gpio_configure[0][12] ),
    .A2(_3974_),
    .B1(_4264_),
    .C1(_3689_),
    .X(_4265_));
 sky130_fd_sc_hd__a21o_1 _8703_ (.A1(_1525_),
    .A2(net1476),
    .B1(_3600_),
    .X(_4266_));
 sky130_fd_sc_hd__o22a_1 _8704_ (.A1(\serial_data_staging_2[12] ),
    .A2(_3603_),
    .B1(_4265_),
    .B2(_4266_),
    .X(_0804_));
 sky130_fd_sc_hd__nand2_1 _8705_ (.A(net1502),
    .B(_1523_),
    .Y(_4267_));
 sky130_fd_sc_hd__nand2_1 _8706_ (.A(_1539_),
    .B(net1532),
    .Y(_4268_));
 sky130_fd_sc_hd__o21a_1 _8707_ (.A1(_1539_),
    .A2(_1523_),
    .B1(net1448),
    .X(_4269_));
 sky130_fd_sc_hd__a31o_1 _8708_ (.A1(net326),
    .A2(_4267_),
    .A3(_4268_),
    .B1(_4269_),
    .X(_0805_));
 sky130_fd_sc_hd__and2_1 _8709_ (.A(\wbbd_state[1] ),
    .B(net501),
    .X(_4270_));
 sky130_fd_sc_hd__buf_2 _8710_ (.A(_4270_),
    .X(_4271_));
 sky130_fd_sc_hd__mux2_1 _8711_ (.A0(net343),
    .A1(_1426_),
    .S(_4271_),
    .X(_4272_));
 sky130_fd_sc_hd__clkbuf_1 _8712_ (.A(_4272_),
    .X(_0806_));
 sky130_fd_sc_hd__mux2_1 _8713_ (.A0(net344),
    .A1(_1352_),
    .S(_4271_),
    .X(_4273_));
 sky130_fd_sc_hd__clkbuf_1 _8714_ (.A(_4273_),
    .X(_0807_));
 sky130_fd_sc_hd__mux2_1 _8715_ (.A0(net345),
    .A1(_1285_),
    .S(_4271_),
    .X(_4274_));
 sky130_fd_sc_hd__clkbuf_1 _8716_ (.A(_4274_),
    .X(_0808_));
 sky130_fd_sc_hd__mux2_1 _8717_ (.A0(net346),
    .A1(_1221_),
    .S(_4271_),
    .X(_4275_));
 sky130_fd_sc_hd__clkbuf_1 _8718_ (.A(_4275_),
    .X(_0809_));
 sky130_fd_sc_hd__mux2_2 _8719_ (.A0(net347),
    .A1(clknet_1_1__leaf__1160_),
    .S(_4271_),
    .X(_4276_));
 sky130_fd_sc_hd__buf_1 _8720_ (.A(_4276_),
    .X(_0810_));
 sky130_fd_sc_hd__mux2_1 _8721_ (.A0(net348),
    .A1(_1062_),
    .S(_4271_),
    .X(_4277_));
 sky130_fd_sc_hd__clkbuf_1 _8722_ (.A(_4277_),
    .X(_0811_));
 sky130_fd_sc_hd__mux2_1 _8723_ (.A0(net350),
    .A1(_1022_),
    .S(_4271_),
    .X(_4278_));
 sky130_fd_sc_hd__clkbuf_1 _8724_ (.A(_4278_),
    .X(_0812_));
 sky130_fd_sc_hd__mux2_1 _8725_ (.A0(net351),
    .A1(_0982_),
    .S(_4271_),
    .X(_4279_));
 sky130_fd_sc_hd__clkbuf_1 _8726_ (.A(_4279_),
    .X(_0813_));
 sky130_fd_sc_hd__nor3_4 _8727_ (.A(\wbbd_state[8] ),
    .B(\wbbd_state[7] ),
    .C(\wbbd_state[9] ),
    .Y(_4280_));
 sky130_fd_sc_hd__a22o_1 _8728_ (.A1(_1536_),
    .A2(net171),
    .B1(net164),
    .B2(_4280_),
    .X(_4281_));
 sky130_fd_sc_hd__a221o_1 _8729_ (.A1(_1538_),
    .A2(net180),
    .B1(net194),
    .B2(_1537_),
    .C1(_4281_),
    .X(_4282_));
 sky130_fd_sc_hd__a21boi_1 _8730_ (.A1(net202),
    .A2(net198),
    .B1_N(\wbbd_state[8] ),
    .Y(_4283_));
 sky130_fd_sc_hd__nand2_1 _8731_ (.A(net200),
    .B(net202),
    .Y(_4284_));
 sky130_fd_sc_hd__nand2_1 _8732_ (.A(net202),
    .B(net199),
    .Y(_4285_));
 sky130_fd_sc_hd__a22o_1 _8733_ (.A1(\wbbd_state[9] ),
    .A2(_4284_),
    .B1(_4285_),
    .B2(\wbbd_state[7] ),
    .X(_4286_));
 sky130_fd_sc_hd__a21bo_1 _8734_ (.A1(net202),
    .A2(net197),
    .B1_N(\wbbd_state[5] ),
    .X(_4287_));
 sky130_fd_sc_hd__or4b_1 _8735_ (.A(_2533_),
    .B(_4283_),
    .C(_4286_),
    .D_N(_4287_),
    .X(_4288_));
 sky130_fd_sc_hd__buf_2 _8736_ (.A(_4288_),
    .X(_4289_));
 sky130_fd_sc_hd__mux2_1 _8737_ (.A0(_4282_),
    .A1(net1559),
    .S(_4289_),
    .X(_4290_));
 sky130_fd_sc_hd__clkbuf_1 _8738_ (.A(_4290_),
    .X(_0814_));
 sky130_fd_sc_hd__a22o_1 _8739_ (.A1(_1538_),
    .A2(net181),
    .B1(net195),
    .B2(_1537_),
    .X(_4291_));
 sky130_fd_sc_hd__a221o_1 _8740_ (.A1(_1536_),
    .A2(net172),
    .B1(net175),
    .B2(_4280_),
    .C1(_4291_),
    .X(_4292_));
 sky130_fd_sc_hd__mux2_1 _8741_ (.A0(_4292_),
    .A1(net574),
    .S(_4289_),
    .X(_4293_));
 sky130_fd_sc_hd__clkbuf_1 _8742_ (.A(_4293_),
    .X(_0815_));
 sky130_fd_sc_hd__a22o_1 _8743_ (.A1(_1538_),
    .A2(net182),
    .B1(net165),
    .B2(_1537_),
    .X(_4294_));
 sky130_fd_sc_hd__a221o_1 _8744_ (.A1(_1536_),
    .A2(net173),
    .B1(net186),
    .B2(_4280_),
    .C1(_4294_),
    .X(_4295_));
 sky130_fd_sc_hd__mux2_1 _8745_ (.A0(_4295_),
    .A1(net1558),
    .S(_4289_),
    .X(_4296_));
 sky130_fd_sc_hd__clkbuf_1 _8746_ (.A(_4296_),
    .X(_0816_));
 sky130_fd_sc_hd__a22o_1 _8747_ (.A1(_1538_),
    .A2(net183),
    .B1(net166),
    .B2(_1537_),
    .X(_4297_));
 sky130_fd_sc_hd__a221o_1 _8748_ (.A1(_1536_),
    .A2(net174),
    .B1(net189),
    .B2(_4280_),
    .C1(_4297_),
    .X(_4298_));
 sky130_fd_sc_hd__mux2_1 _8749_ (.A0(_4298_),
    .A1(net1563),
    .S(_4289_),
    .X(_4299_));
 sky130_fd_sc_hd__clkbuf_1 _8750_ (.A(_4299_),
    .X(_0817_));
 sky130_fd_sc_hd__a22o_1 _8751_ (.A1(_1538_),
    .A2(net184),
    .B1(net167),
    .B2(_1537_),
    .X(_4300_));
 sky130_fd_sc_hd__a221o_1 _8752_ (.A1(_1536_),
    .A2(net176),
    .B1(net190),
    .B2(_4280_),
    .C1(_4300_),
    .X(_4301_));
 sky130_fd_sc_hd__mux2_1 _8753_ (.A0(_4301_),
    .A1(net618),
    .S(_4289_),
    .X(_4302_));
 sky130_fd_sc_hd__clkbuf_1 _8754_ (.A(_4302_),
    .X(_0818_));
 sky130_fd_sc_hd__a22o_1 _8755_ (.A1(_1538_),
    .A2(net185),
    .B1(net168),
    .B2(_1537_),
    .X(_4303_));
 sky130_fd_sc_hd__a221o_1 _8756_ (.A1(_1536_),
    .A2(net177),
    .B1(net191),
    .B2(_4280_),
    .C1(_4303_),
    .X(_4304_));
 sky130_fd_sc_hd__mux2_1 _8757_ (.A0(_4304_),
    .A1(net1564),
    .S(_4289_),
    .X(_4305_));
 sky130_fd_sc_hd__clkbuf_1 _8758_ (.A(_4305_),
    .X(_0819_));
 sky130_fd_sc_hd__a22o_1 _8759_ (.A1(\wbbd_state[7] ),
    .A2(net178),
    .B1(net169),
    .B2(_1537_),
    .X(_4306_));
 sky130_fd_sc_hd__a221o_1 _8760_ (.A1(_1538_),
    .A2(net187),
    .B1(net192),
    .B2(_4280_),
    .C1(_4306_),
    .X(_4307_));
 sky130_fd_sc_hd__mux2_1 _8761_ (.A0(_4307_),
    .A1(net1533),
    .S(_4289_),
    .X(_4308_));
 sky130_fd_sc_hd__clkbuf_1 _8762_ (.A(_4308_),
    .X(_0820_));
 sky130_fd_sc_hd__a22o_1 _8763_ (.A1(\wbbd_state[9] ),
    .A2(net188),
    .B1(net170),
    .B2(net1521),
    .X(_4309_));
 sky130_fd_sc_hd__a221o_1 _8764_ (.A1(_1536_),
    .A2(net179),
    .B1(net193),
    .B2(_4280_),
    .C1(net1522),
    .X(_4310_));
 sky130_fd_sc_hd__mux2_1 _8765_ (.A0(_4310_),
    .A1(\wbbd_data[7] ),
    .S(_4289_),
    .X(_4311_));
 sky130_fd_sc_hd__clkbuf_1 _8766_ (.A(net1523),
    .X(_0821_));
 sky130_fd_sc_hd__o211a_2 _8767_ (.A1(clknet_1_1__leaf_wbbd_sck),
    .A2(_1946_),
    .B1(_2533_),
    .C1(_1540_),
    .X(_0822_));
 sky130_fd_sc_hd__a22o_1 _8768_ (.A1(_1538_),
    .A2(net200),
    .B1(net199),
    .B2(_1536_),
    .X(_4312_));
 sky130_fd_sc_hd__a21o_1 _8769_ (.A1(_1537_),
    .A2(net198),
    .B1(_4312_),
    .X(_4313_));
 sky130_fd_sc_hd__a32o_1 _8770_ (.A1(_1540_),
    .A2(_4280_),
    .A3(_4287_),
    .B1(_4313_),
    .B2(net202),
    .X(_4314_));
 sky130_fd_sc_hd__o31a_1 _8771_ (.A1(net609),
    .A2(net1498),
    .A3(_1949_),
    .B1(_4314_),
    .X(_0823_));
 sky130_fd_sc_hd__dfrtp_4 _8772_ (.CLK(clknet_leaf_67_csclk),
    .D(_0065_),
    .RESET_B(net427),
    .Q(\gpio_configure[26][8] ));
 sky130_fd_sc_hd__dfrtp_4 _8773_ (.CLK(clknet_leaf_61_csclk),
    .D(_0066_),
    .RESET_B(net438),
    .Q(\gpio_configure[26][9] ));
 sky130_fd_sc_hd__dfstp_2 _8774_ (.CLK(clknet_leaf_61_csclk),
    .D(_0067_),
    .SET_B(net438),
    .Q(\gpio_configure[26][10] ));
 sky130_fd_sc_hd__dfrtp_4 _8775_ (.CLK(clknet_leaf_63_csclk),
    .D(_0068_),
    .RESET_B(net438),
    .Q(\gpio_configure[26][11] ));
 sky130_fd_sc_hd__dfrtp_4 _8776_ (.CLK(clknet_leaf_67_csclk),
    .D(_0069_),
    .RESET_B(net430),
    .Q(\gpio_configure[26][12] ));
 sky130_fd_sc_hd__dfrtn_1 _8777_ (.CLK_N(clknet_2_2_0_mgmt_gpio_in[4]),
    .D(_0070_),
    .RESET_B(_0019_),
    .Q(\hkspi.wrstb ));
 sky130_fd_sc_hd__dfrtp_1 _8778_ (.CLK(clknet_2_0_0_mgmt_gpio_in[4]),
    .D(_0071_),
    .RESET_B(_0020_),
    .Q(\hkspi.pre_pass_thru_user ));
 sky130_fd_sc_hd__dfstp_1 _8779_ (.CLK(net505),
    .D(_0018_),
    .SET_B(_0021_),
    .Q(\hkspi.sdoenb ));
 sky130_fd_sc_hd__dfrtp_2 _8780_ (.CLK(clknet_2_0_0_mgmt_gpio_in[4]),
    .D(_0072_),
    .RESET_B(_0023_),
    .Q(\hkspi.pre_pass_thru_mgmt ));
 sky130_fd_sc_hd__dfrtp_1 _8781_ (.CLK(clknet_2_3_0_mgmt_gpio_in[4]),
    .D(_0073_),
    .RESET_B(_0024_),
    .Q(\hkspi.odata[1] ));
 sky130_fd_sc_hd__dfrtp_1 _8782_ (.CLK(clknet_2_3_0_mgmt_gpio_in[4]),
    .D(_0074_),
    .RESET_B(_0025_),
    .Q(\hkspi.odata[2] ));
 sky130_fd_sc_hd__dfrtp_1 _8783_ (.CLK(clknet_2_3_0_mgmt_gpio_in[4]),
    .D(_0075_),
    .RESET_B(_0026_),
    .Q(\hkspi.odata[3] ));
 sky130_fd_sc_hd__dfrtp_1 _8784_ (.CLK(clknet_2_3_0_mgmt_gpio_in[4]),
    .D(_0076_),
    .RESET_B(_0027_),
    .Q(\hkspi.odata[4] ));
 sky130_fd_sc_hd__dfrtp_1 _8785_ (.CLK(clknet_2_3_0_mgmt_gpio_in[4]),
    .D(_0077_),
    .RESET_B(_0028_),
    .Q(\hkspi.odata[5] ));
 sky130_fd_sc_hd__dfrtp_1 _8786_ (.CLK(clknet_2_3_0_mgmt_gpio_in[4]),
    .D(_0078_),
    .RESET_B(_0029_),
    .Q(\hkspi.odata[6] ));
 sky130_fd_sc_hd__dfrtp_1 _8787_ (.CLK(clknet_2_3_0_mgmt_gpio_in[4]),
    .D(_0079_),
    .RESET_B(_0030_),
    .Q(\hkspi.odata[7] ));
 sky130_fd_sc_hd__dfrtp_1 _8788_ (.CLK(clknet_2_1_0_mgmt_gpio_in[4]),
    .D(_0080_),
    .RESET_B(_0031_),
    .Q(\hkspi.fixed[0] ));
 sky130_fd_sc_hd__dfrtp_1 _8789_ (.CLK(clknet_2_0_0_mgmt_gpio_in[4]),
    .D(_0081_),
    .RESET_B(_0032_),
    .Q(\hkspi.fixed[1] ));
 sky130_fd_sc_hd__dfrtp_1 _8790_ (.CLK(clknet_2_1_0_mgmt_gpio_in[4]),
    .D(net1472),
    .RESET_B(_0033_),
    .Q(\hkspi.fixed[2] ));
 sky130_fd_sc_hd__dfrtp_1 _8791_ (.CLK(clknet_2_1_0_mgmt_gpio_in[4]),
    .D(_0083_),
    .RESET_B(_0034_),
    .Q(\hkspi.readmode ));
 sky130_fd_sc_hd__dfrtp_1 _8792_ (.CLK(clknet_2_0_0_mgmt_gpio_in[4]),
    .D(_0084_),
    .RESET_B(_0035_),
    .Q(\hkspi.writemode ));
 sky130_fd_sc_hd__dfrtp_1 _8793_ (.CLK(clknet_2_0_0_mgmt_gpio_in[4]),
    .D(_0085_),
    .RESET_B(_0036_),
    .Q(\hkspi.rdstb ));
 sky130_fd_sc_hd__dfrtp_4 _8794_ (.CLK(clknet_2_1_0_mgmt_gpio_in[4]),
    .D(net1458),
    .RESET_B(_0037_),
    .Q(\hkspi.pass_thru_mgmt ));
 sky130_fd_sc_hd__dfrtp_4 _8795_ (.CLK(clknet_2_1_0_mgmt_gpio_in[4]),
    .D(_0087_),
    .RESET_B(_0038_),
    .Q(\hkspi.pass_thru_mgmt_delay ));
 sky130_fd_sc_hd__dfrtp_4 _8796_ (.CLK(clknet_2_0_0_mgmt_gpio_in[4]),
    .D(_0088_),
    .RESET_B(_0039_),
    .Q(\hkspi.pass_thru_user ));
 sky130_fd_sc_hd__dfrtp_4 _8797_ (.CLK(clknet_2_1_0_mgmt_gpio_in[4]),
    .D(_0089_),
    .RESET_B(_0040_),
    .Q(\hkspi.pass_thru_user_delay ));
 sky130_fd_sc_hd__dfrtp_4 _8798_ (.CLK(clknet_2_0_0_mgmt_gpio_in[4]),
    .D(_0090_),
    .RESET_B(_0041_),
    .Q(\hkspi.addr[0] ));
 sky130_fd_sc_hd__dfrtp_2 _8799_ (.CLK(clknet_2_1_0_mgmt_gpio_in[4]),
    .D(_0091_),
    .RESET_B(_0042_),
    .Q(\hkspi.addr[1] ));
 sky130_fd_sc_hd__dfrtp_1 _8800_ (.CLK(clknet_2_1_0_mgmt_gpio_in[4]),
    .D(_0092_),
    .RESET_B(_0043_),
    .Q(\hkspi.addr[2] ));
 sky130_fd_sc_hd__dfrtp_1 _8801_ (.CLK(clknet_2_1_0_mgmt_gpio_in[4]),
    .D(_0093_),
    .RESET_B(_0044_),
    .Q(\hkspi.addr[3] ));
 sky130_fd_sc_hd__dfrtp_1 _8802_ (.CLK(clknet_2_1_0_mgmt_gpio_in[4]),
    .D(_0094_),
    .RESET_B(_0045_),
    .Q(\hkspi.addr[4] ));
 sky130_fd_sc_hd__dfrtp_1 _8803_ (.CLK(clknet_2_1_0_mgmt_gpio_in[4]),
    .D(_0095_),
    .RESET_B(_0046_),
    .Q(\hkspi.addr[5] ));
 sky130_fd_sc_hd__dfrtp_1 _8804_ (.CLK(clknet_2_1_0_mgmt_gpio_in[4]),
    .D(_0096_),
    .RESET_B(_0047_),
    .Q(\hkspi.addr[6] ));
 sky130_fd_sc_hd__dfrtp_1 _8805_ (.CLK(clknet_2_1_0_mgmt_gpio_in[4]),
    .D(_0097_),
    .RESET_B(_0048_),
    .Q(\hkspi.addr[7] ));
 sky130_fd_sc_hd__dfrtp_1 _8806_ (.CLK(clknet_2_1_0_mgmt_gpio_in[4]),
    .D(_0098_),
    .RESET_B(_0049_),
    .Q(\hkspi.count[0] ));
 sky130_fd_sc_hd__dfrtp_2 _8807_ (.CLK(clknet_2_0_0_mgmt_gpio_in[4]),
    .D(_0099_),
    .RESET_B(_0050_),
    .Q(\hkspi.count[1] ));
 sky130_fd_sc_hd__dfrtp_4 _8808_ (.CLK(clknet_2_1_0_mgmt_gpio_in[4]),
    .D(_0100_),
    .RESET_B(_0051_),
    .Q(\hkspi.count[2] ));
 sky130_fd_sc_hd__dfstp_1 _8809_ (.CLK(clknet_leaf_79_csclk),
    .D(_0101_),
    .SET_B(net414),
    .Q(net298));
 sky130_fd_sc_hd__dfstp_2 _8810_ (.CLK(clknet_leaf_67_csclk),
    .D(_0102_),
    .SET_B(net427),
    .Q(net299));
 sky130_fd_sc_hd__dfstp_2 _8811_ (.CLK(clknet_leaf_78_csclk),
    .D(_0103_),
    .SET_B(net427),
    .Q(net275));
 sky130_fd_sc_hd__dfstp_2 _8812_ (.CLK(clknet_leaf_68_csclk),
    .D(_0104_),
    .SET_B(net427),
    .Q(net276));
 sky130_fd_sc_hd__dfrtp_2 _8813_ (.CLK(clknet_leaf_67_csclk),
    .D(_0105_),
    .RESET_B(net428),
    .Q(net277));
 sky130_fd_sc_hd__dfstp_2 _8814_ (.CLK(clknet_leaf_80_csclk),
    .D(_0106_),
    .SET_B(net411),
    .Q(net278));
 sky130_fd_sc_hd__dfstp_2 _8815_ (.CLK(clknet_leaf_80_csclk),
    .D(_0107_),
    .SET_B(net411),
    .Q(net279));
 sky130_fd_sc_hd__dfstp_2 _8816_ (.CLK(clknet_leaf_80_csclk),
    .D(_0108_),
    .SET_B(net411),
    .Q(net280));
 sky130_fd_sc_hd__dfstp_1 _8817_ (.CLK(clknet_leaf_78_csclk),
    .D(_0109_),
    .SET_B(net414),
    .Q(net274));
 sky130_fd_sc_hd__dfstp_2 _8818_ (.CLK(clknet_leaf_67_csclk),
    .D(_0110_),
    .SET_B(net430),
    .Q(net285));
 sky130_fd_sc_hd__dfstp_1 _8819_ (.CLK(clknet_leaf_78_csclk),
    .D(_0111_),
    .SET_B(net414),
    .Q(net292));
 sky130_fd_sc_hd__dfstp_2 _8820_ (.CLK(clknet_leaf_67_csclk),
    .D(_0112_),
    .SET_B(net430),
    .Q(net293));
 sky130_fd_sc_hd__dfstp_2 _8821_ (.CLK(clknet_leaf_67_csclk),
    .D(_0113_),
    .SET_B(net430),
    .Q(net294));
 sky130_fd_sc_hd__dfstp_1 _8822_ (.CLK(clknet_leaf_80_csclk),
    .D(_0114_),
    .SET_B(net412),
    .Q(net295));
 sky130_fd_sc_hd__dfstp_2 _8823_ (.CLK(clknet_leaf_80_csclk),
    .D(_0115_),
    .SET_B(net412),
    .Q(net296));
 sky130_fd_sc_hd__dfstp_1 _8824_ (.CLK(clknet_leaf_80_csclk),
    .D(_0116_),
    .SET_B(net412),
    .Q(net297));
 sky130_fd_sc_hd__dfstp_1 _8825_ (.CLK(clknet_leaf_68_csclk),
    .D(_0117_),
    .SET_B(net427),
    .Q(net290));
 sky130_fd_sc_hd__dfstp_1 _8826_ (.CLK(clknet_leaf_68_csclk),
    .D(_0118_),
    .SET_B(net427),
    .Q(net291));
 sky130_fd_sc_hd__dfstp_1 _8827_ (.CLK(clknet_2_1_0_mgmt_gpio_in[4]),
    .D(net1515),
    .SET_B(_0052_),
    .Q(\hkspi.state[0] ));
 sky130_fd_sc_hd__dfrtp_1 _8828_ (.CLK(clknet_2_0_0_mgmt_gpio_in[4]),
    .D(net1456),
    .RESET_B(_0053_),
    .Q(\hkspi.state[1] ));
 sky130_fd_sc_hd__dfrtp_4 _8829_ (.CLK(clknet_2_0_0_mgmt_gpio_in[4]),
    .D(_0006_),
    .RESET_B(_0054_),
    .Q(\hkspi.state[2] ));
 sky130_fd_sc_hd__dfrtp_4 _8830_ (.CLK(clknet_2_0_0_mgmt_gpio_in[4]),
    .D(net1501),
    .RESET_B(_0055_),
    .Q(\hkspi.state[3] ));
 sky130_fd_sc_hd__dfrtp_1 _8831_ (.CLK(clknet_2_0_0_mgmt_gpio_in[4]),
    .D(_0008_),
    .RESET_B(_0056_),
    .Q(\hkspi.state[4] ));
 sky130_fd_sc_hd__dfrtp_1 _8832_ (.CLK(clknet_leaf_39_csclk),
    .D(_0119_),
    .RESET_B(net493),
    .Q(\mgmt_gpio_data_buf[16] ));
 sky130_fd_sc_hd__dfrtp_1 _8833_ (.CLK(clknet_leaf_37_csclk),
    .D(_0120_),
    .RESET_B(net493),
    .Q(\mgmt_gpio_data_buf[17] ));
 sky130_fd_sc_hd__dfrtp_1 _8834_ (.CLK(clknet_leaf_37_csclk),
    .D(_0121_),
    .RESET_B(net494),
    .Q(\mgmt_gpio_data_buf[18] ));
 sky130_fd_sc_hd__dfrtp_1 _8835_ (.CLK(clknet_leaf_37_csclk),
    .D(_0122_),
    .RESET_B(net494),
    .Q(\mgmt_gpio_data_buf[19] ));
 sky130_fd_sc_hd__dfrtp_1 _8836_ (.CLK(clknet_leaf_30_csclk),
    .D(_0123_),
    .RESET_B(net477),
    .Q(\mgmt_gpio_data_buf[20] ));
 sky130_fd_sc_hd__dfrtp_1 _8837_ (.CLK(clknet_leaf_29_csclk),
    .D(_0124_),
    .RESET_B(net477),
    .Q(\mgmt_gpio_data_buf[21] ));
 sky130_fd_sc_hd__dfrtp_1 _8838_ (.CLK(clknet_leaf_29_csclk),
    .D(_0125_),
    .RESET_B(net477),
    .Q(\mgmt_gpio_data_buf[22] ));
 sky130_fd_sc_hd__dfrtp_1 _8839_ (.CLK(clknet_leaf_31_csclk),
    .D(_0126_),
    .RESET_B(net481),
    .Q(\mgmt_gpio_data_buf[23] ));
 sky130_fd_sc_hd__dfrtp_1 _8840_ (.CLK(clknet_leaf_39_csclk),
    .D(_0127_),
    .RESET_B(net486),
    .Q(\mgmt_gpio_data_buf[8] ));
 sky130_fd_sc_hd__dfrtp_1 _8841_ (.CLK(clknet_leaf_37_csclk),
    .D(_0128_),
    .RESET_B(net493),
    .Q(\mgmt_gpio_data_buf[9] ));
 sky130_fd_sc_hd__dfrtp_1 _8842_ (.CLK(clknet_leaf_39_csclk),
    .D(_0129_),
    .RESET_B(net486),
    .Q(\mgmt_gpio_data_buf[10] ));
 sky130_fd_sc_hd__dfrtp_1 _8843_ (.CLK(clknet_leaf_37_csclk),
    .D(_0130_),
    .RESET_B(net493),
    .Q(\mgmt_gpio_data_buf[11] ));
 sky130_fd_sc_hd__dfrtp_1 _8844_ (.CLK(clknet_leaf_38_csclk),
    .D(_0131_),
    .RESET_B(net493),
    .Q(\mgmt_gpio_data_buf[12] ));
 sky130_fd_sc_hd__dfrtp_1 _8845_ (.CLK(clknet_leaf_37_csclk),
    .D(_0132_),
    .RESET_B(net489),
    .Q(\mgmt_gpio_data_buf[13] ));
 sky130_fd_sc_hd__dfrtp_1 _8846_ (.CLK(clknet_leaf_37_csclk),
    .D(_0133_),
    .RESET_B(net493),
    .Q(\mgmt_gpio_data_buf[14] ));
 sky130_fd_sc_hd__dfrtp_1 _8847_ (.CLK(clknet_leaf_37_csclk),
    .D(_0134_),
    .RESET_B(net491),
    .Q(\mgmt_gpio_data_buf[15] ));
 sky130_fd_sc_hd__dfrtp_4 _8848_ (.CLK(clknet_leaf_64_csclk),
    .D(_0135_),
    .RESET_B(net443),
    .Q(\gpio_configure[0][8] ));
 sky130_fd_sc_hd__dfrtp_4 _8849_ (.CLK(clknet_leaf_58_csclk),
    .D(_0136_),
    .RESET_B(net447),
    .Q(\gpio_configure[0][9] ));
 sky130_fd_sc_hd__dfrtp_4 _8850_ (.CLK(clknet_leaf_58_csclk),
    .D(_0137_),
    .RESET_B(net447),
    .Q(\gpio_configure[0][10] ));
 sky130_fd_sc_hd__dfstp_2 _8851_ (.CLK(clknet_leaf_58_csclk),
    .D(_0138_),
    .SET_B(net447),
    .Q(\gpio_configure[0][11] ));
 sky130_fd_sc_hd__dfstp_1 _8852_ (.CLK(clknet_leaf_64_csclk),
    .D(_0139_),
    .SET_B(net444),
    .Q(\gpio_configure[0][12] ));
 sky130_fd_sc_hd__dfrtp_4 _8853_ (.CLK(clknet_leaf_63_csclk),
    .D(_0140_),
    .RESET_B(net443),
    .Q(\gpio_configure[1][8] ));
 sky130_fd_sc_hd__dfrtp_4 _8854_ (.CLK(clknet_leaf_58_csclk),
    .D(_0141_),
    .RESET_B(net445),
    .Q(\gpio_configure[1][9] ));
 sky130_fd_sc_hd__dfrtp_4 _8855_ (.CLK(clknet_leaf_58_csclk),
    .D(_0142_),
    .RESET_B(net445),
    .Q(\gpio_configure[1][10] ));
 sky130_fd_sc_hd__dfstp_1 _8856_ (.CLK(clknet_leaf_58_csclk),
    .D(_0143_),
    .SET_B(net445),
    .Q(\gpio_configure[1][11] ));
 sky130_fd_sc_hd__dfstp_2 _8857_ (.CLK(clknet_leaf_63_csclk),
    .D(_0144_),
    .SET_B(net443),
    .Q(\gpio_configure[1][12] ));
 sky130_fd_sc_hd__dfrtp_4 _8858_ (.CLK(clknet_leaf_69_csclk),
    .D(_0145_),
    .RESET_B(net434),
    .Q(\gpio_configure[4][8] ));
 sky130_fd_sc_hd__dfrtp_4 _8859_ (.CLK(clknet_leaf_63_csclk),
    .D(_0146_),
    .RESET_B(net443),
    .Q(\gpio_configure[4][9] ));
 sky130_fd_sc_hd__dfstp_2 _8860_ (.CLK(clknet_leaf_63_csclk),
    .D(_0147_),
    .SET_B(net443),
    .Q(\gpio_configure[4][10] ));
 sky130_fd_sc_hd__dfrtp_4 _8861_ (.CLK(clknet_leaf_63_csclk),
    .D(_0148_),
    .RESET_B(net443),
    .Q(\gpio_configure[4][11] ));
 sky130_fd_sc_hd__dfrtp_2 _8862_ (.CLK(clknet_leaf_69_csclk),
    .D(_0149_),
    .RESET_B(net433),
    .Q(\gpio_configure[4][12] ));
 sky130_fd_sc_hd__dfrtp_4 _8863_ (.CLK(clknet_leaf_27_csclk),
    .D(_0150_),
    .RESET_B(net471),
    .Q(\gpio_configure[10][8] ));
 sky130_fd_sc_hd__dfrtp_4 _8864_ (.CLK(clknet_leaf_35_csclk),
    .D(_0151_),
    .RESET_B(net484),
    .Q(\gpio_configure[10][9] ));
 sky130_fd_sc_hd__dfstp_2 _8865_ (.CLK(clknet_leaf_35_csclk),
    .D(_0152_),
    .SET_B(net489),
    .Q(\gpio_configure[10][10] ));
 sky130_fd_sc_hd__dfrtp_4 _8866_ (.CLK(clknet_leaf_41_csclk),
    .D(_0153_),
    .RESET_B(net485),
    .Q(\gpio_configure[10][11] ));
 sky130_fd_sc_hd__dfrtp_4 _8867_ (.CLK(clknet_leaf_28_csclk),
    .D(_0154_),
    .RESET_B(net471),
    .Q(\gpio_configure[10][12] ));
 sky130_fd_sc_hd__dfrtp_4 _8868_ (.CLK(clknet_leaf_27_csclk),
    .D(_0155_),
    .RESET_B(net471),
    .Q(\gpio_configure[11][8] ));
 sky130_fd_sc_hd__dfrtp_4 _8869_ (.CLK(clknet_leaf_40_csclk),
    .D(_0156_),
    .RESET_B(net486),
    .Q(\gpio_configure[11][9] ));
 sky130_fd_sc_hd__dfstp_2 _8870_ (.CLK(clknet_leaf_40_csclk),
    .D(_0157_),
    .SET_B(net486),
    .Q(\gpio_configure[11][10] ));
 sky130_fd_sc_hd__dfrtp_4 _8871_ (.CLK(clknet_leaf_40_csclk),
    .D(_0158_),
    .RESET_B(net488),
    .Q(\gpio_configure[11][11] ));
 sky130_fd_sc_hd__dfrtp_4 _8872_ (.CLK(clknet_leaf_25_csclk),
    .D(_0159_),
    .RESET_B(net474),
    .Q(\gpio_configure[11][12] ));
 sky130_fd_sc_hd__dfrtp_4 _8873_ (.CLK(clknet_leaf_26_csclk),
    .D(_0160_),
    .RESET_B(net471),
    .Q(\gpio_configure[12][8] ));
 sky130_fd_sc_hd__dfrtp_2 _8874_ (.CLK(clknet_leaf_41_csclk),
    .D(_0161_),
    .RESET_B(net486),
    .Q(\gpio_configure[12][9] ));
 sky130_fd_sc_hd__dfstp_1 _8875_ (.CLK(clknet_leaf_41_csclk),
    .D(_0162_),
    .SET_B(net485),
    .Q(\gpio_configure[12][10] ));
 sky130_fd_sc_hd__dfrtp_4 _8876_ (.CLK(clknet_leaf_41_csclk),
    .D(_0163_),
    .RESET_B(net486),
    .Q(\gpio_configure[12][11] ));
 sky130_fd_sc_hd__dfrtp_4 _8877_ (.CLK(clknet_leaf_26_csclk),
    .D(_0164_),
    .RESET_B(net471),
    .Q(\gpio_configure[12][12] ));
 sky130_fd_sc_hd__dfrtp_4 _8878_ (.CLK(clknet_leaf_70_csclk),
    .D(_0165_),
    .RESET_B(net433),
    .Q(\gpio_configure[13][8] ));
 sky130_fd_sc_hd__dfrtp_4 _8879_ (.CLK(clknet_leaf_58_csclk),
    .D(_0166_),
    .RESET_B(net447),
    .Q(\gpio_configure[13][9] ));
 sky130_fd_sc_hd__dfstp_2 _8880_ (.CLK(clknet_leaf_57_csclk),
    .D(_0167_),
    .SET_B(net447),
    .Q(\gpio_configure[13][10] ));
 sky130_fd_sc_hd__dfrtp_4 _8881_ (.CLK(clknet_leaf_58_csclk),
    .D(_0168_),
    .RESET_B(net444),
    .Q(\gpio_configure[13][11] ));
 sky130_fd_sc_hd__dfrtp_1 _8882_ (.CLK(clknet_leaf_70_csclk),
    .D(_0169_),
    .RESET_B(net433),
    .Q(\gpio_configure[13][12] ));
 sky130_fd_sc_hd__dfrtp_4 _8883_ (.CLK(clknet_leaf_33_csclk),
    .D(_0170_),
    .RESET_B(net473),
    .Q(\gpio_configure[14][8] ));
 sky130_fd_sc_hd__dfrtp_2 _8884_ (.CLK(clknet_leaf_34_csclk),
    .D(_0171_),
    .RESET_B(net484),
    .Q(\gpio_configure[14][9] ));
 sky130_fd_sc_hd__dfstp_1 _8885_ (.CLK(clknet_leaf_34_csclk),
    .D(_0172_),
    .SET_B(net484),
    .Q(\gpio_configure[14][10] ));
 sky130_fd_sc_hd__dfrtp_4 _8886_ (.CLK(clknet_leaf_34_csclk),
    .D(_0173_),
    .RESET_B(net484),
    .Q(\gpio_configure[14][11] ));
 sky130_fd_sc_hd__dfrtp_4 _8887_ (.CLK(clknet_leaf_33_csclk),
    .D(_0174_),
    .RESET_B(net473),
    .Q(\gpio_configure[14][12] ));
 sky130_fd_sc_hd__dfrtp_2 _8888_ (.CLK(clknet_leaf_57_csclk),
    .D(_0175_),
    .RESET_B(net444),
    .Q(\gpio_configure[15][8] ));
 sky130_fd_sc_hd__dfrtp_4 _8889_ (.CLK(clknet_leaf_57_csclk),
    .D(_0176_),
    .RESET_B(net453),
    .Q(\gpio_configure[15][9] ));
 sky130_fd_sc_hd__dfstp_2 _8890_ (.CLK(clknet_leaf_57_csclk),
    .D(_0177_),
    .SET_B(net451),
    .Q(\gpio_configure[15][10] ));
 sky130_fd_sc_hd__dfrtp_1 _8891_ (.CLK(clknet_leaf_57_csclk),
    .D(_0178_),
    .RESET_B(net453),
    .Q(\gpio_configure[15][11] ));
 sky130_fd_sc_hd__dfrtp_4 _8892_ (.CLK(clknet_leaf_57_csclk),
    .D(_0179_),
    .RESET_B(net444),
    .Q(\gpio_configure[15][12] ));
 sky130_fd_sc_hd__dfrtp_1 _8893_ (.CLK(clknet_leaf_67_csclk),
    .D(_0180_),
    .RESET_B(net430),
    .Q(\gpio_configure[37][8] ));
 sky130_fd_sc_hd__dfrtp_4 _8894_ (.CLK(clknet_leaf_63_csclk),
    .D(_0181_),
    .RESET_B(net432),
    .Q(\gpio_configure[37][9] ));
 sky130_fd_sc_hd__dfrtp_4 _8895_ (.CLK(clknet_leaf_66_csclk),
    .D(_0182_),
    .RESET_B(net432),
    .Q(\gpio_configure[37][10] ));
 sky130_fd_sc_hd__dfstp_1 _8896_ (.CLK(clknet_leaf_66_csclk),
    .D(_0183_),
    .SET_B(net432),
    .Q(\gpio_configure[37][11] ));
 sky130_fd_sc_hd__dfstp_1 _8897_ (.CLK(clknet_leaf_67_csclk),
    .D(_0184_),
    .SET_B(net430),
    .Q(\gpio_configure[37][12] ));
 sky130_fd_sc_hd__dfrtp_4 _8898_ (.CLK(clknet_leaf_66_csclk),
    .D(_0185_),
    .RESET_B(net436),
    .Q(\gpio_configure[35][8] ));
 sky130_fd_sc_hd__dfrtp_4 _8899_ (.CLK(clknet_leaf_62_csclk),
    .D(_0186_),
    .RESET_B(net436),
    .Q(\gpio_configure[35][9] ));
 sky130_fd_sc_hd__dfstp_2 _8900_ (.CLK(clknet_leaf_62_csclk),
    .D(_0187_),
    .SET_B(net438),
    .Q(\gpio_configure[35][10] ));
 sky130_fd_sc_hd__dfrtp_2 _8901_ (.CLK(clknet_leaf_63_csclk),
    .D(_0188_),
    .RESET_B(net438),
    .Q(\gpio_configure[35][11] ));
 sky130_fd_sc_hd__dfrtp_4 _8902_ (.CLK(clknet_leaf_62_csclk),
    .D(_0189_),
    .RESET_B(net436),
    .Q(\gpio_configure[35][12] ));
 sky130_fd_sc_hd__dfrtp_4 _8903_ (.CLK(clknet_leaf_62_csclk),
    .D(_0190_),
    .RESET_B(net436),
    .Q(\gpio_configure[17][8] ));
 sky130_fd_sc_hd__dfrtp_4 _8904_ (.CLK(clknet_leaf_63_csclk),
    .D(_0191_),
    .RESET_B(net438),
    .Q(\gpio_configure[17][9] ));
 sky130_fd_sc_hd__dfstp_2 _8905_ (.CLK(clknet_leaf_62_csclk),
    .D(_0192_),
    .SET_B(net436),
    .Q(\gpio_configure[17][10] ));
 sky130_fd_sc_hd__dfrtp_4 _8906_ (.CLK(clknet_leaf_62_csclk),
    .D(_0193_),
    .RESET_B(net436),
    .Q(\gpio_configure[17][11] ));
 sky130_fd_sc_hd__dfrtp_4 _8907_ (.CLK(clknet_leaf_62_csclk),
    .D(_0194_),
    .RESET_B(net436),
    .Q(\gpio_configure[17][12] ));
 sky130_fd_sc_hd__dfrtp_1 _8908_ (.CLK(clknet_leaf_69_csclk),
    .D(_0195_),
    .RESET_B(net429),
    .Q(\gpio_configure[34][8] ));
 sky130_fd_sc_hd__dfrtp_1 _8909_ (.CLK(clknet_leaf_53_csclk),
    .D(_0196_),
    .RESET_B(net469),
    .Q(\gpio_configure[34][9] ));
 sky130_fd_sc_hd__dfstp_1 _8910_ (.CLK(clknet_leaf_63_csclk),
    .D(_0197_),
    .SET_B(net438),
    .Q(\gpio_configure[34][10] ));
 sky130_fd_sc_hd__dfrtp_1 _8911_ (.CLK(clknet_leaf_57_csclk),
    .D(_0198_),
    .RESET_B(net453),
    .Q(\gpio_configure[34][11] ));
 sky130_fd_sc_hd__dfrtp_4 _8912_ (.CLK(clknet_leaf_48_csclk),
    .D(_0199_),
    .RESET_B(net450),
    .Q(\gpio_configure[34][12] ));
 sky130_fd_sc_hd__dfrtp_4 _8913_ (.CLK(clknet_leaf_30_csclk),
    .D(_0200_),
    .RESET_B(net478),
    .Q(\gpio_configure[18][8] ));
 sky130_fd_sc_hd__dfrtp_4 _8914_ (.CLK(clknet_leaf_37_csclk),
    .D(_0201_),
    .RESET_B(net492),
    .Q(\gpio_configure[18][9] ));
 sky130_fd_sc_hd__dfstp_1 _8915_ (.CLK(clknet_leaf_37_csclk),
    .D(_0202_),
    .SET_B(net492),
    .Q(\gpio_configure[18][10] ));
 sky130_fd_sc_hd__dfrtp_4 _8916_ (.CLK(clknet_leaf_35_csclk),
    .D(_0203_),
    .RESET_B(net490),
    .Q(\gpio_configure[18][11] ));
 sky130_fd_sc_hd__dfrtp_4 _8917_ (.CLK(clknet_leaf_33_csclk),
    .D(_0204_),
    .RESET_B(net474),
    .Q(\gpio_configure[18][12] ));
 sky130_fd_sc_hd__dfrtp_2 _8918_ (.CLK(clknet_leaf_70_csclk),
    .D(_0205_),
    .RESET_B(net434),
    .Q(\gpio_configure[33][8] ));
 sky130_fd_sc_hd__dfrtp_4 _8919_ (.CLK(clknet_leaf_57_csclk),
    .D(_0206_),
    .RESET_B(net444),
    .Q(\gpio_configure[33][9] ));
 sky130_fd_sc_hd__dfstp_2 _8920_ (.CLK(clknet_leaf_58_csclk),
    .D(_0207_),
    .SET_B(net444),
    .Q(\gpio_configure[33][10] ));
 sky130_fd_sc_hd__dfrtp_1 _8921_ (.CLK(clknet_leaf_58_csclk),
    .D(_0208_),
    .RESET_B(net444),
    .Q(\gpio_configure[33][11] ));
 sky130_fd_sc_hd__dfrtp_1 _8922_ (.CLK(clknet_leaf_70_csclk),
    .D(_0209_),
    .RESET_B(net433),
    .Q(\gpio_configure[33][12] ));
 sky130_fd_sc_hd__dfrtp_4 _8923_ (.CLK(clknet_leaf_28_csclk),
    .D(_0210_),
    .RESET_B(net475),
    .Q(\gpio_configure[19][8] ));
 sky130_fd_sc_hd__dfrtp_4 _8924_ (.CLK(clknet_leaf_35_csclk),
    .D(_0211_),
    .RESET_B(net489),
    .Q(\gpio_configure[19][9] ));
 sky130_fd_sc_hd__dfstp_2 _8925_ (.CLK(clknet_leaf_34_csclk),
    .D(_0212_),
    .SET_B(net489),
    .Q(\gpio_configure[19][10] ));
 sky130_fd_sc_hd__dfrtp_4 _8926_ (.CLK(clknet_leaf_35_csclk),
    .D(_0213_),
    .RESET_B(net489),
    .Q(\gpio_configure[19][11] ));
 sky130_fd_sc_hd__dfrtp_4 _8927_ (.CLK(clknet_leaf_28_csclk),
    .D(_0214_),
    .RESET_B(net475),
    .Q(\gpio_configure[19][12] ));
 sky130_fd_sc_hd__dfrtp_1 _8928_ (.CLK(clknet_leaf_67_csclk),
    .D(_0215_),
    .RESET_B(net432),
    .Q(\gpio_configure[32][8] ));
 sky130_fd_sc_hd__dfrtp_1 _8929_ (.CLK(clknet_leaf_66_csclk),
    .D(_0216_),
    .RESET_B(net438),
    .Q(\gpio_configure[32][9] ));
 sky130_fd_sc_hd__dfstp_1 _8930_ (.CLK(clknet_leaf_63_csclk),
    .D(_0217_),
    .SET_B(net439),
    .Q(\gpio_configure[32][10] ));
 sky130_fd_sc_hd__dfrtp_1 _8931_ (.CLK(clknet_leaf_63_csclk),
    .D(_0218_),
    .RESET_B(net438),
    .Q(\gpio_configure[32][11] ));
 sky130_fd_sc_hd__dfrtp_1 _8932_ (.CLK(clknet_leaf_67_csclk),
    .D(_0219_),
    .RESET_B(net432),
    .Q(\gpio_configure[32][12] ));
 sky130_fd_sc_hd__dfrtp_4 _8933_ (.CLK(clknet_leaf_28_csclk),
    .D(_0220_),
    .RESET_B(net476),
    .Q(\gpio_configure[20][8] ));
 sky130_fd_sc_hd__dfrtp_4 _8934_ (.CLK(clknet_leaf_35_csclk),
    .D(_0221_),
    .RESET_B(net490),
    .Q(\gpio_configure[20][9] ));
 sky130_fd_sc_hd__dfstp_4 _8935_ (.CLK(clknet_leaf_35_csclk),
    .D(_0222_),
    .SET_B(net490),
    .Q(\gpio_configure[20][10] ));
 sky130_fd_sc_hd__dfrtp_4 _8936_ (.CLK(clknet_leaf_35_csclk),
    .D(_0223_),
    .RESET_B(net490),
    .Q(\gpio_configure[20][11] ));
 sky130_fd_sc_hd__dfrtp_4 _8937_ (.CLK(clknet_leaf_26_csclk),
    .D(_0224_),
    .RESET_B(net472),
    .Q(\gpio_configure[20][12] ));
 sky130_fd_sc_hd__dfrtp_4 _8938_ (.CLK(clknet_leaf_70_csclk),
    .D(_0225_),
    .RESET_B(net433),
    .Q(\gpio_configure[31][8] ));
 sky130_fd_sc_hd__dfrtp_4 _8939_ (.CLK(clknet_leaf_60_csclk),
    .D(_0226_),
    .RESET_B(net445),
    .Q(\gpio_configure[31][9] ));
 sky130_fd_sc_hd__dfstp_4 _8940_ (.CLK(clknet_leaf_59_csclk),
    .D(_0227_),
    .SET_B(net445),
    .Q(\gpio_configure[31][10] ));
 sky130_fd_sc_hd__dfrtp_2 _8941_ (.CLK(clknet_leaf_59_csclk),
    .D(_0228_),
    .RESET_B(net445),
    .Q(\gpio_configure[31][11] ));
 sky130_fd_sc_hd__dfrtp_2 _8942_ (.CLK(clknet_leaf_65_csclk),
    .D(_0229_),
    .RESET_B(net433),
    .Q(\gpio_configure[31][12] ));
 sky130_fd_sc_hd__dfrtp_4 _8943_ (.CLK(clknet_leaf_57_csclk),
    .D(_0230_),
    .RESET_B(net444),
    .Q(\gpio_configure[21][8] ));
 sky130_fd_sc_hd__dfrtp_2 _8944_ (.CLK(clknet_leaf_43_csclk),
    .D(_0231_),
    .RESET_B(net469),
    .Q(\gpio_configure[21][9] ));
 sky130_fd_sc_hd__dfstp_1 _8945_ (.CLK(clknet_leaf_55_csclk),
    .D(_0232_),
    .SET_B(net454),
    .Q(\gpio_configure[21][10] ));
 sky130_fd_sc_hd__dfrtp_1 _8946_ (.CLK(clknet_leaf_57_csclk),
    .D(_0233_),
    .RESET_B(net453),
    .Q(\gpio_configure[21][11] ));
 sky130_fd_sc_hd__dfrtp_4 _8947_ (.CLK(clknet_leaf_55_csclk),
    .D(_0234_),
    .RESET_B(net454),
    .Q(\gpio_configure[21][12] ));
 sky130_fd_sc_hd__dfrtp_4 _8948_ (.CLK(clknet_leaf_28_csclk),
    .D(_0235_),
    .RESET_B(net476),
    .Q(\gpio_configure[30][8] ));
 sky130_fd_sc_hd__dfrtp_4 _8949_ (.CLK(clknet_leaf_34_csclk),
    .D(_0236_),
    .RESET_B(net485),
    .Q(\gpio_configure[30][9] ));
 sky130_fd_sc_hd__dfstp_2 _8950_ (.CLK(clknet_leaf_36_csclk),
    .D(_0237_),
    .SET_B(net489),
    .Q(\gpio_configure[30][10] ));
 sky130_fd_sc_hd__dfrtp_4 _8951_ (.CLK(clknet_leaf_35_csclk),
    .D(_0238_),
    .RESET_B(net489),
    .Q(\gpio_configure[30][11] ));
 sky130_fd_sc_hd__dfrtp_4 _8952_ (.CLK(clknet_leaf_28_csclk),
    .D(_0239_),
    .RESET_B(net476),
    .Q(\gpio_configure[30][12] ));
 sky130_fd_sc_hd__dfrtp_1 _8953_ (.CLK(clknet_leaf_49_csclk),
    .D(_0240_),
    .RESET_B(net450),
    .Q(\gpio_configure[22][8] ));
 sky130_fd_sc_hd__dfrtp_1 _8954_ (.CLK(clknet_3_6_0_csclk),
    .D(_0241_),
    .RESET_B(net469),
    .Q(\gpio_configure[22][9] ));
 sky130_fd_sc_hd__dfstp_2 _8955_ (.CLK(clknet_leaf_53_csclk),
    .D(_0242_),
    .SET_B(net455),
    .Q(\gpio_configure[22][10] ));
 sky130_fd_sc_hd__dfrtp_2 _8956_ (.CLK(clknet_leaf_52_csclk),
    .D(_0243_),
    .RESET_B(net455),
    .Q(\gpio_configure[22][11] ));
 sky130_fd_sc_hd__dfrtp_1 _8957_ (.CLK(clknet_leaf_49_csclk),
    .D(_0244_),
    .RESET_B(net450),
    .Q(\gpio_configure[22][12] ));
 sky130_fd_sc_hd__dfrtp_4 _8958_ (.CLK(clknet_leaf_61_csclk),
    .D(_0245_),
    .RESET_B(net436),
    .Q(\gpio_configure[29][8] ));
 sky130_fd_sc_hd__dfrtp_1 _8959_ (.CLK(clknet_leaf_55_csclk),
    .D(_0246_),
    .RESET_B(net454),
    .Q(\gpio_configure[29][9] ));
 sky130_fd_sc_hd__dfstp_1 _8960_ (.CLK(clknet_leaf_55_csclk),
    .D(_0247_),
    .SET_B(net454),
    .Q(\gpio_configure[29][10] ));
 sky130_fd_sc_hd__dfrtp_4 _8961_ (.CLK(clknet_leaf_61_csclk),
    .D(_0248_),
    .RESET_B(net441),
    .Q(\gpio_configure[29][11] ));
 sky130_fd_sc_hd__dfrtp_4 _8962_ (.CLK(clknet_leaf_59_csclk),
    .D(_0249_),
    .RESET_B(net446),
    .Q(\gpio_configure[29][12] ));
 sky130_fd_sc_hd__dfrtp_4 _8963_ (.CLK(clknet_leaf_65_csclk),
    .D(_0250_),
    .RESET_B(net432),
    .Q(\gpio_configure[23][8] ));
 sky130_fd_sc_hd__dfrtp_4 _8964_ (.CLK(clknet_leaf_63_csclk),
    .D(_0251_),
    .RESET_B(net443),
    .Q(\gpio_configure[23][9] ));
 sky130_fd_sc_hd__dfstp_4 _8965_ (.CLK(clknet_leaf_63_csclk),
    .D(_0252_),
    .SET_B(net439),
    .Q(\gpio_configure[23][10] ));
 sky130_fd_sc_hd__dfrtp_4 _8966_ (.CLK(clknet_leaf_63_csclk),
    .D(_0253_),
    .RESET_B(net439),
    .Q(\gpio_configure[23][11] ));
 sky130_fd_sc_hd__dfrtp_2 _8967_ (.CLK(clknet_leaf_65_csclk),
    .D(_0254_),
    .RESET_B(net432),
    .Q(\gpio_configure[23][12] ));
 sky130_fd_sc_hd__dfrtp_4 _8968_ (.CLK(clknet_leaf_28_csclk),
    .D(_0255_),
    .RESET_B(net476),
    .Q(\gpio_configure[28][8] ));
 sky130_fd_sc_hd__dfrtp_4 _8969_ (.CLK(clknet_leaf_36_csclk),
    .D(_0256_),
    .RESET_B(net491),
    .Q(\gpio_configure[28][9] ));
 sky130_fd_sc_hd__dfstp_2 _8970_ (.CLK(clknet_leaf_36_csclk),
    .D(_0257_),
    .SET_B(net492),
    .Q(\gpio_configure[28][10] ));
 sky130_fd_sc_hd__dfrtp_2 _8971_ (.CLK(clknet_leaf_36_csclk),
    .D(_0258_),
    .RESET_B(net491),
    .Q(\gpio_configure[28][11] ));
 sky130_fd_sc_hd__dfrtp_4 _8972_ (.CLK(clknet_leaf_30_csclk),
    .D(_0259_),
    .RESET_B(net478),
    .Q(\gpio_configure[28][12] ));
 sky130_fd_sc_hd__dfrtp_4 _8973_ (.CLK(clknet_leaf_59_csclk),
    .D(_0260_),
    .RESET_B(net447),
    .Q(\gpio_configure[24][8] ));
 sky130_fd_sc_hd__dfrtp_2 _8974_ (.CLK(clknet_leaf_43_csclk),
    .D(_0261_),
    .RESET_B(net469),
    .Q(\gpio_configure[24][9] ));
 sky130_fd_sc_hd__dfstp_2 _8975_ (.CLK(clknet_leaf_43_csclk),
    .D(_0262_),
    .SET_B(net469),
    .Q(\gpio_configure[24][10] ));
 sky130_fd_sc_hd__dfrtp_2 _8976_ (.CLK(clknet_leaf_56_csclk),
    .D(_0263_),
    .RESET_B(net451),
    .Q(\gpio_configure[24][11] ));
 sky130_fd_sc_hd__dfrtp_4 _8977_ (.CLK(clknet_leaf_59_csclk),
    .D(_0264_),
    .RESET_B(net447),
    .Q(\gpio_configure[24][12] ));
 sky130_fd_sc_hd__dfrtp_4 _8978_ (.CLK(clknet_leaf_27_csclk),
    .D(_0265_),
    .RESET_B(net472),
    .Q(\gpio_configure[27][8] ));
 sky130_fd_sc_hd__dfrtp_2 _8979_ (.CLK(clknet_leaf_34_csclk),
    .D(_0266_),
    .RESET_B(net485),
    .Q(\gpio_configure[27][9] ));
 sky130_fd_sc_hd__dfstp_4 _8980_ (.CLK(clknet_leaf_35_csclk),
    .D(_0267_),
    .SET_B(net485),
    .Q(\gpio_configure[27][10] ));
 sky130_fd_sc_hd__dfrtp_4 _8981_ (.CLK(clknet_leaf_34_csclk),
    .D(_0268_),
    .RESET_B(net484),
    .Q(\gpio_configure[27][11] ));
 sky130_fd_sc_hd__dfrtp_4 _8982_ (.CLK(clknet_leaf_26_csclk),
    .D(_0269_),
    .RESET_B(net471),
    .Q(\gpio_configure[27][12] ));
 sky130_fd_sc_hd__dfrtp_2 _8983_ (.CLK(clknet_leaf_70_csclk),
    .D(_0270_),
    .RESET_B(net433),
    .Q(\gpio_configure[25][8] ));
 sky130_fd_sc_hd__dfrtp_4 _8984_ (.CLK(clknet_leaf_58_csclk),
    .D(_0271_),
    .RESET_B(net445),
    .Q(\gpio_configure[25][9] ));
 sky130_fd_sc_hd__dfstp_2 _8985_ (.CLK(clknet_leaf_58_csclk),
    .D(_0272_),
    .SET_B(net445),
    .Q(\gpio_configure[25][10] ));
 sky130_fd_sc_hd__dfrtp_2 _8986_ (.CLK(clknet_leaf_58_csclk),
    .D(_0273_),
    .RESET_B(net446),
    .Q(\gpio_configure[25][11] ));
 sky130_fd_sc_hd__dfrtp_2 _8987_ (.CLK(clknet_leaf_70_csclk),
    .D(_0274_),
    .RESET_B(net433),
    .Q(\gpio_configure[25][12] ));
 sky130_fd_sc_hd__dfrtp_1 _8988_ (.CLK(clknet_leaf_39_csclk),
    .D(net1570),
    .RESET_B(net486),
    .Q(\mgmt_gpio_data[16] ));
 sky130_fd_sc_hd__dfrtp_1 _8989_ (.CLK(clknet_leaf_38_csclk),
    .D(net1568),
    .RESET_B(net493),
    .Q(\mgmt_gpio_data[17] ));
 sky130_fd_sc_hd__dfrtp_1 _8990_ (.CLK(clknet_leaf_38_csclk),
    .D(net1566),
    .RESET_B(net494),
    .Q(\mgmt_gpio_data[18] ));
 sky130_fd_sc_hd__dfrtp_1 _8991_ (.CLK(clknet_leaf_38_csclk),
    .D(net1588),
    .RESET_B(net494),
    .Q(\mgmt_gpio_data[19] ));
 sky130_fd_sc_hd__dfrtp_1 _8992_ (.CLK(clknet_leaf_30_csclk),
    .D(net1586),
    .RESET_B(net478),
    .Q(\mgmt_gpio_data[20] ));
 sky130_fd_sc_hd__dfrtp_1 _8993_ (.CLK(clknet_leaf_29_csclk),
    .D(net1584),
    .RESET_B(net477),
    .Q(\mgmt_gpio_data[21] ));
 sky130_fd_sc_hd__dfrtp_1 _8994_ (.CLK(clknet_leaf_16_csclk),
    .D(net1572),
    .RESET_B(net477),
    .Q(\mgmt_gpio_data[22] ));
 sky130_fd_sc_hd__dfrtp_1 _8995_ (.CLK(clknet_leaf_31_csclk),
    .D(net1590),
    .RESET_B(net481),
    .Q(\mgmt_gpio_data[23] ));
 sky130_fd_sc_hd__dfstp_4 _8996_ (.CLK(clknet_3_2_0_wb_clk_i),
    .D(_0014_),
    .SET_B(net441),
    .Q(\xfer_state[0] ));
 sky130_fd_sc_hd__dfrtp_4 _8997_ (.CLK(clknet_3_2_0_wb_clk_i),
    .D(_0015_),
    .RESET_B(net446),
    .Q(\xfer_state[1] ));
 sky130_fd_sc_hd__dfrtp_1 _8998_ (.CLK(clknet_3_0_0_wb_clk_i),
    .D(_0016_),
    .RESET_B(net446),
    .Q(\xfer_state[2] ));
 sky130_fd_sc_hd__dfrtp_2 _8999_ (.CLK(clknet_3_2_0_wb_clk_i),
    .D(_0017_),
    .RESET_B(net446),
    .Q(\xfer_state[3] ));
 sky130_fd_sc_hd__dfrtp_2 _9000_ (.CLK(clknet_leaf_39_csclk),
    .D(_0283_),
    .RESET_B(net486),
    .Q(\mgmt_gpio_data[8] ));
 sky130_fd_sc_hd__dfrtp_2 _9001_ (.CLK(clknet_leaf_38_csclk),
    .D(net1582),
    .RESET_B(net493),
    .Q(\mgmt_gpio_data[9] ));
 sky130_fd_sc_hd__dfrtp_1 _9002_ (.CLK(clknet_leaf_39_csclk),
    .D(_0285_),
    .RESET_B(net487),
    .Q(\mgmt_gpio_data[10] ));
 sky130_fd_sc_hd__dfrtp_2 _9003_ (.CLK(clknet_leaf_38_csclk),
    .D(_0286_),
    .RESET_B(net493),
    .Q(\mgmt_gpio_data[11] ));
 sky130_fd_sc_hd__dfrtp_1 _9004_ (.CLK(clknet_leaf_38_csclk),
    .D(_0287_),
    .RESET_B(net493),
    .Q(\mgmt_gpio_data[12] ));
 sky130_fd_sc_hd__dfrtp_1 _9005_ (.CLK(clknet_leaf_35_csclk),
    .D(net1576),
    .RESET_B(net490),
    .Q(\mgmt_gpio_data[13] ));
 sky130_fd_sc_hd__dfrtp_1 _9006_ (.CLK(clknet_leaf_38_csclk),
    .D(net1578),
    .RESET_B(net494),
    .Q(\mgmt_gpio_data[14] ));
 sky130_fd_sc_hd__dfrtp_1 _9007_ (.CLK(clknet_leaf_37_csclk),
    .D(net1540),
    .RESET_B(net490),
    .Q(\mgmt_gpio_data[15] ));
 sky130_fd_sc_hd__dfrtp_4 _9008_ (.CLK(clknet_3_2_0_wb_clk_i),
    .D(_0291_),
    .RESET_B(net503),
    .Q(wbbd_busy));
 sky130_fd_sc_hd__dfrtp_1 _9009_ (.CLK(clknet_leaf_4_csclk),
    .D(net1403),
    .RESET_B(net420),
    .Q(\mgmt_gpio_data[0] ));
 sky130_fd_sc_hd__dfrtp_1 _9010_ (.CLK(clknet_leaf_4_csclk),
    .D(net1574),
    .RESET_B(net420),
    .Q(\mgmt_gpio_data[1] ));
 sky130_fd_sc_hd__dfrtp_4 _9011_ (.CLK(clknet_leaf_40_csclk),
    .D(_0294_),
    .RESET_B(net487),
    .Q(\mgmt_gpio_data[2] ));
 sky130_fd_sc_hd__dfrtp_4 _9012_ (.CLK(clknet_leaf_40_csclk),
    .D(_0295_),
    .RESET_B(net488),
    .Q(\mgmt_gpio_data[3] ));
 sky130_fd_sc_hd__dfrtp_1 _9013_ (.CLK(clknet_leaf_40_csclk),
    .D(_0296_),
    .RESET_B(net487),
    .Q(\mgmt_gpio_data[4] ));
 sky130_fd_sc_hd__dfrtp_1 _9014_ (.CLK(clknet_leaf_40_csclk),
    .D(_0297_),
    .RESET_B(net488),
    .Q(\mgmt_gpio_data[5] ));
 sky130_fd_sc_hd__dfrtp_1 _9015_ (.CLK(clknet_leaf_4_csclk),
    .D(net608),
    .RESET_B(net420),
    .Q(\mgmt_gpio_data[6] ));
 sky130_fd_sc_hd__dfrtp_2 _9016_ (.CLK(clknet_leaf_40_csclk),
    .D(_0299_),
    .RESET_B(net487),
    .Q(\mgmt_gpio_data[7] ));
 sky130_fd_sc_hd__dfrtp_1 _9017_ (.CLK(clknet_leaf_31_csclk),
    .D(_0300_),
    .RESET_B(net481),
    .Q(\mgmt_gpio_data[24] ));
 sky130_fd_sc_hd__dfrtp_1 _9018_ (.CLK(clknet_leaf_31_csclk),
    .D(net948),
    .RESET_B(net481),
    .Q(\mgmt_gpio_data[25] ));
 sky130_fd_sc_hd__dfrtp_1 _9019_ (.CLK(clknet_leaf_31_csclk),
    .D(net1030),
    .RESET_B(net481),
    .Q(\mgmt_gpio_data[26] ));
 sky130_fd_sc_hd__dfrtp_1 _9020_ (.CLK(clknet_leaf_36_csclk),
    .D(net898),
    .RESET_B(net491),
    .Q(\mgmt_gpio_data[27] ));
 sky130_fd_sc_hd__dfrtp_1 _9021_ (.CLK(clknet_leaf_36_csclk),
    .D(net660),
    .RESET_B(net491),
    .Q(\mgmt_gpio_data[28] ));
 sky130_fd_sc_hd__dfrtp_1 _9022_ (.CLK(clknet_leaf_36_csclk),
    .D(net1167),
    .RESET_B(net491),
    .Q(\mgmt_gpio_data[29] ));
 sky130_fd_sc_hd__dfrtp_1 _9023_ (.CLK(clknet_leaf_36_csclk),
    .D(net1165),
    .RESET_B(net492),
    .Q(\mgmt_gpio_data[30] ));
 sky130_fd_sc_hd__dfrtp_1 _9024_ (.CLK(clknet_leaf_37_csclk),
    .D(net988),
    .RESET_B(net492),
    .Q(\mgmt_gpio_data[31] ));
 sky130_fd_sc_hd__dfstp_1 _9025_ (.CLK(clknet_3_7_0_wb_clk_i),
    .D(_0009_),
    .SET_B(net499),
    .Q(\wbbd_state[0] ));
 sky130_fd_sc_hd__dfrtp_1 _9026_ (.CLK(clknet_3_7_0_wb_clk_i),
    .D(_0000_),
    .RESET_B(net499),
    .Q(\wbbd_state[1] ));
 sky130_fd_sc_hd__dfrtp_1 _9027_ (.CLK(clknet_3_7_0_wb_clk_i),
    .D(_0001_),
    .RESET_B(net499),
    .Q(\wbbd_state[2] ));
 sky130_fd_sc_hd__dfrtp_1 _9028_ (.CLK(clknet_3_7_0_wb_clk_i),
    .D(_0002_),
    .RESET_B(net499),
    .Q(\wbbd_state[3] ));
 sky130_fd_sc_hd__dfrtp_1 _9029_ (.CLK(clknet_3_7_0_wb_clk_i),
    .D(_0003_),
    .RESET_B(net499),
    .Q(\wbbd_state[4] ));
 sky130_fd_sc_hd__dfrtp_4 _9030_ (.CLK(clknet_3_7_0_wb_clk_i),
    .D(_0010_),
    .RESET_B(net499),
    .Q(\wbbd_state[5] ));
 sky130_fd_sc_hd__dfrtp_1 _9031_ (.CLK(clknet_3_7_0_wb_clk_i),
    .D(net1448),
    .RESET_B(net501),
    .Q(\wbbd_state[6] ));
 sky130_fd_sc_hd__dfrtp_4 _9032_ (.CLK(clknet_3_7_0_wb_clk_i),
    .D(_0011_),
    .RESET_B(net499),
    .Q(\wbbd_state[7] ));
 sky130_fd_sc_hd__dfrtp_4 _9033_ (.CLK(clknet_3_7_0_wb_clk_i),
    .D(_0012_),
    .RESET_B(net499),
    .Q(\wbbd_state[8] ));
 sky130_fd_sc_hd__dfrtp_4 _9034_ (.CLK(clknet_3_7_0_wb_clk_i),
    .D(_0013_),
    .RESET_B(net499),
    .Q(\wbbd_state[9] ));
 sky130_fd_sc_hd__dfrtp_2 _9035_ (.CLK(clknet_leaf_72_csclk),
    .D(_0308_),
    .RESET_B(net450),
    .Q(\gpio_configure[2][8] ));
 sky130_fd_sc_hd__dfrtp_1 _9036_ (.CLK(clknet_leaf_47_csclk),
    .D(_0309_),
    .RESET_B(net467),
    .Q(\gpio_configure[2][9] ));
 sky130_fd_sc_hd__dfstp_1 _9037_ (.CLK(clknet_leaf_50_csclk),
    .D(_0310_),
    .SET_B(net455),
    .Q(\gpio_configure[2][10] ));
 sky130_fd_sc_hd__dfrtp_1 _9038_ (.CLK(clknet_3_3_0_csclk),
    .D(_0311_),
    .RESET_B(net453),
    .Q(\gpio_configure[2][11] ));
 sky130_fd_sc_hd__dfrtp_1 _9039_ (.CLK(clknet_leaf_50_csclk),
    .D(_0312_),
    .RESET_B(net450),
    .Q(\gpio_configure[2][12] ));
 sky130_fd_sc_hd__dfxtp_1 _9040_ (.CLK(clknet_3_5_0_wb_clk_i),
    .D(_0313_),
    .Q(net334));
 sky130_fd_sc_hd__dfxtp_1 _9041_ (.CLK(clknet_3_5_0_wb_clk_i),
    .D(_0314_),
    .Q(net335));
 sky130_fd_sc_hd__dfxtp_1 _9042_ (.CLK(clknet_3_5_0_wb_clk_i),
    .D(_0315_),
    .Q(net336));
 sky130_fd_sc_hd__dfxtp_1 _9043_ (.CLK(clknet_3_5_0_wb_clk_i),
    .D(_0316_),
    .Q(net337));
 sky130_fd_sc_hd__dfxtp_1 _9044_ (.CLK(clknet_3_5_0_wb_clk_i),
    .D(_0317_),
    .Q(net339));
 sky130_fd_sc_hd__dfxtp_1 _9045_ (.CLK(clknet_3_5_0_wb_clk_i),
    .D(_0318_),
    .Q(net340));
 sky130_fd_sc_hd__dfxtp_1 _9046_ (.CLK(clknet_3_5_0_wb_clk_i),
    .D(_0319_),
    .Q(net341));
 sky130_fd_sc_hd__dfxtp_1 _9047_ (.CLK(clknet_3_5_0_wb_clk_i),
    .D(_0320_),
    .Q(net342));
 sky130_fd_sc_hd__dfrtp_4 _9048_ (.CLK(clknet_leaf_69_csclk),
    .D(_0321_),
    .RESET_B(net429),
    .Q(\gpio_configure[3][8] ));
 sky130_fd_sc_hd__dfrtp_4 _9049_ (.CLK(clknet_leaf_63_csclk),
    .D(_0322_),
    .RESET_B(net443),
    .Q(\gpio_configure[3][9] ));
 sky130_fd_sc_hd__dfstp_2 _9050_ (.CLK(clknet_leaf_63_csclk),
    .D(_0323_),
    .SET_B(net443),
    .Q(\gpio_configure[3][10] ));
 sky130_fd_sc_hd__dfrtp_1 _9051_ (.CLK(clknet_leaf_57_csclk),
    .D(_0324_),
    .RESET_B(net453),
    .Q(\gpio_configure[3][11] ));
 sky130_fd_sc_hd__dfrtp_2 _9052_ (.CLK(clknet_leaf_50_csclk),
    .D(_0325_),
    .RESET_B(net450),
    .Q(\gpio_configure[3][12] ));
 sky130_fd_sc_hd__dfxtp_1 _9053_ (.CLK(clknet_3_4_0_wb_clk_i),
    .D(_0326_),
    .Q(net357));
 sky130_fd_sc_hd__dfxtp_1 _9054_ (.CLK(clknet_3_4_0_wb_clk_i),
    .D(_0327_),
    .Q(net358));
 sky130_fd_sc_hd__dfxtp_1 _9055_ (.CLK(clknet_3_4_0_wb_clk_i),
    .D(_0328_),
    .Q(net328));
 sky130_fd_sc_hd__dfxtp_1 _9056_ (.CLK(clknet_3_4_0_wb_clk_i),
    .D(_0329_),
    .Q(net329));
 sky130_fd_sc_hd__dfxtp_1 _9057_ (.CLK(clknet_3_4_0_wb_clk_i),
    .D(_0330_),
    .Q(net330));
 sky130_fd_sc_hd__dfxtp_1 _9058_ (.CLK(clknet_3_5_0_wb_clk_i),
    .D(_0331_),
    .Q(net331));
 sky130_fd_sc_hd__dfxtp_1 _9059_ (.CLK(clknet_3_5_0_wb_clk_i),
    .D(_0332_),
    .Q(net332));
 sky130_fd_sc_hd__dfxtp_1 _9060_ (.CLK(clknet_3_5_0_wb_clk_i),
    .D(_0333_),
    .Q(net333));
 sky130_fd_sc_hd__dfxtp_1 _9061_ (.CLK(clknet_3_4_0_wb_clk_i),
    .D(_0334_),
    .Q(net327));
 sky130_fd_sc_hd__dfxtp_1 _9062_ (.CLK(clknet_3_4_0_wb_clk_i),
    .D(_0335_),
    .Q(net338));
 sky130_fd_sc_hd__dfxtp_1 _9063_ (.CLK(clknet_3_4_0_wb_clk_i),
    .D(_0336_),
    .Q(net349));
 sky130_fd_sc_hd__dfxtp_1 _9064_ (.CLK(clknet_3_4_0_wb_clk_i),
    .D(_0337_),
    .Q(net352));
 sky130_fd_sc_hd__dfxtp_1 _9065_ (.CLK(clknet_3_4_0_wb_clk_i),
    .D(_0338_),
    .Q(net353));
 sky130_fd_sc_hd__dfxtp_1 _9066_ (.CLK(clknet_3_4_0_wb_clk_i),
    .D(_0339_),
    .Q(net354));
 sky130_fd_sc_hd__dfxtp_1 _9067_ (.CLK(clknet_3_4_0_wb_clk_i),
    .D(_0340_),
    .Q(net355));
 sky130_fd_sc_hd__dfxtp_1 _9068_ (.CLK(clknet_3_4_0_wb_clk_i),
    .D(_0341_),
    .Q(net356));
 sky130_fd_sc_hd__dfrtp_2 _9069_ (.CLK(clknet_leaf_69_csclk),
    .D(_0342_),
    .RESET_B(net434),
    .Q(\gpio_configure[5][8] ));
 sky130_fd_sc_hd__dfrtp_4 _9070_ (.CLK(clknet_leaf_60_csclk),
    .D(_0343_),
    .RESET_B(net441),
    .Q(\gpio_configure[5][9] ));
 sky130_fd_sc_hd__dfstp_4 _9071_ (.CLK(clknet_leaf_60_csclk),
    .D(_0344_),
    .SET_B(net445),
    .Q(\gpio_configure[5][10] ));
 sky130_fd_sc_hd__dfrtp_2 _9072_ (.CLK(clknet_leaf_58_csclk),
    .D(_0345_),
    .RESET_B(net445),
    .Q(\gpio_configure[5][11] ));
 sky130_fd_sc_hd__dfrtp_2 _9073_ (.CLK(clknet_leaf_65_csclk),
    .D(_0346_),
    .RESET_B(net433),
    .Q(\gpio_configure[5][12] ));
 sky130_fd_sc_hd__dfrtp_4 _9074_ (.CLK(clknet_leaf_67_csclk),
    .D(_0347_),
    .RESET_B(net428),
    .Q(\gpio_configure[6][8] ));
 sky130_fd_sc_hd__dfrtp_4 _9075_ (.CLK(clknet_leaf_61_csclk),
    .D(_0348_),
    .RESET_B(net436),
    .Q(\gpio_configure[6][9] ));
 sky130_fd_sc_hd__dfstp_4 _9076_ (.CLK(clknet_leaf_61_csclk),
    .D(_0349_),
    .SET_B(net437),
    .Q(\gpio_configure[6][10] ));
 sky130_fd_sc_hd__dfrtp_4 _9077_ (.CLK(clknet_leaf_61_csclk),
    .D(_0350_),
    .RESET_B(net437),
    .Q(\gpio_configure[6][11] ));
 sky130_fd_sc_hd__dfrtp_4 _9078_ (.CLK(clknet_leaf_67_csclk),
    .D(_0351_),
    .RESET_B(net430),
    .Q(\gpio_configure[6][12] ));
 sky130_fd_sc_hd__dfrtp_4 _9079_ (.CLK(clknet_leaf_61_csclk),
    .D(_0352_),
    .RESET_B(net440),
    .Q(\gpio_configure[7][8] ));
 sky130_fd_sc_hd__dfrtp_4 _9080_ (.CLK(clknet_leaf_61_csclk),
    .D(_0353_),
    .RESET_B(net440),
    .Q(\gpio_configure[7][9] ));
 sky130_fd_sc_hd__dfstp_2 _9081_ (.CLK(clknet_leaf_60_csclk),
    .D(_0354_),
    .SET_B(net441),
    .Q(\gpio_configure[7][10] ));
 sky130_fd_sc_hd__dfrtp_4 _9082_ (.CLK(clknet_leaf_61_csclk),
    .D(_0355_),
    .RESET_B(net439),
    .Q(\gpio_configure[7][11] ));
 sky130_fd_sc_hd__dfrtp_4 _9083_ (.CLK(clknet_leaf_61_csclk),
    .D(_0356_),
    .RESET_B(net441),
    .Q(\gpio_configure[7][12] ));
 sky130_fd_sc_hd__dfrtp_4 _9084_ (.CLK(clknet_leaf_58_csclk),
    .D(_0357_),
    .RESET_B(net447),
    .Q(\gpio_configure[8][8] ));
 sky130_fd_sc_hd__dfrtp_2 _9085_ (.CLK(clknet_leaf_55_csclk),
    .D(_0358_),
    .RESET_B(net455),
    .Q(\gpio_configure[8][9] ));
 sky130_fd_sc_hd__dfstp_2 _9086_ (.CLK(clknet_leaf_55_csclk),
    .D(_0359_),
    .SET_B(net455),
    .Q(\gpio_configure[8][10] ));
 sky130_fd_sc_hd__dfrtp_2 _9087_ (.CLK(clknet_leaf_59_csclk),
    .D(_0360_),
    .RESET_B(net447),
    .Q(\gpio_configure[8][11] ));
 sky130_fd_sc_hd__dfrtp_4 _9088_ (.CLK(clknet_leaf_55_csclk),
    .D(_0361_),
    .RESET_B(net455),
    .Q(\gpio_configure[8][12] ));
 sky130_fd_sc_hd__dfrtp_2 _9089_ (.CLK(clknet_leaf_70_csclk),
    .D(_0362_),
    .RESET_B(net434),
    .Q(\gpio_configure[9][8] ));
 sky130_fd_sc_hd__dfrtp_4 _9090_ (.CLK(clknet_3_3_0_csclk),
    .D(_0363_),
    .RESET_B(net454),
    .Q(\gpio_configure[9][9] ));
 sky130_fd_sc_hd__dfstp_2 _9091_ (.CLK(clknet_leaf_52_csclk),
    .D(_0364_),
    .SET_B(net455),
    .Q(\gpio_configure[9][10] ));
 sky130_fd_sc_hd__dfrtp_1 _9092_ (.CLK(clknet_leaf_56_csclk),
    .D(_0365_),
    .RESET_B(net451),
    .Q(\gpio_configure[9][11] ));
 sky130_fd_sc_hd__dfrtp_1 _9093_ (.CLK(clknet_leaf_73_csclk),
    .D(_0366_),
    .RESET_B(net450),
    .Q(\gpio_configure[9][12] ));
 sky130_fd_sc_hd__dfrtp_1 _9094_ (.CLK(clknet_leaf_67_csclk),
    .D(_0367_),
    .RESET_B(net428),
    .Q(\gpio_configure[36][8] ));
 sky130_fd_sc_hd__dfrtp_1 _9095_ (.CLK(clknet_leaf_66_csclk),
    .D(_0368_),
    .RESET_B(net430),
    .Q(\gpio_configure[36][9] ));
 sky130_fd_sc_hd__dfrtp_4 _9096_ (.CLK(clknet_leaf_66_csclk),
    .D(_0369_),
    .RESET_B(net431),
    .Q(\gpio_configure[36][10] ));
 sky130_fd_sc_hd__dfstp_1 _9097_ (.CLK(clknet_leaf_66_csclk),
    .D(_0370_),
    .SET_B(net431),
    .Q(\gpio_configure[36][11] ));
 sky130_fd_sc_hd__dfstp_2 _9098_ (.CLK(clknet_leaf_67_csclk),
    .D(_0371_),
    .SET_B(net428),
    .Q(\gpio_configure[36][12] ));
 sky130_fd_sc_hd__dfrtp_4 _9099_ (.CLK(clknet_leaf_66_csclk),
    .D(_0372_),
    .RESET_B(net431),
    .Q(\gpio_configure[16][8] ));
 sky130_fd_sc_hd__dfrtp_4 _9100_ (.CLK(clknet_leaf_62_csclk),
    .D(_0373_),
    .RESET_B(net437),
    .Q(\gpio_configure[16][9] ));
 sky130_fd_sc_hd__dfstp_2 _9101_ (.CLK(clknet_leaf_62_csclk),
    .D(_0374_),
    .SET_B(net437),
    .Q(\gpio_configure[16][10] ));
 sky130_fd_sc_hd__dfrtp_4 _9102_ (.CLK(clknet_leaf_62_csclk),
    .D(_0375_),
    .RESET_B(net436),
    .Q(\gpio_configure[16][11] ));
 sky130_fd_sc_hd__dfrtp_4 _9103_ (.CLK(clknet_leaf_66_csclk),
    .D(_0376_),
    .RESET_B(net431),
    .Q(\gpio_configure[16][12] ));
 sky130_fd_sc_hd__dfrtp_4 _9104_ (.CLK(clknet_3_7_0_wb_clk_i),
    .D(_0377_),
    .RESET_B(net502),
    .Q(\wbbd_addr[0] ));
 sky130_fd_sc_hd__dfrtp_4 _9105_ (.CLK(clknet_3_7_0_wb_clk_i),
    .D(_0378_),
    .RESET_B(net502),
    .Q(\wbbd_addr[1] ));
 sky130_fd_sc_hd__dfrtp_4 _9106_ (.CLK(clknet_3_4_0_wb_clk_i),
    .D(_0379_),
    .RESET_B(net502),
    .Q(\wbbd_addr[2] ));
 sky130_fd_sc_hd__dfrtp_4 _9107_ (.CLK(clknet_3_4_0_wb_clk_i),
    .D(_0380_),
    .RESET_B(net503),
    .Q(\wbbd_addr[3] ));
 sky130_fd_sc_hd__dfrtp_4 _9108_ (.CLK(clknet_3_4_0_wb_clk_i),
    .D(_0381_),
    .RESET_B(net503),
    .Q(\wbbd_addr[4] ));
 sky130_fd_sc_hd__dfrtp_4 _9109_ (.CLK(clknet_3_4_0_wb_clk_i),
    .D(_0382_),
    .RESET_B(net503),
    .Q(\wbbd_addr[5] ));
 sky130_fd_sc_hd__dfrtp_4 _9110_ (.CLK(clknet_3_4_0_wb_clk_i),
    .D(_0383_),
    .RESET_B(net503),
    .Q(\wbbd_addr[6] ));
 sky130_fd_sc_hd__dfrtn_1 _9111_ (.CLK_N(clknet_2_2_0_mgmt_gpio_in[4]),
    .D(_0384_),
    .RESET_B(_0057_),
    .Q(\hkspi.ldata[0] ));
 sky130_fd_sc_hd__dfrtn_1 _9112_ (.CLK_N(clknet_2_2_0_mgmt_gpio_in[4]),
    .D(_0385_),
    .RESET_B(_0058_),
    .Q(\hkspi.ldata[1] ));
 sky130_fd_sc_hd__dfrtn_1 _9113_ (.CLK_N(clknet_2_2_0_mgmt_gpio_in[4]),
    .D(_0386_),
    .RESET_B(_0059_),
    .Q(\hkspi.ldata[2] ));
 sky130_fd_sc_hd__dfrtn_1 _9114_ (.CLK_N(clknet_2_2_0_mgmt_gpio_in[4]),
    .D(_0387_),
    .RESET_B(_0060_),
    .Q(\hkspi.ldata[3] ));
 sky130_fd_sc_hd__dfrtn_1 _9115_ (.CLK_N(clknet_2_2_0_mgmt_gpio_in[4]),
    .D(_0388_),
    .RESET_B(_0061_),
    .Q(\hkspi.ldata[4] ));
 sky130_fd_sc_hd__dfrtn_1 _9116_ (.CLK_N(clknet_2_2_0_mgmt_gpio_in[4]),
    .D(_0389_),
    .RESET_B(_0062_),
    .Q(\hkspi.ldata[5] ));
 sky130_fd_sc_hd__dfrtn_1 _9117_ (.CLK_N(clknet_2_2_0_mgmt_gpio_in[4]),
    .D(_0390_),
    .RESET_B(_0063_),
    .Q(\hkspi.ldata[6] ));
 sky130_fd_sc_hd__dfrtn_1 _9118_ (.CLK_N(clknet_2_2_0_mgmt_gpio_in[4]),
    .D(_0391_),
    .RESET_B(_0064_),
    .Q(\hkspi.SDO ));
 sky130_fd_sc_hd__dfrtp_2 _9119_ (.CLK(clknet_leaf_84_csclk),
    .D(_0392_),
    .RESET_B(net404),
    .Q(net270));
 sky130_fd_sc_hd__dfstp_1 _9120_ (.CLK(clknet_leaf_84_csclk),
    .D(_0393_),
    .SET_B(net404),
    .Q(net264));
 sky130_fd_sc_hd__dfrtp_2 _9121_ (.CLK(clknet_leaf_83_csclk),
    .D(_0394_),
    .RESET_B(net404),
    .Q(net265));
 sky130_fd_sc_hd__dfrtp_4 _9122_ (.CLK(clknet_leaf_83_csclk),
    .D(_0395_),
    .RESET_B(net404),
    .Q(net266));
 sky130_fd_sc_hd__dfstp_2 _9123_ (.CLK(clknet_leaf_83_csclk),
    .D(_0396_),
    .SET_B(net404),
    .Q(net267));
 sky130_fd_sc_hd__dfrtp_4 _9124_ (.CLK(clknet_leaf_83_csclk),
    .D(_0397_),
    .RESET_B(net404),
    .Q(net268));
 sky130_fd_sc_hd__dfrtp_2 _9125_ (.CLK(clknet_leaf_83_csclk),
    .D(_0398_),
    .RESET_B(net405),
    .Q(net269));
 sky130_fd_sc_hd__dfrtp_4 _9126_ (.CLK(clknet_leaf_83_csclk),
    .D(_0399_),
    .RESET_B(net405),
    .Q(net271));
 sky130_fd_sc_hd__dfstp_2 _9127_ (.CLK(clknet_leaf_83_csclk),
    .D(_0400_),
    .SET_B(net405),
    .Q(net272));
 sky130_fd_sc_hd__dfrtp_4 _9128_ (.CLK(clknet_leaf_83_csclk),
    .D(_0401_),
    .RESET_B(net405),
    .Q(net273));
 sky130_fd_sc_hd__dfrtp_4 _9129_ (.CLK(clknet_leaf_80_csclk),
    .D(_0402_),
    .RESET_B(net411),
    .Q(net260));
 sky130_fd_sc_hd__dfstp_2 _9130_ (.CLK(clknet_leaf_80_csclk),
    .D(_0403_),
    .SET_B(net411),
    .Q(net261));
 sky130_fd_sc_hd__dfrtp_1 _9131_ (.CLK(clknet_leaf_80_csclk),
    .D(_0404_),
    .RESET_B(net411),
    .Q(net262));
 sky130_fd_sc_hd__dfstp_1 _9132_ (.CLK(clknet_leaf_68_csclk),
    .D(_0405_),
    .SET_B(net427),
    .Q(net281));
 sky130_fd_sc_hd__dfstp_1 _9133_ (.CLK(clknet_leaf_67_csclk),
    .D(_0406_),
    .SET_B(net428),
    .Q(net282));
 sky130_fd_sc_hd__dfstp_2 _9134_ (.CLK(clknet_leaf_78_csclk),
    .D(_0407_),
    .SET_B(net414),
    .Q(net283));
 sky130_fd_sc_hd__dfstp_2 _9135_ (.CLK(clknet_leaf_66_csclk),
    .D(_0408_),
    .SET_B(net430),
    .Q(net284));
 sky130_fd_sc_hd__dfstp_2 _9136_ (.CLK(clknet_leaf_78_csclk),
    .D(_0409_),
    .SET_B(net414),
    .Q(net286));
 sky130_fd_sc_hd__dfstp_2 _9137_ (.CLK(clknet_leaf_79_csclk),
    .D(_0410_),
    .SET_B(net412),
    .Q(net287));
 sky130_fd_sc_hd__dfstp_2 _9138_ (.CLK(clknet_leaf_79_csclk),
    .D(_0411_),
    .SET_B(net412),
    .Q(net288));
 sky130_fd_sc_hd__dfstp_1 _9139_ (.CLK(clknet_leaf_79_csclk),
    .D(_0412_),
    .SET_B(net412),
    .Q(net289));
 sky130_fd_sc_hd__dfstp_1 _9140_ (.CLK(clknet_leaf_68_csclk),
    .D(_0413_),
    .SET_B(net427),
    .Q(net263));
 sky130_fd_sc_hd__dfrtp_4 _9141_ (.CLK(clknet_leaf_60_csclk),
    .D(_0414_),
    .RESET_B(net440),
    .Q(net300));
 sky130_fd_sc_hd__dfrtp_2 _9142_ (.CLK(clknet_leaf_60_csclk),
    .D(net1580),
    .RESET_B(net440),
    .Q(net301));
 sky130_fd_sc_hd__dfrtp_4 _9143_ (.CLK(clknet_leaf_61_csclk),
    .D(_0416_),
    .RESET_B(net437),
    .Q(net302));
 sky130_fd_sc_hd__dfrtp_4 _9144_ (.CLK(clknet_leaf_61_csclk),
    .D(_0417_),
    .RESET_B(net440),
    .Q(net303));
 sky130_fd_sc_hd__dfrtp_4 _9145_ (.CLK(clknet_leaf_85_csclk),
    .D(_0418_),
    .RESET_B(net408),
    .Q(net324));
 sky130_fd_sc_hd__dfstp_2 _9146_ (.CLK(clknet_leaf_85_csclk),
    .D(_0419_),
    .SET_B(net408),
    .Q(net325));
 sky130_fd_sc_hd__dfrtp_4 _9147_ (.CLK(clknet_leaf_84_csclk),
    .D(_0420_),
    .RESET_B(net407),
    .Q(net316));
 sky130_fd_sc_hd__dfrtp_4 _9148_ (.CLK(clknet_leaf_84_csclk),
    .D(_0421_),
    .RESET_B(net407),
    .Q(net317));
 sky130_fd_sc_hd__dfrtp_4 _9149_ (.CLK(clknet_leaf_83_csclk),
    .D(_0422_),
    .RESET_B(net404),
    .Q(net318));
 sky130_fd_sc_hd__dfrtp_4 _9150_ (.CLK(clknet_leaf_84_csclk),
    .D(_0423_),
    .RESET_B(net407),
    .Q(net319));
 sky130_fd_sc_hd__dfrtp_4 _9151_ (.CLK(clknet_leaf_84_csclk),
    .D(_0424_),
    .RESET_B(net404),
    .Q(net320));
 sky130_fd_sc_hd__dfrtp_4 _9152_ (.CLK(clknet_leaf_84_csclk),
    .D(_0425_),
    .RESET_B(net404),
    .Q(net321));
 sky130_fd_sc_hd__dfrtp_4 _9153_ (.CLK(clknet_leaf_84_csclk),
    .D(_0426_),
    .RESET_B(net407),
    .Q(net322));
 sky130_fd_sc_hd__dfrtp_4 _9154_ (.CLK(clknet_leaf_84_csclk),
    .D(_0427_),
    .RESET_B(net406),
    .Q(net323));
 sky130_fd_sc_hd__dfrtp_1 _9155_ (.CLK(clknet_leaf_85_csclk),
    .D(net1416),
    .RESET_B(net408),
    .Q(reset_reg));
 sky130_fd_sc_hd__dfrtp_4 _9156_ (.CLK(clknet_leaf_77_csclk),
    .D(net940),
    .RESET_B(net415),
    .Q(net204));
 sky130_fd_sc_hd__dfrtp_4 _9157_ (.CLK(clknet_leaf_61_csclk),
    .D(_0430_),
    .RESET_B(net440),
    .Q(serial_bb_clock));
 sky130_fd_sc_hd__dfrtp_1 _9158_ (.CLK(clknet_leaf_61_csclk),
    .D(_0431_),
    .RESET_B(net440),
    .Q(serial_bb_load));
 sky130_fd_sc_hd__dfrtp_1 _9159_ (.CLK(clknet_leaf_60_csclk),
    .D(_0432_),
    .RESET_B(net440),
    .Q(serial_bb_resetn));
 sky130_fd_sc_hd__dfrtp_1 _9160_ (.CLK(clknet_leaf_60_csclk),
    .D(net1096),
    .RESET_B(net442),
    .Q(serial_bb_data_1));
 sky130_fd_sc_hd__dfrtp_1 _9161_ (.CLK(clknet_leaf_60_csclk),
    .D(net1135),
    .RESET_B(net442),
    .Q(serial_bb_data_2));
 sky130_fd_sc_hd__dfrtp_4 _9162_ (.CLK(clknet_leaf_61_csclk),
    .D(_0435_),
    .RESET_B(net440),
    .Q(serial_bb_enable));
 sky130_fd_sc_hd__dfrtp_4 _9163_ (.CLK(clknet_leaf_77_csclk),
    .D(net1196),
    .RESET_B(net415),
    .Q(serial_xfer));
 sky130_fd_sc_hd__dfrtp_4 _9164_ (.CLK(clknet_leaf_86_csclk),
    .D(_0437_),
    .RESET_B(net408),
    .Q(hkspi_disable));
 sky130_fd_sc_hd__dfrtp_4 _9165_ (.CLK(clknet_leaf_42_csclk),
    .D(_0438_),
    .RESET_B(net484),
    .Q(clk1_output_dest));
 sky130_fd_sc_hd__dfrtp_2 _9166_ (.CLK(clknet_leaf_42_csclk),
    .D(_0439_),
    .RESET_B(net484),
    .Q(clk2_output_dest));
 sky130_fd_sc_hd__dfrtp_1 _9167_ (.CLK(clknet_leaf_42_csclk),
    .D(_0440_),
    .RESET_B(net484),
    .Q(trap_output_dest));
 sky130_fd_sc_hd__dfrtp_4 _9168_ (.CLK(clknet_leaf_85_csclk),
    .D(_0441_),
    .RESET_B(net408),
    .Q(irq_1_inputsrc));
 sky130_fd_sc_hd__dfrtp_4 _9169_ (.CLK(clknet_leaf_85_csclk),
    .D(_0442_),
    .RESET_B(net408),
    .Q(irq_2_inputsrc));
 sky130_fd_sc_hd__dfrtp_1 _9170_ (.CLK(clknet_leaf_4_csclk),
    .D(net1440),
    .RESET_B(net420),
    .Q(\mgmt_gpio_data[32] ));
 sky130_fd_sc_hd__dfrtp_1 _9171_ (.CLK(clknet_leaf_14_csclk),
    .D(net653),
    .RESET_B(net459),
    .Q(\mgmt_gpio_data[33] ));
 sky130_fd_sc_hd__dfrtp_1 _9172_ (.CLK(clknet_leaf_37_csclk),
    .D(net923),
    .RESET_B(net494),
    .Q(\mgmt_gpio_data[34] ));
 sky130_fd_sc_hd__dfrtp_1 _9173_ (.CLK(clknet_leaf_14_csclk),
    .D(net967),
    .RESET_B(net459),
    .Q(\mgmt_gpio_data[35] ));
 sky130_fd_sc_hd__dfrtp_1 _9174_ (.CLK(clknet_leaf_16_csclk),
    .D(net788),
    .RESET_B(net466),
    .Q(\mgmt_gpio_data[36] ));
 sky130_fd_sc_hd__dfrtp_1 _9175_ (.CLK(clknet_leaf_16_csclk),
    .D(net1325),
    .RESET_B(net466),
    .Q(\mgmt_gpio_data[37] ));
 sky130_fd_sc_hd__dfrtp_1 _9176_ (.CLK(clknet_leaf_4_csclk),
    .D(_0449_),
    .RESET_B(net420),
    .Q(\mgmt_gpio_data_buf[0] ));
 sky130_fd_sc_hd__dfrtp_1 _9177_ (.CLK(clknet_leaf_4_csclk),
    .D(_0450_),
    .RESET_B(net420),
    .Q(\mgmt_gpio_data_buf[1] ));
 sky130_fd_sc_hd__dfrtp_1 _9178_ (.CLK(clknet_leaf_39_csclk),
    .D(_0451_),
    .RESET_B(net487),
    .Q(\mgmt_gpio_data_buf[2] ));
 sky130_fd_sc_hd__dfrtp_1 _9179_ (.CLK(clknet_leaf_40_csclk),
    .D(_0452_),
    .RESET_B(net488),
    .Q(\mgmt_gpio_data_buf[3] ));
 sky130_fd_sc_hd__dfrtp_1 _9180_ (.CLK(clknet_leaf_40_csclk),
    .D(net613),
    .RESET_B(net486),
    .Q(\mgmt_gpio_data_buf[4] ));
 sky130_fd_sc_hd__dfrtp_1 _9181_ (.CLK(clknet_leaf_40_csclk),
    .D(_0454_),
    .RESET_B(net487),
    .Q(\mgmt_gpio_data_buf[5] ));
 sky130_fd_sc_hd__dfrtp_1 _9182_ (.CLK(clknet_leaf_4_csclk),
    .D(_0455_),
    .RESET_B(net420),
    .Q(\mgmt_gpio_data_buf[6] ));
 sky130_fd_sc_hd__dfrtp_1 _9183_ (.CLK(clknet_leaf_41_csclk),
    .D(_0456_),
    .RESET_B(net486),
    .Q(\mgmt_gpio_data_buf[7] ));
 sky130_fd_sc_hd__dfstp_2 _9184_ (.CLK(clknet_leaf_63_csclk),
    .D(_0457_),
    .SET_B(net443),
    .Q(\gpio_configure[0][0] ));
 sky130_fd_sc_hd__dfstp_1 _9185_ (.CLK(clknet_leaf_65_csclk),
    .D(_0458_),
    .SET_B(net433),
    .Q(\gpio_configure[0][1] ));
 sky130_fd_sc_hd__dfrtp_1 _9186_ (.CLK(clknet_leaf_73_csclk),
    .D(_0459_),
    .RESET_B(net456),
    .Q(\gpio_configure[0][2] ));
 sky130_fd_sc_hd__dfrtp_4 _9187_ (.CLK(clknet_leaf_50_csclk),
    .D(_0460_),
    .RESET_B(net456),
    .Q(\gpio_configure[0][3] ));
 sky130_fd_sc_hd__dfrtp_4 _9188_ (.CLK(clknet_leaf_71_csclk),
    .D(_0461_),
    .RESET_B(net450),
    .Q(\gpio_configure[0][4] ));
 sky130_fd_sc_hd__dfrtp_2 _9189_ (.CLK(clknet_leaf_81_csclk),
    .D(_0462_),
    .RESET_B(net416),
    .Q(\gpio_configure[0][5] ));
 sky130_fd_sc_hd__dfrtp_4 _9190_ (.CLK(clknet_leaf_75_csclk),
    .D(_0463_),
    .RESET_B(net425),
    .Q(\gpio_configure[0][6] ));
 sky130_fd_sc_hd__dfrtp_1 _9191_ (.CLK(clknet_leaf_81_csclk),
    .D(_0464_),
    .RESET_B(net416),
    .Q(\gpio_configure[0][7] ));
 sky130_fd_sc_hd__dfstp_1 _9192_ (.CLK(clknet_leaf_7_csclk),
    .D(_0465_),
    .SET_B(net422),
    .Q(\gpio_configure[1][0] ));
 sky130_fd_sc_hd__dfstp_1 _9193_ (.CLK(clknet_leaf_46_csclk),
    .D(_0466_),
    .SET_B(net467),
    .Q(\gpio_configure[1][1] ));
 sky130_fd_sc_hd__dfrtp_2 _9194_ (.CLK(clknet_leaf_73_csclk),
    .D(_0467_),
    .RESET_B(net456),
    .Q(\gpio_configure[1][2] ));
 sky130_fd_sc_hd__dfrtp_1 _9195_ (.CLK(clknet_leaf_46_csclk),
    .D(_0468_),
    .RESET_B(net467),
    .Q(\gpio_configure[1][3] ));
 sky130_fd_sc_hd__dfrtp_1 _9196_ (.CLK(clknet_leaf_21_csclk),
    .D(_0469_),
    .RESET_B(net461),
    .Q(\gpio_configure[1][4] ));
 sky130_fd_sc_hd__dfrtp_1 _9197_ (.CLK(clknet_leaf_12_csclk),
    .D(_0470_),
    .RESET_B(net458),
    .Q(\gpio_configure[1][5] ));
 sky130_fd_sc_hd__dfrtp_2 _9198_ (.CLK(clknet_leaf_0_csclk),
    .D(_0471_),
    .RESET_B(net409),
    .Q(\gpio_configure[1][6] ));
 sky130_fd_sc_hd__dfrtp_2 _9199_ (.CLK(clknet_leaf_0_csclk),
    .D(_0472_),
    .RESET_B(net409),
    .Q(\gpio_configure[1][7] ));
 sky130_fd_sc_hd__dfstp_1 _9200_ (.CLK(clknet_leaf_5_csclk),
    .D(_0473_),
    .SET_B(net422),
    .Q(\gpio_configure[2][0] ));
 sky130_fd_sc_hd__dfstp_1 _9201_ (.CLK(clknet_leaf_25_csclk),
    .D(_0474_),
    .SET_B(net473),
    .Q(\gpio_configure[2][1] ));
 sky130_fd_sc_hd__dfrtp_2 _9202_ (.CLK(clknet_leaf_18_csclk),
    .D(_0475_),
    .RESET_B(net463),
    .Q(\gpio_configure[2][2] ));
 sky130_fd_sc_hd__dfrtp_4 _9203_ (.CLK(clknet_leaf_71_csclk),
    .D(_0476_),
    .RESET_B(net434),
    .Q(\gpio_configure[2][3] ));
 sky130_fd_sc_hd__dfrtp_4 _9204_ (.CLK(clknet_leaf_74_csclk),
    .D(_0477_),
    .RESET_B(net425),
    .Q(\gpio_configure[2][4] ));
 sky130_fd_sc_hd__dfrtp_1 _9205_ (.CLK(clknet_leaf_5_csclk),
    .D(_0478_),
    .RESET_B(net423),
    .Q(\gpio_configure[2][5] ));
 sky130_fd_sc_hd__dfrtp_1 _9206_ (.CLK(clknet_leaf_0_csclk),
    .D(_0479_),
    .RESET_B(net409),
    .Q(\gpio_configure[2][6] ));
 sky130_fd_sc_hd__dfrtp_1 _9207_ (.CLK(clknet_leaf_0_csclk),
    .D(_0480_),
    .RESET_B(net419),
    .Q(\gpio_configure[2][7] ));
 sky130_fd_sc_hd__dfstp_1 _9208_ (.CLK(clknet_leaf_1_csclk),
    .D(_0481_),
    .SET_B(net418),
    .Q(\gpio_configure[3][0] ));
 sky130_fd_sc_hd__dfstp_1 _9209_ (.CLK(clknet_leaf_47_csclk),
    .D(_0482_),
    .SET_B(net467),
    .Q(\gpio_configure[3][1] ));
 sky130_fd_sc_hd__dfrtp_1 _9210_ (.CLK(clknet_3_4_0_csclk),
    .D(_0483_),
    .RESET_B(net467),
    .Q(\gpio_configure[3][2] ));
 sky130_fd_sc_hd__dfrtp_4 _9211_ (.CLK(clknet_leaf_48_csclk),
    .D(_0484_),
    .RESET_B(net467),
    .Q(\gpio_configure[3][3] ));
 sky130_fd_sc_hd__dfrtp_4 _9212_ (.CLK(clknet_leaf_85_csclk),
    .D(_0485_),
    .RESET_B(net408),
    .Q(\gpio_configure[3][4] ));
 sky130_fd_sc_hd__dfrtp_4 _9213_ (.CLK(clknet_leaf_0_csclk),
    .D(_0486_),
    .RESET_B(net419),
    .Q(\gpio_configure[3][5] ));
 sky130_fd_sc_hd__dfrtp_4 _9214_ (.CLK(clknet_leaf_85_csclk),
    .D(_0487_),
    .RESET_B(net408),
    .Q(\gpio_configure[3][6] ));
 sky130_fd_sc_hd__dfrtp_2 _9215_ (.CLK(clknet_leaf_86_csclk),
    .D(_0488_),
    .RESET_B(net409),
    .Q(\gpio_configure[3][7] ));
 sky130_fd_sc_hd__dfstp_2 _9216_ (.CLK(clknet_leaf_86_csclk),
    .D(_0489_),
    .SET_B(net409),
    .Q(\gpio_configure[4][0] ));
 sky130_fd_sc_hd__dfstp_2 _9217_ (.CLK(clknet_leaf_49_csclk),
    .D(_0490_),
    .SET_B(net456),
    .Q(\gpio_configure[4][1] ));
 sky130_fd_sc_hd__dfrtp_4 _9218_ (.CLK(clknet_leaf_68_csclk),
    .D(_0491_),
    .RESET_B(net429),
    .Q(\gpio_configure[4][2] ));
 sky130_fd_sc_hd__dfrtp_4 _9219_ (.CLK(clknet_leaf_47_csclk),
    .D(_0492_),
    .RESET_B(net469),
    .Q(\gpio_configure[4][3] ));
 sky130_fd_sc_hd__dfrtp_4 _9220_ (.CLK(clknet_leaf_77_csclk),
    .D(_0493_),
    .RESET_B(net415),
    .Q(\gpio_configure[4][4] ));
 sky130_fd_sc_hd__dfrtp_4 _9221_ (.CLK(clknet_leaf_82_csclk),
    .D(_0494_),
    .RESET_B(net406),
    .Q(\gpio_configure[4][5] ));
 sky130_fd_sc_hd__dfrtp_2 _9222_ (.CLK(clknet_leaf_82_csclk),
    .D(_0495_),
    .RESET_B(net409),
    .Q(\gpio_configure[4][6] ));
 sky130_fd_sc_hd__dfrtp_2 _9223_ (.CLK(clknet_leaf_83_csclk),
    .D(_0496_),
    .RESET_B(net406),
    .Q(\gpio_configure[4][7] ));
 sky130_fd_sc_hd__dfstp_1 _9224_ (.CLK(clknet_leaf_7_csclk),
    .D(_0497_),
    .SET_B(net419),
    .Q(\gpio_configure[5][0] ));
 sky130_fd_sc_hd__dfstp_1 _9225_ (.CLK(clknet_leaf_26_csclk),
    .D(_0498_),
    .SET_B(net471),
    .Q(\gpio_configure[5][1] ));
 sky130_fd_sc_hd__dfrtp_4 _9226_ (.CLK(clknet_leaf_27_csclk),
    .D(_0499_),
    .RESET_B(net472),
    .Q(\gpio_configure[5][2] ));
 sky130_fd_sc_hd__dfrtp_4 _9227_ (.CLK(clknet_leaf_48_csclk),
    .D(_0500_),
    .RESET_B(net467),
    .Q(\gpio_configure[5][3] ));
 sky130_fd_sc_hd__dfrtp_4 _9228_ (.CLK(clknet_leaf_77_csclk),
    .D(_0501_),
    .RESET_B(net415),
    .Q(\gpio_configure[5][4] ));
 sky130_fd_sc_hd__dfrtp_1 _9229_ (.CLK(clknet_leaf_12_csclk),
    .D(_0502_),
    .RESET_B(net458),
    .Q(\gpio_configure[5][5] ));
 sky130_fd_sc_hd__dfrtp_1 _9230_ (.CLK(clknet_leaf_0_csclk),
    .D(_0503_),
    .RESET_B(net419),
    .Q(\gpio_configure[5][6] ));
 sky130_fd_sc_hd__dfrtp_1 _9231_ (.CLK(clknet_leaf_0_csclk),
    .D(_0504_),
    .RESET_B(net419),
    .Q(\gpio_configure[5][7] ));
 sky130_fd_sc_hd__dfstp_2 _9232_ (.CLK(clknet_leaf_0_csclk),
    .D(_0505_),
    .SET_B(net419),
    .Q(\gpio_configure[6][0] ));
 sky130_fd_sc_hd__dfstp_2 _9233_ (.CLK(clknet_leaf_25_csclk),
    .D(_0506_),
    .SET_B(net473),
    .Q(\gpio_configure[6][1] ));
 sky130_fd_sc_hd__dfrtp_4 _9234_ (.CLK(clknet_leaf_27_csclk),
    .D(_0507_),
    .RESET_B(net471),
    .Q(\gpio_configure[6][2] ));
 sky130_fd_sc_hd__dfrtp_4 _9235_ (.CLK(clknet_leaf_34_csclk),
    .D(_0508_),
    .RESET_B(net484),
    .Q(\gpio_configure[6][3] ));
 sky130_fd_sc_hd__dfrtp_4 _9236_ (.CLK(clknet_leaf_18_csclk),
    .D(_0509_),
    .RESET_B(net463),
    .Q(\gpio_configure[6][4] ));
 sky130_fd_sc_hd__dfrtp_1 _9237_ (.CLK(clknet_leaf_11_csclk),
    .D(_0510_),
    .RESET_B(net460),
    .Q(\gpio_configure[6][5] ));
 sky130_fd_sc_hd__dfrtp_1 _9238_ (.CLK(clknet_leaf_7_csclk),
    .D(_0511_),
    .RESET_B(net419),
    .Q(\gpio_configure[6][6] ));
 sky130_fd_sc_hd__dfrtp_1 _9239_ (.CLK(clknet_leaf_1_csclk),
    .D(_0512_),
    .RESET_B(net419),
    .Q(\gpio_configure[6][7] ));
 sky130_fd_sc_hd__dfstp_2 _9240_ (.CLK(clknet_leaf_5_csclk),
    .D(_0513_),
    .SET_B(net420),
    .Q(\gpio_configure[7][0] ));
 sky130_fd_sc_hd__dfstp_1 _9241_ (.CLK(clknet_leaf_49_csclk),
    .D(_0514_),
    .SET_B(net467),
    .Q(\gpio_configure[7][1] ));
 sky130_fd_sc_hd__dfrtp_4 _9242_ (.CLK(clknet_leaf_68_csclk),
    .D(_0515_),
    .RESET_B(net429),
    .Q(\gpio_configure[7][2] ));
 sky130_fd_sc_hd__dfrtp_4 _9243_ (.CLK(clknet_leaf_43_csclk),
    .D(_0516_),
    .RESET_B(net469),
    .Q(\gpio_configure[7][3] ));
 sky130_fd_sc_hd__dfrtp_2 _9244_ (.CLK(clknet_leaf_13_csclk),
    .D(_0517_),
    .RESET_B(net459),
    .Q(\gpio_configure[7][4] ));
 sky130_fd_sc_hd__dfrtp_4 _9245_ (.CLK(clknet_leaf_82_csclk),
    .D(_0518_),
    .RESET_B(net406),
    .Q(\gpio_configure[7][5] ));
 sky130_fd_sc_hd__dfrtp_1 _9246_ (.CLK(clknet_leaf_0_csclk),
    .D(_0519_),
    .RESET_B(net419),
    .Q(\gpio_configure[7][6] ));
 sky130_fd_sc_hd__dfrtp_2 _9247_ (.CLK(clknet_leaf_1_csclk),
    .D(_0520_),
    .RESET_B(net418),
    .Q(\gpio_configure[7][7] ));
 sky130_fd_sc_hd__dfstp_2 _9248_ (.CLK(clknet_leaf_78_csclk),
    .D(_0521_),
    .SET_B(net415),
    .Q(\gpio_configure[8][0] ));
 sky130_fd_sc_hd__dfstp_2 _9249_ (.CLK(clknet_leaf_33_csclk),
    .D(_0522_),
    .SET_B(net474),
    .Q(\gpio_configure[8][1] ));
 sky130_fd_sc_hd__dfrtp_1 _9250_ (.CLK(clknet_leaf_23_csclk),
    .D(_0523_),
    .RESET_B(net467),
    .Q(\gpio_configure[8][2] ));
 sky130_fd_sc_hd__dfrtp_4 _9251_ (.CLK(clknet_leaf_41_csclk),
    .D(_0524_),
    .RESET_B(net485),
    .Q(\gpio_configure[8][3] ));
 sky130_fd_sc_hd__dfrtp_1 _9252_ (.CLK(clknet_leaf_17_csclk),
    .D(_0525_),
    .RESET_B(net463),
    .Q(\gpio_configure[8][4] ));
 sky130_fd_sc_hd__dfrtp_4 _9253_ (.CLK(clknet_leaf_80_csclk),
    .D(_0526_),
    .RESET_B(net411),
    .Q(\gpio_configure[8][5] ));
 sky130_fd_sc_hd__dfrtp_4 _9254_ (.CLK(clknet_leaf_80_csclk),
    .D(_0527_),
    .RESET_B(net411),
    .Q(\gpio_configure[8][6] ));
 sky130_fd_sc_hd__dfrtp_2 _9255_ (.CLK(clknet_leaf_81_csclk),
    .D(_0528_),
    .RESET_B(net416),
    .Q(\gpio_configure[8][7] ));
 sky130_fd_sc_hd__dfstp_2 _9256_ (.CLK(clknet_leaf_18_csclk),
    .D(_0529_),
    .SET_B(net463),
    .Q(\gpio_configure[9][0] ));
 sky130_fd_sc_hd__dfstp_2 _9257_ (.CLK(clknet_leaf_25_csclk),
    .D(_0530_),
    .SET_B(net473),
    .Q(\gpio_configure[9][1] ));
 sky130_fd_sc_hd__dfrtp_1 _9258_ (.CLK(clknet_leaf_27_csclk),
    .D(_0531_),
    .RESET_B(net471),
    .Q(\gpio_configure[9][2] ));
 sky130_fd_sc_hd__dfrtp_4 _9259_ (.CLK(clknet_leaf_25_csclk),
    .D(_0532_),
    .RESET_B(net473),
    .Q(\gpio_configure[9][3] ));
 sky130_fd_sc_hd__dfrtp_1 _9260_ (.CLK(clknet_leaf_18_csclk),
    .D(_0533_),
    .RESET_B(net463),
    .Q(\gpio_configure[9][4] ));
 sky130_fd_sc_hd__dfrtp_4 _9261_ (.CLK(clknet_leaf_19_csclk),
    .D(_0534_),
    .RESET_B(net460),
    .Q(\gpio_configure[9][5] ));
 sky130_fd_sc_hd__dfrtp_4 _9262_ (.CLK(clknet_leaf_19_csclk),
    .D(_0535_),
    .RESET_B(net460),
    .Q(\gpio_configure[9][6] ));
 sky130_fd_sc_hd__dfrtp_4 _9263_ (.CLK(clknet_leaf_19_csclk),
    .D(_0536_),
    .RESET_B(net464),
    .Q(\gpio_configure[9][7] ));
 sky130_fd_sc_hd__dfstp_1 _9264_ (.CLK(clknet_leaf_20_csclk),
    .D(_0537_),
    .SET_B(net462),
    .Q(\gpio_configure[10][0] ));
 sky130_fd_sc_hd__dfstp_2 _9265_ (.CLK(clknet_leaf_25_csclk),
    .D(_0538_),
    .SET_B(net473),
    .Q(\gpio_configure[10][1] ));
 sky130_fd_sc_hd__dfrtp_1 _9266_ (.CLK(clknet_leaf_27_csclk),
    .D(_0539_),
    .RESET_B(net472),
    .Q(\gpio_configure[10][2] ));
 sky130_fd_sc_hd__dfrtp_4 _9267_ (.CLK(clknet_leaf_34_csclk),
    .D(_0540_),
    .RESET_B(net484),
    .Q(\gpio_configure[10][3] ));
 sky130_fd_sc_hd__dfrtp_4 _9268_ (.CLK(clknet_leaf_17_csclk),
    .D(_0541_),
    .RESET_B(net463),
    .Q(\gpio_configure[10][4] ));
 sky130_fd_sc_hd__dfrtp_1 _9269_ (.CLK(clknet_leaf_11_csclk),
    .D(_0542_),
    .RESET_B(net460),
    .Q(\gpio_configure[10][5] ));
 sky130_fd_sc_hd__dfrtp_4 _9270_ (.CLK(clknet_leaf_11_csclk),
    .D(_0543_),
    .RESET_B(net460),
    .Q(\gpio_configure[10][6] ));
 sky130_fd_sc_hd__dfrtp_2 _9271_ (.CLK(clknet_leaf_11_csclk),
    .D(_0544_),
    .RESET_B(net460),
    .Q(\gpio_configure[10][7] ));
 sky130_fd_sc_hd__dfstp_2 _9272_ (.CLK(clknet_leaf_7_csclk),
    .D(_0545_),
    .SET_B(net421),
    .Q(\gpio_configure[11][0] ));
 sky130_fd_sc_hd__dfstp_1 _9273_ (.CLK(clknet_leaf_24_csclk),
    .D(_0546_),
    .SET_B(net467),
    .Q(\gpio_configure[11][1] ));
 sky130_fd_sc_hd__dfrtp_1 _9274_ (.CLK(clknet_leaf_23_csclk),
    .D(_0547_),
    .RESET_B(net468),
    .Q(\gpio_configure[11][2] ));
 sky130_fd_sc_hd__dfrtp_4 _9275_ (.CLK(clknet_leaf_45_csclk),
    .D(_0548_),
    .RESET_B(net468),
    .Q(\gpio_configure[11][3] ));
 sky130_fd_sc_hd__dfrtp_4 _9276_ (.CLK(clknet_leaf_21_csclk),
    .D(_0549_),
    .RESET_B(net462),
    .Q(\gpio_configure[11][4] ));
 sky130_fd_sc_hd__dfrtp_1 _9277_ (.CLK(clknet_leaf_13_csclk),
    .D(_0550_),
    .RESET_B(net458),
    .Q(\gpio_configure[11][5] ));
 sky130_fd_sc_hd__dfrtp_2 _9278_ (.CLK(clknet_leaf_1_csclk),
    .D(_0551_),
    .RESET_B(net426),
    .Q(\gpio_configure[11][6] ));
 sky130_fd_sc_hd__dfrtp_2 _9279_ (.CLK(clknet_leaf_3_csclk),
    .D(_0552_),
    .RESET_B(net417),
    .Q(\gpio_configure[11][7] ));
 sky130_fd_sc_hd__dfstp_1 _9280_ (.CLK(clknet_leaf_18_csclk),
    .D(_0553_),
    .SET_B(net463),
    .Q(\gpio_configure[12][0] ));
 sky130_fd_sc_hd__dfstp_2 _9281_ (.CLK(clknet_leaf_25_csclk),
    .D(_0554_),
    .SET_B(net474),
    .Q(\gpio_configure[12][1] ));
 sky130_fd_sc_hd__dfrtp_1 _9282_ (.CLK(clknet_leaf_27_csclk),
    .D(_0555_),
    .RESET_B(net472),
    .Q(\gpio_configure[12][2] ));
 sky130_fd_sc_hd__dfrtp_4 _9283_ (.CLK(clknet_leaf_34_csclk),
    .D(_0556_),
    .RESET_B(net473),
    .Q(\gpio_configure[12][3] ));
 sky130_fd_sc_hd__dfrtp_1 _9284_ (.CLK(clknet_leaf_18_csclk),
    .D(_0557_),
    .RESET_B(net463),
    .Q(\gpio_configure[12][4] ));
 sky130_fd_sc_hd__dfrtp_1 _9285_ (.CLK(clknet_leaf_19_csclk),
    .D(_0558_),
    .RESET_B(net464),
    .Q(\gpio_configure[12][5] ));
 sky130_fd_sc_hd__dfrtp_4 _9286_ (.CLK(clknet_leaf_19_csclk),
    .D(_0559_),
    .RESET_B(net464),
    .Q(\gpio_configure[12][6] ));
 sky130_fd_sc_hd__dfrtp_1 _9287_ (.CLK(clknet_leaf_19_csclk),
    .D(_0560_),
    .RESET_B(net464),
    .Q(\gpio_configure[12][7] ));
 sky130_fd_sc_hd__dfstp_1 _9288_ (.CLK(clknet_leaf_75_csclk),
    .D(_0561_),
    .SET_B(net425),
    .Q(\gpio_configure[13][0] ));
 sky130_fd_sc_hd__dfstp_1 _9289_ (.CLK(clknet_leaf_24_csclk),
    .D(_0562_),
    .SET_B(net468),
    .Q(\gpio_configure[13][1] ));
 sky130_fd_sc_hd__dfrtp_1 _9290_ (.CLK(clknet_leaf_23_csclk),
    .D(_0563_),
    .RESET_B(net468),
    .Q(\gpio_configure[13][2] ));
 sky130_fd_sc_hd__dfrtp_4 _9291_ (.CLK(clknet_leaf_45_csclk),
    .D(_0564_),
    .RESET_B(net468),
    .Q(\gpio_configure[13][3] ));
 sky130_fd_sc_hd__dfrtp_2 _9292_ (.CLK(clknet_leaf_20_csclk),
    .D(_0565_),
    .RESET_B(net462),
    .Q(\gpio_configure[13][4] ));
 sky130_fd_sc_hd__dfrtp_1 _9293_ (.CLK(clknet_leaf_13_csclk),
    .D(_0566_),
    .RESET_B(net458),
    .Q(\gpio_configure[13][5] ));
 sky130_fd_sc_hd__dfrtp_4 _9294_ (.CLK(clknet_leaf_5_csclk),
    .D(_0567_),
    .RESET_B(net422),
    .Q(\gpio_configure[13][6] ));
 sky130_fd_sc_hd__dfrtp_2 _9295_ (.CLK(clknet_leaf_1_csclk),
    .D(_0568_),
    .RESET_B(net417),
    .Q(\gpio_configure[13][7] ));
 sky130_fd_sc_hd__dfstp_2 _9296_ (.CLK(clknet_leaf_18_csclk),
    .D(_0569_),
    .SET_B(net463),
    .Q(\gpio_configure[14][0] ));
 sky130_fd_sc_hd__dfstp_2 _9297_ (.CLK(clknet_leaf_32_csclk),
    .D(_0570_),
    .SET_B(net479),
    .Q(\gpio_configure[14][1] ));
 sky130_fd_sc_hd__dfrtp_4 _9298_ (.CLK(clknet_leaf_28_csclk),
    .D(_0571_),
    .RESET_B(net475),
    .Q(\gpio_configure[14][2] ));
 sky130_fd_sc_hd__dfrtp_4 _9299_ (.CLK(clknet_leaf_32_csclk),
    .D(_0572_),
    .RESET_B(net479),
    .Q(\gpio_configure[14][3] ));
 sky130_fd_sc_hd__dfrtp_2 _9300_ (.CLK(clknet_leaf_17_csclk),
    .D(_0573_),
    .RESET_B(net465),
    .Q(\gpio_configure[14][4] ));
 sky130_fd_sc_hd__dfrtp_1 _9301_ (.CLK(clknet_leaf_19_csclk),
    .D(_0574_),
    .RESET_B(net460),
    .Q(\gpio_configure[14][5] ));
 sky130_fd_sc_hd__dfrtp_4 _9302_ (.CLK(clknet_leaf_19_csclk),
    .D(_0575_),
    .RESET_B(net464),
    .Q(\gpio_configure[14][6] ));
 sky130_fd_sc_hd__dfrtp_4 _9303_ (.CLK(clknet_3_5_0_csclk),
    .D(_0576_),
    .RESET_B(net464),
    .Q(\gpio_configure[14][7] ));
 sky130_fd_sc_hd__dfstp_2 _9304_ (.CLK(clknet_leaf_4_csclk),
    .D(_0577_),
    .SET_B(net420),
    .Q(\gpio_configure[15][0] ));
 sky130_fd_sc_hd__dfstp_2 _9305_ (.CLK(clknet_leaf_24_csclk),
    .D(_0578_),
    .SET_B(net468),
    .Q(\gpio_configure[15][1] ));
 sky130_fd_sc_hd__dfrtp_4 _9306_ (.CLK(clknet_leaf_29_csclk),
    .D(_0579_),
    .RESET_B(net475),
    .Q(\gpio_configure[15][2] ));
 sky130_fd_sc_hd__dfrtp_4 _9307_ (.CLK(clknet_leaf_32_csclk),
    .D(_0580_),
    .RESET_B(net489),
    .Q(\gpio_configure[15][3] ));
 sky130_fd_sc_hd__dfrtp_4 _9308_ (.CLK(clknet_leaf_17_csclk),
    .D(_0581_),
    .RESET_B(net465),
    .Q(\gpio_configure[15][4] ));
 sky130_fd_sc_hd__dfrtp_1 _9309_ (.CLK(clknet_leaf_12_csclk),
    .D(_0582_),
    .RESET_B(net458),
    .Q(\gpio_configure[15][5] ));
 sky130_fd_sc_hd__dfrtp_2 _9310_ (.CLK(clknet_leaf_1_csclk),
    .D(_0583_),
    .RESET_B(net419),
    .Q(\gpio_configure[15][6] ));
 sky130_fd_sc_hd__dfrtp_2 _9311_ (.CLK(clknet_leaf_1_csclk),
    .D(_0584_),
    .RESET_B(net417),
    .Q(\gpio_configure[15][7] ));
 sky130_fd_sc_hd__dfstp_1 _9312_ (.CLK(clknet_leaf_9_csclk),
    .D(_0585_),
    .SET_B(net461),
    .Q(\gpio_configure[16][0] ));
 sky130_fd_sc_hd__dfstp_2 _9313_ (.CLK(clknet_leaf_33_csclk),
    .D(_0586_),
    .SET_B(net474),
    .Q(\gpio_configure[16][1] ));
 sky130_fd_sc_hd__dfrtp_4 _9314_ (.CLK(clknet_leaf_77_csclk),
    .D(_0587_),
    .RESET_B(net429),
    .Q(\gpio_configure[16][2] ));
 sky130_fd_sc_hd__dfrtp_4 _9315_ (.CLK(clknet_leaf_26_csclk),
    .D(_0588_),
    .RESET_B(net474),
    .Q(\gpio_configure[16][3] ));
 sky130_fd_sc_hd__dfrtp_2 _9316_ (.CLK(clknet_leaf_17_csclk),
    .D(_0589_),
    .RESET_B(net464),
    .Q(\gpio_configure[16][4] ));
 sky130_fd_sc_hd__dfrtp_4 _9317_ (.CLK(clknet_leaf_79_csclk),
    .D(_0590_),
    .RESET_B(net413),
    .Q(\gpio_configure[16][5] ));
 sky130_fd_sc_hd__dfrtp_4 _9318_ (.CLK(clknet_leaf_81_csclk),
    .D(_0591_),
    .RESET_B(net413),
    .Q(\gpio_configure[16][6] ));
 sky130_fd_sc_hd__dfrtp_1 _9319_ (.CLK(clknet_leaf_76_csclk),
    .D(_0592_),
    .RESET_B(net425),
    .Q(\gpio_configure[16][7] ));
 sky130_fd_sc_hd__dfstp_2 _9320_ (.CLK(clknet_leaf_18_csclk),
    .D(_0593_),
    .SET_B(net464),
    .Q(\gpio_configure[17][0] ));
 sky130_fd_sc_hd__dfstp_1 _9321_ (.CLK(clknet_leaf_32_csclk),
    .D(_0594_),
    .SET_B(net479),
    .Q(\gpio_configure[17][1] ));
 sky130_fd_sc_hd__dfrtp_4 _9322_ (.CLK(clknet_leaf_29_csclk),
    .D(_0595_),
    .RESET_B(net475),
    .Q(\gpio_configure[17][2] ));
 sky130_fd_sc_hd__dfrtp_4 _9323_ (.CLK(clknet_leaf_32_csclk),
    .D(_0596_),
    .RESET_B(net489),
    .Q(\gpio_configure[17][3] ));
 sky130_fd_sc_hd__dfrtp_4 _9324_ (.CLK(clknet_leaf_17_csclk),
    .D(_0597_),
    .RESET_B(net465),
    .Q(\gpio_configure[17][4] ));
 sky130_fd_sc_hd__dfrtp_1 _9325_ (.CLK(clknet_leaf_19_csclk),
    .D(_0598_),
    .RESET_B(net460),
    .Q(\gpio_configure[17][5] ));
 sky130_fd_sc_hd__dfrtp_4 _9326_ (.CLK(clknet_leaf_6_csclk),
    .D(_0599_),
    .RESET_B(net423),
    .Q(\gpio_configure[17][6] ));
 sky130_fd_sc_hd__dfrtp_4 _9327_ (.CLK(clknet_leaf_6_csclk),
    .D(_0600_),
    .RESET_B(net423),
    .Q(\gpio_configure[17][7] ));
 sky130_fd_sc_hd__dfstp_2 _9328_ (.CLK(clknet_leaf_18_csclk),
    .D(_0601_),
    .SET_B(net463),
    .Q(\gpio_configure[18][0] ));
 sky130_fd_sc_hd__dfstp_1 _9329_ (.CLK(clknet_leaf_32_csclk),
    .D(_0602_),
    .SET_B(net479),
    .Q(\gpio_configure[18][1] ));
 sky130_fd_sc_hd__dfrtp_4 _9330_ (.CLK(clknet_leaf_29_csclk),
    .D(_0603_),
    .RESET_B(net477),
    .Q(\gpio_configure[18][2] ));
 sky130_fd_sc_hd__dfrtp_4 _9331_ (.CLK(clknet_leaf_36_csclk),
    .D(_0604_),
    .RESET_B(net491),
    .Q(\gpio_configure[18][3] ));
 sky130_fd_sc_hd__dfrtp_4 _9332_ (.CLK(clknet_leaf_16_csclk),
    .D(_0605_),
    .RESET_B(net466),
    .Q(\gpio_configure[18][4] ));
 sky130_fd_sc_hd__dfrtp_1 _9333_ (.CLK(clknet_leaf_20_csclk),
    .D(_0606_),
    .RESET_B(net460),
    .Q(\gpio_configure[18][5] ));
 sky130_fd_sc_hd__dfrtp_1 _9334_ (.CLK(clknet_leaf_6_csclk),
    .D(_0607_),
    .RESET_B(net423),
    .Q(\gpio_configure[18][6] ));
 sky130_fd_sc_hd__dfrtp_1 _9335_ (.CLK(clknet_leaf_6_csclk),
    .D(_0608_),
    .RESET_B(net422),
    .Q(\gpio_configure[18][7] ));
 sky130_fd_sc_hd__dfstp_2 _9336_ (.CLK(clknet_leaf_1_csclk),
    .D(_0609_),
    .SET_B(net417),
    .Q(\gpio_configure[19][0] ));
 sky130_fd_sc_hd__dfstp_2 _9337_ (.CLK(clknet_leaf_25_csclk),
    .D(_0610_),
    .SET_B(net473),
    .Q(\gpio_configure[19][1] ));
 sky130_fd_sc_hd__dfrtp_4 _9338_ (.CLK(clknet_leaf_29_csclk),
    .D(_0611_),
    .RESET_B(net478),
    .Q(\gpio_configure[19][2] ));
 sky130_fd_sc_hd__dfrtp_4 _9339_ (.CLK(clknet_leaf_31_csclk),
    .D(_0612_),
    .RESET_B(net481),
    .Q(\gpio_configure[19][3] ));
 sky130_fd_sc_hd__dfrtp_4 _9340_ (.CLK(clknet_leaf_16_csclk),
    .D(_0613_),
    .RESET_B(net466),
    .Q(\gpio_configure[19][4] ));
 sky130_fd_sc_hd__dfrtp_2 _9341_ (.CLK(clknet_leaf_12_csclk),
    .D(_0614_),
    .RESET_B(net458),
    .Q(\gpio_configure[19][5] ));
 sky130_fd_sc_hd__dfrtp_2 _9342_ (.CLK(clknet_leaf_1_csclk),
    .D(_0615_),
    .RESET_B(net417),
    .Q(\gpio_configure[19][6] ));
 sky130_fd_sc_hd__dfrtp_2 _9343_ (.CLK(clknet_leaf_3_csclk),
    .D(_0616_),
    .RESET_B(net418),
    .Q(\gpio_configure[19][7] ));
 sky130_fd_sc_hd__dfstp_1 _9344_ (.CLK(clknet_leaf_9_csclk),
    .D(_0617_),
    .SET_B(net425),
    .Q(\gpio_configure[20][0] ));
 sky130_fd_sc_hd__dfstp_2 _9345_ (.CLK(clknet_leaf_33_csclk),
    .D(_0618_),
    .SET_B(net479),
    .Q(\gpio_configure[20][1] ));
 sky130_fd_sc_hd__dfrtp_4 _9346_ (.CLK(clknet_leaf_29_csclk),
    .D(_0619_),
    .RESET_B(net477),
    .Q(\gpio_configure[20][2] ));
 sky130_fd_sc_hd__dfrtp_4 _9347_ (.CLK(clknet_leaf_30_csclk),
    .D(_0620_),
    .RESET_B(net478),
    .Q(\gpio_configure[20][3] ));
 sky130_fd_sc_hd__dfrtp_4 _9348_ (.CLK(clknet_leaf_29_csclk),
    .D(_0621_),
    .RESET_B(net466),
    .Q(\gpio_configure[20][4] ));
 sky130_fd_sc_hd__dfrtp_1 _9349_ (.CLK(clknet_leaf_11_csclk),
    .D(_0622_),
    .RESET_B(net461),
    .Q(\gpio_configure[20][5] ));
 sky130_fd_sc_hd__dfrtp_4 _9350_ (.CLK(clknet_leaf_5_csclk),
    .D(_0623_),
    .RESET_B(net422),
    .Q(\gpio_configure[20][6] ));
 sky130_fd_sc_hd__dfrtp_1 _9351_ (.CLK(clknet_leaf_5_csclk),
    .D(_0624_),
    .RESET_B(net422),
    .Q(\gpio_configure[20][7] ));
 sky130_fd_sc_hd__dfstp_2 _9352_ (.CLK(clknet_leaf_9_csclk),
    .D(_0625_),
    .SET_B(net425),
    .Q(\gpio_configure[21][0] ));
 sky130_fd_sc_hd__dfstp_4 _9353_ (.CLK(clknet_leaf_30_csclk),
    .D(_0626_),
    .SET_B(net479),
    .Q(\gpio_configure[21][1] ));
 sky130_fd_sc_hd__dfrtp_4 _9354_ (.CLK(clknet_leaf_29_csclk),
    .D(_0627_),
    .RESET_B(net477),
    .Q(\gpio_configure[21][2] ));
 sky130_fd_sc_hd__dfrtp_4 _9355_ (.CLK(clknet_leaf_31_csclk),
    .D(_0628_),
    .RESET_B(net478),
    .Q(\gpio_configure[21][3] ));
 sky130_fd_sc_hd__dfrtp_4 _9356_ (.CLK(clknet_leaf_16_csclk),
    .D(_0629_),
    .RESET_B(net466),
    .Q(\gpio_configure[21][4] ));
 sky130_fd_sc_hd__dfrtp_1 _9357_ (.CLK(clknet_leaf_11_csclk),
    .D(_0630_),
    .RESET_B(net460),
    .Q(\gpio_configure[21][5] ));
 sky130_fd_sc_hd__dfrtp_2 _9358_ (.CLK(clknet_leaf_6_csclk),
    .D(_0631_),
    .RESET_B(net422),
    .Q(\gpio_configure[21][6] ));
 sky130_fd_sc_hd__dfrtp_1 _9359_ (.CLK(clknet_3_1_0_csclk),
    .D(_0632_),
    .RESET_B(net422),
    .Q(\gpio_configure[21][7] ));
 sky130_fd_sc_hd__dfstp_1 _9360_ (.CLK(clknet_leaf_9_csclk),
    .D(_0633_),
    .SET_B(net425),
    .Q(\gpio_configure[22][0] ));
 sky130_fd_sc_hd__dfstp_2 _9361_ (.CLK(clknet_leaf_31_csclk),
    .D(_0634_),
    .SET_B(net479),
    .Q(\gpio_configure[22][1] ));
 sky130_fd_sc_hd__dfrtp_4 _9362_ (.CLK(clknet_leaf_29_csclk),
    .D(_0635_),
    .RESET_B(net477),
    .Q(\gpio_configure[22][2] ));
 sky130_fd_sc_hd__dfrtp_4 _9363_ (.CLK(clknet_leaf_30_csclk),
    .D(_0636_),
    .RESET_B(net481),
    .Q(\gpio_configure[22][3] ));
 sky130_fd_sc_hd__dfrtp_4 _9364_ (.CLK(clknet_leaf_16_csclk),
    .D(_0637_),
    .RESET_B(net466),
    .Q(\gpio_configure[22][4] ));
 sky130_fd_sc_hd__dfrtp_4 _9365_ (.CLK(clknet_leaf_10_csclk),
    .D(_0638_),
    .RESET_B(net461),
    .Q(\gpio_configure[22][5] ));
 sky130_fd_sc_hd__dfrtp_2 _9366_ (.CLK(clknet_leaf_6_csclk),
    .D(_0639_),
    .RESET_B(net422),
    .Q(\gpio_configure[22][6] ));
 sky130_fd_sc_hd__dfrtp_2 _9367_ (.CLK(clknet_leaf_6_csclk),
    .D(_0640_),
    .RESET_B(net422),
    .Q(\gpio_configure[22][7] ));
 sky130_fd_sc_hd__dfstp_2 _9368_ (.CLK(clknet_leaf_9_csclk),
    .D(_0641_),
    .SET_B(net425),
    .Q(\gpio_configure[23][0] ));
 sky130_fd_sc_hd__dfstp_2 _9369_ (.CLK(clknet_leaf_31_csclk),
    .D(_0642_),
    .SET_B(net481),
    .Q(\gpio_configure[23][1] ));
 sky130_fd_sc_hd__dfrtp_2 _9370_ (.CLK(clknet_leaf_29_csclk),
    .D(_0643_),
    .RESET_B(net477),
    .Q(\gpio_configure[23][2] ));
 sky130_fd_sc_hd__dfrtp_4 _9371_ (.CLK(clknet_leaf_31_csclk),
    .D(_0644_),
    .RESET_B(net481),
    .Q(\gpio_configure[23][3] ));
 sky130_fd_sc_hd__dfrtp_4 _9372_ (.CLK(clknet_leaf_16_csclk),
    .D(_0645_),
    .RESET_B(net465),
    .Q(\gpio_configure[23][4] ));
 sky130_fd_sc_hd__dfrtp_4 _9373_ (.CLK(clknet_leaf_12_csclk),
    .D(_0646_),
    .RESET_B(net458),
    .Q(\gpio_configure[23][5] ));
 sky130_fd_sc_hd__dfrtp_4 _9374_ (.CLK(clknet_leaf_5_csclk),
    .D(_0647_),
    .RESET_B(net423),
    .Q(\gpio_configure[23][6] ));
 sky130_fd_sc_hd__dfrtp_2 _9375_ (.CLK(clknet_leaf_5_csclk),
    .D(_0648_),
    .RESET_B(net423),
    .Q(\gpio_configure[23][7] ));
 sky130_fd_sc_hd__dfstp_1 _9376_ (.CLK(clknet_leaf_76_csclk),
    .D(_0649_),
    .SET_B(net416),
    .Q(\gpio_configure[24][0] ));
 sky130_fd_sc_hd__dfstp_1 _9377_ (.CLK(clknet_leaf_25_csclk),
    .D(_0650_),
    .SET_B(net473),
    .Q(\gpio_configure[24][1] ));
 sky130_fd_sc_hd__dfrtp_2 _9378_ (.CLK(clknet_leaf_27_csclk),
    .D(_0651_),
    .RESET_B(net471),
    .Q(\gpio_configure[24][2] ));
 sky130_fd_sc_hd__dfrtp_4 _9379_ (.CLK(clknet_leaf_32_csclk),
    .D(_0652_),
    .RESET_B(net480),
    .Q(\gpio_configure[24][3] ));
 sky130_fd_sc_hd__dfrtp_2 _9380_ (.CLK(clknet_leaf_17_csclk),
    .D(_0653_),
    .RESET_B(net464),
    .Q(\gpio_configure[24][4] ));
 sky130_fd_sc_hd__dfrtp_1 _9381_ (.CLK(clknet_leaf_11_csclk),
    .D(_0654_),
    .RESET_B(net461),
    .Q(\gpio_configure[24][5] ));
 sky130_fd_sc_hd__dfrtp_4 _9382_ (.CLK(clknet_leaf_86_csclk),
    .D(_0655_),
    .RESET_B(net409),
    .Q(\gpio_configure[24][6] ));
 sky130_fd_sc_hd__dfrtp_2 _9383_ (.CLK(clknet_leaf_86_csclk),
    .D(_0656_),
    .RESET_B(net409),
    .Q(\gpio_configure[24][7] ));
 sky130_fd_sc_hd__dfstp_2 _9384_ (.CLK(clknet_leaf_3_csclk),
    .D(_0657_),
    .SET_B(net417),
    .Q(\gpio_configure[25][0] ));
 sky130_fd_sc_hd__dfstp_2 _9385_ (.CLK(clknet_leaf_30_csclk),
    .D(_0658_),
    .SET_B(net479),
    .Q(\gpio_configure[25][1] ));
 sky130_fd_sc_hd__dfrtp_4 _9386_ (.CLK(clknet_leaf_28_csclk),
    .D(_0659_),
    .RESET_B(net476),
    .Q(\gpio_configure[25][2] ));
 sky130_fd_sc_hd__dfrtp_4 _9387_ (.CLK(clknet_leaf_31_csclk),
    .D(_0660_),
    .RESET_B(net482),
    .Q(\gpio_configure[25][3] ));
 sky130_fd_sc_hd__dfrtp_4 _9388_ (.CLK(clknet_leaf_16_csclk),
    .D(_0661_),
    .RESET_B(net466),
    .Q(\gpio_configure[25][4] ));
 sky130_fd_sc_hd__dfrtp_4 _9389_ (.CLK(clknet_leaf_12_csclk),
    .D(_0662_),
    .RESET_B(net458),
    .Q(\gpio_configure[25][5] ));
 sky130_fd_sc_hd__dfrtp_2 _9390_ (.CLK(clknet_leaf_1_csclk),
    .D(_0663_),
    .RESET_B(net418),
    .Q(\gpio_configure[25][6] ));
 sky130_fd_sc_hd__dfrtp_2 _9391_ (.CLK(clknet_leaf_2_csclk),
    .D(_0664_),
    .RESET_B(net418),
    .Q(\gpio_configure[25][7] ));
 sky130_fd_sc_hd__dfstp_1 _9392_ (.CLK(clknet_leaf_74_csclk),
    .D(_0665_),
    .SET_B(net425),
    .Q(\gpio_configure[26][0] ));
 sky130_fd_sc_hd__dfstp_2 _9393_ (.CLK(clknet_leaf_30_csclk),
    .D(_0666_),
    .SET_B(net476),
    .Q(\gpio_configure[26][1] ));
 sky130_fd_sc_hd__dfrtp_4 _9394_ (.CLK(clknet_leaf_3_csclk),
    .D(_0667_),
    .RESET_B(net417),
    .Q(\gpio_configure[26][2] ));
 sky130_fd_sc_hd__dfrtp_4 _9395_ (.CLK(clknet_leaf_31_csclk),
    .D(_0668_),
    .RESET_B(net480),
    .Q(\gpio_configure[26][3] ));
 sky130_fd_sc_hd__dfrtp_4 _9396_ (.CLK(clknet_leaf_17_csclk),
    .D(_0669_),
    .RESET_B(net465),
    .Q(\gpio_configure[26][4] ));
 sky130_fd_sc_hd__dfrtp_1 _9397_ (.CLK(clknet_leaf_10_csclk),
    .D(_0670_),
    .RESET_B(net461),
    .Q(\gpio_configure[26][5] ));
 sky130_fd_sc_hd__dfrtp_2 _9398_ (.CLK(clknet_leaf_1_csclk),
    .D(_0671_),
    .RESET_B(net418),
    .Q(\gpio_configure[26][6] ));
 sky130_fd_sc_hd__dfrtp_2 _9399_ (.CLK(clknet_leaf_2_csclk),
    .D(_0672_),
    .RESET_B(net417),
    .Q(\gpio_configure[26][7] ));
 sky130_fd_sc_hd__dfstp_1 _9400_ (.CLK(clknet_leaf_9_csclk),
    .D(_0673_),
    .SET_B(net425),
    .Q(\gpio_configure[27][0] ));
 sky130_fd_sc_hd__dfstp_4 _9401_ (.CLK(clknet_leaf_30_csclk),
    .D(_0674_),
    .SET_B(net479),
    .Q(\gpio_configure[27][1] ));
 sky130_fd_sc_hd__dfrtp_4 _9402_ (.CLK(clknet_leaf_28_csclk),
    .D(_0675_),
    .RESET_B(net475),
    .Q(\gpio_configure[27][2] ));
 sky130_fd_sc_hd__dfrtp_4 _9403_ (.CLK(clknet_leaf_36_csclk),
    .D(_0676_),
    .RESET_B(net482),
    .Q(\gpio_configure[27][3] ));
 sky130_fd_sc_hd__dfrtp_4 _9404_ (.CLK(clknet_leaf_17_csclk),
    .D(_0677_),
    .RESET_B(net465),
    .Q(\gpio_configure[27][4] ));
 sky130_fd_sc_hd__dfrtp_2 _9405_ (.CLK(clknet_leaf_12_csclk),
    .D(_0678_),
    .RESET_B(net458),
    .Q(\gpio_configure[27][5] ));
 sky130_fd_sc_hd__dfrtp_4 _9406_ (.CLK(clknet_leaf_5_csclk),
    .D(_0679_),
    .RESET_B(net423),
    .Q(\gpio_configure[27][6] ));
 sky130_fd_sc_hd__dfrtp_2 _9407_ (.CLK(clknet_leaf_5_csclk),
    .D(_0680_),
    .RESET_B(net423),
    .Q(\gpio_configure[27][7] ));
 sky130_fd_sc_hd__dfstp_2 _9408_ (.CLK(clknet_leaf_4_csclk),
    .D(_0681_),
    .SET_B(net420),
    .Q(\gpio_configure[28][0] ));
 sky130_fd_sc_hd__dfstp_4 _9409_ (.CLK(clknet_leaf_32_csclk),
    .D(_0682_),
    .SET_B(net480),
    .Q(\gpio_configure[28][1] ));
 sky130_fd_sc_hd__dfrtp_1 _9410_ (.CLK(clknet_leaf_28_csclk),
    .D(_0683_),
    .RESET_B(net475),
    .Q(\gpio_configure[28][2] ));
 sky130_fd_sc_hd__dfrtp_4 _9411_ (.CLK(clknet_leaf_31_csclk),
    .D(_0684_),
    .RESET_B(net480),
    .Q(\gpio_configure[28][3] ));
 sky130_fd_sc_hd__dfrtp_4 _9412_ (.CLK(clknet_leaf_16_csclk),
    .D(_0685_),
    .RESET_B(net465),
    .Q(\gpio_configure[28][4] ));
 sky130_fd_sc_hd__dfrtp_1 _9413_ (.CLK(clknet_leaf_13_csclk),
    .D(_0686_),
    .RESET_B(net458),
    .Q(\gpio_configure[28][5] ));
 sky130_fd_sc_hd__dfrtp_4 _9414_ (.CLK(clknet_leaf_3_csclk),
    .D(_0687_),
    .RESET_B(net421),
    .Q(\gpio_configure[28][6] ));
 sky130_fd_sc_hd__dfrtp_1 _9415_ (.CLK(clknet_leaf_5_csclk),
    .D(_0688_),
    .RESET_B(net424),
    .Q(\gpio_configure[28][7] ));
 sky130_fd_sc_hd__dfstp_2 _9416_ (.CLK(clknet_leaf_9_csclk),
    .D(_0689_),
    .SET_B(net426),
    .Q(\gpio_configure[29][0] ));
 sky130_fd_sc_hd__dfstp_1 _9417_ (.CLK(clknet_leaf_32_csclk),
    .D(_0690_),
    .SET_B(net479),
    .Q(\gpio_configure[29][1] ));
 sky130_fd_sc_hd__dfrtp_1 _9418_ (.CLK(clknet_leaf_27_csclk),
    .D(_0691_),
    .RESET_B(net475),
    .Q(\gpio_configure[29][2] ));
 sky130_fd_sc_hd__dfrtp_4 _9419_ (.CLK(clknet_leaf_36_csclk),
    .D(_0692_),
    .RESET_B(net491),
    .Q(\gpio_configure[29][3] ));
 sky130_fd_sc_hd__dfrtp_2 _9420_ (.CLK(clknet_leaf_17_csclk),
    .D(_0693_),
    .RESET_B(net465),
    .Q(\gpio_configure[29][4] ));
 sky130_fd_sc_hd__dfrtp_1 _9421_ (.CLK(clknet_leaf_11_csclk),
    .D(_0694_),
    .RESET_B(net461),
    .Q(\gpio_configure[29][5] ));
 sky130_fd_sc_hd__dfrtp_4 _9422_ (.CLK(clknet_leaf_4_csclk),
    .D(_0695_),
    .RESET_B(net421),
    .Q(\gpio_configure[29][6] ));
 sky130_fd_sc_hd__dfrtp_1 _9423_ (.CLK(clknet_leaf_5_csclk),
    .D(_0696_),
    .RESET_B(net421),
    .Q(\gpio_configure[29][7] ));
 sky130_fd_sc_hd__dfstp_2 _9424_ (.CLK(clknet_leaf_3_csclk),
    .D(_0697_),
    .SET_B(net417),
    .Q(\gpio_configure[30][0] ));
 sky130_fd_sc_hd__dfstp_4 _9425_ (.CLK(clknet_leaf_30_csclk),
    .D(_0698_),
    .SET_B(net476),
    .Q(\gpio_configure[30][1] ));
 sky130_fd_sc_hd__dfrtp_2 _9426_ (.CLK(clknet_leaf_28_csclk),
    .D(_0699_),
    .RESET_B(net475),
    .Q(\gpio_configure[30][2] ));
 sky130_fd_sc_hd__dfrtp_4 _9427_ (.CLK(clknet_leaf_30_csclk),
    .D(_0700_),
    .RESET_B(net478),
    .Q(\gpio_configure[30][3] ));
 sky130_fd_sc_hd__dfrtp_4 _9428_ (.CLK(clknet_leaf_16_csclk),
    .D(_0701_),
    .RESET_B(net465),
    .Q(\gpio_configure[30][4] ));
 sky130_fd_sc_hd__dfrtp_4 _9429_ (.CLK(clknet_leaf_10_csclk),
    .D(_0702_),
    .RESET_B(net461),
    .Q(\gpio_configure[30][5] ));
 sky130_fd_sc_hd__dfrtp_4 _9430_ (.CLK(clknet_leaf_3_csclk),
    .D(_0703_),
    .RESET_B(net421),
    .Q(\gpio_configure[30][6] ));
 sky130_fd_sc_hd__dfrtp_1 _9431_ (.CLK(clknet_leaf_3_csclk),
    .D(_0704_),
    .RESET_B(net421),
    .Q(\gpio_configure[30][7] ));
 sky130_fd_sc_hd__dfstp_1 _9432_ (.CLK(clknet_leaf_72_csclk),
    .D(_0705_),
    .SET_B(net450),
    .Q(\gpio_configure[31][0] ));
 sky130_fd_sc_hd__dfstp_4 _9433_ (.CLK(clknet_leaf_31_csclk),
    .D(_0706_),
    .SET_B(net481),
    .Q(\gpio_configure[31][1] ));
 sky130_fd_sc_hd__dfrtp_4 _9434_ (.CLK(clknet_leaf_72_csclk),
    .D(_0707_),
    .RESET_B(net450),
    .Q(\gpio_configure[31][2] ));
 sky130_fd_sc_hd__dfrtp_4 _9435_ (.CLK(clknet_leaf_31_csclk),
    .D(_0708_),
    .RESET_B(net491),
    .Q(\gpio_configure[31][3] ));
 sky130_fd_sc_hd__dfrtp_1 _9436_ (.CLK(clknet_leaf_20_csclk),
    .D(_0709_),
    .RESET_B(net462),
    .Q(\gpio_configure[31][4] ));
 sky130_fd_sc_hd__dfrtp_4 _9437_ (.CLK(clknet_leaf_0_csclk),
    .D(_0710_),
    .RESET_B(net410),
    .Q(\gpio_configure[31][5] ));
 sky130_fd_sc_hd__dfrtp_4 _9438_ (.CLK(clknet_leaf_82_csclk),
    .D(_0711_),
    .RESET_B(net409),
    .Q(\gpio_configure[31][6] ));
 sky130_fd_sc_hd__dfrtp_2 _9439_ (.CLK(clknet_leaf_82_csclk),
    .D(_0712_),
    .RESET_B(net409),
    .Q(\gpio_configure[31][7] ));
 sky130_fd_sc_hd__dfstp_1 _9440_ (.CLK(clknet_leaf_79_csclk),
    .D(_0713_),
    .SET_B(net414),
    .Q(\gpio_configure[32][0] ));
 sky130_fd_sc_hd__dfstp_1 _9441_ (.CLK(clknet_leaf_65_csclk),
    .D(_0714_),
    .SET_B(net432),
    .Q(\gpio_configure[32][1] ));
 sky130_fd_sc_hd__dfrtp_1 _9442_ (.CLK(clknet_leaf_62_csclk),
    .D(_0715_),
    .RESET_B(net438),
    .Q(\gpio_configure[32][2] ));
 sky130_fd_sc_hd__dfrtp_4 _9443_ (.CLK(clknet_leaf_32_csclk),
    .D(net554),
    .RESET_B(net489),
    .Q(\gpio_configure[32][3] ));
 sky130_fd_sc_hd__dfrtp_2 _9444_ (.CLK(clknet_leaf_67_csclk),
    .D(_0717_),
    .RESET_B(net429),
    .Q(\gpio_configure[32][4] ));
 sky130_fd_sc_hd__dfrtp_1 _9445_ (.CLK(clknet_leaf_83_csclk),
    .D(_0718_),
    .RESET_B(net411),
    .Q(\gpio_configure[32][5] ));
 sky130_fd_sc_hd__dfrtp_1 _9446_ (.CLK(clknet_leaf_81_csclk),
    .D(_0719_),
    .RESET_B(net413),
    .Q(\gpio_configure[32][6] ));
 sky130_fd_sc_hd__dfrtp_1 _9447_ (.CLK(clknet_leaf_81_csclk),
    .D(_0720_),
    .RESET_B(net413),
    .Q(\gpio_configure[32][7] ));
 sky130_fd_sc_hd__dfstp_2 _9448_ (.CLK(clknet_leaf_78_csclk),
    .D(_0721_),
    .SET_B(net414),
    .Q(\gpio_configure[33][0] ));
 sky130_fd_sc_hd__dfstp_1 _9449_ (.CLK(clknet_leaf_33_csclk),
    .D(_0722_),
    .SET_B(net474),
    .Q(\gpio_configure[33][1] ));
 sky130_fd_sc_hd__dfrtp_4 _9450_ (.CLK(clknet_leaf_68_csclk),
    .D(_0723_),
    .RESET_B(net427),
    .Q(\gpio_configure[33][2] ));
 sky130_fd_sc_hd__dfrtp_4 _9451_ (.CLK(clknet_leaf_32_csclk),
    .D(_0724_),
    .RESET_B(net480),
    .Q(\gpio_configure[33][3] ));
 sky130_fd_sc_hd__dfrtp_4 _9452_ (.CLK(clknet_leaf_77_csclk),
    .D(_0725_),
    .RESET_B(net416),
    .Q(\gpio_configure[33][4] ));
 sky130_fd_sc_hd__dfrtp_1 _9453_ (.CLK(clknet_leaf_10_csclk),
    .D(_0726_),
    .RESET_B(net461),
    .Q(\gpio_configure[33][5] ));
 sky130_fd_sc_hd__dfrtp_2 _9454_ (.CLK(clknet_leaf_85_csclk),
    .D(_0727_),
    .RESET_B(net408),
    .Q(\gpio_configure[33][6] ));
 sky130_fd_sc_hd__dfrtp_1 _9455_ (.CLK(clknet_leaf_3_csclk),
    .D(_0728_),
    .RESET_B(net421),
    .Q(\gpio_configure[33][7] ));
 sky130_fd_sc_hd__dfstp_2 _9456_ (.CLK(clknet_leaf_84_csclk),
    .D(_0729_),
    .SET_B(net404),
    .Q(\gpio_configure[34][0] ));
 sky130_fd_sc_hd__dfstp_1 _9457_ (.CLK(clknet_leaf_66_csclk),
    .D(_0730_),
    .SET_B(net430),
    .Q(\gpio_configure[34][1] ));
 sky130_fd_sc_hd__dfrtp_1 _9458_ (.CLK(clknet_leaf_68_csclk),
    .D(_0731_),
    .RESET_B(net427),
    .Q(\gpio_configure[34][2] ));
 sky130_fd_sc_hd__dfrtp_4 _9459_ (.CLK(clknet_leaf_32_csclk),
    .D(_0732_),
    .RESET_B(net491),
    .Q(\gpio_configure[34][3] ));
 sky130_fd_sc_hd__dfrtp_4 _9460_ (.CLK(clknet_leaf_78_csclk),
    .D(_0733_),
    .RESET_B(net414),
    .Q(\gpio_configure[34][4] ));
 sky130_fd_sc_hd__dfrtp_1 _9461_ (.CLK(clknet_leaf_5_csclk),
    .D(_0734_),
    .RESET_B(net423),
    .Q(\gpio_configure[34][5] ));
 sky130_fd_sc_hd__dfrtp_1 _9462_ (.CLK(clknet_leaf_85_csclk),
    .D(_0735_),
    .RESET_B(net408),
    .Q(\gpio_configure[34][6] ));
 sky130_fd_sc_hd__dfrtp_1 _9463_ (.CLK(clknet_leaf_2_csclk),
    .D(_0736_),
    .RESET_B(net410),
    .Q(\gpio_configure[34][7] ));
 sky130_fd_sc_hd__dfstp_1 _9464_ (.CLK(clknet_leaf_4_csclk),
    .D(_0737_),
    .SET_B(net421),
    .Q(\gpio_configure[35][0] ));
 sky130_fd_sc_hd__dfstp_1 _9465_ (.CLK(clknet_leaf_26_csclk),
    .D(_0738_),
    .SET_B(net472),
    .Q(\gpio_configure[35][1] ));
 sky130_fd_sc_hd__dfrtp_2 _9466_ (.CLK(clknet_leaf_27_csclk),
    .D(_0739_),
    .RESET_B(net475),
    .Q(\gpio_configure[35][2] ));
 sky130_fd_sc_hd__dfrtp_4 _9467_ (.CLK(clknet_leaf_28_csclk),
    .D(_0740_),
    .RESET_B(net476),
    .Q(\gpio_configure[35][3] ));
 sky130_fd_sc_hd__dfrtp_4 _9468_ (.CLK(clknet_leaf_16_csclk),
    .D(_0741_),
    .RESET_B(net465),
    .Q(\gpio_configure[35][4] ));
 sky130_fd_sc_hd__dfrtp_1 _9469_ (.CLK(clknet_leaf_12_csclk),
    .D(_0742_),
    .RESET_B(net459),
    .Q(\gpio_configure[35][5] ));
 sky130_fd_sc_hd__dfrtp_2 _9470_ (.CLK(clknet_leaf_3_csclk),
    .D(_0743_),
    .RESET_B(net421),
    .Q(\gpio_configure[35][6] ));
 sky130_fd_sc_hd__dfrtp_1 _9471_ (.CLK(clknet_leaf_3_csclk),
    .D(_0744_),
    .RESET_B(net421),
    .Q(\gpio_configure[35][7] ));
 sky130_fd_sc_hd__dfstp_2 _9472_ (.CLK(clknet_leaf_78_csclk),
    .D(_0745_),
    .SET_B(net414),
    .Q(\gpio_configure[36][0] ));
 sky130_fd_sc_hd__dfstp_1 _9473_ (.CLK(clknet_leaf_66_csclk),
    .D(_0746_),
    .SET_B(net431),
    .Q(\gpio_configure[36][1] ));
 sky130_fd_sc_hd__dfrtp_1 _9474_ (.CLK(clknet_leaf_68_csclk),
    .D(_0747_),
    .RESET_B(net429),
    .Q(\gpio_configure[36][2] ));
 sky130_fd_sc_hd__dfrtp_4 _9475_ (.CLK(clknet_leaf_31_csclk),
    .D(_0748_),
    .RESET_B(net482),
    .Q(\gpio_configure[36][3] ));
 sky130_fd_sc_hd__dfrtp_1 _9476_ (.CLK(clknet_leaf_78_csclk),
    .D(_0749_),
    .RESET_B(net414),
    .Q(\gpio_configure[36][4] ));
 sky130_fd_sc_hd__dfrtp_1 _9477_ (.CLK(clknet_leaf_82_csclk),
    .D(_0750_),
    .RESET_B(net406),
    .Q(\gpio_configure[36][5] ));
 sky130_fd_sc_hd__dfrtp_1 _9478_ (.CLK(clknet_leaf_83_csclk),
    .D(_0751_),
    .RESET_B(net405),
    .Q(\gpio_configure[36][6] ));
 sky130_fd_sc_hd__dfrtp_1 _9479_ (.CLK(clknet_leaf_83_csclk),
    .D(_0752_),
    .RESET_B(net405),
    .Q(\gpio_configure[36][7] ));
 sky130_fd_sc_hd__dfstp_1 _9480_ (.CLK(clknet_leaf_79_csclk),
    .D(_0753_),
    .SET_B(net415),
    .Q(\gpio_configure[37][0] ));
 sky130_fd_sc_hd__dfstp_1 _9481_ (.CLK(clknet_leaf_65_csclk),
    .D(_0754_),
    .SET_B(net435),
    .Q(\gpio_configure[37][1] ));
 sky130_fd_sc_hd__dfrtp_1 _9482_ (.CLK(clknet_leaf_65_csclk),
    .D(_0755_),
    .RESET_B(net435),
    .Q(\gpio_configure[37][2] ));
 sky130_fd_sc_hd__dfrtp_4 _9483_ (.CLK(clknet_leaf_25_csclk),
    .D(_0756_),
    .RESET_B(net474),
    .Q(\gpio_configure[37][3] ));
 sky130_fd_sc_hd__dfrtp_4 _9484_ (.CLK(clknet_leaf_67_csclk),
    .D(_0757_),
    .RESET_B(net429),
    .Q(\gpio_configure[37][4] ));
 sky130_fd_sc_hd__dfrtp_1 _9485_ (.CLK(clknet_leaf_83_csclk),
    .D(_0758_),
    .RESET_B(net413),
    .Q(\gpio_configure[37][5] ));
 sky130_fd_sc_hd__dfrtp_1 _9486_ (.CLK(clknet_leaf_81_csclk),
    .D(_0759_),
    .RESET_B(net416),
    .Q(\gpio_configure[37][6] ));
 sky130_fd_sc_hd__dfrtp_1 _9487_ (.CLK(clknet_leaf_80_csclk),
    .D(_0760_),
    .RESET_B(net411),
    .Q(\gpio_configure[37][7] ));
 sky130_fd_sc_hd__dfrtp_2 _9488_ (.CLK(clknet_3_3_0_wb_clk_i),
    .D(_0761_),
    .RESET_B(net440),
    .Q(\xfer_count[0] ));
 sky130_fd_sc_hd__dfrtp_2 _9489_ (.CLK(clknet_3_2_0_wb_clk_i),
    .D(_0762_),
    .RESET_B(net442),
    .Q(\xfer_count[1] ));
 sky130_fd_sc_hd__dfrtp_1 _9490_ (.CLK(clknet_3_0_0_wb_clk_i),
    .D(_0763_),
    .RESET_B(net441),
    .Q(\xfer_count[2] ));
 sky130_fd_sc_hd__dfrtp_1 _9491_ (.CLK(clknet_3_2_0_wb_clk_i),
    .D(_0764_),
    .RESET_B(net441),
    .Q(\xfer_count[3] ));
 sky130_fd_sc_hd__dfrtp_4 _9492_ (.CLK(clknet_3_1_0_wb_clk_i),
    .D(_0765_),
    .RESET_B(net469),
    .Q(\pad_count_1[0] ));
 sky130_fd_sc_hd__dfstp_2 _9493_ (.CLK(clknet_3_1_0_wb_clk_i),
    .D(_0766_),
    .SET_B(net469),
    .Q(\pad_count_1[1] ));
 sky130_fd_sc_hd__dfrtp_2 _9494_ (.CLK(clknet_3_1_0_wb_clk_i),
    .D(_0767_),
    .RESET_B(net469),
    .Q(\pad_count_1[2] ));
 sky130_fd_sc_hd__dfrtp_4 _9495_ (.CLK(clknet_3_1_0_wb_clk_i),
    .D(_0768_),
    .RESET_B(net470),
    .Q(\pad_count_1[3] ));
 sky130_fd_sc_hd__dfstp_4 _9496_ (.CLK(clknet_3_1_0_wb_clk_i),
    .D(_0769_),
    .SET_B(net470),
    .Q(\pad_count_1[4] ));
 sky130_fd_sc_hd__dfstp_1 _9497_ (.CLK(net508),
    .D(_0770_),
    .SET_B(net488),
    .Q(\pad_count_2[0] ));
 sky130_fd_sc_hd__dfstp_1 _9498_ (.CLK(net508),
    .D(_0771_),
    .SET_B(net488),
    .Q(\pad_count_2[1] ));
 sky130_fd_sc_hd__dfrtp_2 _9499_ (.CLK(net508),
    .D(_0772_),
    .RESET_B(net470),
    .Q(\pad_count_2[2] ));
 sky130_fd_sc_hd__dfrtp_2 _9500_ (.CLK(net508),
    .D(_0773_),
    .RESET_B(net470),
    .Q(\pad_count_2[3] ));
 sky130_fd_sc_hd__dfstp_2 _9501_ (.CLK(net508),
    .D(_0774_),
    .SET_B(net470),
    .Q(\pad_count_2[4] ));
 sky130_fd_sc_hd__dfrtp_2 _9502_ (.CLK(clknet_3_1_0_wb_clk_i),
    .D(_0775_),
    .RESET_B(net470),
    .Q(\pad_count_2[5] ));
 sky130_fd_sc_hd__dfrtp_1 _9503_ (.CLK(clknet_3_2_0_wb_clk_i),
    .D(net504),
    .RESET_B(net441),
    .Q(serial_resetn_pre));
 sky130_fd_sc_hd__dfrtp_1 _9504_ (.CLK(clknet_3_3_0_wb_clk_i),
    .D(_0776_),
    .RESET_B(net441),
    .Q(serial_clock_pre));
 sky130_fd_sc_hd__dfrtp_1 _9505_ (.CLK(clknet_3_3_0_wb_clk_i),
    .D(net1451),
    .RESET_B(net442),
    .Q(serial_load_pre));
 sky130_fd_sc_hd__dfrtp_1 _9506_ (.CLK(clknet_3_3_0_wb_clk_i),
    .D(_0778_),
    .RESET_B(net442),
    .Q(serial_busy));
 sky130_fd_sc_hd__dfrtp_1 _9507_ (.CLK(clknet_3_0_0_wb_clk_i),
    .D(_0779_),
    .RESET_B(net454),
    .Q(\serial_data_staging_1[0] ));
 sky130_fd_sc_hd__dfrtp_1 _9508_ (.CLK(clknet_3_1_0_wb_clk_i),
    .D(net1454),
    .RESET_B(net454),
    .Q(\serial_data_staging_1[1] ));
 sky130_fd_sc_hd__dfrtp_1 _9509_ (.CLK(clknet_3_1_0_wb_clk_i),
    .D(_0781_),
    .RESET_B(net454),
    .Q(\serial_data_staging_1[2] ));
 sky130_fd_sc_hd__dfrtp_1 _9510_ (.CLK(clknet_3_0_0_wb_clk_i),
    .D(net1481),
    .RESET_B(net454),
    .Q(\serial_data_staging_1[3] ));
 sky130_fd_sc_hd__dfrtp_1 _9511_ (.CLK(clknet_3_0_0_wb_clk_i),
    .D(_0783_),
    .RESET_B(net451),
    .Q(\serial_data_staging_1[4] ));
 sky130_fd_sc_hd__dfrtp_1 _9512_ (.CLK(clknet_3_0_0_wb_clk_i),
    .D(_0784_),
    .RESET_B(net451),
    .Q(\serial_data_staging_1[5] ));
 sky130_fd_sc_hd__dfrtp_1 _9513_ (.CLK(clknet_3_0_0_wb_clk_i),
    .D(net1483),
    .RESET_B(net452),
    .Q(\serial_data_staging_1[6] ));
 sky130_fd_sc_hd__dfrtp_1 _9514_ (.CLK(clknet_3_0_0_wb_clk_i),
    .D(_0786_),
    .RESET_B(net452),
    .Q(\serial_data_staging_1[7] ));
 sky130_fd_sc_hd__dfrtp_1 _9515_ (.CLK(clknet_3_0_0_wb_clk_i),
    .D(_0787_),
    .RESET_B(net452),
    .Q(\serial_data_staging_1[8] ));
 sky130_fd_sc_hd__dfrtp_1 _9516_ (.CLK(clknet_3_0_0_wb_clk_i),
    .D(net1485),
    .RESET_B(net452),
    .Q(\serial_data_staging_1[9] ));
 sky130_fd_sc_hd__dfrtp_1 _9517_ (.CLK(clknet_3_0_0_wb_clk_i),
    .D(_0789_),
    .RESET_B(net452),
    .Q(\serial_data_staging_1[10] ));
 sky130_fd_sc_hd__dfrtp_1 _9518_ (.CLK(clknet_3_0_0_wb_clk_i),
    .D(net1492),
    .RESET_B(net452),
    .Q(\serial_data_staging_1[11] ));
 sky130_fd_sc_hd__dfrtp_1 _9519_ (.CLK(clknet_3_3_0_wb_clk_i),
    .D(net1494),
    .RESET_B(net446),
    .Q(\serial_data_staging_1[12] ));
 sky130_fd_sc_hd__dfrtp_1 _9520_ (.CLK(clknet_3_1_0_wb_clk_i),
    .D(_0792_),
    .RESET_B(net454),
    .Q(\serial_data_staging_2[0] ));
 sky130_fd_sc_hd__dfrtp_1 _9521_ (.CLK(clknet_3_3_0_wb_clk_i),
    .D(_0793_),
    .RESET_B(net451),
    .Q(\serial_data_staging_2[1] ));
 sky130_fd_sc_hd__dfrtp_1 _9522_ (.CLK(clknet_3_3_0_wb_clk_i),
    .D(net1475),
    .RESET_B(net451),
    .Q(\serial_data_staging_2[2] ));
 sky130_fd_sc_hd__dfrtp_1 _9523_ (.CLK(clknet_3_3_0_wb_clk_i),
    .D(_0795_),
    .RESET_B(net451),
    .Q(\serial_data_staging_2[3] ));
 sky130_fd_sc_hd__dfrtp_1 _9524_ (.CLK(clknet_3_3_0_wb_clk_i),
    .D(net1461),
    .RESET_B(net451),
    .Q(\serial_data_staging_2[4] ));
 sky130_fd_sc_hd__dfrtp_1 _9525_ (.CLK(clknet_3_3_0_wb_clk_i),
    .D(_0797_),
    .RESET_B(net451),
    .Q(\serial_data_staging_2[5] ));
 sky130_fd_sc_hd__dfrtp_1 _9526_ (.CLK(clknet_3_3_0_wb_clk_i),
    .D(_0798_),
    .RESET_B(net447),
    .Q(\serial_data_staging_2[6] ));
 sky130_fd_sc_hd__dfrtp_1 _9527_ (.CLK(clknet_3_3_0_wb_clk_i),
    .D(net1497),
    .RESET_B(net448),
    .Q(\serial_data_staging_2[7] ));
 sky130_fd_sc_hd__dfrtp_1 _9528_ (.CLK(clknet_3_2_0_wb_clk_i),
    .D(net1466),
    .RESET_B(net448),
    .Q(\serial_data_staging_2[8] ));
 sky130_fd_sc_hd__dfrtp_1 _9529_ (.CLK(clknet_3_3_0_wb_clk_i),
    .D(_0801_),
    .RESET_B(net448),
    .Q(\serial_data_staging_2[9] ));
 sky130_fd_sc_hd__dfrtp_1 _9530_ (.CLK(clknet_3_0_0_wb_clk_i),
    .D(_0802_),
    .RESET_B(net448),
    .Q(\serial_data_staging_2[10] ));
 sky130_fd_sc_hd__dfrtp_1 _9531_ (.CLK(clknet_3_0_0_wb_clk_i),
    .D(net1477),
    .RESET_B(net446),
    .Q(\serial_data_staging_2[11] ));
 sky130_fd_sc_hd__dfrtp_1 _9532_ (.CLK(clknet_3_2_0_wb_clk_i),
    .D(net1504),
    .RESET_B(net446),
    .Q(\serial_data_staging_2[12] ));
 sky130_fd_sc_hd__dfrtp_4 _9533_ (.CLK(clknet_3_7_0_wb_clk_i),
    .D(_0805_),
    .RESET_B(net501),
    .Q(net326));
 sky130_fd_sc_hd__dfxtp_1 _9534_ (.CLK(clknet_3_5_0_wb_clk_i),
    .D(_0806_),
    .Q(net343));
 sky130_fd_sc_hd__dfxtp_1 _9535_ (.CLK(clknet_3_5_0_wb_clk_i),
    .D(_0807_),
    .Q(net344));
 sky130_fd_sc_hd__dfxtp_1 _9536_ (.CLK(clknet_3_5_0_wb_clk_i),
    .D(_0808_),
    .Q(net345));
 sky130_fd_sc_hd__dfxtp_1 _9537_ (.CLK(clknet_3_5_0_wb_clk_i),
    .D(_0809_),
    .Q(net346));
 sky130_fd_sc_hd__dfxtp_1 _9538_ (.CLK(clknet_3_5_0_wb_clk_i),
    .D(_0810_),
    .Q(net347));
 sky130_fd_sc_hd__dfxtp_1 _9539_ (.CLK(clknet_3_5_0_wb_clk_i),
    .D(_0811_),
    .Q(net348));
 sky130_fd_sc_hd__dfxtp_1 _9540_ (.CLK(clknet_3_5_0_wb_clk_i),
    .D(_0812_),
    .Q(net350));
 sky130_fd_sc_hd__dfxtp_1 _9541_ (.CLK(clknet_3_5_0_wb_clk_i),
    .D(_0813_),
    .Q(net351));
 sky130_fd_sc_hd__dfrtp_1 _9542_ (.CLK(net507),
    .D(_0814_),
    .RESET_B(net499),
    .Q(\wbbd_data[0] ));
 sky130_fd_sc_hd__dfrtp_1 _9543_ (.CLK(clknet_3_7_0_wb_clk_i),
    .D(_0815_),
    .RESET_B(net500),
    .Q(\wbbd_data[1] ));
 sky130_fd_sc_hd__dfrtp_1 _9544_ (.CLK(net507),
    .D(_0816_),
    .RESET_B(net500),
    .Q(\wbbd_data[2] ));
 sky130_fd_sc_hd__dfrtp_1 _9545_ (.CLK(net507),
    .D(_0817_),
    .RESET_B(net500),
    .Q(\wbbd_data[3] ));
 sky130_fd_sc_hd__dfrtp_1 _9546_ (.CLK(clknet_3_7_0_wb_clk_i),
    .D(_0818_),
    .RESET_B(net500),
    .Q(\wbbd_data[4] ));
 sky130_fd_sc_hd__dfrtp_1 _9547_ (.CLK(net507),
    .D(_0819_),
    .RESET_B(net501),
    .Q(\wbbd_data[5] ));
 sky130_fd_sc_hd__dfrtp_1 _9548_ (.CLK(clknet_3_7_0_wb_clk_i),
    .D(_0820_),
    .RESET_B(net500),
    .Q(\wbbd_data[6] ));
 sky130_fd_sc_hd__dfrtp_1 _9549_ (.CLK(net507),
    .D(_0821_),
    .RESET_B(net500),
    .Q(\wbbd_data[7] ));
 sky130_fd_sc_hd__dfrtp_2 _9550_ (.CLK(net507),
    .D(_0822_),
    .RESET_B(net501),
    .Q(wbbd_sck));
 sky130_fd_sc_hd__dfrtp_1 _9551_ (.CLK(clknet_3_7_0_wb_clk_i),
    .D(_0823_),
    .RESET_B(net501),
    .Q(wbbd_write));
 sky130_fd_sc_hd__inv_2 _5235__1 (.A(clknet_2_2_0_mgmt_gpio_in[4]),
    .Y(net505));
 sky130_fd_sc_hd__clkbuf_2 _9553_ (.A(net87),
    .X(net257));
 sky130_fd_sc_hd__clkbuf_1 _9554_ (.A(net65),
    .X(net314));
 sky130_fd_sc_hd__clkbuf_1 _9555_ (.A(net66),
    .X(net315));
 sky130_fd_sc_hd__ebufn_8 _9556_ (.A(\mgmt_gpio_data[2] ),
    .TE_B(_4315_),
    .Z(mgmt_gpio_out[2]));
 sky130_fd_sc_hd__ebufn_8 _9557_ (.A(\mgmt_gpio_data[3] ),
    .TE_B(_4316_),
    .Z(mgmt_gpio_out[3]));
 sky130_fd_sc_hd__ebufn_8 _9558_ (.A(\mgmt_gpio_data[4] ),
    .TE_B(_4317_),
    .Z(mgmt_gpio_out[4]));
 sky130_fd_sc_hd__ebufn_8 _9559_ (.A(\mgmt_gpio_data[5] ),
    .TE_B(_4318_),
    .Z(mgmt_gpio_out[5]));
 sky130_fd_sc_hd__ebufn_8 _9560_ (.A(\mgmt_gpio_out_pre[6] ),
    .TE_B(_4319_),
    .Z(mgmt_gpio_out[6]));
 sky130_fd_sc_hd__ebufn_8 _9561_ (.A(\mgmt_gpio_data[7] ),
    .TE_B(_4320_),
    .Z(mgmt_gpio_out[7]));
 sky130_fd_sc_hd__ebufn_8 _9562_ (.A(\mgmt_gpio_out_pre[8] ),
    .TE_B(_4321_),
    .Z(mgmt_gpio_out[8]));
 sky130_fd_sc_hd__ebufn_2 _9563_ (.A(\mgmt_gpio_out_pre[9] ),
    .TE_B(_4322_),
    .Z(mgmt_gpio_out[9]));
 sky130_fd_sc_hd__ebufn_8 _9564_ (.A(\mgmt_gpio_out_pre[10] ),
    .TE_B(_4323_),
    .Z(mgmt_gpio_out[10]));
 sky130_fd_sc_hd__ebufn_8 _9565_ (.A(\mgmt_gpio_data[11] ),
    .TE_B(_4324_),
    .Z(mgmt_gpio_out[11]));
 sky130_fd_sc_hd__ebufn_8 _9566_ (.A(\mgmt_gpio_data[12] ),
    .TE_B(_4325_),
    .Z(mgmt_gpio_out[12]));
 sky130_fd_sc_hd__ebufn_8 _9567_ (.A(\mgmt_gpio_out_pre[13] ),
    .TE_B(_4326_),
    .Z(mgmt_gpio_out[13]));
 sky130_fd_sc_hd__ebufn_8 _9568_ (.A(\mgmt_gpio_out_pre[14] ),
    .TE_B(_4327_),
    .Z(mgmt_gpio_out[14]));
 sky130_fd_sc_hd__ebufn_2 _9569_ (.A(\mgmt_gpio_out_pre[15] ),
    .TE_B(_4328_),
    .Z(mgmt_gpio_out[15]));
 sky130_fd_sc_hd__ebufn_8 _9570_ (.A(\mgmt_gpio_data[16] ),
    .TE_B(_4329_),
    .Z(mgmt_gpio_out[16]));
 sky130_fd_sc_hd__ebufn_8 _9571_ (.A(\mgmt_gpio_data[17] ),
    .TE_B(_4330_),
    .Z(mgmt_gpio_out[17]));
 sky130_fd_sc_hd__ebufn_8 _9572_ (.A(\mgmt_gpio_data[18] ),
    .TE_B(_4331_),
    .Z(mgmt_gpio_out[18]));
 sky130_fd_sc_hd__ebufn_8 _9573_ (.A(\mgmt_gpio_data[19] ),
    .TE_B(_4332_),
    .Z(mgmt_gpio_out[19]));
 sky130_fd_sc_hd__ebufn_8 _9574_ (.A(\mgmt_gpio_data[20] ),
    .TE_B(_4333_),
    .Z(mgmt_gpio_out[20]));
 sky130_fd_sc_hd__ebufn_8 _9575_ (.A(\mgmt_gpio_data[21] ),
    .TE_B(_4334_),
    .Z(mgmt_gpio_out[21]));
 sky130_fd_sc_hd__ebufn_8 _9576_ (.A(\mgmt_gpio_data[22] ),
    .TE_B(_4335_),
    .Z(mgmt_gpio_out[22]));
 sky130_fd_sc_hd__ebufn_8 _9577_ (.A(\mgmt_gpio_data[23] ),
    .TE_B(_4336_),
    .Z(mgmt_gpio_out[23]));
 sky130_fd_sc_hd__ebufn_8 _9578_ (.A(\mgmt_gpio_data[24] ),
    .TE_B(_4337_),
    .Z(mgmt_gpio_out[24]));
 sky130_fd_sc_hd__ebufn_8 _9579_ (.A(\mgmt_gpio_data[25] ),
    .TE_B(_4338_),
    .Z(mgmt_gpio_out[25]));
 sky130_fd_sc_hd__ebufn_8 _9580_ (.A(\mgmt_gpio_data[26] ),
    .TE_B(_4339_),
    .Z(mgmt_gpio_out[26]));
 sky130_fd_sc_hd__ebufn_8 _9581_ (.A(\mgmt_gpio_data[27] ),
    .TE_B(_4340_),
    .Z(mgmt_gpio_out[27]));
 sky130_fd_sc_hd__ebufn_8 _9582_ (.A(\mgmt_gpio_data[28] ),
    .TE_B(_4341_),
    .Z(mgmt_gpio_out[28]));
 sky130_fd_sc_hd__ebufn_8 _9583_ (.A(\mgmt_gpio_data[29] ),
    .TE_B(_4342_),
    .Z(mgmt_gpio_out[29]));
 sky130_fd_sc_hd__ebufn_8 _9584_ (.A(\mgmt_gpio_data[30] ),
    .TE_B(_4343_),
    .Z(mgmt_gpio_out[30]));
 sky130_fd_sc_hd__ebufn_8 _9585_ (.A(\mgmt_gpio_data[31] ),
    .TE_B(_4344_),
    .Z(mgmt_gpio_out[31]));
 sky130_fd_sc_hd__ebufn_8 _9586_ (.A(\mgmt_gpio_out_pre[32] ),
    .TE_B(_4345_),
    .Z(mgmt_gpio_out[32]));
 sky130_fd_sc_hd__ebufn_8 _9587_ (.A(\mgmt_gpio_out_pre[33] ),
    .TE_B(_4346_),
    .Z(mgmt_gpio_out[33]));
 sky130_fd_sc_hd__ebufn_8 _9588_ (.A(\mgmt_gpio_data[34] ),
    .TE_B(_4347_),
    .Z(mgmt_gpio_out[34]));
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_28 ();
 sky130_fd_sc_hd__decap_3 PHY_29 ();
 sky130_fd_sc_hd__decap_3 PHY_30 ();
 sky130_fd_sc_hd__decap_3 PHY_31 ();
 sky130_fd_sc_hd__decap_3 PHY_32 ();
 sky130_fd_sc_hd__decap_3 PHY_33 ();
 sky130_fd_sc_hd__decap_3 PHY_34 ();
 sky130_fd_sc_hd__decap_3 PHY_35 ();
 sky130_fd_sc_hd__decap_3 PHY_36 ();
 sky130_fd_sc_hd__decap_3 PHY_37 ();
 sky130_fd_sc_hd__decap_3 PHY_38 ();
 sky130_fd_sc_hd__decap_3 PHY_39 ();
 sky130_fd_sc_hd__decap_3 PHY_40 ();
 sky130_fd_sc_hd__decap_3 PHY_41 ();
 sky130_fd_sc_hd__decap_3 PHY_42 ();
 sky130_fd_sc_hd__decap_3 PHY_43 ();
 sky130_fd_sc_hd__decap_3 PHY_44 ();
 sky130_fd_sc_hd__decap_3 PHY_45 ();
 sky130_fd_sc_hd__decap_3 PHY_46 ();
 sky130_fd_sc_hd__decap_3 PHY_47 ();
 sky130_fd_sc_hd__decap_3 PHY_48 ();
 sky130_fd_sc_hd__decap_3 PHY_49 ();
 sky130_fd_sc_hd__decap_3 PHY_50 ();
 sky130_fd_sc_hd__decap_3 PHY_51 ();
 sky130_fd_sc_hd__decap_3 PHY_52 ();
 sky130_fd_sc_hd__decap_3 PHY_53 ();
 sky130_fd_sc_hd__decap_3 PHY_54 ();
 sky130_fd_sc_hd__decap_3 PHY_55 ();
 sky130_fd_sc_hd__decap_3 PHY_56 ();
 sky130_fd_sc_hd__decap_3 PHY_57 ();
 sky130_fd_sc_hd__decap_3 PHY_58 ();
 sky130_fd_sc_hd__decap_3 PHY_59 ();
 sky130_fd_sc_hd__decap_3 PHY_60 ();
 sky130_fd_sc_hd__decap_3 PHY_61 ();
 sky130_fd_sc_hd__decap_3 PHY_62 ();
 sky130_fd_sc_hd__decap_3 PHY_63 ();
 sky130_fd_sc_hd__decap_3 PHY_64 ();
 sky130_fd_sc_hd__decap_3 PHY_65 ();
 sky130_fd_sc_hd__decap_3 PHY_66 ();
 sky130_fd_sc_hd__decap_3 PHY_67 ();
 sky130_fd_sc_hd__decap_3 PHY_68 ();
 sky130_fd_sc_hd__decap_3 PHY_69 ();
 sky130_fd_sc_hd__decap_3 PHY_70 ();
 sky130_fd_sc_hd__decap_3 PHY_71 ();
 sky130_fd_sc_hd__decap_3 PHY_72 ();
 sky130_fd_sc_hd__decap_3 PHY_73 ();
 sky130_fd_sc_hd__decap_3 PHY_74 ();
 sky130_fd_sc_hd__decap_3 PHY_75 ();
 sky130_fd_sc_hd__decap_3 PHY_76 ();
 sky130_fd_sc_hd__decap_3 PHY_77 ();
 sky130_fd_sc_hd__decap_3 PHY_78 ();
 sky130_fd_sc_hd__decap_3 PHY_79 ();
 sky130_fd_sc_hd__decap_3 PHY_80 ();
 sky130_fd_sc_hd__decap_3 PHY_81 ();
 sky130_fd_sc_hd__decap_3 PHY_82 ();
 sky130_fd_sc_hd__decap_3 PHY_83 ();
 sky130_fd_sc_hd__decap_3 PHY_84 ();
 sky130_fd_sc_hd__decap_3 PHY_85 ();
 sky130_fd_sc_hd__decap_3 PHY_86 ();
 sky130_fd_sc_hd__decap_3 PHY_87 ();
 sky130_fd_sc_hd__decap_3 PHY_88 ();
 sky130_fd_sc_hd__decap_3 PHY_89 ();
 sky130_fd_sc_hd__decap_3 PHY_90 ();
 sky130_fd_sc_hd__decap_3 PHY_91 ();
 sky130_fd_sc_hd__decap_3 PHY_92 ();
 sky130_fd_sc_hd__decap_3 PHY_93 ();
 sky130_fd_sc_hd__decap_3 PHY_94 ();
 sky130_fd_sc_hd__decap_3 PHY_95 ();
 sky130_fd_sc_hd__decap_3 PHY_96 ();
 sky130_fd_sc_hd__decap_3 PHY_97 ();
 sky130_fd_sc_hd__decap_3 PHY_98 ();
 sky130_fd_sc_hd__decap_3 PHY_99 ();
 sky130_fd_sc_hd__decap_3 PHY_100 ();
 sky130_fd_sc_hd__decap_3 PHY_101 ();
 sky130_fd_sc_hd__decap_3 PHY_102 ();
 sky130_fd_sc_hd__decap_3 PHY_103 ();
 sky130_fd_sc_hd__decap_3 PHY_104 ();
 sky130_fd_sc_hd__decap_3 PHY_105 ();
 sky130_fd_sc_hd__decap_3 PHY_106 ();
 sky130_fd_sc_hd__decap_3 PHY_107 ();
 sky130_fd_sc_hd__decap_3 PHY_108 ();
 sky130_fd_sc_hd__decap_3 PHY_109 ();
 sky130_fd_sc_hd__decap_3 PHY_110 ();
 sky130_fd_sc_hd__decap_3 PHY_111 ();
 sky130_fd_sc_hd__decap_3 PHY_112 ();
 sky130_fd_sc_hd__decap_3 PHY_113 ();
 sky130_fd_sc_hd__decap_3 PHY_114 ();
 sky130_fd_sc_hd__decap_3 PHY_115 ();
 sky130_fd_sc_hd__decap_3 PHY_116 ();
 sky130_fd_sc_hd__decap_3 PHY_117 ();
 sky130_fd_sc_hd__decap_3 PHY_118 ();
 sky130_fd_sc_hd__decap_3 PHY_119 ();
 sky130_fd_sc_hd__decap_3 PHY_120 ();
 sky130_fd_sc_hd__decap_3 PHY_121 ();
 sky130_fd_sc_hd__decap_3 PHY_122 ();
 sky130_fd_sc_hd__decap_3 PHY_123 ();
 sky130_fd_sc_hd__decap_3 PHY_124 ();
 sky130_fd_sc_hd__decap_3 PHY_125 ();
 sky130_fd_sc_hd__decap_3 PHY_126 ();
 sky130_fd_sc_hd__decap_3 PHY_127 ();
 sky130_fd_sc_hd__decap_3 PHY_128 ();
 sky130_fd_sc_hd__decap_3 PHY_129 ();
 sky130_fd_sc_hd__decap_3 PHY_130 ();
 sky130_fd_sc_hd__decap_3 PHY_131 ();
 sky130_fd_sc_hd__decap_3 PHY_132 ();
 sky130_fd_sc_hd__decap_3 PHY_133 ();
 sky130_fd_sc_hd__decap_3 PHY_134 ();
 sky130_fd_sc_hd__decap_3 PHY_135 ();
 sky130_fd_sc_hd__decap_3 PHY_136 ();
 sky130_fd_sc_hd__decap_3 PHY_137 ();
 sky130_fd_sc_hd__decap_3 PHY_138 ();
 sky130_fd_sc_hd__decap_3 PHY_139 ();
 sky130_fd_sc_hd__decap_3 PHY_140 ();
 sky130_fd_sc_hd__decap_3 PHY_141 ();
 sky130_fd_sc_hd__decap_3 PHY_142 ();
 sky130_fd_sc_hd__decap_3 PHY_143 ();
 sky130_fd_sc_hd__decap_3 PHY_144 ();
 sky130_fd_sc_hd__decap_3 PHY_145 ();
 sky130_fd_sc_hd__decap_3 PHY_146 ();
 sky130_fd_sc_hd__decap_3 PHY_147 ();
 sky130_fd_sc_hd__decap_3 PHY_148 ();
 sky130_fd_sc_hd__decap_3 PHY_149 ();
 sky130_fd_sc_hd__decap_3 PHY_150 ();
 sky130_fd_sc_hd__decap_3 PHY_151 ();
 sky130_fd_sc_hd__decap_3 PHY_152 ();
 sky130_fd_sc_hd__decap_3 PHY_153 ();
 sky130_fd_sc_hd__decap_3 PHY_154 ();
 sky130_fd_sc_hd__decap_3 PHY_155 ();
 sky130_fd_sc_hd__decap_3 PHY_156 ();
 sky130_fd_sc_hd__decap_3 PHY_157 ();
 sky130_fd_sc_hd__decap_3 PHY_158 ();
 sky130_fd_sc_hd__decap_3 PHY_159 ();
 sky130_fd_sc_hd__decap_3 PHY_160 ();
 sky130_fd_sc_hd__decap_3 PHY_161 ();
 sky130_fd_sc_hd__decap_3 PHY_162 ();
 sky130_fd_sc_hd__decap_3 PHY_163 ();
 sky130_fd_sc_hd__decap_3 PHY_164 ();
 sky130_fd_sc_hd__decap_3 PHY_165 ();
 sky130_fd_sc_hd__decap_3 PHY_166 ();
 sky130_fd_sc_hd__decap_3 PHY_167 ();
 sky130_fd_sc_hd__decap_3 PHY_168 ();
 sky130_fd_sc_hd__decap_3 PHY_169 ();
 sky130_fd_sc_hd__decap_3 PHY_170 ();
 sky130_fd_sc_hd__decap_3 PHY_171 ();
 sky130_fd_sc_hd__decap_3 PHY_172 ();
 sky130_fd_sc_hd__decap_3 PHY_173 ();
 sky130_fd_sc_hd__decap_3 PHY_174 ();
 sky130_fd_sc_hd__decap_3 PHY_175 ();
 sky130_fd_sc_hd__decap_3 PHY_176 ();
 sky130_fd_sc_hd__decap_3 PHY_177 ();
 sky130_fd_sc_hd__decap_3 PHY_178 ();
 sky130_fd_sc_hd__decap_3 PHY_179 ();
 sky130_fd_sc_hd__decap_3 PHY_180 ();
 sky130_fd_sc_hd__decap_3 PHY_181 ();
 sky130_fd_sc_hd__decap_3 PHY_182 ();
 sky130_fd_sc_hd__decap_3 PHY_183 ();
 sky130_fd_sc_hd__decap_3 PHY_184 ();
 sky130_fd_sc_hd__decap_3 PHY_185 ();
 sky130_fd_sc_hd__decap_3 PHY_186 ();
 sky130_fd_sc_hd__decap_3 PHY_187 ();
 sky130_fd_sc_hd__decap_3 PHY_188 ();
 sky130_fd_sc_hd__decap_3 PHY_189 ();
 sky130_fd_sc_hd__decap_3 PHY_190 ();
 sky130_fd_sc_hd__decap_3 PHY_191 ();
 sky130_fd_sc_hd__decap_3 PHY_192 ();
 sky130_fd_sc_hd__decap_3 PHY_193 ();
 sky130_fd_sc_hd__decap_3 PHY_194 ();
 sky130_fd_sc_hd__decap_3 PHY_195 ();
 sky130_fd_sc_hd__decap_3 PHY_196 ();
 sky130_fd_sc_hd__decap_3 PHY_197 ();
 sky130_fd_sc_hd__decap_3 PHY_198 ();
 sky130_fd_sc_hd__decap_3 PHY_199 ();
 sky130_fd_sc_hd__decap_3 PHY_200 ();
 sky130_fd_sc_hd__decap_3 PHY_201 ();
 sky130_fd_sc_hd__decap_3 PHY_202 ();
 sky130_fd_sc_hd__decap_3 PHY_203 ();
 sky130_fd_sc_hd__decap_3 PHY_204 ();
 sky130_fd_sc_hd__decap_3 PHY_205 ();
 sky130_fd_sc_hd__decap_3 PHY_206 ();
 sky130_fd_sc_hd__decap_3 PHY_207 ();
 sky130_fd_sc_hd__decap_3 PHY_208 ();
 sky130_fd_sc_hd__decap_3 PHY_209 ();
 sky130_fd_sc_hd__decap_3 PHY_210 ();
 sky130_fd_sc_hd__decap_3 PHY_211 ();
 sky130_fd_sc_hd__decap_3 PHY_212 ();
 sky130_fd_sc_hd__decap_3 PHY_213 ();
 sky130_fd_sc_hd__decap_3 PHY_214 ();
 sky130_fd_sc_hd__decap_3 PHY_215 ();
 sky130_fd_sc_hd__decap_3 PHY_216 ();
 sky130_fd_sc_hd__decap_3 PHY_217 ();
 sky130_fd_sc_hd__decap_3 PHY_218 ();
 sky130_fd_sc_hd__decap_3 PHY_219 ();
 sky130_fd_sc_hd__decap_3 PHY_220 ();
 sky130_fd_sc_hd__decap_3 PHY_221 ();
 sky130_fd_sc_hd__decap_3 PHY_222 ();
 sky130_fd_sc_hd__decap_3 PHY_223 ();
 sky130_fd_sc_hd__decap_3 PHY_224 ();
 sky130_fd_sc_hd__decap_3 PHY_225 ();
 sky130_fd_sc_hd__decap_3 PHY_226 ();
 sky130_fd_sc_hd__decap_3 PHY_227 ();
 sky130_fd_sc_hd__decap_3 PHY_228 ();
 sky130_fd_sc_hd__decap_3 PHY_229 ();
 sky130_fd_sc_hd__decap_3 PHY_230 ();
 sky130_fd_sc_hd__decap_3 PHY_231 ();
 sky130_fd_sc_hd__decap_3 PHY_232 ();
 sky130_fd_sc_hd__decap_3 PHY_233 ();
 sky130_fd_sc_hd__decap_3 PHY_234 ();
 sky130_fd_sc_hd__decap_3 PHY_235 ();
 sky130_fd_sc_hd__decap_3 PHY_236 ();
 sky130_fd_sc_hd__decap_3 PHY_237 ();
 sky130_fd_sc_hd__decap_3 PHY_238 ();
 sky130_fd_sc_hd__decap_3 PHY_239 ();
 sky130_fd_sc_hd__decap_3 PHY_240 ();
 sky130_fd_sc_hd__decap_3 PHY_241 ();
 sky130_fd_sc_hd__decap_3 PHY_242 ();
 sky130_fd_sc_hd__decap_3 PHY_243 ();
 sky130_fd_sc_hd__decap_3 PHY_244 ();
 sky130_fd_sc_hd__decap_3 PHY_245 ();
 sky130_fd_sc_hd__decap_3 PHY_246 ();
 sky130_fd_sc_hd__decap_3 PHY_247 ();
 sky130_fd_sc_hd__decap_3 PHY_248 ();
 sky130_fd_sc_hd__decap_3 PHY_249 ();
 sky130_fd_sc_hd__decap_3 PHY_250 ();
 sky130_fd_sc_hd__decap_3 PHY_251 ();
 sky130_fd_sc_hd__decap_3 PHY_252 ();
 sky130_fd_sc_hd__decap_3 PHY_253 ();
 sky130_fd_sc_hd__decap_3 PHY_254 ();
 sky130_fd_sc_hd__decap_3 PHY_255 ();
 sky130_fd_sc_hd__decap_3 PHY_256 ();
 sky130_fd_sc_hd__decap_3 PHY_257 ();
 sky130_fd_sc_hd__decap_3 PHY_258 ();
 sky130_fd_sc_hd__decap_3 PHY_259 ();
 sky130_fd_sc_hd__decap_3 PHY_260 ();
 sky130_fd_sc_hd__decap_3 PHY_261 ();
 sky130_fd_sc_hd__decap_3 PHY_262 ();
 sky130_fd_sc_hd__decap_3 PHY_263 ();
 sky130_fd_sc_hd__decap_3 PHY_264 ();
 sky130_fd_sc_hd__decap_3 PHY_265 ();
 sky130_fd_sc_hd__decap_3 PHY_266 ();
 sky130_fd_sc_hd__decap_3 PHY_267 ();
 sky130_fd_sc_hd__decap_3 PHY_268 ();
 sky130_fd_sc_hd__decap_3 PHY_269 ();
 sky130_fd_sc_hd__decap_3 PHY_270 ();
 sky130_fd_sc_hd__decap_3 PHY_271 ();
 sky130_fd_sc_hd__decap_3 PHY_272 ();
 sky130_fd_sc_hd__decap_3 PHY_273 ();
 sky130_fd_sc_hd__decap_3 PHY_274 ();
 sky130_fd_sc_hd__decap_3 PHY_275 ();
 sky130_fd_sc_hd__decap_3 PHY_276 ();
 sky130_fd_sc_hd__decap_3 PHY_277 ();
 sky130_fd_sc_hd__decap_3 PHY_278 ();
 sky130_fd_sc_hd__decap_3 PHY_279 ();
 sky130_fd_sc_hd__decap_3 PHY_280 ();
 sky130_fd_sc_hd__decap_3 PHY_281 ();
 sky130_fd_sc_hd__decap_3 PHY_282 ();
 sky130_fd_sc_hd__decap_3 PHY_283 ();
 sky130_fd_sc_hd__decap_3 PHY_284 ();
 sky130_fd_sc_hd__decap_3 PHY_285 ();
 sky130_fd_sc_hd__decap_3 PHY_286 ();
 sky130_fd_sc_hd__decap_3 PHY_287 ();
 sky130_fd_sc_hd__decap_3 PHY_288 ();
 sky130_fd_sc_hd__decap_3 PHY_289 ();
 sky130_fd_sc_hd__decap_3 PHY_290 ();
 sky130_fd_sc_hd__decap_3 PHY_291 ();
 sky130_fd_sc_hd__decap_3 PHY_292 ();
 sky130_fd_sc_hd__decap_3 PHY_293 ();
 sky130_fd_sc_hd__decap_3 PHY_294 ();
 sky130_fd_sc_hd__decap_3 PHY_295 ();
 sky130_fd_sc_hd__decap_3 PHY_296 ();
 sky130_fd_sc_hd__decap_3 PHY_297 ();
 sky130_fd_sc_hd__decap_3 PHY_298 ();
 sky130_fd_sc_hd__decap_3 PHY_299 ();
 sky130_fd_sc_hd__decap_3 PHY_300 ();
 sky130_fd_sc_hd__decap_3 PHY_301 ();
 sky130_fd_sc_hd__decap_3 PHY_302 ();
 sky130_fd_sc_hd__decap_3 PHY_303 ();
 sky130_fd_sc_hd__decap_3 PHY_304 ();
 sky130_fd_sc_hd__decap_3 PHY_305 ();
 sky130_fd_sc_hd__decap_3 PHY_306 ();
 sky130_fd_sc_hd__decap_3 PHY_307 ();
 sky130_fd_sc_hd__decap_3 PHY_308 ();
 sky130_fd_sc_hd__decap_3 PHY_309 ();
 sky130_fd_sc_hd__decap_3 PHY_310 ();
 sky130_fd_sc_hd__decap_3 PHY_311 ();
 sky130_fd_sc_hd__decap_3 PHY_312 ();
 sky130_fd_sc_hd__decap_3 PHY_313 ();
 sky130_fd_sc_hd__decap_3 PHY_314 ();
 sky130_fd_sc_hd__decap_3 PHY_315 ();
 sky130_fd_sc_hd__decap_3 PHY_316 ();
 sky130_fd_sc_hd__decap_3 PHY_317 ();
 sky130_fd_sc_hd__decap_3 PHY_318 ();
 sky130_fd_sc_hd__decap_3 PHY_319 ();
 sky130_fd_sc_hd__decap_3 PHY_320 ();
 sky130_fd_sc_hd__decap_3 PHY_321 ();
 sky130_fd_sc_hd__decap_3 PHY_322 ();
 sky130_fd_sc_hd__decap_3 PHY_323 ();
 sky130_fd_sc_hd__decap_3 PHY_324 ();
 sky130_fd_sc_hd__decap_3 PHY_325 ();
 sky130_fd_sc_hd__decap_3 PHY_326 ();
 sky130_fd_sc_hd__decap_3 PHY_327 ();
 sky130_fd_sc_hd__decap_3 PHY_328 ();
 sky130_fd_sc_hd__decap_3 PHY_329 ();
 sky130_fd_sc_hd__decap_3 PHY_330 ();
 sky130_fd_sc_hd__decap_3 PHY_331 ();
 sky130_fd_sc_hd__decap_3 PHY_332 ();
 sky130_fd_sc_hd__decap_3 PHY_333 ();
 sky130_fd_sc_hd__decap_3 PHY_334 ();
 sky130_fd_sc_hd__decap_3 PHY_335 ();
 sky130_fd_sc_hd__decap_3 PHY_336 ();
 sky130_fd_sc_hd__decap_3 PHY_337 ();
 sky130_fd_sc_hd__decap_3 PHY_338 ();
 sky130_fd_sc_hd__decap_3 PHY_339 ();
 sky130_fd_sc_hd__decap_3 PHY_340 ();
 sky130_fd_sc_hd__decap_3 PHY_341 ();
 sky130_fd_sc_hd__decap_3 PHY_342 ();
 sky130_fd_sc_hd__decap_3 PHY_343 ();
 sky130_fd_sc_hd__decap_3 PHY_344 ();
 sky130_fd_sc_hd__decap_3 PHY_345 ();
 sky130_fd_sc_hd__decap_3 PHY_346 ();
 sky130_fd_sc_hd__decap_3 PHY_347 ();
 sky130_fd_sc_hd__decap_3 PHY_348 ();
 sky130_fd_sc_hd__decap_3 PHY_349 ();
 sky130_fd_sc_hd__decap_3 PHY_350 ();
 sky130_fd_sc_hd__decap_3 PHY_351 ();
 sky130_fd_sc_hd__decap_3 PHY_352 ();
 sky130_fd_sc_hd__decap_3 PHY_353 ();
 sky130_fd_sc_hd__decap_3 PHY_354 ();
 sky130_fd_sc_hd__decap_3 PHY_355 ();
 sky130_fd_sc_hd__decap_3 PHY_356 ();
 sky130_fd_sc_hd__decap_3 PHY_357 ();
 sky130_fd_sc_hd__decap_3 PHY_358 ();
 sky130_fd_sc_hd__decap_3 PHY_359 ();
 sky130_fd_sc_hd__decap_3 PHY_360 ();
 sky130_fd_sc_hd__decap_3 PHY_361 ();
 sky130_fd_sc_hd__decap_3 PHY_362 ();
 sky130_fd_sc_hd__decap_3 PHY_363 ();
 sky130_fd_sc_hd__decap_3 PHY_364 ();
 sky130_fd_sc_hd__decap_3 PHY_365 ();
 sky130_fd_sc_hd__decap_3 PHY_366 ();
 sky130_fd_sc_hd__decap_3 PHY_367 ();
 sky130_fd_sc_hd__decap_3 PHY_368 ();
 sky130_fd_sc_hd__decap_3 PHY_369 ();
 sky130_fd_sc_hd__decap_3 PHY_370 ();
 sky130_fd_sc_hd__decap_3 PHY_371 ();
 sky130_fd_sc_hd__decap_3 PHY_372 ();
 sky130_fd_sc_hd__decap_3 PHY_373 ();
 sky130_fd_sc_hd__decap_3 PHY_374 ();
 sky130_fd_sc_hd__decap_3 PHY_375 ();
 sky130_fd_sc_hd__decap_3 PHY_376 ();
 sky130_fd_sc_hd__decap_3 PHY_377 ();
 sky130_fd_sc_hd__decap_3 PHY_378 ();
 sky130_fd_sc_hd__decap_3 PHY_379 ();
 sky130_fd_sc_hd__decap_3 PHY_380 ();
 sky130_fd_sc_hd__decap_3 PHY_381 ();
 sky130_fd_sc_hd__decap_3 PHY_382 ();
 sky130_fd_sc_hd__decap_3 PHY_383 ();
 sky130_fd_sc_hd__decap_3 PHY_384 ();
 sky130_fd_sc_hd__decap_3 PHY_385 ();
 sky130_fd_sc_hd__decap_3 PHY_386 ();
 sky130_fd_sc_hd__decap_3 PHY_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3033 ();
 sky130_fd_sc_hd__clkbuf_1 input99 (.A(sram_ro_data[15]),
    .X(net99));
 sky130_fd_sc_hd__dlymetal6s2s_1 input98 (.A(sram_ro_data[14]),
    .X(net98));
 sky130_fd_sc_hd__clkbuf_1 input97 (.A(sram_ro_data[13]),
    .X(net97));
 sky130_fd_sc_hd__dlymetal6s2s_1 input96 (.A(sram_ro_data[12]),
    .X(net96));
 sky130_fd_sc_hd__clkbuf_2 input95 (.A(sram_ro_data[11]),
    .X(net95));
 sky130_fd_sc_hd__clkbuf_2 input94 (.A(sram_ro_data[10]),
    .X(net94));
 sky130_fd_sc_hd__clkbuf_2 input93 (.A(sram_ro_data[0]),
    .X(net93));
 sky130_fd_sc_hd__clkbuf_2 input92 (.A(spimemio_flash_io3_oeb),
    .X(net92));
 sky130_fd_sc_hd__dlymetal6s2s_1 input91 (.A(spimemio_flash_io3_do),
    .X(net91));
 sky130_fd_sc_hd__clkbuf_2 input90 (.A(spimemio_flash_io2_oeb),
    .X(net90));
 sky130_fd_sc_hd__dlymetal6s2s_1 input89 (.A(spimemio_flash_io2_do),
    .X(net89));
 sky130_fd_sc_hd__buf_2 input88 (.A(spimemio_flash_io1_oeb),
    .X(net88));
 sky130_fd_sc_hd__clkbuf_4 input87 (.A(spimemio_flash_io1_do),
    .X(net87));
 sky130_fd_sc_hd__buf_2 input86 (.A(spimemio_flash_io0_oeb),
    .X(net86));
 sky130_fd_sc_hd__buf_2 input85 (.A(spimemio_flash_io0_do),
    .X(net85));
 sky130_fd_sc_hd__buf_2 input84 (.A(spimemio_flash_csb),
    .X(net84));
 sky130_fd_sc_hd__buf_2 input83 (.A(spimemio_flash_clk),
    .X(net83));
 sky130_fd_sc_hd__clkbuf_1 input82 (.A(spi_sdoenb),
    .X(net82));
 sky130_fd_sc_hd__clkbuf_1 input81 (.A(spi_sdo),
    .X(net81));
 sky130_fd_sc_hd__clkbuf_1 input80 (.A(spi_sck),
    .X(net80));
 sky130_fd_sc_hd__clkbuf_4 input79 (.A(spi_enabled),
    .X(net79));
 sky130_fd_sc_hd__clkbuf_1 input78 (.A(spi_csb),
    .X(net78));
 sky130_fd_sc_hd__clkbuf_1 input77 (.A(ser_tx),
    .X(net77));
 sky130_fd_sc_hd__buf_4 input76 (.A(qspi_enabled),
    .X(net76));
 sky130_fd_sc_hd__buf_2 input75 (.A(porb),
    .X(net75));
 sky130_fd_sc_hd__clkbuf_1 input74 (.A(pad_flash_io1_di),
    .X(net74));
 sky130_fd_sc_hd__dlymetal6s2s_1 input73 (.A(pad_flash_io0_di),
    .X(net73));
 sky130_fd_sc_hd__clkbuf_1 input72 (.A(mgmt_gpio_in[9]),
    .X(net72));
 sky130_fd_sc_hd__dlymetal6s2s_1 input71 (.A(mgmt_gpio_in[8]),
    .X(net71));
 sky130_fd_sc_hd__buf_2 input70 (.A(mgmt_gpio_in[7]),
    .X(net70));
 sky130_fd_sc_hd__buf_2 input69 (.A(mgmt_gpio_in[6]),
    .X(net69));
 sky130_fd_sc_hd__clkbuf_4 input68 (.A(mgmt_gpio_in[5]),
    .X(net68));
 sky130_fd_sc_hd__buf_6 input67 (.A(mgmt_gpio_in[3]),
    .X(net67));
 sky130_fd_sc_hd__buf_4 input66 (.A(mgmt_gpio_in[37]),
    .X(net66));
 sky130_fd_sc_hd__buf_4 input65 (.A(mgmt_gpio_in[36]),
    .X(net65));
 sky130_fd_sc_hd__clkbuf_4 input64 (.A(mgmt_gpio_in[35]),
    .X(net64));
 sky130_fd_sc_hd__buf_4 input63 (.A(mgmt_gpio_in[34]),
    .X(net63));
 sky130_fd_sc_hd__clkbuf_2 input62 (.A(mgmt_gpio_in[33]),
    .X(net62));
 sky130_fd_sc_hd__clkbuf_2 input61 (.A(mgmt_gpio_in[32]),
    .X(net61));
 sky130_fd_sc_hd__buf_4 input60 (.A(mgmt_gpio_in[31]),
    .X(net60));
 sky130_fd_sc_hd__buf_4 input59 (.A(mgmt_gpio_in[30]),
    .X(net59));
 sky130_fd_sc_hd__clkbuf_4 input58 (.A(mgmt_gpio_in[2]),
    .X(net58));
 sky130_fd_sc_hd__buf_2 input57 (.A(mgmt_gpio_in[29]),
    .X(net57));
 sky130_fd_sc_hd__dlymetal6s2s_1 input56 (.A(mgmt_gpio_in[28]),
    .X(net56));
 sky130_fd_sc_hd__dlymetal6s2s_1 input55 (.A(mgmt_gpio_in[27]),
    .X(net55));
 sky130_fd_sc_hd__clkbuf_2 input54 (.A(mgmt_gpio_in[26]),
    .X(net54));
 sky130_fd_sc_hd__clkbuf_4 input53 (.A(mgmt_gpio_in[25]),
    .X(net53));
 sky130_fd_sc_hd__dlymetal6s2s_1 input52 (.A(mgmt_gpio_in[24]),
    .X(net52));
 sky130_fd_sc_hd__clkbuf_4 input51 (.A(mgmt_gpio_in[23]),
    .X(net51));
 sky130_fd_sc_hd__clkbuf_4 input50 (.A(mgmt_gpio_in[22]),
    .X(net50));
 sky130_fd_sc_hd__buf_2 input49 (.A(mgmt_gpio_in[21]),
    .X(net49));
 sky130_fd_sc_hd__clkbuf_2 input48 (.A(mgmt_gpio_in[20]),
    .X(net48));
 sky130_fd_sc_hd__buf_2 input47 (.A(mgmt_gpio_in[1]),
    .X(net47));
 sky130_fd_sc_hd__buf_2 input46 (.A(mgmt_gpio_in[19]),
    .X(net46));
 sky130_fd_sc_hd__buf_2 input45 (.A(mgmt_gpio_in[18]),
    .X(net45));
 sky130_fd_sc_hd__clkbuf_2 input44 (.A(mgmt_gpio_in[17]),
    .X(net44));
 sky130_fd_sc_hd__clkbuf_4 input43 (.A(mgmt_gpio_in[16]),
    .X(net43));
 sky130_fd_sc_hd__clkbuf_4 input42 (.A(mgmt_gpio_in[15]),
    .X(net42));
 sky130_fd_sc_hd__clkbuf_4 input41 (.A(mgmt_gpio_in[14]),
    .X(net41));
 sky130_fd_sc_hd__buf_2 input40 (.A(mgmt_gpio_in[13]),
    .X(net40));
 sky130_fd_sc_hd__clkbuf_8 input39 (.A(mgmt_gpio_in[12]),
    .X(net39));
 sky130_fd_sc_hd__clkbuf_4 input38 (.A(mgmt_gpio_in[11]),
    .X(net38));
 sky130_fd_sc_hd__clkbuf_1 input37 (.A(mgmt_gpio_in[10]),
    .X(net37));
 sky130_fd_sc_hd__clkbuf_4 input36 (.A(mgmt_gpio_in[0]),
    .X(net36));
 sky130_fd_sc_hd__clkbuf_1 input35 (.A(mask_rev_in[9]),
    .X(net35));
 sky130_fd_sc_hd__clkbuf_1 input34 (.A(mask_rev_in[8]),
    .X(net34));
 sky130_fd_sc_hd__clkbuf_2 input33 (.A(mask_rev_in[7]),
    .X(net33));
 sky130_fd_sc_hd__clkbuf_1 input32 (.A(mask_rev_in[6]),
    .X(net32));
 sky130_fd_sc_hd__dlymetal6s2s_1 input31 (.A(mask_rev_in[5]),
    .X(net31));
 sky130_fd_sc_hd__clkbuf_1 input30 (.A(mask_rev_in[4]),
    .X(net30));
 sky130_fd_sc_hd__clkbuf_2 input29 (.A(mask_rev_in[3]),
    .X(net29));
 sky130_fd_sc_hd__clkbuf_4 input28 (.A(mask_rev_in[31]),
    .X(net28));
 sky130_fd_sc_hd__dlymetal6s2s_1 input27 (.A(mask_rev_in[30]),
    .X(net27));
 sky130_fd_sc_hd__clkbuf_1 input26 (.A(mask_rev_in[2]),
    .X(net26));
 sky130_fd_sc_hd__clkbuf_2 input25 (.A(mask_rev_in[29]),
    .X(net25));
 sky130_fd_sc_hd__dlymetal6s2s_1 input24 (.A(mask_rev_in[28]),
    .X(net24));
 sky130_fd_sc_hd__clkbuf_1 input23 (.A(mask_rev_in[27]),
    .X(net23));
 sky130_fd_sc_hd__dlymetal6s2s_1 input22 (.A(mask_rev_in[26]),
    .X(net22));
 sky130_fd_sc_hd__clkbuf_4 input21 (.A(mask_rev_in[25]),
    .X(net21));
 sky130_fd_sc_hd__clkbuf_2 input20 (.A(mask_rev_in[24]),
    .X(net20));
 sky130_fd_sc_hd__clkbuf_2 input19 (.A(mask_rev_in[23]),
    .X(net19));
 sky130_fd_sc_hd__buf_2 input18 (.A(mask_rev_in[22]),
    .X(net18));
 sky130_fd_sc_hd__buf_2 input17 (.A(mask_rev_in[21]),
    .X(net17));
 sky130_fd_sc_hd__dlymetal6s2s_1 input16 (.A(mask_rev_in[20]),
    .X(net16));
 sky130_fd_sc_hd__clkbuf_2 input15 (.A(mask_rev_in[1]),
    .X(net15));
 sky130_fd_sc_hd__clkbuf_1 input14 (.A(mask_rev_in[19]),
    .X(net14));
 sky130_fd_sc_hd__clkbuf_1 input13 (.A(mask_rev_in[18]),
    .X(net13));
 sky130_fd_sc_hd__clkbuf_1 input12 (.A(mask_rev_in[17]),
    .X(net12));
 sky130_fd_sc_hd__clkbuf_1 input11 (.A(mask_rev_in[16]),
    .X(net11));
 sky130_fd_sc_hd__clkbuf_2 input10 (.A(mask_rev_in[15]),
    .X(net10));
 sky130_fd_sc_hd__clkbuf_2 input9 (.A(mask_rev_in[14]),
    .X(net9));
 sky130_fd_sc_hd__dlymetal6s2s_1 input8 (.A(mask_rev_in[13]),
    .X(net8));
 sky130_fd_sc_hd__clkbuf_1 input7 (.A(mask_rev_in[12]),
    .X(net7));
 sky130_fd_sc_hd__clkbuf_1 input6 (.A(mask_rev_in[11]),
    .X(net6));
 sky130_fd_sc_hd__clkbuf_1 input5 (.A(mask_rev_in[10]),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_1 input4 (.A(mask_rev_in[0]),
    .X(net4));
 sky130_fd_sc_hd__clkbuf_1 input3 (.A(debug_out),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_1 input2 (.A(debug_oeb),
    .X(net2));
 sky130_fd_sc_hd__dlymetal6s2s_1 input1 (.A(debug_mode),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_1 input100 (.A(sram_ro_data[16]),
    .X(net100));
 sky130_fd_sc_hd__dlymetal6s2s_1 input101 (.A(sram_ro_data[17]),
    .X(net101));
 sky130_fd_sc_hd__buf_2 input102 (.A(sram_ro_data[18]),
    .X(net102));
 sky130_fd_sc_hd__clkbuf_2 input103 (.A(sram_ro_data[19]),
    .X(net103));
 sky130_fd_sc_hd__clkbuf_4 input104 (.A(sram_ro_data[1]),
    .X(net104));
 sky130_fd_sc_hd__clkbuf_2 input105 (.A(sram_ro_data[20]),
    .X(net105));
 sky130_fd_sc_hd__clkbuf_1 input106 (.A(sram_ro_data[21]),
    .X(net106));
 sky130_fd_sc_hd__clkbuf_1 input107 (.A(sram_ro_data[22]),
    .X(net107));
 sky130_fd_sc_hd__clkbuf_1 input108 (.A(sram_ro_data[23]),
    .X(net108));
 sky130_fd_sc_hd__clkbuf_2 input109 (.A(sram_ro_data[24]),
    .X(net109));
 sky130_fd_sc_hd__buf_2 input110 (.A(sram_ro_data[25]),
    .X(net110));
 sky130_fd_sc_hd__clkbuf_2 input111 (.A(sram_ro_data[26]),
    .X(net111));
 sky130_fd_sc_hd__clkbuf_2 input112 (.A(sram_ro_data[27]),
    .X(net112));
 sky130_fd_sc_hd__clkbuf_2 input113 (.A(sram_ro_data[28]),
    .X(net113));
 sky130_fd_sc_hd__clkbuf_2 input114 (.A(sram_ro_data[29]),
    .X(net114));
 sky130_fd_sc_hd__clkbuf_2 input115 (.A(sram_ro_data[2]),
    .X(net115));
 sky130_fd_sc_hd__dlymetal6s2s_1 input116 (.A(sram_ro_data[30]),
    .X(net116));
 sky130_fd_sc_hd__clkbuf_1 input117 (.A(sram_ro_data[31]),
    .X(net117));
 sky130_fd_sc_hd__clkbuf_2 input118 (.A(sram_ro_data[3]),
    .X(net118));
 sky130_fd_sc_hd__clkbuf_2 input119 (.A(sram_ro_data[4]),
    .X(net119));
 sky130_fd_sc_hd__clkbuf_1 input120 (.A(sram_ro_data[5]),
    .X(net120));
 sky130_fd_sc_hd__clkbuf_1 input121 (.A(sram_ro_data[6]),
    .X(net121));
 sky130_fd_sc_hd__clkbuf_1 input122 (.A(sram_ro_data[7]),
    .X(net122));
 sky130_fd_sc_hd__clkbuf_2 input123 (.A(sram_ro_data[8]),
    .X(net123));
 sky130_fd_sc_hd__clkbuf_2 input124 (.A(sram_ro_data[9]),
    .X(net124));
 sky130_fd_sc_hd__buf_4 input125 (.A(trap),
    .X(net125));
 sky130_fd_sc_hd__clkbuf_1 input126 (.A(uart_enabled),
    .X(net126));
 sky130_fd_sc_hd__clkbuf_2 input127 (.A(usr1_vcc_pwrgood),
    .X(net127));
 sky130_fd_sc_hd__clkbuf_2 input128 (.A(usr1_vdd_pwrgood),
    .X(net128));
 sky130_fd_sc_hd__clkbuf_4 input129 (.A(usr2_vcc_pwrgood),
    .X(net129));
 sky130_fd_sc_hd__clkbuf_4 input130 (.A(usr2_vdd_pwrgood),
    .X(net130));
 sky130_fd_sc_hd__clkbuf_4 input131 (.A(wb_adr_i[0]),
    .X(net131));
 sky130_fd_sc_hd__clkbuf_1 input132 (.A(wb_adr_i[10]),
    .X(net132));
 sky130_fd_sc_hd__clkbuf_1 input133 (.A(wb_adr_i[11]),
    .X(net133));
 sky130_fd_sc_hd__clkbuf_1 input134 (.A(wb_adr_i[12]),
    .X(net134));
 sky130_fd_sc_hd__clkbuf_1 input135 (.A(wb_adr_i[13]),
    .X(net135));
 sky130_fd_sc_hd__clkbuf_1 input136 (.A(wb_adr_i[14]),
    .X(net136));
 sky130_fd_sc_hd__clkbuf_1 input137 (.A(wb_adr_i[15]),
    .X(net137));
 sky130_fd_sc_hd__clkbuf_1 input138 (.A(wb_adr_i[16]),
    .X(net138));
 sky130_fd_sc_hd__clkbuf_1 input139 (.A(wb_adr_i[17]),
    .X(net139));
 sky130_fd_sc_hd__clkbuf_1 input140 (.A(wb_adr_i[18]),
    .X(net140));
 sky130_fd_sc_hd__clkbuf_1 input141 (.A(wb_adr_i[19]),
    .X(net141));
 sky130_fd_sc_hd__clkbuf_2 input142 (.A(wb_adr_i[1]),
    .X(net142));
 sky130_fd_sc_hd__clkbuf_1 input143 (.A(wb_adr_i[20]),
    .X(net143));
 sky130_fd_sc_hd__clkbuf_2 input144 (.A(wb_adr_i[21]),
    .X(net144));
 sky130_fd_sc_hd__clkbuf_1 input145 (.A(wb_adr_i[22]),
    .X(net145));
 sky130_fd_sc_hd__clkbuf_1 input146 (.A(wb_adr_i[23]),
    .X(net146));
 sky130_fd_sc_hd__clkbuf_1 input147 (.A(wb_adr_i[24]),
    .X(net147));
 sky130_fd_sc_hd__clkbuf_1 input148 (.A(wb_adr_i[25]),
    .X(net148));
 sky130_fd_sc_hd__clkbuf_1 input149 (.A(wb_adr_i[26]),
    .X(net149));
 sky130_fd_sc_hd__clkbuf_1 input150 (.A(wb_adr_i[27]),
    .X(net150));
 sky130_fd_sc_hd__clkbuf_1 input151 (.A(wb_adr_i[28]),
    .X(net151));
 sky130_fd_sc_hd__clkbuf_1 input152 (.A(wb_adr_i[29]),
    .X(net152));
 sky130_fd_sc_hd__dlymetal6s2s_1 input153 (.A(wb_adr_i[2]),
    .X(net153));
 sky130_fd_sc_hd__clkbuf_1 input154 (.A(wb_adr_i[30]),
    .X(net154));
 sky130_fd_sc_hd__clkbuf_1 input155 (.A(wb_adr_i[31]),
    .X(net155));
 sky130_fd_sc_hd__clkbuf_4 input156 (.A(wb_adr_i[3]),
    .X(net156));
 sky130_fd_sc_hd__buf_4 input157 (.A(wb_adr_i[4]),
    .X(net157));
 sky130_fd_sc_hd__buf_2 input158 (.A(wb_adr_i[5]),
    .X(net158));
 sky130_fd_sc_hd__clkbuf_1 input159 (.A(wb_adr_i[6]),
    .X(net159));
 sky130_fd_sc_hd__buf_2 input160 (.A(wb_adr_i[7]),
    .X(net160));
 sky130_fd_sc_hd__clkbuf_1 input161 (.A(wb_adr_i[8]),
    .X(net161));
 sky130_fd_sc_hd__clkbuf_1 input162 (.A(wb_adr_i[9]),
    .X(net162));
 sky130_fd_sc_hd__clkbuf_1 input163 (.A(wb_cyc_i),
    .X(net163));
 sky130_fd_sc_hd__clkbuf_1 input164 (.A(wb_dat_i[0]),
    .X(net164));
 sky130_fd_sc_hd__clkbuf_1 input165 (.A(wb_dat_i[10]),
    .X(net165));
 sky130_fd_sc_hd__clkbuf_1 input166 (.A(wb_dat_i[11]),
    .X(net166));
 sky130_fd_sc_hd__clkbuf_1 input167 (.A(wb_dat_i[12]),
    .X(net167));
 sky130_fd_sc_hd__clkbuf_1 input168 (.A(wb_dat_i[13]),
    .X(net168));
 sky130_fd_sc_hd__clkbuf_1 input169 (.A(wb_dat_i[14]),
    .X(net169));
 sky130_fd_sc_hd__clkbuf_1 input170 (.A(wb_dat_i[15]),
    .X(net170));
 sky130_fd_sc_hd__clkbuf_1 input171 (.A(wb_dat_i[16]),
    .X(net171));
 sky130_fd_sc_hd__clkbuf_1 input172 (.A(wb_dat_i[17]),
    .X(net172));
 sky130_fd_sc_hd__clkbuf_1 input173 (.A(wb_dat_i[18]),
    .X(net173));
 sky130_fd_sc_hd__clkbuf_1 input174 (.A(wb_dat_i[19]),
    .X(net174));
 sky130_fd_sc_hd__clkbuf_1 input175 (.A(wb_dat_i[1]),
    .X(net175));
 sky130_fd_sc_hd__clkbuf_1 input176 (.A(wb_dat_i[20]),
    .X(net176));
 sky130_fd_sc_hd__clkbuf_1 input177 (.A(wb_dat_i[21]),
    .X(net177));
 sky130_fd_sc_hd__clkbuf_1 input178 (.A(wb_dat_i[22]),
    .X(net178));
 sky130_fd_sc_hd__clkbuf_1 input179 (.A(wb_dat_i[23]),
    .X(net179));
 sky130_fd_sc_hd__clkbuf_1 input180 (.A(wb_dat_i[24]),
    .X(net180));
 sky130_fd_sc_hd__clkbuf_1 input181 (.A(wb_dat_i[25]),
    .X(net181));
 sky130_fd_sc_hd__clkbuf_1 input182 (.A(wb_dat_i[26]),
    .X(net182));
 sky130_fd_sc_hd__clkbuf_1 input183 (.A(wb_dat_i[27]),
    .X(net183));
 sky130_fd_sc_hd__clkbuf_1 input184 (.A(wb_dat_i[28]),
    .X(net184));
 sky130_fd_sc_hd__clkbuf_1 input185 (.A(wb_dat_i[29]),
    .X(net185));
 sky130_fd_sc_hd__clkbuf_1 input186 (.A(wb_dat_i[2]),
    .X(net186));
 sky130_fd_sc_hd__clkbuf_1 input187 (.A(wb_dat_i[30]),
    .X(net187));
 sky130_fd_sc_hd__clkbuf_1 input188 (.A(wb_dat_i[31]),
    .X(net188));
 sky130_fd_sc_hd__clkbuf_1 input189 (.A(wb_dat_i[3]),
    .X(net189));
 sky130_fd_sc_hd__clkbuf_1 input190 (.A(wb_dat_i[4]),
    .X(net190));
 sky130_fd_sc_hd__clkbuf_1 input191 (.A(wb_dat_i[5]),
    .X(net191));
 sky130_fd_sc_hd__clkbuf_1 input192 (.A(wb_dat_i[6]),
    .X(net192));
 sky130_fd_sc_hd__clkbuf_1 input193 (.A(wb_dat_i[7]),
    .X(net193));
 sky130_fd_sc_hd__clkbuf_1 input194 (.A(wb_dat_i[8]),
    .X(net194));
 sky130_fd_sc_hd__clkbuf_1 input195 (.A(wb_dat_i[9]),
    .X(net195));
 sky130_fd_sc_hd__clkbuf_2 input196 (.A(wb_rstn_i),
    .X(net196));
 sky130_fd_sc_hd__clkbuf_1 input197 (.A(wb_sel_i[0]),
    .X(net197));
 sky130_fd_sc_hd__clkbuf_1 input198 (.A(wb_sel_i[1]),
    .X(net198));
 sky130_fd_sc_hd__clkbuf_1 input199 (.A(wb_sel_i[2]),
    .X(net199));
 sky130_fd_sc_hd__clkbuf_1 input200 (.A(wb_sel_i[3]),
    .X(net200));
 sky130_fd_sc_hd__buf_2 input201 (.A(wb_stb_i),
    .X(net201));
 sky130_fd_sc_hd__clkbuf_2 input202 (.A(wb_we_i),
    .X(net202));
 sky130_fd_sc_hd__buf_12 output203 (.A(net203),
    .X(debug_in));
 sky130_fd_sc_hd__buf_12 output204 (.A(net204),
    .X(irq[0]));
 sky130_fd_sc_hd__buf_12 output205 (.A(net205),
    .X(irq[1]));
 sky130_fd_sc_hd__buf_12 output206 (.A(net206),
    .X(irq[2]));
 sky130_fd_sc_hd__buf_12 output207 (.A(net207),
    .X(mgmt_gpio_oeb[0]));
 sky130_fd_sc_hd__buf_12 output208 (.A(net208),
    .X(mgmt_gpio_oeb[10]));
 sky130_fd_sc_hd__buf_12 output209 (.A(net209),
    .X(mgmt_gpio_oeb[11]));
 sky130_fd_sc_hd__buf_12 output210 (.A(net210),
    .X(mgmt_gpio_oeb[12]));
 sky130_fd_sc_hd__buf_12 output211 (.A(net211),
    .X(mgmt_gpio_oeb[13]));
 sky130_fd_sc_hd__buf_12 output212 (.A(net212),
    .X(mgmt_gpio_oeb[14]));
 sky130_fd_sc_hd__buf_12 output213 (.A(net213),
    .X(mgmt_gpio_oeb[15]));
 sky130_fd_sc_hd__buf_12 output214 (.A(net214),
    .X(mgmt_gpio_oeb[16]));
 sky130_fd_sc_hd__buf_12 output215 (.A(net215),
    .X(mgmt_gpio_oeb[17]));
 sky130_fd_sc_hd__buf_12 output216 (.A(net216),
    .X(mgmt_gpio_oeb[18]));
 sky130_fd_sc_hd__buf_12 output217 (.A(net217),
    .X(mgmt_gpio_oeb[19]));
 sky130_fd_sc_hd__buf_12 output218 (.A(net218),
    .X(mgmt_gpio_oeb[1]));
 sky130_fd_sc_hd__buf_12 output219 (.A(net219),
    .X(mgmt_gpio_oeb[20]));
 sky130_fd_sc_hd__buf_12 output220 (.A(net220),
    .X(mgmt_gpio_oeb[21]));
 sky130_fd_sc_hd__buf_12 output221 (.A(net221),
    .X(mgmt_gpio_oeb[22]));
 sky130_fd_sc_hd__buf_12 output222 (.A(net222),
    .X(mgmt_gpio_oeb[23]));
 sky130_fd_sc_hd__buf_12 output223 (.A(net223),
    .X(mgmt_gpio_oeb[24]));
 sky130_fd_sc_hd__buf_12 output224 (.A(net224),
    .X(mgmt_gpio_oeb[25]));
 sky130_fd_sc_hd__buf_12 output225 (.A(net225),
    .X(mgmt_gpio_oeb[26]));
 sky130_fd_sc_hd__buf_12 output226 (.A(net226),
    .X(mgmt_gpio_oeb[27]));
 sky130_fd_sc_hd__buf_12 output227 (.A(net227),
    .X(mgmt_gpio_oeb[28]));
 sky130_fd_sc_hd__buf_12 output228 (.A(net228),
    .X(mgmt_gpio_oeb[29]));
 sky130_fd_sc_hd__buf_12 output229 (.A(net229),
    .X(mgmt_gpio_oeb[2]));
 sky130_fd_sc_hd__buf_12 output230 (.A(net230),
    .X(mgmt_gpio_oeb[30]));
 sky130_fd_sc_hd__buf_12 output231 (.A(net231),
    .X(mgmt_gpio_oeb[31]));
 sky130_fd_sc_hd__buf_12 output232 (.A(net232),
    .X(mgmt_gpio_oeb[32]));
 sky130_fd_sc_hd__buf_12 output233 (.A(net233),
    .X(mgmt_gpio_oeb[33]));
 sky130_fd_sc_hd__buf_12 output234 (.A(net234),
    .X(mgmt_gpio_oeb[34]));
 sky130_fd_sc_hd__buf_12 output235 (.A(net235),
    .X(mgmt_gpio_oeb[35]));
 sky130_fd_sc_hd__buf_12 output236 (.A(net236),
    .X(mgmt_gpio_oeb[36]));
 sky130_fd_sc_hd__buf_12 output237 (.A(net237),
    .X(mgmt_gpio_oeb[37]));
 sky130_fd_sc_hd__buf_12 output238 (.A(net238),
    .X(mgmt_gpio_oeb[3]));
 sky130_fd_sc_hd__buf_12 output239 (.A(net239),
    .X(mgmt_gpio_oeb[4]));
 sky130_fd_sc_hd__buf_12 output240 (.A(net240),
    .X(mgmt_gpio_oeb[5]));
 sky130_fd_sc_hd__buf_12 output241 (.A(net241),
    .X(mgmt_gpio_oeb[6]));
 sky130_fd_sc_hd__buf_12 output242 (.A(net242),
    .X(mgmt_gpio_oeb[7]));
 sky130_fd_sc_hd__buf_12 output243 (.A(net243),
    .X(mgmt_gpio_oeb[8]));
 sky130_fd_sc_hd__buf_12 output244 (.A(net244),
    .X(mgmt_gpio_oeb[9]));
 sky130_fd_sc_hd__buf_12 output245 (.A(net245),
    .X(mgmt_gpio_out[0]));
 sky130_fd_sc_hd__buf_12 output246 (.A(net246),
    .X(mgmt_gpio_out[1]));
 sky130_fd_sc_hd__buf_12 output247 (.A(net247),
    .X(mgmt_gpio_out[35]));
 sky130_fd_sc_hd__buf_12 output248 (.A(net248),
    .X(mgmt_gpio_out[36]));
 sky130_fd_sc_hd__buf_12 output249 (.A(net249),
    .X(mgmt_gpio_out[37]));
 sky130_fd_sc_hd__clkbuf_1 output250 (.A(net250),
    .X(pad_flash_clk));
 sky130_fd_sc_hd__buf_12 output251 (.A(net251),
    .X(pad_flash_clk_oeb));
 sky130_fd_sc_hd__buf_12 output252 (.A(net252),
    .X(pad_flash_csb));
 sky130_fd_sc_hd__buf_12 output253 (.A(net253),
    .X(pad_flash_csb_oeb));
 sky130_fd_sc_hd__buf_12 output254 (.A(net254),
    .X(pad_flash_io0_do));
 sky130_fd_sc_hd__buf_12 output255 (.A(net255),
    .X(pad_flash_io0_ieb));
 sky130_fd_sc_hd__buf_12 output256 (.A(net256),
    .X(pad_flash_io0_oeb));
 sky130_fd_sc_hd__buf_12 output257 (.A(net257),
    .X(pad_flash_io1_do));
 sky130_fd_sc_hd__buf_12 output258 (.A(net258),
    .X(pad_flash_io1_ieb));
 sky130_fd_sc_hd__buf_12 output259 (.A(net259),
    .X(pad_flash_io1_oeb));
 sky130_fd_sc_hd__buf_12 output260 (.A(net260),
    .X(pll90_sel[0]));
 sky130_fd_sc_hd__buf_12 output261 (.A(net261),
    .X(pll90_sel[1]));
 sky130_fd_sc_hd__buf_12 output262 (.A(net262),
    .X(pll90_sel[2]));
 sky130_fd_sc_hd__buf_12 output263 (.A(net263),
    .X(pll_bypass));
 sky130_fd_sc_hd__buf_12 output264 (.A(net264),
    .X(pll_dco_ena));
 sky130_fd_sc_hd__buf_12 output265 (.A(net265),
    .X(pll_div[0]));
 sky130_fd_sc_hd__buf_12 output266 (.A(net266),
    .X(pll_div[1]));
 sky130_fd_sc_hd__buf_12 output267 (.A(net267),
    .X(pll_div[2]));
 sky130_fd_sc_hd__buf_12 output268 (.A(net268),
    .X(pll_div[3]));
 sky130_fd_sc_hd__buf_12 output269 (.A(net269),
    .X(pll_div[4]));
 sky130_fd_sc_hd__buf_12 output270 (.A(net270),
    .X(pll_ena));
 sky130_fd_sc_hd__buf_12 output271 (.A(net271),
    .X(pll_sel[0]));
 sky130_fd_sc_hd__buf_12 output272 (.A(net272),
    .X(pll_sel[1]));
 sky130_fd_sc_hd__buf_12 output273 (.A(net273),
    .X(pll_sel[2]));
 sky130_fd_sc_hd__buf_12 output274 (.A(net274),
    .X(pll_trim[0]));
 sky130_fd_sc_hd__buf_12 output275 (.A(net275),
    .X(pll_trim[10]));
 sky130_fd_sc_hd__buf_12 output276 (.A(net276),
    .X(pll_trim[11]));
 sky130_fd_sc_hd__buf_12 output277 (.A(net277),
    .X(pll_trim[12]));
 sky130_fd_sc_hd__buf_12 output278 (.A(net278),
    .X(pll_trim[13]));
 sky130_fd_sc_hd__buf_12 output279 (.A(net279),
    .X(pll_trim[14]));
 sky130_fd_sc_hd__buf_12 output280 (.A(net280),
    .X(pll_trim[15]));
 sky130_fd_sc_hd__buf_12 output281 (.A(net281),
    .X(pll_trim[16]));
 sky130_fd_sc_hd__buf_12 output282 (.A(net282),
    .X(pll_trim[17]));
 sky130_fd_sc_hd__buf_12 output283 (.A(net283),
    .X(pll_trim[18]));
 sky130_fd_sc_hd__buf_12 output284 (.A(net284),
    .X(pll_trim[19]));
 sky130_fd_sc_hd__buf_12 output285 (.A(net285),
    .X(pll_trim[1]));
 sky130_fd_sc_hd__buf_12 output286 (.A(net286),
    .X(pll_trim[20]));
 sky130_fd_sc_hd__buf_12 output287 (.A(net287),
    .X(pll_trim[21]));
 sky130_fd_sc_hd__buf_12 output288 (.A(net288),
    .X(pll_trim[22]));
 sky130_fd_sc_hd__buf_12 output289 (.A(net289),
    .X(pll_trim[23]));
 sky130_fd_sc_hd__buf_12 output290 (.A(net290),
    .X(pll_trim[24]));
 sky130_fd_sc_hd__buf_12 output291 (.A(net291),
    .X(pll_trim[25]));
 sky130_fd_sc_hd__buf_12 output292 (.A(net292),
    .X(pll_trim[2]));
 sky130_fd_sc_hd__buf_12 output293 (.A(net293),
    .X(pll_trim[3]));
 sky130_fd_sc_hd__buf_12 output294 (.A(net294),
    .X(pll_trim[4]));
 sky130_fd_sc_hd__buf_12 output295 (.A(net295),
    .X(pll_trim[5]));
 sky130_fd_sc_hd__buf_12 output296 (.A(net296),
    .X(pll_trim[6]));
 sky130_fd_sc_hd__buf_12 output297 (.A(net297),
    .X(pll_trim[7]));
 sky130_fd_sc_hd__buf_12 output298 (.A(net298),
    .X(pll_trim[8]));
 sky130_fd_sc_hd__buf_12 output299 (.A(net299),
    .X(pll_trim[9]));
 sky130_fd_sc_hd__buf_12 output300 (.A(net300),
    .X(pwr_ctrl_out[0]));
 sky130_fd_sc_hd__buf_12 output301 (.A(net301),
    .X(pwr_ctrl_out[1]));
 sky130_fd_sc_hd__buf_12 output302 (.A(net302),
    .X(pwr_ctrl_out[2]));
 sky130_fd_sc_hd__buf_12 output303 (.A(net303),
    .X(pwr_ctrl_out[3]));
 sky130_fd_sc_hd__buf_12 output304 (.A(net304),
    .X(reset));
 sky130_fd_sc_hd__buf_12 output305 (.A(net305),
    .X(ser_rx));
 sky130_fd_sc_hd__buf_12 output306 (.A(net306),
    .X(serial_clock));
 sky130_fd_sc_hd__buf_12 output307 (.A(net307),
    .X(serial_data_1));
 sky130_fd_sc_hd__buf_12 output308 (.A(net308),
    .X(serial_data_2));
 sky130_fd_sc_hd__buf_12 output309 (.A(net309),
    .X(serial_load));
 sky130_fd_sc_hd__buf_12 output310 (.A(net310),
    .X(serial_resetn));
 sky130_fd_sc_hd__buf_12 output311 (.A(net311),
    .X(spi_sdi));
 sky130_fd_sc_hd__buf_12 output312 (.A(net312),
    .X(spimemio_flash_io0_di));
 sky130_fd_sc_hd__buf_12 output313 (.A(net313),
    .X(spimemio_flash_io1_di));
 sky130_fd_sc_hd__buf_12 output314 (.A(net314),
    .X(spimemio_flash_io2_di));
 sky130_fd_sc_hd__buf_12 output315 (.A(net315),
    .X(spimemio_flash_io3_di));
 sky130_fd_sc_hd__buf_12 output316 (.A(net316),
    .X(sram_ro_addr[0]));
 sky130_fd_sc_hd__buf_12 output317 (.A(net317),
    .X(sram_ro_addr[1]));
 sky130_fd_sc_hd__buf_12 output318 (.A(net318),
    .X(sram_ro_addr[2]));
 sky130_fd_sc_hd__buf_12 output319 (.A(net319),
    .X(sram_ro_addr[3]));
 sky130_fd_sc_hd__buf_12 output320 (.A(net320),
    .X(sram_ro_addr[4]));
 sky130_fd_sc_hd__buf_12 output321 (.A(net321),
    .X(sram_ro_addr[5]));
 sky130_fd_sc_hd__buf_12 output322 (.A(net322),
    .X(sram_ro_addr[6]));
 sky130_fd_sc_hd__buf_12 output323 (.A(net323),
    .X(sram_ro_addr[7]));
 sky130_fd_sc_hd__buf_12 output324 (.A(net324),
    .X(sram_ro_clk));
 sky130_fd_sc_hd__buf_12 output325 (.A(net325),
    .X(sram_ro_csb));
 sky130_fd_sc_hd__buf_12 output326 (.A(net326),
    .X(wb_ack_o));
 sky130_fd_sc_hd__buf_12 output327 (.A(net327),
    .X(wb_dat_o[0]));
 sky130_fd_sc_hd__buf_12 output328 (.A(net328),
    .X(wb_dat_o[10]));
 sky130_fd_sc_hd__buf_12 output329 (.A(net329),
    .X(wb_dat_o[11]));
 sky130_fd_sc_hd__buf_12 output330 (.A(net330),
    .X(wb_dat_o[12]));
 sky130_fd_sc_hd__buf_12 output331 (.A(net331),
    .X(wb_dat_o[13]));
 sky130_fd_sc_hd__buf_12 output332 (.A(net332),
    .X(wb_dat_o[14]));
 sky130_fd_sc_hd__buf_12 output333 (.A(net333),
    .X(wb_dat_o[15]));
 sky130_fd_sc_hd__buf_12 output334 (.A(net334),
    .X(wb_dat_o[16]));
 sky130_fd_sc_hd__buf_12 output335 (.A(net335),
    .X(wb_dat_o[17]));
 sky130_fd_sc_hd__buf_12 output336 (.A(net336),
    .X(wb_dat_o[18]));
 sky130_fd_sc_hd__buf_12 output337 (.A(net337),
    .X(wb_dat_o[19]));
 sky130_fd_sc_hd__buf_12 output338 (.A(net338),
    .X(wb_dat_o[1]));
 sky130_fd_sc_hd__buf_12 output339 (.A(net339),
    .X(wb_dat_o[20]));
 sky130_fd_sc_hd__buf_12 output340 (.A(net340),
    .X(wb_dat_o[21]));
 sky130_fd_sc_hd__buf_12 output341 (.A(net341),
    .X(wb_dat_o[22]));
 sky130_fd_sc_hd__buf_12 output342 (.A(net342),
    .X(wb_dat_o[23]));
 sky130_fd_sc_hd__buf_12 output343 (.A(net343),
    .X(wb_dat_o[24]));
 sky130_fd_sc_hd__buf_12 output344 (.A(net344),
    .X(wb_dat_o[25]));
 sky130_fd_sc_hd__buf_12 output345 (.A(net345),
    .X(wb_dat_o[26]));
 sky130_fd_sc_hd__buf_12 output346 (.A(net346),
    .X(wb_dat_o[27]));
 sky130_fd_sc_hd__buf_12 output347 (.A(net347),
    .X(wb_dat_o[28]));
 sky130_fd_sc_hd__buf_12 output348 (.A(net348),
    .X(wb_dat_o[29]));
 sky130_fd_sc_hd__buf_12 output349 (.A(net349),
    .X(wb_dat_o[2]));
 sky130_fd_sc_hd__buf_12 output350 (.A(net350),
    .X(wb_dat_o[30]));
 sky130_fd_sc_hd__buf_12 output351 (.A(net351),
    .X(wb_dat_o[31]));
 sky130_fd_sc_hd__buf_12 output352 (.A(net352),
    .X(wb_dat_o[3]));
 sky130_fd_sc_hd__buf_12 output353 (.A(net353),
    .X(wb_dat_o[4]));
 sky130_fd_sc_hd__buf_12 output354 (.A(net354),
    .X(wb_dat_o[5]));
 sky130_fd_sc_hd__buf_12 output355 (.A(net355),
    .X(wb_dat_o[6]));
 sky130_fd_sc_hd__buf_12 output356 (.A(net356),
    .X(wb_dat_o[7]));
 sky130_fd_sc_hd__buf_12 output357 (.A(net357),
    .X(wb_dat_o[8]));
 sky130_fd_sc_hd__buf_12 output358 (.A(net358),
    .X(wb_dat_o[9]));
 sky130_fd_sc_hd__buf_6 max_cap359 (.A(_0957_),
    .X(net359));
 sky130_fd_sc_hd__buf_8 max_cap360 (.A(_0953_),
    .X(net360));
 sky130_fd_sc_hd__buf_8 max_cap361 (.A(_0934_),
    .X(net361));
 sky130_fd_sc_hd__buf_6 max_cap362 (.A(_0933_),
    .X(net362));
 sky130_fd_sc_hd__buf_8 max_cap363 (.A(_0929_),
    .X(net363));
 sky130_fd_sc_hd__buf_8 max_cap364 (.A(_0925_),
    .X(net364));
 sky130_fd_sc_hd__buf_8 max_cap365 (.A(_0902_),
    .X(net365));
 sky130_fd_sc_hd__buf_8 max_cap366 (.A(_0884_),
    .X(net366));
 sky130_fd_sc_hd__clkbuf_1 wire367 (.A(net368),
    .X(net367));
 sky130_fd_sc_hd__clkbuf_1 wire368 (.A(net369),
    .X(net368));
 sky130_fd_sc_hd__clkbuf_1 wire369 (.A(_2601_),
    .X(net369));
 sky130_fd_sc_hd__buf_8 max_cap370 (.A(_1056_),
    .X(net370));
 sky130_fd_sc_hd__buf_8 max_cap371 (.A(_0976_),
    .X(net371));
 sky130_fd_sc_hd__buf_8 max_cap372 (.A(_0966_),
    .X(net372));
 sky130_fd_sc_hd__buf_6 wire373 (.A(_0960_),
    .X(net373));
 sky130_fd_sc_hd__buf_8 max_cap374 (.A(_0939_),
    .X(net374));
 sky130_fd_sc_hd__buf_6 wire375 (.A(_0932_),
    .X(net375));
 sky130_fd_sc_hd__buf_8 max_cap376 (.A(_0930_),
    .X(net376));
 sky130_fd_sc_hd__buf_6 max_cap377 (.A(_0924_),
    .X(net377));
 sky130_fd_sc_hd__buf_6 max_cap378 (.A(_0923_),
    .X(net378));
 sky130_fd_sc_hd__buf_6 max_cap379 (.A(_0922_),
    .X(net379));
 sky130_fd_sc_hd__buf_8 max_cap380 (.A(_0920_),
    .X(net380));
 sky130_fd_sc_hd__buf_8 max_cap381 (.A(_0913_),
    .X(net381));
 sky130_fd_sc_hd__buf_8 wire382 (.A(_0903_),
    .X(net382));
 sky130_fd_sc_hd__buf_8 max_cap383 (.A(_0899_),
    .X(net383));
 sky130_fd_sc_hd__buf_6 max_cap384 (.A(_0894_),
    .X(net384));
 sky130_fd_sc_hd__buf_8 max_cap385 (.A(_0891_),
    .X(net385));
 sky130_fd_sc_hd__buf_8 max_cap386 (.A(_0889_),
    .X(net386));
 sky130_fd_sc_hd__buf_6 max_cap387 (.A(_0882_),
    .X(net387));
 sky130_fd_sc_hd__buf_6 max_cap388 (.A(_0959_),
    .X(net388));
 sky130_fd_sc_hd__buf_6 max_cap389 (.A(_0949_),
    .X(net389));
 sky130_fd_sc_hd__buf_8 wire390 (.A(_0914_),
    .X(net390));
 sky130_fd_sc_hd__buf_8 max_cap391 (.A(_0912_),
    .X(net391));
 sky130_fd_sc_hd__buf_8 max_cap392 (.A(_0864_),
    .X(net392));
 sky130_fd_sc_hd__clkbuf_2 wire393 (.A(_3940_),
    .X(net393));
 sky130_fd_sc_hd__clkbuf_2 max_cap394 (.A(_2288_),
    .X(net394));
 sky130_fd_sc_hd__clkbuf_2 max_cap395 (.A(_2164_),
    .X(net395));
 sky130_fd_sc_hd__clkbuf_4 wire396 (.A(_1586_),
    .X(net396));
 sky130_fd_sc_hd__buf_4 max_cap397 (.A(net548),
    .X(net397));
 sky130_fd_sc_hd__buf_4 max_cap398 (.A(_0858_),
    .X(net398));
 sky130_fd_sc_hd__buf_4 max_cap399 (.A(_0849_),
    .X(net399));
 sky130_fd_sc_hd__buf_4 max_cap400 (.A(_0844_),
    .X(net400));
 sky130_fd_sc_hd__clkbuf_1 max_cap401 (.A(_1484_),
    .X(net401));
 sky130_fd_sc_hd__clkbuf_2 max_cap402 (.A(_0983_),
    .X(net402));
 sky130_fd_sc_hd__buf_2 max_cap403 (.A(net523),
    .X(net403));
 sky130_fd_sc_hd__clkbuf_4 fanout404 (.A(net406),
    .X(net404));
 sky130_fd_sc_hd__clkbuf_2 fanout405 (.A(net406),
    .X(net405));
 sky130_fd_sc_hd__buf_2 fanout406 (.A(net407),
    .X(net406));
 sky130_fd_sc_hd__clkbuf_2 fanout407 (.A(net410),
    .X(net407));
 sky130_fd_sc_hd__clkbuf_4 fanout408 (.A(net410),
    .X(net408));
 sky130_fd_sc_hd__clkbuf_4 fanout409 (.A(net410),
    .X(net409));
 sky130_fd_sc_hd__buf_2 fanout410 (.A(net457),
    .X(net410));
 sky130_fd_sc_hd__clkbuf_4 fanout411 (.A(net413),
    .X(net411));
 sky130_fd_sc_hd__clkbuf_2 fanout412 (.A(net413),
    .X(net412));
 sky130_fd_sc_hd__buf_2 fanout413 (.A(net416),
    .X(net413));
 sky130_fd_sc_hd__clkbuf_4 fanout414 (.A(net415),
    .X(net414));
 sky130_fd_sc_hd__buf_2 fanout415 (.A(net416),
    .X(net415));
 sky130_fd_sc_hd__clkbuf_4 fanout416 (.A(net457),
    .X(net416));
 sky130_fd_sc_hd__clkbuf_4 fanout417 (.A(net418),
    .X(net417));
 sky130_fd_sc_hd__clkbuf_4 fanout418 (.A(net426),
    .X(net418));
 sky130_fd_sc_hd__clkbuf_4 fanout419 (.A(net426),
    .X(net419));
 sky130_fd_sc_hd__clkbuf_4 fanout420 (.A(net424),
    .X(net420));
 sky130_fd_sc_hd__clkbuf_4 fanout421 (.A(net424),
    .X(net421));
 sky130_fd_sc_hd__clkbuf_4 fanout422 (.A(net424),
    .X(net422));
 sky130_fd_sc_hd__clkbuf_4 fanout423 (.A(net424),
    .X(net423));
 sky130_fd_sc_hd__clkbuf_2 fanout424 (.A(net426),
    .X(net424));
 sky130_fd_sc_hd__buf_4 fanout425 (.A(net426),
    .X(net425));
 sky130_fd_sc_hd__clkbuf_4 fanout426 (.A(net457),
    .X(net426));
 sky130_fd_sc_hd__clkbuf_4 fanout427 (.A(net429),
    .X(net427));
 sky130_fd_sc_hd__clkbuf_2 fanout428 (.A(net429),
    .X(net428));
 sky130_fd_sc_hd__clkbuf_4 fanout429 (.A(net435),
    .X(net429));
 sky130_fd_sc_hd__clkbuf_4 fanout430 (.A(net432),
    .X(net430));
 sky130_fd_sc_hd__clkbuf_2 fanout431 (.A(net432),
    .X(net431));
 sky130_fd_sc_hd__buf_4 fanout432 (.A(net435),
    .X(net432));
 sky130_fd_sc_hd__clkbuf_4 fanout433 (.A(net434),
    .X(net433));
 sky130_fd_sc_hd__buf_2 fanout434 (.A(net435),
    .X(net434));
 sky130_fd_sc_hd__buf_2 fanout435 (.A(net457),
    .X(net435));
 sky130_fd_sc_hd__clkbuf_4 fanout436 (.A(net439),
    .X(net436));
 sky130_fd_sc_hd__clkbuf_2 fanout437 (.A(net439),
    .X(net437));
 sky130_fd_sc_hd__clkbuf_4 fanout438 (.A(net439),
    .X(net438));
 sky130_fd_sc_hd__buf_2 fanout439 (.A(net449),
    .X(net439));
 sky130_fd_sc_hd__clkbuf_4 fanout440 (.A(net441),
    .X(net440));
 sky130_fd_sc_hd__buf_4 fanout441 (.A(net449),
    .X(net441));
 sky130_fd_sc_hd__clkbuf_2 fanout442 (.A(net449),
    .X(net442));
 sky130_fd_sc_hd__clkbuf_4 fanout443 (.A(net449),
    .X(net443));
 sky130_fd_sc_hd__clkbuf_4 fanout444 (.A(net449),
    .X(net444));
 sky130_fd_sc_hd__clkbuf_4 fanout445 (.A(net446),
    .X(net445));
 sky130_fd_sc_hd__clkbuf_4 fanout446 (.A(net448),
    .X(net446));
 sky130_fd_sc_hd__clkbuf_4 fanout447 (.A(net448),
    .X(net447));
 sky130_fd_sc_hd__buf_2 fanout448 (.A(net449),
    .X(net448));
 sky130_fd_sc_hd__buf_2 fanout449 (.A(net457),
    .X(net449));
 sky130_fd_sc_hd__buf_4 fanout450 (.A(net456),
    .X(net450));
 sky130_fd_sc_hd__buf_4 fanout451 (.A(net453),
    .X(net451));
 sky130_fd_sc_hd__clkbuf_2 fanout452 (.A(net453),
    .X(net452));
 sky130_fd_sc_hd__clkbuf_4 fanout453 (.A(net456),
    .X(net453));
 sky130_fd_sc_hd__clkbuf_4 fanout454 (.A(net455),
    .X(net454));
 sky130_fd_sc_hd__clkbuf_4 fanout455 (.A(net456),
    .X(net455));
 sky130_fd_sc_hd__buf_4 fanout456 (.A(net457),
    .X(net456));
 sky130_fd_sc_hd__buf_4 fanout457 (.A(net75),
    .X(net457));
 sky130_fd_sc_hd__clkbuf_4 fanout458 (.A(net459),
    .X(net458));
 sky130_fd_sc_hd__clkbuf_2 fanout459 (.A(net462),
    .X(net459));
 sky130_fd_sc_hd__clkbuf_4 fanout460 (.A(net461),
    .X(net460));
 sky130_fd_sc_hd__buf_4 fanout461 (.A(net462),
    .X(net461));
 sky130_fd_sc_hd__clkbuf_4 fanout462 (.A(net498),
    .X(net462));
 sky130_fd_sc_hd__clkbuf_4 fanout463 (.A(net464),
    .X(net463));
 sky130_fd_sc_hd__clkbuf_4 fanout464 (.A(net498),
    .X(net464));
 sky130_fd_sc_hd__clkbuf_4 fanout465 (.A(net498),
    .X(net465));
 sky130_fd_sc_hd__buf_2 fanout466 (.A(net498),
    .X(net466));
 sky130_fd_sc_hd__buf_4 fanout467 (.A(net497),
    .X(net467));
 sky130_fd_sc_hd__buf_2 fanout468 (.A(net497),
    .X(net468));
 sky130_fd_sc_hd__buf_4 fanout469 (.A(net497),
    .X(net469));
 sky130_fd_sc_hd__clkbuf_2 fanout470 (.A(net497),
    .X(net470));
 sky130_fd_sc_hd__buf_4 fanout471 (.A(net496),
    .X(net471));
 sky130_fd_sc_hd__buf_2 fanout472 (.A(net496),
    .X(net472));
 sky130_fd_sc_hd__clkbuf_4 fanout473 (.A(net474),
    .X(net473));
 sky130_fd_sc_hd__clkbuf_4 fanout474 (.A(net496),
    .X(net474));
 sky130_fd_sc_hd__clkbuf_4 fanout475 (.A(net483),
    .X(net475));
 sky130_fd_sc_hd__clkbuf_4 fanout476 (.A(net483),
    .X(net476));
 sky130_fd_sc_hd__clkbuf_4 fanout477 (.A(net483),
    .X(net477));
 sky130_fd_sc_hd__buf_2 fanout478 (.A(net483),
    .X(net478));
 sky130_fd_sc_hd__clkbuf_4 fanout479 (.A(net482),
    .X(net479));
 sky130_fd_sc_hd__clkbuf_2 fanout480 (.A(net482),
    .X(net480));
 sky130_fd_sc_hd__clkbuf_4 fanout481 (.A(net482),
    .X(net481));
 sky130_fd_sc_hd__buf_2 fanout482 (.A(net483),
    .X(net482));
 sky130_fd_sc_hd__clkbuf_2 fanout483 (.A(net496),
    .X(net483));
 sky130_fd_sc_hd__buf_4 fanout484 (.A(net496),
    .X(net484));
 sky130_fd_sc_hd__buf_2 fanout485 (.A(net496),
    .X(net485));
 sky130_fd_sc_hd__clkbuf_4 fanout486 (.A(net488),
    .X(net486));
 sky130_fd_sc_hd__clkbuf_2 fanout487 (.A(net488),
    .X(net487));
 sky130_fd_sc_hd__buf_2 fanout488 (.A(net496),
    .X(net488));
 sky130_fd_sc_hd__clkbuf_4 fanout489 (.A(net495),
    .X(net489));
 sky130_fd_sc_hd__clkbuf_2 fanout490 (.A(net495),
    .X(net490));
 sky130_fd_sc_hd__clkbuf_4 fanout491 (.A(net495),
    .X(net491));
 sky130_fd_sc_hd__clkbuf_2 fanout492 (.A(net495),
    .X(net492));
 sky130_fd_sc_hd__clkbuf_4 fanout493 (.A(net494),
    .X(net493));
 sky130_fd_sc_hd__buf_2 fanout494 (.A(net495),
    .X(net494));
 sky130_fd_sc_hd__clkbuf_2 fanout495 (.A(net496),
    .X(net495));
 sky130_fd_sc_hd__clkbuf_4 fanout496 (.A(net497),
    .X(net496));
 sky130_fd_sc_hd__clkbuf_4 fanout497 (.A(net498),
    .X(net497));
 sky130_fd_sc_hd__buf_4 fanout498 (.A(net75),
    .X(net498));
 sky130_fd_sc_hd__clkbuf_4 fanout499 (.A(net501),
    .X(net499));
 sky130_fd_sc_hd__clkbuf_2 fanout500 (.A(net501),
    .X(net500));
 sky130_fd_sc_hd__buf_2 fanout501 (.A(net502),
    .X(net501));
 sky130_fd_sc_hd__clkbuf_4 fanout502 (.A(net503),
    .X(net502));
 sky130_fd_sc_hd__buf_4 fanout503 (.A(net196),
    .X(net503));
 sky130_fd_sc_hd__conb_1 _9503__504 (.HI(net504));
 sky130_fd_sc_hd__inv_2 net499_2 (.A(clknet_2_3_0_mgmt_gpio_in[4]),
    .Y(net506));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_1_0_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_1_0_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_1_0_1_wb_clk_i (.A(clknet_1_0_0_wb_clk_i),
    .X(clknet_1_0_1_wb_clk_i));
 sky130_fd_sc_hd__buf_8 clkbuf_1_1_0_wb_clk_i (.A(net509),
    .X(clknet_1_1_0_wb_clk_i));
 sky130_fd_sc_hd__buf_8 clkbuf_1_1_1_wb_clk_i (.A(clknet_1_1_0_wb_clk_i),
    .X(clknet_1_1_1_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_2_0_0_wb_clk_i (.A(clknet_1_0_1_wb_clk_i),
    .X(clknet_2_0_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_2_1_0_wb_clk_i (.A(clknet_1_0_1_wb_clk_i),
    .X(clknet_2_1_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_2_2_0_wb_clk_i (.A(clknet_1_1_1_wb_clk_i),
    .X(clknet_2_2_0_wb_clk_i));
 sky130_fd_sc_hd__buf_8 clkbuf_2_3_0_wb_clk_i (.A(clknet_1_1_1_wb_clk_i),
    .X(clknet_2_3_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_0_0_wb_clk_i (.A(clknet_2_0_0_wb_clk_i),
    .X(clknet_3_0_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_1_0_wb_clk_i (.A(clknet_2_0_0_wb_clk_i),
    .X(clknet_3_1_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_2_0_wb_clk_i (.A(clknet_2_1_0_wb_clk_i),
    .X(clknet_3_2_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_3_0_wb_clk_i (.A(clknet_2_1_0_wb_clk_i),
    .X(clknet_3_3_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_4_0_wb_clk_i (.A(clknet_2_2_0_wb_clk_i),
    .X(clknet_3_4_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_5_0_wb_clk_i (.A(clknet_2_2_0_wb_clk_i),
    .X(clknet_3_5_0_wb_clk_i));
 sky130_fd_sc_hd__buf_12 clkbuf_3_6_0_wb_clk_i (.A(clknet_2_3_0_wb_clk_i),
    .X(clknet_3_6_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_7_0_wb_clk_i (.A(clknet_2_3_0_wb_clk_i),
    .X(clknet_3_7_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_mgmt_gpio_in[4]  (.A(mgmt_gpio_in[4]),
    .X(clknet_0_mgmt_gpio_in[4]));
 sky130_fd_sc_hd__clkbuf_8 \clkbuf_1_0_0_mgmt_gpio_in[4]  (.A(clknet_0_mgmt_gpio_in[4]),
    .X(clknet_1_0_0_mgmt_gpio_in[4]));
 sky130_fd_sc_hd__clkbuf_8 \clkbuf_1_1_0_mgmt_gpio_in[4]  (.A(clknet_0_mgmt_gpio_in[4]),
    .X(clknet_1_1_0_mgmt_gpio_in[4]));
 sky130_fd_sc_hd__clkbuf_8 \clkbuf_2_0_0_mgmt_gpio_in[4]  (.A(clknet_1_0_0_mgmt_gpio_in[4]),
    .X(clknet_2_0_0_mgmt_gpio_in[4]));
 sky130_fd_sc_hd__clkbuf_8 \clkbuf_2_1_0_mgmt_gpio_in[4]  (.A(clknet_1_0_0_mgmt_gpio_in[4]),
    .X(clknet_2_1_0_mgmt_gpio_in[4]));
 sky130_fd_sc_hd__clkbuf_8 \clkbuf_2_2_0_mgmt_gpio_in[4]  (.A(clknet_1_1_0_mgmt_gpio_in[4]),
    .X(clknet_2_2_0_mgmt_gpio_in[4]));
 sky130_fd_sc_hd__clkbuf_8 \clkbuf_2_3_0_mgmt_gpio_in[4]  (.A(clknet_1_1_0_mgmt_gpio_in[4]),
    .X(clknet_2_3_0_mgmt_gpio_in[4]));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_0_csclk (.A(clknet_3_1_0_csclk),
    .X(clknet_leaf_0_csclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_1_csclk (.A(clknet_3_1_0_csclk),
    .X(clknet_leaf_1_csclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_2_csclk (.A(clknet_3_1_0_csclk),
    .X(clknet_leaf_2_csclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_3_csclk (.A(clknet_3_1_0_csclk),
    .X(clknet_leaf_3_csclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_4_csclk (.A(clknet_3_1_0_csclk),
    .X(clknet_leaf_4_csclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_5_csclk (.A(clknet_3_1_0_csclk),
    .X(clknet_leaf_5_csclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_6_csclk (.A(clknet_3_1_0_csclk),
    .X(clknet_leaf_6_csclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_7_csclk (.A(clknet_3_1_0_csclk),
    .X(clknet_leaf_7_csclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_9_csclk (.A(clknet_3_1_0_csclk),
    .X(clknet_leaf_9_csclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_10_csclk (.A(clknet_3_4_0_csclk),
    .X(clknet_leaf_10_csclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_11_csclk (.A(clknet_3_4_0_csclk),
    .X(clknet_leaf_11_csclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_12_csclk (.A(clknet_3_4_0_csclk),
    .X(clknet_leaf_12_csclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_13_csclk (.A(clknet_3_4_0_csclk),
    .X(clknet_leaf_13_csclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_14_csclk (.A(clknet_opt_1_0_csclk),
    .X(clknet_leaf_14_csclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_16_csclk (.A(clknet_3_5_0_csclk),
    .X(clknet_leaf_16_csclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_17_csclk (.A(clknet_3_5_0_csclk),
    .X(clknet_leaf_17_csclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_18_csclk (.A(clknet_3_5_0_csclk),
    .X(clknet_leaf_18_csclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_19_csclk (.A(clknet_3_5_0_csclk),
    .X(clknet_leaf_19_csclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_20_csclk (.A(clknet_3_4_0_csclk),
    .X(clknet_leaf_20_csclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_21_csclk (.A(clknet_3_4_0_csclk),
    .X(clknet_leaf_21_csclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_23_csclk (.A(clknet_3_4_0_csclk),
    .X(clknet_leaf_23_csclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_24_csclk (.A(clknet_3_5_0_csclk),
    .X(clknet_leaf_24_csclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_25_csclk (.A(clknet_3_7_0_csclk),
    .X(clknet_leaf_25_csclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_26_csclk (.A(clknet_3_7_0_csclk),
    .X(clknet_leaf_26_csclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_27_csclk (.A(clknet_3_5_0_csclk),
    .X(clknet_leaf_27_csclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_28_csclk (.A(clknet_3_7_0_csclk),
    .X(clknet_leaf_28_csclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_29_csclk (.A(clknet_3_5_0_csclk),
    .X(clknet_leaf_29_csclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_30_csclk (.A(clknet_3_7_0_csclk),
    .X(clknet_leaf_30_csclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_31_csclk (.A(clknet_3_7_0_csclk),
    .X(clknet_leaf_31_csclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_32_csclk (.A(clknet_3_7_0_csclk),
    .X(clknet_leaf_32_csclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_33_csclk (.A(clknet_3_7_0_csclk),
    .X(clknet_leaf_33_csclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_34_csclk (.A(clknet_3_7_0_csclk),
    .X(clknet_leaf_34_csclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_35_csclk (.A(clknet_3_7_0_csclk),
    .X(clknet_leaf_35_csclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_36_csclk (.A(clknet_3_7_0_csclk),
    .X(clknet_leaf_36_csclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_37_csclk (.A(clknet_3_7_0_csclk),
    .X(clknet_leaf_37_csclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_38_csclk (.A(clknet_3_7_0_csclk),
    .X(clknet_leaf_38_csclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_39_csclk (.A(clknet_3_7_0_csclk),
    .X(clknet_leaf_39_csclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_40_csclk (.A(clknet_3_7_0_csclk),
    .X(clknet_leaf_40_csclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_41_csclk (.A(clknet_3_7_0_csclk),
    .X(clknet_leaf_41_csclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_42_csclk (.A(clknet_3_6_0_csclk),
    .X(clknet_leaf_42_csclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_43_csclk (.A(clknet_3_6_0_csclk),
    .X(clknet_leaf_43_csclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_45_csclk (.A(clknet_3_6_0_csclk),
    .X(clknet_leaf_45_csclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_46_csclk (.A(clknet_3_6_0_csclk),
    .X(clknet_leaf_46_csclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_47_csclk (.A(clknet_3_6_0_csclk),
    .X(clknet_leaf_47_csclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_48_csclk (.A(clknet_3_6_0_csclk),
    .X(clknet_leaf_48_csclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_49_csclk (.A(clknet_3_6_0_csclk),
    .X(clknet_leaf_49_csclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_50_csclk (.A(clknet_3_3_0_csclk),
    .X(clknet_leaf_50_csclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_52_csclk (.A(clknet_3_3_0_csclk),
    .X(clknet_leaf_52_csclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_53_csclk (.A(clknet_3_6_0_csclk),
    .X(clknet_leaf_53_csclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_55_csclk (.A(clknet_opt_2_0_csclk),
    .X(clknet_leaf_55_csclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_56_csclk (.A(clknet_3_3_0_csclk),
    .X(clknet_leaf_56_csclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_57_csclk (.A(clknet_3_3_0_csclk),
    .X(clknet_leaf_57_csclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_58_csclk (.A(clknet_3_2_0_csclk),
    .X(clknet_leaf_58_csclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_59_csclk (.A(clknet_3_2_0_csclk),
    .X(clknet_leaf_59_csclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_60_csclk (.A(clknet_3_2_0_csclk),
    .X(clknet_leaf_60_csclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_61_csclk (.A(clknet_3_2_0_csclk),
    .X(clknet_leaf_61_csclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_62_csclk (.A(clknet_3_2_0_csclk),
    .X(clknet_leaf_62_csclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_63_csclk (.A(clknet_3_2_0_csclk),
    .X(clknet_leaf_63_csclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_64_csclk (.A(clknet_3_3_0_csclk),
    .X(clknet_leaf_64_csclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_65_csclk (.A(clknet_3_2_0_csclk),
    .X(clknet_leaf_65_csclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_66_csclk (.A(clknet_3_2_0_csclk),
    .X(clknet_leaf_66_csclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_67_csclk (.A(clknet_3_2_0_csclk),
    .X(clknet_leaf_67_csclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_68_csclk (.A(clknet_3_2_0_csclk),
    .X(clknet_leaf_68_csclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_69_csclk (.A(clknet_3_2_0_csclk),
    .X(clknet_leaf_69_csclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_70_csclk (.A(clknet_3_2_0_csclk),
    .X(clknet_leaf_70_csclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_71_csclk (.A(clknet_3_3_0_csclk),
    .X(clknet_leaf_71_csclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_72_csclk (.A(clknet_3_3_0_csclk),
    .X(clknet_leaf_72_csclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_73_csclk (.A(clknet_3_3_0_csclk),
    .X(clknet_leaf_73_csclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_74_csclk (.A(clknet_3_1_0_csclk),
    .X(clknet_leaf_74_csclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_75_csclk (.A(clknet_3_1_0_csclk),
    .X(clknet_leaf_75_csclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_76_csclk (.A(clknet_3_0_0_csclk),
    .X(clknet_leaf_76_csclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_77_csclk (.A(clknet_3_2_0_csclk),
    .X(clknet_leaf_77_csclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_78_csclk (.A(clknet_3_2_0_csclk),
    .X(clknet_leaf_78_csclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_79_csclk (.A(clknet_3_0_0_csclk),
    .X(clknet_leaf_79_csclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_80_csclk (.A(clknet_3_0_0_csclk),
    .X(clknet_leaf_80_csclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_81_csclk (.A(clknet_3_0_0_csclk),
    .X(clknet_leaf_81_csclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_82_csclk (.A(clknet_3_0_0_csclk),
    .X(clknet_leaf_82_csclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_83_csclk (.A(clknet_3_0_0_csclk),
    .X(clknet_leaf_83_csclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_84_csclk (.A(clknet_3_0_0_csclk),
    .X(clknet_leaf_84_csclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_85_csclk (.A(clknet_3_0_0_csclk),
    .X(clknet_leaf_85_csclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_86_csclk (.A(clknet_3_0_0_csclk),
    .X(clknet_leaf_86_csclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_csclk (.A(csclk),
    .X(clknet_0_csclk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_1_0_0_csclk (.A(clknet_0_csclk),
    .X(clknet_1_0_0_csclk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_1_0_1_csclk (.A(clknet_1_0_0_csclk),
    .X(clknet_1_0_1_csclk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_1_1_0_csclk (.A(clknet_0_csclk),
    .X(clknet_1_1_0_csclk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_1_1_1_csclk (.A(clknet_1_1_0_csclk),
    .X(clknet_1_1_1_csclk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_2_0_0_csclk (.A(clknet_1_0_1_csclk),
    .X(clknet_2_0_0_csclk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_2_1_0_csclk (.A(clknet_1_0_1_csclk),
    .X(clknet_2_1_0_csclk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_2_2_0_csclk (.A(clknet_1_1_1_csclk),
    .X(clknet_2_2_0_csclk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_2_3_0_csclk (.A(clknet_1_1_1_csclk),
    .X(clknet_2_3_0_csclk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_0_0_csclk (.A(clknet_2_0_0_csclk),
    .X(clknet_3_0_0_csclk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_1_0_csclk (.A(clknet_2_0_0_csclk),
    .X(clknet_3_1_0_csclk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_2_0_csclk (.A(clknet_2_1_0_csclk),
    .X(clknet_3_2_0_csclk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_3_0_csclk (.A(clknet_2_1_0_csclk),
    .X(clknet_3_3_0_csclk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_4_0_csclk (.A(clknet_2_2_0_csclk),
    .X(clknet_3_4_0_csclk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_5_0_csclk (.A(clknet_2_2_0_csclk),
    .X(clknet_3_5_0_csclk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_6_0_csclk (.A(clknet_2_3_0_csclk),
    .X(clknet_3_6_0_csclk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_7_0_csclk (.A(clknet_2_3_0_csclk),
    .X(clknet_3_7_0_csclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_opt_1_0_csclk (.A(clknet_3_4_0_csclk),
    .X(clknet_opt_1_0_csclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_opt_2_0_csclk (.A(clknet_3_6_0_csclk),
    .X(clknet_opt_2_0_csclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__1160_ (.A(_1160_),
    .X(clknet_0__1160_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__1160_ (.A(clknet_0__1160_),
    .X(clknet_1_0__leaf__1160_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__1160_ (.A(clknet_0__1160_),
    .X(clknet_1_1__leaf__1160_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_wbbd_sck (.A(wbbd_sck),
    .X(clknet_0_wbbd_sck));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_wbbd_sck (.A(clknet_0_wbbd_sck),
    .X(clknet_1_0__leaf_wbbd_sck));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_wbbd_sck (.A(clknet_0_wbbd_sck),
    .X(clknet_1_1__leaf_wbbd_sck));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer1 (.A(clknet_3_6_0_wb_clk_i),
    .X(net507));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer2 (.A(clknet_3_6_0_wb_clk_i),
    .X(net508));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4 (.A(\hkspi.odata[7] ),
    .X(net510));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5 (.A(net1542),
    .X(net511));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6 (.A(_1927_),
    .X(net512));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7 (.A(net582),
    .X(net513));
 sky130_fd_sc_hd__dlygate4sd3_1 hold8 (.A(\hkspi.addr[1] ),
    .X(net514));
 sky130_fd_sc_hd__dlygate4sd3_1 hold9 (.A(_0845_),
    .X(net515));
 sky130_fd_sc_hd__dlygate4sd3_1 hold10 (.A(_0846_),
    .X(net516));
 sky130_fd_sc_hd__dlygate4sd3_1 hold11 (.A(\hkspi.odata[2] ),
    .X(net517));
 sky130_fd_sc_hd__dlygate4sd3_1 hold12 (.A(net1064),
    .X(net518));
 sky130_fd_sc_hd__dlygate4sd3_1 hold13 (.A(_1955_),
    .X(net519));
 sky130_fd_sc_hd__dlygate4sd3_1 hold14 (.A(\hkspi.odata[5] ),
    .X(net520));
 sky130_fd_sc_hd__dlygate4sd3_1 hold15 (.A(net1554),
    .X(net521));
 sky130_fd_sc_hd__dlygate4sd3_1 hold16 (.A(_1940_),
    .X(net522));
 sky130_fd_sc_hd__dlygate4sd3_1 hold17 (.A(\hkspi.wrstb ),
    .X(net523));
 sky130_fd_sc_hd__dlygate4sd3_1 hold18 (.A(net403),
    .X(net524));
 sky130_fd_sc_hd__dlygate4sd3_1 hold19 (.A(_1600_),
    .X(net525));
 sky130_fd_sc_hd__dlygate4sd3_1 hold20 (.A(_1601_),
    .X(net526));
 sky130_fd_sc_hd__dlygate4sd3_1 hold21 (.A(_1912_),
    .X(net527));
 sky130_fd_sc_hd__dlygate4sd3_1 hold22 (.A(net600),
    .X(net528));
 sky130_fd_sc_hd__dlygate4sd3_1 hold23 (.A(net1668),
    .X(net529));
 sky130_fd_sc_hd__dlygate4sd3_1 hold24 (.A(_1617_),
    .X(net530));
 sky130_fd_sc_hd__dlygate4sd3_1 hold25 (.A(_1921_),
    .X(net531));
 sky130_fd_sc_hd__dlygate4sd3_1 hold26 (.A(net1560),
    .X(net532));
 sky130_fd_sc_hd__dlygate4sd3_1 hold27 (.A(_1674_),
    .X(net533));
 sky130_fd_sc_hd__dlygate4sd3_1 hold28 (.A(_1942_),
    .X(net534));
 sky130_fd_sc_hd__dlygate4sd3_1 hold29 (.A(\hkspi.addr[6] ),
    .X(net535));
 sky130_fd_sc_hd__dlygate4sd3_1 hold30 (.A(_0827_),
    .X(net536));
 sky130_fd_sc_hd__dlygate4sd3_1 hold31 (.A(_0861_),
    .X(net537));
 sky130_fd_sc_hd__dlygate4sd3_1 hold32 (.A(_0907_),
    .X(net538));
 sky130_fd_sc_hd__buf_12 hold33 (.A(_0908_),
    .X(net539));
 sky130_fd_sc_hd__dlygate4sd3_1 hold34 (.A(_1959_),
    .X(net540));
 sky130_fd_sc_hd__dlygate4sd3_1 hold35 (.A(net591),
    .X(net541));
 sky130_fd_sc_hd__dlygate4sd3_1 hold36 (.A(\hkspi.odata[1] ),
    .X(net542));
 sky130_fd_sc_hd__dlygate4sd3_1 hold37 (.A(net575),
    .X(net543));
 sky130_fd_sc_hd__dlygate4sd3_1 hold38 (.A(_1932_),
    .X(net544));
 sky130_fd_sc_hd__dlygate4sd3_1 hold39 (.A(\hkspi.addr[2] ),
    .X(net545));
 sky130_fd_sc_hd__dlygate4sd3_1 hold40 (.A(_0842_),
    .X(net546));
 sky130_fd_sc_hd__dlygate4sd3_1 hold41 (.A(_0843_),
    .X(net547));
 sky130_fd_sc_hd__dlygate4sd3_1 hold42 (.A(_0892_),
    .X(net548));
 sky130_fd_sc_hd__dlygate4sd3_1 hold43 (.A(_1913_),
    .X(net549));
 sky130_fd_sc_hd__dlygate4sd3_1 hold44 (.A(\hkspi.odata[3] ),
    .X(net550));
 sky130_fd_sc_hd__dlygate4sd3_1 hold45 (.A(net704),
    .X(net551));
 sky130_fd_sc_hd__dlygate4sd3_1 hold46 (.A(_1835_),
    .X(net552));
 sky130_fd_sc_hd__dlygate4sd3_1 hold47 (.A(_3405_),
    .X(net553));
 sky130_fd_sc_hd__dlygate4sd3_1 hold48 (.A(_0716_),
    .X(net554));
 sky130_fd_sc_hd__dlygate4sd3_1 hold49 (.A(net1749),
    .X(net555));
 sky130_fd_sc_hd__dlygate4sd3_1 hold50 (.A(_0836_),
    .X(net556));
 sky130_fd_sc_hd__dlygate4sd3_1 hold51 (.A(_0837_),
    .X(net557));
 sky130_fd_sc_hd__dlygate4sd3_1 hold52 (.A(_0878_),
    .X(net558));
 sky130_fd_sc_hd__dlygate4sd3_1 hold53 (.A(_0887_),
    .X(net559));
 sky130_fd_sc_hd__dlygate4sd3_1 hold54 (.A(_3323_),
    .X(net560));
 sky130_fd_sc_hd__dlygate4sd3_1 hold55 (.A(\hkspi.addr[5] ),
    .X(net561));
 sky130_fd_sc_hd__dlygate4sd3_1 hold56 (.A(_0828_),
    .X(net562));
 sky130_fd_sc_hd__dlygate4sd3_1 hold57 (.A(_0830_),
    .X(net563));
 sky130_fd_sc_hd__dlygate4sd3_1 hold58 (.A(_0831_),
    .X(net564));
 sky130_fd_sc_hd__dlygate4sd3_1 hold59 (.A(_0866_),
    .X(net565));
 sky130_fd_sc_hd__dlygate4sd3_1 hold60 (.A(_0867_),
    .X(net566));
 sky130_fd_sc_hd__dlygate4sd3_1 hold61 (.A(_3245_),
    .X(net567));
 sky130_fd_sc_hd__dlygate4sd3_1 hold62 (.A(\wbbd_addr[3] ),
    .X(net568));
 sky130_fd_sc_hd__dlygate4sd3_1 hold63 (.A(_0841_),
    .X(net569));
 sky130_fd_sc_hd__dlygate4sd3_1 hold64 (.A(_0869_),
    .X(net570));
 sky130_fd_sc_hd__dlygate4sd3_1 hold65 (.A(_3030_),
    .X(net571));
 sky130_fd_sc_hd__dlygate4sd3_1 hold66 (.A(net1764),
    .X(net572));
 sky130_fd_sc_hd__dlygate4sd3_1 hold67 (.A(_3172_),
    .X(net573));
 sky130_fd_sc_hd__dlygate4sd3_1 hold68 (.A(\wbbd_data[1] ),
    .X(net574));
 sky130_fd_sc_hd__dlygate4sd3_1 hold69 (.A(_1605_),
    .X(net575));
 sky130_fd_sc_hd__dlygate4sd3_1 hold70 (.A(_1953_),
    .X(net576));
 sky130_fd_sc_hd__dlygate4sd3_1 hold71 (.A(\gpio_configure[16][11] ),
    .X(net577));
 sky130_fd_sc_hd__dlygate4sd3_1 hold72 (.A(_2065_),
    .X(net578));
 sky130_fd_sc_hd__dlygate4sd3_1 hold73 (.A(wbbd_busy),
    .X(net579));
 sky130_fd_sc_hd__dlygate4sd3_1 hold74 (.A(_0824_),
    .X(net580));
 sky130_fd_sc_hd__dlygate4sd3_1 hold75 (.A(_3314_),
    .X(net581));
 sky130_fd_sc_hd__dlygate4sd3_1 hold76 (.A(\hkspi.addr[0] ),
    .X(net582));
 sky130_fd_sc_hd__dlygate4sd3_1 hold77 (.A(net513),
    .X(net583));
 sky130_fd_sc_hd__dlygate4sd3_1 hold78 (.A(_3305_),
    .X(net584));
 sky130_fd_sc_hd__dlygate4sd3_1 hold79 (.A(_3023_),
    .X(net585));
 sky130_fd_sc_hd__dlygate4sd3_1 hold80 (.A(\hkspi.addr[4] ),
    .X(net586));
 sky130_fd_sc_hd__dlygate4sd3_1 hold81 (.A(_0833_),
    .X(net587));
 sky130_fd_sc_hd__dlygate4sd3_1 hold82 (.A(_0834_),
    .X(net588));
 sky130_fd_sc_hd__dlygate4sd3_1 hold83 (.A(_0862_),
    .X(net589));
 sky130_fd_sc_hd__dlygate4sd3_1 hold84 (.A(_3342_),
    .X(net590));
 sky130_fd_sc_hd__dlygate4sd3_1 hold85 (.A(\wbbd_addr[0] ),
    .X(net591));
 sky130_fd_sc_hd__dlygate4sd3_1 hold86 (.A(_3391_),
    .X(net592));
 sky130_fd_sc_hd__dlygate4sd3_1 hold87 (.A(_3393_),
    .X(net593));
 sky130_fd_sc_hd__dlygate4sd3_1 hold88 (.A(\gpio_configure[29][1] ),
    .X(net594));
 sky130_fd_sc_hd__dlygate4sd3_1 hold89 (.A(_3375_),
    .X(net595));
 sky130_fd_sc_hd__dlygate4sd3_1 hold90 (.A(\gpio_configure[25][1] ),
    .X(net596));
 sky130_fd_sc_hd__dlygate4sd3_1 hold91 (.A(_3335_),
    .X(net597));
 sky130_fd_sc_hd__dlygate4sd3_1 hold92 (.A(\gpio_configure[27][1] ),
    .X(net598));
 sky130_fd_sc_hd__dlygate4sd3_1 hold93 (.A(_3357_),
    .X(net599));
 sky130_fd_sc_hd__dlygate4sd3_1 hold94 (.A(\hkspi.state[3] ),
    .X(net600));
 sky130_fd_sc_hd__dlygate4sd3_1 hold95 (.A(_3382_),
    .X(net601));
 sky130_fd_sc_hd__dlygate4sd3_1 hold96 (.A(\gpio_configure[28][1] ),
    .X(net602));
 sky130_fd_sc_hd__dlygate4sd3_1 hold97 (.A(_3366_),
    .X(net603));
 sky130_fd_sc_hd__dlygate4sd3_1 hold98 (.A(\wbbd_addr[1] ),
    .X(net604));
 sky130_fd_sc_hd__dlygate4sd3_1 hold99 (.A(_3295_),
    .X(net605));
 sky130_fd_sc_hd__dlygate4sd3_1 hold100 (.A(_3298_),
    .X(net606));
 sky130_fd_sc_hd__dlygate4sd3_1 hold101 (.A(_1964_),
    .X(net607));
 sky130_fd_sc_hd__dlygate4sd3_1 hold102 (.A(_0298_),
    .X(net608));
 sky130_fd_sc_hd__dlygate4sd3_1 hold103 (.A(wbbd_write),
    .X(net609));
 sky130_fd_sc_hd__dlygate4sd3_1 hold104 (.A(_1599_),
    .X(net610));
 sky130_fd_sc_hd__dlygate4sd3_1 hold105 (.A(_1700_),
    .X(net611));
 sky130_fd_sc_hd__dlygate4sd3_1 hold106 (.A(_3082_),
    .X(net612));
 sky130_fd_sc_hd__dlygate4sd3_1 hold107 (.A(_0453_),
    .X(net613));
 sky130_fd_sc_hd__dlygate4sd3_1 hold108 (.A(\gpio_configure[8][1] ),
    .X(net614));
 sky130_fd_sc_hd__dlygate4sd3_1 hold109 (.A(\gpio_configure[16][1] ),
    .X(net615));
 sky130_fd_sc_hd__dlygate4sd3_1 hold110 (.A(\mgmt_gpio_data_buf[20] ),
    .X(net616));
 sky130_fd_sc_hd__dlygate4sd3_1 hold111 (.A(_1707_),
    .X(net617));
 sky130_fd_sc_hd__dlygate4sd3_1 hold112 (.A(\wbbd_data[4] ),
    .X(net618));
 sky130_fd_sc_hd__dlygate4sd3_1 hold113 (.A(_1751_),
    .X(net619));
 sky130_fd_sc_hd__dlygate4sd3_1 hold114 (.A(\gpio_configure[24][1] ),
    .X(net620));
 sky130_fd_sc_hd__dlygate4sd3_1 hold115 (.A(\gpio_configure[6][1] ),
    .X(net621));
 sky130_fd_sc_hd__dlygate4sd3_1 hold116 (.A(_3148_),
    .X(net622));
 sky130_fd_sc_hd__dlygate4sd3_1 hold117 (.A(\gpio_configure[32][4] ),
    .X(net623));
 sky130_fd_sc_hd__dlygate4sd3_1 hold118 (.A(_3406_),
    .X(net624));
 sky130_fd_sc_hd__dlygate4sd3_1 hold119 (.A(\gpio_configure[9][1] ),
    .X(net625));
 sky130_fd_sc_hd__dlygate4sd3_1 hold120 (.A(_3179_),
    .X(net626));
 sky130_fd_sc_hd__dlygate4sd3_1 hold121 (.A(\gpio_configure[19][12] ),
    .X(net627));
 sky130_fd_sc_hd__dlygate4sd3_1 hold122 (.A(_1829_),
    .X(net628));
 sky130_fd_sc_hd__dlygate4sd3_1 hold123 (.A(\gpio_configure[30][12] ),
    .X(net629));
 sky130_fd_sc_hd__dlygate4sd3_1 hold124 (.A(_1864_),
    .X(net630));
 sky130_fd_sc_hd__dlygate4sd3_1 hold125 (.A(\gpio_configure[17][1] ),
    .X(net631));
 sky130_fd_sc_hd__dlygate4sd3_1 hold126 (.A(_3257_),
    .X(net632));
 sky130_fd_sc_hd__dlygate4sd3_1 hold127 (.A(\gpio_configure[18][1] ),
    .X(net633));
 sky130_fd_sc_hd__dlygate4sd3_1 hold128 (.A(_3267_),
    .X(net634));
 sky130_fd_sc_hd__dlygate4sd3_1 hold129 (.A(\gpio_configure[28][12] ),
    .X(net635));
 sky130_fd_sc_hd__dlygate4sd3_1 hold130 (.A(_1890_),
    .X(net636));
 sky130_fd_sc_hd__dlygate4sd3_1 hold131 (.A(\gpio_configure[26][12] ),
    .X(net637));
 sky130_fd_sc_hd__dlygate4sd3_1 hold132 (.A(_1619_),
    .X(net638));
 sky130_fd_sc_hd__dlygate4sd3_1 hold133 (.A(\gpio_configure[14][1] ),
    .X(net639));
 sky130_fd_sc_hd__dlygate4sd3_1 hold134 (.A(\gpio_configure[5][1] ),
    .X(net640));
 sky130_fd_sc_hd__dlygate4sd3_1 hold135 (.A(\gpio_configure[2][1] ),
    .X(net641));
 sky130_fd_sc_hd__dlygate4sd3_1 hold136 (.A(_3107_),
    .X(net642));
 sky130_fd_sc_hd__dlygate4sd3_1 hold137 (.A(\mgmt_gpio_data_buf[12] ),
    .X(net643));
 sky130_fd_sc_hd__dlygate4sd3_1 hold138 (.A(_1720_),
    .X(net644));
 sky130_fd_sc_hd__dlygate4sd3_1 hold139 (.A(\gpio_configure[6][12] ),
    .X(net645));
 sky130_fd_sc_hd__dlygate4sd3_1 hold140 (.A(_2035_),
    .X(net646));
 sky130_fd_sc_hd__dlygate4sd3_1 hold141 (.A(\gpio_configure[11][12] ),
    .X(net647));
 sky130_fd_sc_hd__dlygate4sd3_1 hold142 (.A(_1757_),
    .X(net648));
 sky130_fd_sc_hd__dlygate4sd3_1 hold143 (.A(\gpio_configure[12][1] ),
    .X(net649));
 sky130_fd_sc_hd__dlygate4sd3_1 hold144 (.A(\gpio_configure[10][1] ),
    .X(net650));
 sky130_fd_sc_hd__dlygate4sd3_1 hold145 (.A(_3189_),
    .X(net651));
 sky130_fd_sc_hd__dlygate4sd3_1 hold146 (.A(_3071_),
    .X(net652));
 sky130_fd_sc_hd__dlygate4sd3_1 hold147 (.A(_0444_),
    .X(net653));
 sky130_fd_sc_hd__dlygate4sd3_1 hold148 (.A(\gpio_configure[19][1] ),
    .X(net654));
 sky130_fd_sc_hd__dlygate4sd3_1 hold149 (.A(\gpio_configure[12][12] ),
    .X(net655));
 sky130_fd_sc_hd__dlygate4sd3_1 hold150 (.A(_1763_),
    .X(net656));
 sky130_fd_sc_hd__dlygate4sd3_1 hold151 (.A(serial_bb_clock),
    .X(net657));
 sky130_fd_sc_hd__dlygate4sd3_1 hold152 (.A(_3051_),
    .X(net658));
 sky130_fd_sc_hd__dlygate4sd3_1 hold153 (.A(_1973_),
    .X(net659));
 sky130_fd_sc_hd__dlygate4sd3_1 hold154 (.A(_0304_),
    .X(net660));
 sky130_fd_sc_hd__dlygate4sd3_1 hold155 (.A(\gpio_configure[36][12] ),
    .X(net661));
 sky130_fd_sc_hd__dlygate4sd3_1 hold156 (.A(_2060_),
    .X(net662));
 sky130_fd_sc_hd__dlygate4sd3_1 hold157 (.A(\gpio_configure[14][12] ),
    .X(net663));
 sky130_fd_sc_hd__dlygate4sd3_1 hold158 (.A(_1775_),
    .X(net664));
 sky130_fd_sc_hd__dlygate4sd3_1 hold159 (.A(\gpio_configure[16][12] ),
    .X(net665));
 sky130_fd_sc_hd__dlygate4sd3_1 hold160 (.A(_2066_),
    .X(net666));
 sky130_fd_sc_hd__dlygate4sd3_1 hold161 (.A(\gpio_configure[20][1] ),
    .X(net667));
 sky130_fd_sc_hd__dlygate4sd3_1 hold162 (.A(\gpio_configure[18][12] ),
    .X(net668));
 sky130_fd_sc_hd__dlygate4sd3_1 hold163 (.A(_1817_),
    .X(net669));
 sky130_fd_sc_hd__dlygate4sd3_1 hold164 (.A(_3024_),
    .X(net670));
 sky130_fd_sc_hd__dlygate4sd3_1 hold165 (.A(\gpio_configure[4][4] ),
    .X(net671));
 sky130_fd_sc_hd__dlygate4sd3_1 hold166 (.A(_3132_),
    .X(net672));
 sky130_fd_sc_hd__dlygate4sd3_1 hold167 (.A(\gpio_configure[5][4] ),
    .X(net673));
 sky130_fd_sc_hd__dlygate4sd3_1 hold168 (.A(_3141_),
    .X(net674));
 sky130_fd_sc_hd__dlygate4sd3_1 hold169 (.A(\gpio_configure[35][12] ),
    .X(net675));
 sky130_fd_sc_hd__dlygate4sd3_1 hold170 (.A(_1794_),
    .X(net676));
 sky130_fd_sc_hd__dlygate4sd3_1 hold171 (.A(\gpio_configure[20][12] ),
    .X(net677));
 sky130_fd_sc_hd__dlygate4sd3_1 hold172 (.A(_1845_),
    .X(net678));
 sky130_fd_sc_hd__dlygate4sd3_1 hold173 (.A(\gpio_configure[27][12] ),
    .X(net679));
 sky130_fd_sc_hd__dlygate4sd3_1 hold174 (.A(_1902_),
    .X(net680));
 sky130_fd_sc_hd__dlygate4sd3_1 hold175 (.A(\gpio_configure[32][1] ),
    .X(net681));
 sky130_fd_sc_hd__dlygate4sd3_1 hold176 (.A(\gpio_configure[34][5] ),
    .X(net682));
 sky130_fd_sc_hd__dlygate4sd3_1 hold177 (.A(_3425_),
    .X(net683));
 sky130_fd_sc_hd__dlygate4sd3_1 hold178 (.A(\gpio_configure[31][5] ),
    .X(net684));
 sky130_fd_sc_hd__dlygate4sd3_1 hold179 (.A(_3397_),
    .X(net685));
 sky130_fd_sc_hd__dlygate4sd3_1 hold180 (.A(\gpio_configure[3][5] ),
    .X(net686));
 sky130_fd_sc_hd__dlygate4sd3_1 hold181 (.A(_3124_),
    .X(net687));
 sky130_fd_sc_hd__dlygate4sd3_1 hold182 (.A(\mgmt_gpio_data_buf[1] ),
    .X(net688));
 sky130_fd_sc_hd__dlygate4sd3_1 hold183 (.A(_3079_),
    .X(net689));
 sky130_fd_sc_hd__dlygate4sd3_1 hold184 (.A(\gpio_configure[34][4] ),
    .X(net690));
 sky130_fd_sc_hd__dlygate4sd3_1 hold185 (.A(_3424_),
    .X(net691));
 sky130_fd_sc_hd__dlygate4sd3_1 hold186 (.A(\gpio_configure[4][12] ),
    .X(net692));
 sky130_fd_sc_hd__dlygate4sd3_1 hold187 (.A(_1745_),
    .X(net693));
 sky130_fd_sc_hd__dlygate4sd3_1 hold188 (.A(\gpio_configure[29][6] ),
    .X(net694));
 sky130_fd_sc_hd__dlygate4sd3_1 hold189 (.A(_3380_),
    .X(net695));
 sky130_fd_sc_hd__dlygate4sd3_1 hold190 (.A(\gpio_configure[36][4] ),
    .X(net696));
 sky130_fd_sc_hd__dlygate4sd3_1 hold191 (.A(_3442_),
    .X(net697));
 sky130_fd_sc_hd__dlygate4sd3_1 hold192 (.A(\gpio_configure[33][4] ),
    .X(net698));
 sky130_fd_sc_hd__dlygate4sd3_1 hold193 (.A(_3415_),
    .X(net699));
 sky130_fd_sc_hd__dlygate4sd3_1 hold194 (.A(\gpio_configure[35][6] ),
    .X(net700));
 sky130_fd_sc_hd__dlygate4sd3_1 hold195 (.A(_3435_),
    .X(net701));
 sky130_fd_sc_hd__dlygate4sd3_1 hold196 (.A(net1728),
    .X(net702));
 sky130_fd_sc_hd__dlygate4sd3_1 hold197 (.A(\wbbd_data[3] ),
    .X(net703));
 sky130_fd_sc_hd__dlygate4sd3_1 hold198 (.A(_1613_),
    .X(net704));
 sky130_fd_sc_hd__dlygate4sd3_1 hold199 (.A(_1957_),
    .X(net705));
 sky130_fd_sc_hd__dlygate4sd3_1 hold200 (.A(net1719),
    .X(net706));
 sky130_fd_sc_hd__dlygate4sd3_1 hold201 (.A(\gpio_configure[28][6] ),
    .X(net707));
 sky130_fd_sc_hd__dlygate4sd3_1 hold202 (.A(_3371_),
    .X(net708));
 sky130_fd_sc_hd__dlygate4sd3_1 hold203 (.A(net1790),
    .X(net709));
 sky130_fd_sc_hd__dlygate4sd3_1 hold204 (.A(net1608),
    .X(net710));
 sky130_fd_sc_hd__dlygate4sd3_1 hold205 (.A(\gpio_configure[0][7] ),
    .X(net711));
 sky130_fd_sc_hd__dlygate4sd3_1 hold206 (.A(_3095_),
    .X(net712));
 sky130_fd_sc_hd__dlygate4sd3_1 hold207 (.A(\gpio_configure[8][7] ),
    .X(net713));
 sky130_fd_sc_hd__dlygate4sd3_1 hold208 (.A(_3176_),
    .X(net714));
 sky130_fd_sc_hd__dlygate4sd3_1 hold209 (.A(\gpio_configure[32][7] ),
    .X(net715));
 sky130_fd_sc_hd__dlygate4sd3_1 hold210 (.A(_3409_),
    .X(net716));
 sky130_fd_sc_hd__dlygate4sd3_1 hold211 (.A(net1635),
    .X(net717));
 sky130_fd_sc_hd__dlygate4sd3_1 hold212 (.A(\gpio_configure[29][5] ),
    .X(net718));
 sky130_fd_sc_hd__dlygate4sd3_1 hold213 (.A(_3379_),
    .X(net719));
 sky130_fd_sc_hd__dlygate4sd3_1 hold214 (.A(\gpio_configure[2][4] ),
    .X(net720));
 sky130_fd_sc_hd__dlygate4sd3_1 hold215 (.A(_3110_),
    .X(net721));
 sky130_fd_sc_hd__dlygate4sd3_1 hold216 (.A(\gpio_configure[10][5] ),
    .X(net722));
 sky130_fd_sc_hd__dlygate4sd3_1 hold217 (.A(_3193_),
    .X(net723));
 sky130_fd_sc_hd__dlygate4sd3_1 hold218 (.A(\gpio_configure[6][5] ),
    .X(net724));
 sky130_fd_sc_hd__dlygate4sd3_1 hold219 (.A(_3152_),
    .X(net725));
 sky130_fd_sc_hd__dlygate4sd3_1 hold220 (.A(\gpio_configure[35][5] ),
    .X(net726));
 sky130_fd_sc_hd__dlygate4sd3_1 hold221 (.A(_3434_),
    .X(net727));
 sky130_fd_sc_hd__dlygate4sd3_1 hold222 (.A(\gpio_configure[5][5] ),
    .X(net728));
 sky130_fd_sc_hd__dlygate4sd3_1 hold223 (.A(_3142_),
    .X(net729));
 sky130_fd_sc_hd__dlygate4sd3_1 hold224 (.A(net1641),
    .X(net730));
 sky130_fd_sc_hd__dlygate4sd3_1 hold225 (.A(\gpio_configure[27][5] ),
    .X(net731));
 sky130_fd_sc_hd__dlygate4sd3_1 hold226 (.A(_3361_),
    .X(net732));
 sky130_fd_sc_hd__dlygate4sd3_1 hold227 (.A(net1714),
    .X(net733));
 sky130_fd_sc_hd__dlygate4sd3_1 hold228 (.A(_3027_),
    .X(net734));
 sky130_fd_sc_hd__dlygate4sd3_1 hold229 (.A(\gpio_configure[25][5] ),
    .X(net735));
 sky130_fd_sc_hd__dlygate4sd3_1 hold230 (.A(_3339_),
    .X(net736));
 sky130_fd_sc_hd__dlygate4sd3_1 hold231 (.A(\gpio_configure[15][5] ),
    .X(net737));
 sky130_fd_sc_hd__dlygate4sd3_1 hold232 (.A(_3242_),
    .X(net738));
 sky130_fd_sc_hd__dlygate4sd3_1 hold233 (.A(\gpio_configure[21][5] ),
    .X(net739));
 sky130_fd_sc_hd__dlygate4sd3_1 hold234 (.A(_3302_),
    .X(net740));
 sky130_fd_sc_hd__dlygate4sd3_1 hold235 (.A(net1643),
    .X(net741));
 sky130_fd_sc_hd__dlygate4sd3_1 hold236 (.A(\gpio_configure[20][5] ),
    .X(net742));
 sky130_fd_sc_hd__dlygate4sd3_1 hold237 (.A(_3292_),
    .X(net743));
 sky130_fd_sc_hd__dlygate4sd3_1 hold238 (.A(\gpio_configure[19][5] ),
    .X(net744));
 sky130_fd_sc_hd__dlygate4sd3_1 hold239 (.A(_3283_),
    .X(net745));
 sky130_fd_sc_hd__dlygate4sd3_1 hold240 (.A(\gpio_configure[19][4] ),
    .X(net746));
 sky130_fd_sc_hd__dlygate4sd3_1 hold241 (.A(net1601),
    .X(net747));
 sky130_fd_sc_hd__dlygate4sd3_1 hold242 (.A(\gpio_configure[4][1] ),
    .X(net748));
 sky130_fd_sc_hd__dlygate4sd3_1 hold243 (.A(_3129_),
    .X(net749));
 sky130_fd_sc_hd__dlygate4sd3_1 hold244 (.A(\gpio_configure[33][5] ),
    .X(net750));
 sky130_fd_sc_hd__dlygate4sd3_1 hold245 (.A(_3416_),
    .X(net751));
 sky130_fd_sc_hd__dlygate4sd3_1 hold246 (.A(\gpio_configure[36][6] ),
    .X(net752));
 sky130_fd_sc_hd__dlygate4sd3_1 hold247 (.A(_3444_),
    .X(net753));
 sky130_fd_sc_hd__dlygate4sd3_1 hold248 (.A(\gpio_configure[22][5] ),
    .X(net754));
 sky130_fd_sc_hd__dlygate4sd3_1 hold249 (.A(_3311_),
    .X(net755));
 sky130_fd_sc_hd__dlygate4sd3_1 hold250 (.A(\gpio_configure[28][5] ),
    .X(net756));
 sky130_fd_sc_hd__dlygate4sd3_1 hold251 (.A(_3370_),
    .X(net757));
 sky130_fd_sc_hd__dlygate4sd3_1 hold252 (.A(\gpio_configure[30][5] ),
    .X(net758));
 sky130_fd_sc_hd__dlygate4sd3_1 hold253 (.A(_3388_),
    .X(net759));
 sky130_fd_sc_hd__dlygate4sd3_1 hold254 (.A(\gpio_configure[25][4] ),
    .X(net760));
 sky130_fd_sc_hd__dlygate4sd3_1 hold255 (.A(_3338_),
    .X(net761));
 sky130_fd_sc_hd__dlygate4sd3_1 hold256 (.A(\gpio_configure[36][5] ),
    .X(net762));
 sky130_fd_sc_hd__dlygate4sd3_1 hold257 (.A(_3443_),
    .X(net763));
 sky130_fd_sc_hd__dlygate4sd3_1 hold258 (.A(\gpio_configure[21][4] ),
    .X(net764));
 sky130_fd_sc_hd__dlygate4sd3_1 hold259 (.A(net1599),
    .X(net765));
 sky130_fd_sc_hd__dlygate4sd3_1 hold260 (.A(\gpio_configure[4][5] ),
    .X(net766));
 sky130_fd_sc_hd__dlygate4sd3_1 hold261 (.A(_3133_),
    .X(net767));
 sky130_fd_sc_hd__dlygate4sd3_1 hold262 (.A(\gpio_configure[18][5] ),
    .X(net768));
 sky130_fd_sc_hd__dlygate4sd3_1 hold263 (.A(_3271_),
    .X(net769));
 sky130_fd_sc_hd__dlygate4sd3_1 hold264 (.A(\gpio_configure[22][4] ),
    .X(net770));
 sky130_fd_sc_hd__dlygate4sd3_1 hold265 (.A(\gpio_configure[7][5] ),
    .X(net771));
 sky130_fd_sc_hd__dlygate4sd3_1 hold266 (.A(_3164_),
    .X(net772));
 sky130_fd_sc_hd__dlygate4sd3_1 hold267 (.A(\gpio_configure[20][4] ),
    .X(net773));
 sky130_fd_sc_hd__dlygate4sd3_1 hold268 (.A(\gpio_configure[7][1] ),
    .X(net774));
 sky130_fd_sc_hd__dlygate4sd3_1 hold269 (.A(_3160_),
    .X(net775));
 sky130_fd_sc_hd__dlygate4sd3_1 hold270 (.A(net1672),
    .X(net776));
 sky130_fd_sc_hd__dlygate4sd3_1 hold271 (.A(\gpio_configure[13][5] ),
    .X(net777));
 sky130_fd_sc_hd__dlygate4sd3_1 hold272 (.A(_3220_),
    .X(net778));
 sky130_fd_sc_hd__dlygate4sd3_1 hold273 (.A(\gpio_configure[11][5] ),
    .X(net779));
 sky130_fd_sc_hd__dlygate4sd3_1 hold274 (.A(_3202_),
    .X(net780));
 sky130_fd_sc_hd__dlygate4sd3_1 hold275 (.A(\gpio_configure[37][5] ),
    .X(net781));
 sky130_fd_sc_hd__dlygate4sd3_1 hold276 (.A(_3452_),
    .X(net782));
 sky130_fd_sc_hd__dlygate4sd3_1 hold277 (.A(\gpio_configure[10][4] ),
    .X(net783));
 sky130_fd_sc_hd__dlygate4sd3_1 hold278 (.A(_3192_),
    .X(net784));
 sky130_fd_sc_hd__dlygate4sd3_1 hold279 (.A(\gpio_configure[12][5] ),
    .X(net785));
 sky130_fd_sc_hd__dlygate4sd3_1 hold280 (.A(_3211_),
    .X(net786));
 sky130_fd_sc_hd__dlygate4sd3_1 hold281 (.A(_3074_),
    .X(net787));
 sky130_fd_sc_hd__dlygate4sd3_1 hold282 (.A(_0447_),
    .X(net788));
 sky130_fd_sc_hd__dlygate4sd3_1 hold283 (.A(\gpio_configure[18][4] ),
    .X(net789));
 sky130_fd_sc_hd__dlygate4sd3_1 hold284 (.A(_3270_),
    .X(net790));
 sky130_fd_sc_hd__dlygate4sd3_1 hold285 (.A(net1647),
    .X(net791));
 sky130_fd_sc_hd__dlygate4sd3_1 hold286 (.A(\gpio_configure[3][4] ),
    .X(net792));
 sky130_fd_sc_hd__dlygate4sd3_1 hold287 (.A(_3122_),
    .X(net793));
 sky130_fd_sc_hd__dlygate4sd3_1 hold288 (.A(net1701),
    .X(net794));
 sky130_fd_sc_hd__dlygate4sd3_1 hold289 (.A(\gpio_configure[6][4] ),
    .X(net795));
 sky130_fd_sc_hd__dlygate4sd3_1 hold290 (.A(_3151_),
    .X(net796));
 sky130_fd_sc_hd__dlygate4sd3_1 hold291 (.A(\gpio_configure[32][5] ),
    .X(net797));
 sky130_fd_sc_hd__dlygate4sd3_1 hold292 (.A(_3407_),
    .X(net798));
 sky130_fd_sc_hd__dlygate4sd3_1 hold293 (.A(\gpio_configure[8][5] ),
    .X(net799));
 sky130_fd_sc_hd__dlygate4sd3_1 hold294 (.A(_3174_),
    .X(net800));
 sky130_fd_sc_hd__dlygate4sd3_1 hold295 (.A(\gpio_configure[3][1] ),
    .X(net801));
 sky130_fd_sc_hd__dlygate4sd3_1 hold296 (.A(_3116_),
    .X(net802));
 sky130_fd_sc_hd__dlygate4sd3_1 hold297 (.A(\gpio_configure[9][5] ),
    .X(net803));
 sky130_fd_sc_hd__dlygate4sd3_1 hold298 (.A(_3183_),
    .X(net804));
 sky130_fd_sc_hd__dlygate4sd3_1 hold299 (.A(\gpio_configure[33][6] ),
    .X(net805));
 sky130_fd_sc_hd__dlygate4sd3_1 hold300 (.A(_3417_),
    .X(net806));
 sky130_fd_sc_hd__dlygate4sd3_1 hold301 (.A(\gpio_configure[17][5] ),
    .X(net807));
 sky130_fd_sc_hd__dlygate4sd3_1 hold302 (.A(_3261_),
    .X(net808));
 sky130_fd_sc_hd__dlygate4sd3_1 hold303 (.A(\gpio_configure[17][4] ),
    .X(net809));
 sky130_fd_sc_hd__dlygate4sd3_1 hold304 (.A(_3260_),
    .X(net810));
 sky130_fd_sc_hd__dlygate4sd3_1 hold305 (.A(\gpio_configure[24][5] ),
    .X(net811));
 sky130_fd_sc_hd__dlygate4sd3_1 hold306 (.A(_3330_),
    .X(net812));
 sky130_fd_sc_hd__dlygate4sd3_1 hold307 (.A(\gpio_configure[7][4] ),
    .X(net813));
 sky130_fd_sc_hd__dlygate4sd3_1 hold308 (.A(_3163_),
    .X(net814));
 sky130_fd_sc_hd__dlygate4sd3_1 hold309 (.A(net1624),
    .X(net815));
 sky130_fd_sc_hd__dlygate4sd3_1 hold310 (.A(net1603),
    .X(net816));
 sky130_fd_sc_hd__dlygate4sd3_1 hold311 (.A(\gpio_configure[14][5] ),
    .X(net817));
 sky130_fd_sc_hd__dlygate4sd3_1 hold312 (.A(_3233_),
    .X(net818));
 sky130_fd_sc_hd__dlygate4sd3_1 hold313 (.A(_1676_),
    .X(net819));
 sky130_fd_sc_hd__dlygate4sd3_1 hold314 (.A(\gpio_configure[9][4] ),
    .X(net820));
 sky130_fd_sc_hd__dlygate4sd3_1 hold315 (.A(_3182_),
    .X(net821));
 sky130_fd_sc_hd__dlygate4sd3_1 hold316 (.A(\gpio_configure[1][1] ),
    .X(net822));
 sky130_fd_sc_hd__dlygate4sd3_1 hold317 (.A(_3098_),
    .X(net823));
 sky130_fd_sc_hd__dlygate4sd3_1 hold318 (.A(\gpio_configure[11][4] ),
    .X(net824));
 sky130_fd_sc_hd__dlygate4sd3_1 hold319 (.A(_3201_),
    .X(net825));
 sky130_fd_sc_hd__dlygate4sd3_1 hold320 (.A(\gpio_configure[37][6] ),
    .X(net826));
 sky130_fd_sc_hd__dlygate4sd3_1 hold321 (.A(_3453_),
    .X(net827));
 sky130_fd_sc_hd__dlygate4sd3_1 hold322 (.A(\gpio_configure[0][6] ),
    .X(net828));
 sky130_fd_sc_hd__dlygate4sd3_1 hold323 (.A(_3094_),
    .X(net829));
 sky130_fd_sc_hd__dlygate4sd3_1 hold324 (.A(\gpio_configure[34][6] ),
    .X(net830));
 sky130_fd_sc_hd__dlygate4sd3_1 hold325 (.A(_3426_),
    .X(net831));
 sky130_fd_sc_hd__dlygate4sd3_1 hold326 (.A(net1679),
    .X(net832));
 sky130_fd_sc_hd__dlygate4sd3_1 hold327 (.A(_3043_),
    .X(net833));
 sky130_fd_sc_hd__dlygate4sd3_1 hold328 (.A(\gpio_configure[34][12] ),
    .X(net834));
 sky130_fd_sc_hd__dlygate4sd3_1 hold329 (.A(_1808_),
    .X(net835));
 sky130_fd_sc_hd__dlygate4sd3_1 hold330 (.A(\gpio_configure[0][5] ),
    .X(net836));
 sky130_fd_sc_hd__dlygate4sd3_1 hold331 (.A(_3093_),
    .X(net837));
 sky130_fd_sc_hd__dlygate4sd3_1 hold332 (.A(\gpio_configure[16][5] ),
    .X(net838));
 sky130_fd_sc_hd__dlygate4sd3_1 hold333 (.A(_3252_),
    .X(net839));
 sky130_fd_sc_hd__dlygate4sd3_1 hold334 (.A(net1612),
    .X(net840));
 sky130_fd_sc_hd__dlygate4sd3_1 hold335 (.A(net1716),
    .X(net841));
 sky130_fd_sc_hd__dlygate4sd3_1 hold336 (.A(net1665),
    .X(net842));
 sky130_fd_sc_hd__dlygate4sd3_1 hold337 (.A(net1619),
    .X(net843));
 sky130_fd_sc_hd__dlygate4sd3_1 hold338 (.A(_1673_),
    .X(net844));
 sky130_fd_sc_hd__dlygate4sd3_1 hold339 (.A(_3025_),
    .X(net845));
 sky130_fd_sc_hd__dlygate4sd3_1 hold340 (.A(_3337_),
    .X(net846));
 sky130_fd_sc_hd__dlygate4sd3_1 hold341 (.A(_3010_),
    .X(net847));
 sky130_fd_sc_hd__dlygate4sd3_1 hold342 (.A(_3281_),
    .X(net848));
 sky130_fd_sc_hd__dlygate4sd3_1 hold343 (.A(_3300_),
    .X(net849));
 sky130_fd_sc_hd__dlygate4sd3_1 hold344 (.A(_3016_),
    .X(net850));
 sky130_fd_sc_hd__dlygate4sd3_1 hold345 (.A(net1687),
    .X(net851));
 sky130_fd_sc_hd__dlygate4sd3_1 hold346 (.A(_3441_),
    .X(net852));
 sky130_fd_sc_hd__dlygate4sd3_1 hold347 (.A(_3259_),
    .X(net853));
 sky130_fd_sc_hd__dlygate4sd3_1 hold348 (.A(_3240_),
    .X(net854));
 sky130_fd_sc_hd__dlygate4sd3_1 hold349 (.A(_3290_),
    .X(net855));
 sky130_fd_sc_hd__dlygate4sd3_1 hold350 (.A(net1731),
    .X(net856));
 sky130_fd_sc_hd__dlygate4sd3_1 hold351 (.A(_3432_),
    .X(net857));
 sky130_fd_sc_hd__dlygate4sd3_1 hold352 (.A(\gpio_configure[1][4] ),
    .X(net858));
 sky130_fd_sc_hd__dlygate4sd3_1 hold353 (.A(_3101_),
    .X(net859));
 sky130_fd_sc_hd__dlygate4sd3_1 hold354 (.A(net1773),
    .X(net860));
 sky130_fd_sc_hd__dlygate4sd3_1 hold355 (.A(net1746),
    .X(net861));
 sky130_fd_sc_hd__dlygate4sd3_1 hold356 (.A(\gpio_configure[3][12] ),
    .X(net862));
 sky130_fd_sc_hd__dlygate4sd3_1 hold357 (.A(_2000_),
    .X(net863));
 sky130_fd_sc_hd__dlygate4sd3_1 hold358 (.A(\gpio_configure[8][6] ),
    .X(net864));
 sky130_fd_sc_hd__dlygate4sd3_1 hold359 (.A(_3175_),
    .X(net865));
 sky130_fd_sc_hd__dlygate4sd3_1 hold360 (.A(\gpio_configure[2][12] ),
    .X(net866));
 sky130_fd_sc_hd__dlygate4sd3_1 hold361 (.A(_1982_),
    .X(net867));
 sky130_fd_sc_hd__dlygate4sd3_1 hold362 (.A(_3423_),
    .X(net868));
 sky130_fd_sc_hd__dlygate4sd3_1 hold363 (.A(\wbbd_addr[2] ),
    .X(net869));
 sky130_fd_sc_hd__dlygate4sd3_1 hold364 (.A(_3414_),
    .X(net870));
 sky130_fd_sc_hd__dlygate4sd3_1 hold365 (.A(_3269_),
    .X(net871));
 sky130_fd_sc_hd__dlygate4sd3_1 hold366 (.A(net1711),
    .X(net872));
 sky130_fd_sc_hd__dlygate4sd3_1 hold367 (.A(\mgmt_gpio_data_buf[11] ),
    .X(net873));
 sky130_fd_sc_hd__dlygate4sd3_1 hold368 (.A(_1719_),
    .X(net874));
 sky130_fd_sc_hd__dlygate4sd3_1 hold369 (.A(_1688_),
    .X(net875));
 sky130_fd_sc_hd__dlygate4sd3_1 hold370 (.A(net1649),
    .X(net876));
 sky130_fd_sc_hd__dlygate4sd3_1 hold371 (.A(_3368_),
    .X(net877));
 sky130_fd_sc_hd__dlygate4sd3_1 hold372 (.A(\gpio_configure[28][4] ),
    .X(net878));
 sky130_fd_sc_hd__dlygate4sd3_1 hold373 (.A(net1696),
    .X(net879));
 sky130_fd_sc_hd__dlygate4sd3_1 hold374 (.A(\mgmt_gpio_data_buf[3] ),
    .X(net880));
 sky130_fd_sc_hd__dlygate4sd3_1 hold375 (.A(_3081_),
    .X(net881));
 sky130_fd_sc_hd__dlygate4sd3_1 hold376 (.A(_3377_),
    .X(net882));
 sky130_fd_sc_hd__dlygate4sd3_1 hold377 (.A(_1690_),
    .X(net883));
 sky130_fd_sc_hd__dlygate4sd3_1 hold378 (.A(net1760),
    .X(net884));
 sky130_fd_sc_hd__dlygate4sd3_1 hold379 (.A(\gpio_configure[32][6] ),
    .X(net885));
 sky130_fd_sc_hd__dlygate4sd3_1 hold380 (.A(_3408_),
    .X(net886));
 sky130_fd_sc_hd__dlygate4sd3_1 hold381 (.A(net1638),
    .X(net887));
 sky130_fd_sc_hd__dlygate4sd3_1 hold382 (.A(_3359_),
    .X(net888));
 sky130_fd_sc_hd__dlygate4sd3_1 hold383 (.A(\mgmt_gpio_data_buf[19] ),
    .X(net889));
 sky130_fd_sc_hd__dlygate4sd3_1 hold384 (.A(_1706_),
    .X(net890));
 sky130_fd_sc_hd__dlygate4sd3_1 hold385 (.A(_3026_),
    .X(net891));
 sky130_fd_sc_hd__dlygate4sd3_1 hold386 (.A(net1735),
    .X(net892));
 sky130_fd_sc_hd__dlygate4sd3_1 hold387 (.A(net1770),
    .X(net893));
 sky130_fd_sc_hd__dlygate4sd3_1 hold388 (.A(\gpio_configure[18][11] ),
    .X(net894));
 sky130_fd_sc_hd__dlygate4sd3_1 hold389 (.A(\gpio_configure[13][1] ),
    .X(net895));
 sky130_fd_sc_hd__dlygate4sd3_1 hold390 (.A(\gpio_configure[30][11] ),
    .X(net896));
 sky130_fd_sc_hd__dlygate4sd3_1 hold391 (.A(_1972_),
    .X(net897));
 sky130_fd_sc_hd__dlygate4sd3_1 hold392 (.A(_0303_),
    .X(net898));
 sky130_fd_sc_hd__dlygate4sd3_1 hold393 (.A(\gpio_configure[11][1] ),
    .X(net899));
 sky130_fd_sc_hd__dlygate4sd3_1 hold394 (.A(\gpio_configure[15][1] ),
    .X(net900));
 sky130_fd_sc_hd__dlygate4sd3_1 hold395 (.A(net1774),
    .X(net901));
 sky130_fd_sc_hd__dlygate4sd3_1 hold396 (.A(\gpio_configure[20][11] ),
    .X(net902));
 sky130_fd_sc_hd__dlygate4sd3_1 hold397 (.A(net1762),
    .X(net903));
 sky130_fd_sc_hd__dlygate4sd3_1 hold398 (.A(net1753),
    .X(net904));
 sky130_fd_sc_hd__dlygate4sd3_1 hold399 (.A(net1675),
    .X(net905));
 sky130_fd_sc_hd__dlygate4sd3_1 hold400 (.A(\gpio_configure[4][11] ),
    .X(net906));
 sky130_fd_sc_hd__dlygate4sd3_1 hold401 (.A(_1744_),
    .X(net907));
 sky130_fd_sc_hd__dlygate4sd3_1 hold402 (.A(\gpio_configure[14][2] ),
    .X(net908));
 sky130_fd_sc_hd__dlygate4sd3_1 hold403 (.A(_3227_),
    .X(net909));
 sky130_fd_sc_hd__dlygate4sd3_1 hold404 (.A(\gpio_configure[28][11] ),
    .X(net910));
 sky130_fd_sc_hd__dlygate4sd3_1 hold405 (.A(net1614),
    .X(net911));
 sky130_fd_sc_hd__dlygate4sd3_1 hold406 (.A(net1771),
    .X(net912));
 sky130_fd_sc_hd__dlygate4sd3_1 hold407 (.A(\gpio_configure[23][11] ),
    .X(net913));
 sky130_fd_sc_hd__dlygate4sd3_1 hold408 (.A(\gpio_configure[25][2] ),
    .X(net914));
 sky130_fd_sc_hd__dlygate4sd3_1 hold409 (.A(_3336_),
    .X(net915));
 sky130_fd_sc_hd__dlygate4sd3_1 hold410 (.A(net1777),
    .X(net916));
 sky130_fd_sc_hd__dlygate4sd3_1 hold411 (.A(\gpio_configure[7][11] ),
    .X(net917));
 sky130_fd_sc_hd__dlygate4sd3_1 hold412 (.A(_2040_),
    .X(net918));
 sky130_fd_sc_hd__dlygate4sd3_1 hold413 (.A(net1782),
    .X(net919));
 sky130_fd_sc_hd__dlygate4sd3_1 hold414 (.A(\gpio_configure[27][2] ),
    .X(net920));
 sky130_fd_sc_hd__dlygate4sd3_1 hold415 (.A(_3358_),
    .X(net921));
 sky130_fd_sc_hd__dlygate4sd3_1 hold416 (.A(_3072_),
    .X(net922));
 sky130_fd_sc_hd__dlygate4sd3_1 hold417 (.A(_0445_),
    .X(net923));
 sky130_fd_sc_hd__dlygate4sd3_1 hold418 (.A(net1646),
    .X(net924));
 sky130_fd_sc_hd__dlygate4sd3_1 hold419 (.A(\gpio_configure[0][11] ),
    .X(net925));
 sky130_fd_sc_hd__dlygate4sd3_1 hold420 (.A(_1729_),
    .X(net926));
 sky130_fd_sc_hd__dlygate4sd3_1 hold421 (.A(net1677),
    .X(net927));
 sky130_fd_sc_hd__dlygate4sd3_1 hold422 (.A(net1737),
    .X(net928));
 sky130_fd_sc_hd__dlygate4sd3_1 hold423 (.A(net1789),
    .X(net929));
 sky130_fd_sc_hd__dlygate4sd3_1 hold424 (.A(_3181_),
    .X(net930));
 sky130_fd_sc_hd__dlygate4sd3_1 hold425 (.A(net1685),
    .X(net931));
 sky130_fd_sc_hd__dlygate4sd3_1 hold426 (.A(\gpio_configure[28][2] ),
    .X(net932));
 sky130_fd_sc_hd__dlygate4sd3_1 hold427 (.A(_3367_),
    .X(net933));
 sky130_fd_sc_hd__dlygate4sd3_1 hold428 (.A(_1686_),
    .X(net934));
 sky130_fd_sc_hd__dlygate4sd3_1 hold429 (.A(_3191_),
    .X(net935));
 sky130_fd_sc_hd__dlygate4sd3_1 hold430 (.A(net1780),
    .X(net936));
 sky130_fd_sc_hd__dlygate4sd3_1 hold431 (.A(\wbbd_data[0] ),
    .X(net937));
 sky130_fd_sc_hd__dlygate4sd3_1 hold432 (.A(_1596_),
    .X(net938));
 sky130_fd_sc_hd__dlygate4sd3_1 hold433 (.A(_1731_),
    .X(net939));
 sky130_fd_sc_hd__dlygate4sd3_1 hold434 (.A(net1695),
    .X(net940));
 sky130_fd_sc_hd__dlygate4sd3_1 hold435 (.A(net1726),
    .X(net941));
 sky130_fd_sc_hd__dlygate4sd3_1 hold436 (.A(net1631),
    .X(net942));
 sky130_fd_sc_hd__dlygate4sd3_1 hold437 (.A(\gpio_configure[1][11] ),
    .X(net943));
 sky130_fd_sc_hd__dlygate4sd3_1 hold438 (.A(_1737_),
    .X(net944));
 sky130_fd_sc_hd__dlygate4sd3_1 hold439 (.A(\gpio_configure[18][9] ),
    .X(net945));
 sky130_fd_sc_hd__dlygate4sd3_1 hold440 (.A(_3150_),
    .X(net946));
 sky130_fd_sc_hd__dlygate4sd3_1 hold441 (.A(_1970_),
    .X(net947));
 sky130_fd_sc_hd__dlygate4sd3_1 hold442 (.A(_0301_),
    .X(net948));
 sky130_fd_sc_hd__dlygate4sd3_1 hold443 (.A(_1667_),
    .X(net949));
 sky130_fd_sc_hd__dlygate4sd3_1 hold444 (.A(net1734),
    .X(net950));
 sky130_fd_sc_hd__dlygate4sd3_1 hold445 (.A(\gpio_configure[6][11] ),
    .X(net951));
 sky130_fd_sc_hd__dlygate4sd3_1 hold446 (.A(_2033_),
    .X(net952));
 sky130_fd_sc_hd__dlygate4sd3_1 hold447 (.A(_1684_),
    .X(net953));
 sky130_fd_sc_hd__dlygate4sd3_1 hold448 (.A(net1659),
    .X(net954));
 sky130_fd_sc_hd__dlygate4sd3_1 hold449 (.A(\gpio_configure[37][11] ),
    .X(net955));
 sky130_fd_sc_hd__dlygate4sd3_1 hold450 (.A(\mgmt_gpio_data_buf[23] ),
    .X(net956));
 sky130_fd_sc_hd__dlygate4sd3_1 hold451 (.A(_1713_),
    .X(net957));
 sky130_fd_sc_hd__dlygate4sd3_1 hold452 (.A(_1663_),
    .X(net958));
 sky130_fd_sc_hd__dlygate4sd3_1 hold453 (.A(net1776),
    .X(net959));
 sky130_fd_sc_hd__dlygate4sd3_1 hold454 (.A(net1663),
    .X(net960));
 sky130_fd_sc_hd__dlygate4sd3_1 hold455 (.A(net1751),
    .X(net961));
 sky130_fd_sc_hd__dlygate4sd3_1 hold456 (.A(\mgmt_gpio_data_buf[18] ),
    .X(net962));
 sky130_fd_sc_hd__dlygate4sd3_1 hold457 (.A(_1705_),
    .X(net963));
 sky130_fd_sc_hd__dlygate4sd3_1 hold458 (.A(\gpio_configure[28][9] ),
    .X(net964));
 sky130_fd_sc_hd__dlygate4sd3_1 hold459 (.A(net1784),
    .X(net965));
 sky130_fd_sc_hd__dlygate4sd3_1 hold460 (.A(_3073_),
    .X(net966));
 sky130_fd_sc_hd__dlygate4sd3_1 hold461 (.A(_0446_),
    .X(net967));
 sky130_fd_sc_hd__dlygate4sd3_1 hold462 (.A(\gpio_configure[26][9] ),
    .X(net968));
 sky130_fd_sc_hd__dlygate4sd3_1 hold463 (.A(\gpio_configure[4][9] ),
    .X(net969));
 sky130_fd_sc_hd__dlygate4sd3_1 hold464 (.A(_1742_),
    .X(net970));
 sky130_fd_sc_hd__dlygate4sd3_1 hold465 (.A(net1781),
    .X(net971));
 sky130_fd_sc_hd__dlygate4sd3_1 hold466 (.A(net1787),
    .X(net972));
 sky130_fd_sc_hd__dlygate4sd3_1 hold467 (.A(net1640),
    .X(net973));
 sky130_fd_sc_hd__dlygate4sd3_1 hold468 (.A(net1660),
    .X(net974));
 sky130_fd_sc_hd__dlygate4sd3_1 hold469 (.A(\mgmt_gpio_data_buf[15] ),
    .X(net975));
 sky130_fd_sc_hd__dlygate4sd3_1 hold470 (.A(_1723_),
    .X(net976));
 sky130_fd_sc_hd__dlygate4sd3_1 hold471 (.A(\mgmt_gpio_data_buf[17] ),
    .X(net977));
 sky130_fd_sc_hd__dlygate4sd3_1 hold472 (.A(_1704_),
    .X(net978));
 sky130_fd_sc_hd__dlygate4sd3_1 hold473 (.A(\gpio_configure[10][10] ),
    .X(net979));
 sky130_fd_sc_hd__dlygate4sd3_1 hold474 (.A(_1749_),
    .X(net980));
 sky130_fd_sc_hd__dlygate4sd3_1 hold475 (.A(\gpio_configure[36][1] ),
    .X(net981));
 sky130_fd_sc_hd__dlygate4sd3_1 hold476 (.A(\gpio_configure[34][1] ),
    .X(net982));
 sky130_fd_sc_hd__dlygate4sd3_1 hold477 (.A(\gpio_configure[0][9] ),
    .X(net983));
 sky130_fd_sc_hd__dlygate4sd3_1 hold478 (.A(_1727_),
    .X(net984));
 sky130_fd_sc_hd__dlygate4sd3_1 hold479 (.A(\gpio_configure[1][9] ),
    .X(net985));
 sky130_fd_sc_hd__dlygate4sd3_1 hold480 (.A(_1735_),
    .X(net986));
 sky130_fd_sc_hd__dlygate4sd3_1 hold481 (.A(_1976_),
    .X(net987));
 sky130_fd_sc_hd__dlygate4sd3_1 hold482 (.A(_0307_),
    .X(net988));
 sky130_fd_sc_hd__dlygate4sd3_1 hold483 (.A(\gpio_configure[7][9] ),
    .X(net989));
 sky130_fd_sc_hd__dlygate4sd3_1 hold484 (.A(_2038_),
    .X(net990));
 sky130_fd_sc_hd__dlygate4sd3_1 hold485 (.A(net1704),
    .X(net991));
 sky130_fd_sc_hd__dlygate4sd3_1 hold486 (.A(\mgmt_gpio_data_buf[2] ),
    .X(net992));
 sky130_fd_sc_hd__dlygate4sd3_1 hold487 (.A(_3080_),
    .X(net993));
 sky130_fd_sc_hd__dlygate4sd3_1 hold488 (.A(\gpio_configure[33][2] ),
    .X(net994));
 sky130_fd_sc_hd__dlygate4sd3_1 hold489 (.A(_3413_),
    .X(net995));
 sky130_fd_sc_hd__dlygate4sd3_1 hold490 (.A(\gpio_configure[36][11] ),
    .X(net996));
 sky130_fd_sc_hd__dlygate4sd3_1 hold491 (.A(\gpio_configure[11][10] ),
    .X(net997));
 sky130_fd_sc_hd__dlygate4sd3_1 hold492 (.A(_1755_),
    .X(net998));
 sky130_fd_sc_hd__dlygate4sd3_1 hold493 (.A(_3021_),
    .X(net999));
 sky130_fd_sc_hd__dlygate4sd3_1 hold494 (.A(net1698),
    .X(net1000));
 sky130_fd_sc_hd__dlygate4sd3_1 hold495 (.A(net1688),
    .X(net1001));
 sky130_fd_sc_hd__dlygate4sd3_1 hold496 (.A(\gpio_configure[36][2] ),
    .X(net1002));
 sky130_fd_sc_hd__dlygate4sd3_1 hold497 (.A(_3440_),
    .X(net1003));
 sky130_fd_sc_hd__dlygate4sd3_1 hold498 (.A(net1700),
    .X(net1004));
 sky130_fd_sc_hd__dlygate4sd3_1 hold499 (.A(\gpio_configure[33][1] ),
    .X(net1005));
 sky130_fd_sc_hd__dlygate4sd3_1 hold500 (.A(net1670),
    .X(net1006));
 sky130_fd_sc_hd__dlygate4sd3_1 hold501 (.A(\gpio_configure[34][10] ),
    .X(net1007));
 sky130_fd_sc_hd__dlygate4sd3_1 hold502 (.A(_1806_),
    .X(net1008));
 sky130_fd_sc_hd__dlygate4sd3_1 hold503 (.A(\gpio_configure[32][2] ),
    .X(net1009));
 sky130_fd_sc_hd__dlygate4sd3_1 hold504 (.A(_3404_),
    .X(net1010));
 sky130_fd_sc_hd__dlygate4sd3_1 hold505 (.A(net1689),
    .X(net1011));
 sky130_fd_sc_hd__dlygate4sd3_1 hold506 (.A(\mgmt_gpio_data_buf[10] ),
    .X(net1012));
 sky130_fd_sc_hd__dlygate4sd3_1 hold507 (.A(_1718_),
    .X(net1013));
 sky130_fd_sc_hd__dlygate4sd3_1 hold508 (.A(\gpio_configure[4][10] ),
    .X(net1014));
 sky130_fd_sc_hd__dlygate4sd3_1 hold509 (.A(_1743_),
    .X(net1015));
 sky130_fd_sc_hd__dlygate4sd3_1 hold510 (.A(\gpio_configure[34][2] ),
    .X(net1016));
 sky130_fd_sc_hd__dlygate4sd3_1 hold511 (.A(_3422_),
    .X(net1017));
 sky130_fd_sc_hd__dlygate4sd3_1 hold512 (.A(\gpio_configure[16][10] ),
    .X(net1018));
 sky130_fd_sc_hd__dlygate4sd3_1 hold513 (.A(_2064_),
    .X(net1019));
 sky130_fd_sc_hd__dlygate4sd3_1 hold514 (.A(\gpio_configure[26][10] ),
    .X(net1020));
 sky130_fd_sc_hd__dlygate4sd3_1 hold515 (.A(_1612_),
    .X(net1021));
 sky130_fd_sc_hd__dlygate4sd3_1 hold516 (.A(net1598),
    .X(net1022));
 sky130_fd_sc_hd__dlygate4sd3_1 hold517 (.A(\gpio_configure[35][1] ),
    .X(net1023));
 sky130_fd_sc_hd__dlygate4sd3_1 hold518 (.A(\mgmt_gpio_data_buf[9] ),
    .X(net1024));
 sky130_fd_sc_hd__dlygate4sd3_1 hold519 (.A(_1717_),
    .X(net1025));
 sky130_fd_sc_hd__dlygate4sd3_1 hold520 (.A(\gpio_configure[15][7] ),
    .X(net1026));
 sky130_fd_sc_hd__dlygate4sd3_1 hold521 (.A(_3244_),
    .X(net1027));
 sky130_fd_sc_hd__dlygate4sd3_1 hold522 (.A(net1722),
    .X(net1028));
 sky130_fd_sc_hd__dlygate4sd3_1 hold523 (.A(_1971_),
    .X(net1029));
 sky130_fd_sc_hd__dlygate4sd3_1 hold524 (.A(_0302_),
    .X(net1030));
 sky130_fd_sc_hd__dlygate4sd3_1 hold525 (.A(net1741),
    .X(net1031));
 sky130_fd_sc_hd__dlygate4sd3_1 hold526 (.A(net1767),
    .X(net1032));
 sky130_fd_sc_hd__dlygate4sd3_1 hold527 (.A(\gpio_configure[7][7] ),
    .X(net1033));
 sky130_fd_sc_hd__dlygate4sd3_1 hold528 (.A(_3166_),
    .X(net1034));
 sky130_fd_sc_hd__dlygate4sd3_1 hold529 (.A(net1636),
    .X(net1035));
 sky130_fd_sc_hd__dlygate4sd3_1 hold530 (.A(\gpio_configure[13][7] ),
    .X(net1036));
 sky130_fd_sc_hd__dlygate4sd3_1 hold531 (.A(_3222_),
    .X(net1037));
 sky130_fd_sc_hd__dlygate4sd3_1 hold532 (.A(net1763),
    .X(net1038));
 sky130_fd_sc_hd__dlygate4sd3_1 hold533 (.A(\gpio_configure[11][7] ),
    .X(net1039));
 sky130_fd_sc_hd__dlygate4sd3_1 hold534 (.A(_3204_),
    .X(net1040));
 sky130_fd_sc_hd__dlygate4sd3_1 hold535 (.A(\gpio_configure[35][10] ),
    .X(net1041));
 sky130_fd_sc_hd__dlygate4sd3_1 hold536 (.A(_1792_),
    .X(net1042));
 sky130_fd_sc_hd__dlygate4sd3_1 hold537 (.A(\gpio_configure[37][1] ),
    .X(net1043));
 sky130_fd_sc_hd__dlygate4sd3_1 hold538 (.A(\gpio_configure[21][10] ),
    .X(net1044));
 sky130_fd_sc_hd__dlygate4sd3_1 hold539 (.A(_1855_),
    .X(net1045));
 sky130_fd_sc_hd__dlygate4sd3_1 hold540 (.A(\gpio_configure[12][10] ),
    .X(net1046));
 sky130_fd_sc_hd__dlygate4sd3_1 hold541 (.A(_1761_),
    .X(net1047));
 sky130_fd_sc_hd__dlygate4sd3_1 hold542 (.A(\gpio_configure[14][10] ),
    .X(net1048));
 sky130_fd_sc_hd__dlygate4sd3_1 hold543 (.A(_1773_),
    .X(net1049));
 sky130_fd_sc_hd__dlygate4sd3_1 hold544 (.A(\gpio_configure[3][9] ),
    .X(net1050));
 sky130_fd_sc_hd__dlygate4sd3_1 hold545 (.A(_1997_),
    .X(net1051));
 sky130_fd_sc_hd__dlygate4sd3_1 hold546 (.A(net1759),
    .X(net1052));
 sky130_fd_sc_hd__dlygate4sd3_1 hold547 (.A(\gpio_configure[7][12] ),
    .X(net1053));
 sky130_fd_sc_hd__dlygate4sd3_1 hold548 (.A(_2041_),
    .X(net1054));
 sky130_fd_sc_hd__dlygate4sd3_1 hold549 (.A(_3022_),
    .X(net1055));
 sky130_fd_sc_hd__dlygate4sd3_1 hold550 (.A(net1778),
    .X(net1056));
 sky130_fd_sc_hd__dlygate4sd3_1 hold551 (.A(\gpio_configure[8][10] ),
    .X(net1057));
 sky130_fd_sc_hd__dlygate4sd3_1 hold552 (.A(_2045_),
    .X(net1058));
 sky130_fd_sc_hd__dlygate4sd3_1 hold553 (.A(net1743),
    .X(net1059));
 sky130_fd_sc_hd__dlygate4sd3_1 hold554 (.A(\gpio_configure[6][9] ),
    .X(net1060));
 sky130_fd_sc_hd__dlygate4sd3_1 hold555 (.A(_2029_),
    .X(net1061));
 sky130_fd_sc_hd__dlygate4sd3_1 hold556 (.A(\gpio_configure[16][9] ),
    .X(net1062));
 sky130_fd_sc_hd__dlygate4sd3_1 hold557 (.A(\wbbd_data[2] ),
    .X(net1063));
 sky130_fd_sc_hd__dlygate4sd3_1 hold558 (.A(_1609_),
    .X(net1064));
 sky130_fd_sc_hd__dlygate4sd3_1 hold559 (.A(_2031_),
    .X(net1065));
 sky130_fd_sc_hd__dlygate4sd3_1 hold560 (.A(\gpio_configure[7][2] ),
    .X(net1066));
 sky130_fd_sc_hd__dlygate4sd3_1 hold561 (.A(_3161_),
    .X(net1067));
 sky130_fd_sc_hd__dlygate4sd3_1 hold562 (.A(\gpio_configure[6][7] ),
    .X(net1068));
 sky130_fd_sc_hd__dlygate4sd3_1 hold563 (.A(_3155_),
    .X(net1069));
 sky130_fd_sc_hd__dlygate4sd3_1 hold564 (.A(\gpio_configure[17][7] ),
    .X(net1070));
 sky130_fd_sc_hd__dlygate4sd3_1 hold565 (.A(_3264_),
    .X(net1071));
 sky130_fd_sc_hd__dlygate4sd3_1 hold566 (.A(net1786),
    .X(net1072));
 sky130_fd_sc_hd__dlygate4sd3_1 hold567 (.A(\mgmt_gpio_data_buf[7] ),
    .X(net1073));
 sky130_fd_sc_hd__dlygate4sd3_1 hold568 (.A(_3085_),
    .X(net1074));
 sky130_fd_sc_hd__dlygate4sd3_1 hold569 (.A(\gpio_configure[29][10] ),
    .X(net1075));
 sky130_fd_sc_hd__dlygate4sd3_1 hold570 (.A(\gpio_configure[4][2] ),
    .X(net1076));
 sky130_fd_sc_hd__dlygate4sd3_1 hold571 (.A(_3130_),
    .X(net1077));
 sky130_fd_sc_hd__dlygate4sd3_1 hold572 (.A(\gpio_configure[18][10] ),
    .X(net1078));
 sky130_fd_sc_hd__dlygate4sd3_1 hold573 (.A(net1709),
    .X(net1079));
 sky130_fd_sc_hd__dlygate4sd3_1 hold574 (.A(\gpio_configure[0][1] ),
    .X(net1080));
 sky130_fd_sc_hd__dlygate4sd3_1 hold575 (.A(_1694_),
    .X(net1081));
 sky130_fd_sc_hd__dlygate4sd3_1 hold576 (.A(net1645),
    .X(net1082));
 sky130_fd_sc_hd__dlygate4sd3_1 hold577 (.A(\gpio_configure[19][10] ),
    .X(net1083));
 sky130_fd_sc_hd__dlygate4sd3_1 hold578 (.A(\gpio_configure[20][10] ),
    .X(net1084));
 sky130_fd_sc_hd__dlygate4sd3_1 hold579 (.A(\gpio_configure[3][10] ),
    .X(net1085));
 sky130_fd_sc_hd__dlygate4sd3_1 hold580 (.A(_1998_),
    .X(net1086));
 sky130_fd_sc_hd__dlygate4sd3_1 hold581 (.A(_1687_),
    .X(net1087));
 sky130_fd_sc_hd__dlygate4sd3_1 hold582 (.A(\gpio_configure[27][10] ),
    .X(net1088));
 sky130_fd_sc_hd__dlygate4sd3_1 hold583 (.A(net1768),
    .X(net1089));
 sky130_fd_sc_hd__dlygate4sd3_1 hold584 (.A(\gpio_configure[23][7] ),
    .X(net1090));
 sky130_fd_sc_hd__dlygate4sd3_1 hold585 (.A(_3322_),
    .X(net1091));
 sky130_fd_sc_hd__dlygate4sd3_1 hold586 (.A(\gpio_configure[28][7] ),
    .X(net1092));
 sky130_fd_sc_hd__dlygate4sd3_1 hold587 (.A(_3372_),
    .X(net1093));
 sky130_fd_sc_hd__dlygate4sd3_1 hold588 (.A(net1633),
    .X(net1094));
 sky130_fd_sc_hd__dlygate4sd3_1 hold589 (.A(_3054_),
    .X(net1095));
 sky130_fd_sc_hd__dlygate4sd3_1 hold590 (.A(_0433_),
    .X(net1096));
 sky130_fd_sc_hd__dlygate4sd3_1 hold591 (.A(net1676),
    .X(net1097));
 sky130_fd_sc_hd__dlygate4sd3_1 hold592 (.A(\gpio_configure[0][10] ),
    .X(net1098));
 sky130_fd_sc_hd__dlygate4sd3_1 hold593 (.A(_1728_),
    .X(net1099));
 sky130_fd_sc_hd__dlygate4sd3_1 hold594 (.A(net1682),
    .X(net1100));
 sky130_fd_sc_hd__dlygate4sd3_1 hold595 (.A(\gpio_configure[20][7] ),
    .X(net1101));
 sky130_fd_sc_hd__dlygate4sd3_1 hold596 (.A(_3294_),
    .X(net1102));
 sky130_fd_sc_hd__dlygate4sd3_1 hold597 (.A(\gpio_configure[30][10] ),
    .X(net1103));
 sky130_fd_sc_hd__dlygate4sd3_1 hold598 (.A(\gpio_configure[19][7] ),
    .X(net1104));
 sky130_fd_sc_hd__dlygate4sd3_1 hold599 (.A(_3285_),
    .X(net1105));
 sky130_fd_sc_hd__dlygate4sd3_1 hold600 (.A(net1739),
    .X(net1106));
 sky130_fd_sc_hd__dlygate4sd3_1 hold601 (.A(\gpio_configure[1][10] ),
    .X(net1107));
 sky130_fd_sc_hd__dlygate4sd3_1 hold602 (.A(_1736_),
    .X(net1108));
 sky130_fd_sc_hd__dlygate4sd3_1 hold603 (.A(\gpio_configure[27][7] ),
    .X(net1109));
 sky130_fd_sc_hd__dlygate4sd3_1 hold604 (.A(_3363_),
    .X(net1110));
 sky130_fd_sc_hd__dlygate4sd3_1 hold605 (.A(\gpio_configure[32][10] ),
    .X(net1111));
 sky130_fd_sc_hd__dlygate4sd3_1 hold606 (.A(\gpio_configure[25][10] ),
    .X(net1112));
 sky130_fd_sc_hd__dlygate4sd3_1 hold607 (.A(\gpio_configure[1][12] ),
    .X(net1113));
 sky130_fd_sc_hd__dlygate4sd3_1 hold608 (.A(_1738_),
    .X(net1114));
 sky130_fd_sc_hd__dlygate4sd3_1 hold609 (.A(net1616),
    .X(net1115));
 sky130_fd_sc_hd__dlygate4sd3_1 hold610 (.A(\gpio_configure[17][10] ),
    .X(net1116));
 sky130_fd_sc_hd__dlygate4sd3_1 hold611 (.A(\mgmt_gpio_data_buf[14] ),
    .X(net1117));
 sky130_fd_sc_hd__dlygate4sd3_1 hold612 (.A(_1722_),
    .X(net1118));
 sky130_fd_sc_hd__dlygate4sd3_1 hold613 (.A(\mgmt_gpio_data_buf[13] ),
    .X(net1119));
 sky130_fd_sc_hd__dlygate4sd3_1 hold614 (.A(_1721_),
    .X(net1120));
 sky130_fd_sc_hd__dlygate4sd3_1 hold615 (.A(\gpio_configure[28][10] ),
    .X(net1121));
 sky130_fd_sc_hd__dlygate4sd3_1 hold616 (.A(net1605),
    .X(net1122));
 sky130_fd_sc_hd__dlygate4sd3_1 hold617 (.A(\gpio_configure[33][10] ),
    .X(net1123));
 sky130_fd_sc_hd__dlygate4sd3_1 hold618 (.A(_1685_),
    .X(net1124));
 sky130_fd_sc_hd__dlygate4sd3_1 hold619 (.A(\gpio_configure[23][10] ),
    .X(net1125));
 sky130_fd_sc_hd__dlygate4sd3_1 hold620 (.A(\gpio_configure[37][12] ),
    .X(net1126));
 sky130_fd_sc_hd__dlygate4sd3_1 hold621 (.A(\gpio_configure[26][2] ),
    .X(net1127));
 sky130_fd_sc_hd__dlygate4sd3_1 hold622 (.A(net1775),
    .X(net1128));
 sky130_fd_sc_hd__dlygate4sd3_1 hold623 (.A(_1665_),
    .X(net1129));
 sky130_fd_sc_hd__dlygate4sd3_1 hold624 (.A(\gpio_configure[5][7] ),
    .X(net1130));
 sky130_fd_sc_hd__dlygate4sd3_1 hold625 (.A(_3145_),
    .X(net1131));
 sky130_fd_sc_hd__dlygate4sd3_1 hold626 (.A(\gpio_configure[2][7] ),
    .X(net1132));
 sky130_fd_sc_hd__dlygate4sd3_1 hold627 (.A(_3113_),
    .X(net1133));
 sky130_fd_sc_hd__dlygate4sd3_1 hold628 (.A(_3055_),
    .X(net1134));
 sky130_fd_sc_hd__dlygate4sd3_1 hold629 (.A(_0434_),
    .X(net1135));
 sky130_fd_sc_hd__dlygate4sd3_1 hold630 (.A(net1653),
    .X(net1136));
 sky130_fd_sc_hd__dlygate4sd3_1 hold631 (.A(\gpio_configure[1][7] ),
    .X(net1137));
 sky130_fd_sc_hd__dlygate4sd3_1 hold632 (.A(_3104_),
    .X(net1138));
 sky130_fd_sc_hd__dlygate4sd3_1 hold633 (.A(\gpio_configure[37][2] ),
    .X(net1139));
 sky130_fd_sc_hd__dlygate4sd3_1 hold634 (.A(_3449_),
    .X(net1140));
 sky130_fd_sc_hd__dlygate4sd3_1 hold635 (.A(net1673),
    .X(net1141));
 sky130_fd_sc_hd__dlygate4sd3_1 hold636 (.A(\gpio_configure[18][7] ),
    .X(net1142));
 sky130_fd_sc_hd__dlygate4sd3_1 hold637 (.A(_3274_),
    .X(net1143));
 sky130_fd_sc_hd__dlygate4sd3_1 hold638 (.A(net1699),
    .X(net1144));
 sky130_fd_sc_hd__dlygate4sd3_1 hold639 (.A(\mgmt_gpio_data_buf[5] ),
    .X(net1145));
 sky130_fd_sc_hd__dlygate4sd3_1 hold640 (.A(_3083_),
    .X(net1146));
 sky130_fd_sc_hd__dlygate4sd3_1 hold641 (.A(net1721),
    .X(net1147));
 sky130_fd_sc_hd__dlygate4sd3_1 hold642 (.A(net1724),
    .X(net1148));
 sky130_fd_sc_hd__dlygate4sd3_1 hold643 (.A(\gpio_configure[29][7] ),
    .X(net1149));
 sky130_fd_sc_hd__dlygate4sd3_1 hold644 (.A(_3381_),
    .X(net1150));
 sky130_fd_sc_hd__dlygate4sd3_1 hold645 (.A(\gpio_configure[5][10] ),
    .X(net1151));
 sky130_fd_sc_hd__dlygate4sd3_1 hold646 (.A(\gpio_configure[22][7] ),
    .X(net1152));
 sky130_fd_sc_hd__dlygate4sd3_1 hold647 (.A(_3313_),
    .X(net1153));
 sky130_fd_sc_hd__dlygate4sd3_1 hold648 (.A(net1630),
    .X(net1154));
 sky130_fd_sc_hd__dlygate4sd3_1 hold649 (.A(\gpio_configure[35][7] ),
    .X(net1155));
 sky130_fd_sc_hd__dlygate4sd3_1 hold650 (.A(_3436_),
    .X(net1156));
 sky130_fd_sc_hd__dlygate4sd3_1 hold651 (.A(\gpio_configure[7][10] ),
    .X(net1157));
 sky130_fd_sc_hd__dlygate4sd3_1 hold652 (.A(_2039_),
    .X(net1158));
 sky130_fd_sc_hd__dlygate4sd3_1 hold653 (.A(\gpio_configure[33][7] ),
    .X(net1159));
 sky130_fd_sc_hd__dlygate4sd3_1 hold654 (.A(_3418_),
    .X(net1160));
 sky130_fd_sc_hd__dlygate4sd3_1 hold655 (.A(\gpio_configure[30][7] ),
    .X(net1161));
 sky130_fd_sc_hd__dlygate4sd3_1 hold656 (.A(_3390_),
    .X(net1162));
 sky130_fd_sc_hd__dlygate4sd3_1 hold657 (.A(net1654),
    .X(net1163));
 sky130_fd_sc_hd__dlygate4sd3_1 hold658 (.A(_1975_),
    .X(net1164));
 sky130_fd_sc_hd__dlygate4sd3_1 hold659 (.A(_0306_),
    .X(net1165));
 sky130_fd_sc_hd__dlygate4sd3_1 hold660 (.A(_1974_),
    .X(net1166));
 sky130_fd_sc_hd__dlygate4sd3_1 hold661 (.A(_0305_),
    .X(net1167));
 sky130_fd_sc_hd__dlygate4sd3_1 hold662 (.A(net1671),
    .X(net1168));
 sky130_fd_sc_hd__dlygate4sd3_1 hold663 (.A(\gpio_configure[31][10] ),
    .X(net1169));
 sky130_fd_sc_hd__dlygate4sd3_1 hold664 (.A(net1658),
    .X(net1170));
 sky130_fd_sc_hd__dlygate4sd3_1 hold665 (.A(\gpio_configure[25][7] ),
    .X(net1171));
 sky130_fd_sc_hd__dlygate4sd3_1 hold666 (.A(_3341_),
    .X(net1172));
 sky130_fd_sc_hd__dlygate4sd3_1 hold667 (.A(net1617),
    .X(net1173));
 sky130_fd_sc_hd__dlygate4sd3_1 hold668 (.A(\gpio_configure[10][7] ),
    .X(net1174));
 sky130_fd_sc_hd__dlygate4sd3_1 hold669 (.A(_3195_),
    .X(net1175));
 sky130_fd_sc_hd__dlygate4sd3_1 hold670 (.A(\gpio_configure[4][7] ),
    .X(net1176));
 sky130_fd_sc_hd__dlygate4sd3_1 hold671 (.A(_3135_),
    .X(net1177));
 sky130_fd_sc_hd__dlygate4sd3_1 hold672 (.A(\gpio_configure[34][11] ),
    .X(net1178));
 sky130_fd_sc_hd__dlygate4sd3_1 hold673 (.A(_1807_),
    .X(net1179));
 sky130_fd_sc_hd__dlygate4sd3_1 hold674 (.A(\gpio_configure[3][11] ),
    .X(net1180));
 sky130_fd_sc_hd__dlygate4sd3_1 hold675 (.A(_1999_),
    .X(net1181));
 sky130_fd_sc_hd__dlygate4sd3_1 hold676 (.A(\gpio_configure[1][6] ),
    .X(net1182));
 sky130_fd_sc_hd__dlygate4sd3_1 hold677 (.A(_3103_),
    .X(net1183));
 sky130_fd_sc_hd__dlygate4sd3_1 hold678 (.A(net1662),
    .X(net1184));
 sky130_fd_sc_hd__dlygate4sd3_1 hold679 (.A(\gpio_configure[2][5] ),
    .X(net1185));
 sky130_fd_sc_hd__dlygate4sd3_1 hold680 (.A(_3111_),
    .X(net1186));
 sky130_fd_sc_hd__dlygate4sd3_1 hold681 (.A(\mgmt_gpio_data_buf[6] ),
    .X(net1187));
 sky130_fd_sc_hd__dlygate4sd3_1 hold682 (.A(_3084_),
    .X(net1188));
 sky130_fd_sc_hd__dlygate4sd3_1 hold683 (.A(\gpio_configure[2][6] ),
    .X(net1189));
 sky130_fd_sc_hd__dlygate4sd3_1 hold684 (.A(_3112_),
    .X(net1190));
 sky130_fd_sc_hd__dlygate4sd3_1 hold685 (.A(\gpio_configure[34][7] ),
    .X(net1191));
 sky130_fd_sc_hd__dlygate4sd3_1 hold686 (.A(_3427_),
    .X(net1192));
 sky130_fd_sc_hd__dlygate4sd3_1 hold687 (.A(net1758),
    .X(net1193));
 sky130_fd_sc_hd__dlygate4sd3_1 hold688 (.A(_3120_),
    .X(net1194));
 sky130_fd_sc_hd__dlygate4sd3_1 hold689 (.A(serial_xfer),
    .X(net1195));
 sky130_fd_sc_hd__dlygate4sd3_1 hold690 (.A(_0436_),
    .X(net1196));
 sky130_fd_sc_hd__dlygate4sd3_1 hold691 (.A(\gpio_configure[9][7] ),
    .X(net1197));
 sky130_fd_sc_hd__dlygate4sd3_1 hold692 (.A(_3185_),
    .X(net1198));
 sky130_fd_sc_hd__dlygate4sd3_1 hold693 (.A(_3131_),
    .X(net1199));
 sky130_fd_sc_hd__dlygate4sd3_1 hold694 (.A(\gpio_configure[12][7] ),
    .X(net1200));
 sky130_fd_sc_hd__dlygate4sd3_1 hold695 (.A(_3213_),
    .X(net1201));
 sky130_fd_sc_hd__dlygate4sd3_1 hold696 (.A(_3009_),
    .X(net1202));
 sky130_fd_sc_hd__dlygate4sd3_1 hold697 (.A(net1788),
    .X(net1203));
 sky130_fd_sc_hd__dlygate4sd3_1 hold698 (.A(_3046_),
    .X(net1204));
 sky130_fd_sc_hd__dlygate4sd3_1 hold699 (.A(net1727),
    .X(net1205));
 sky130_fd_sc_hd__dlygate4sd3_1 hold700 (.A(\gpio_configure[1][3] ),
    .X(net1206));
 sky130_fd_sc_hd__dlygate4sd3_1 hold701 (.A(_3100_),
    .X(net1207));
 sky130_fd_sc_hd__dlygate4sd3_1 hold702 (.A(_3042_),
    .X(net1208));
 sky130_fd_sc_hd__dlygate4sd3_1 hold703 (.A(\gpio_configure[36][7] ),
    .X(net1209));
 sky130_fd_sc_hd__dlygate4sd3_1 hold704 (.A(_3445_),
    .X(net1210));
 sky130_fd_sc_hd__dlygate4sd3_1 hold705 (.A(net1725),
    .X(net1211));
 sky130_fd_sc_hd__dlygate4sd3_1 hold706 (.A(net1744),
    .X(net1212));
 sky130_fd_sc_hd__dlygate4sd3_1 hold707 (.A(\gpio_configure[2][9] ),
    .X(net1213));
 sky130_fd_sc_hd__dlygate4sd3_1 hold708 (.A(_1979_),
    .X(net1214));
 sky130_fd_sc_hd__dlygate4sd3_1 hold709 (.A(_3015_),
    .X(net1215));
 sky130_fd_sc_hd__dlygate4sd3_1 hold710 (.A(net1632),
    .X(net1216));
 sky130_fd_sc_hd__dlygate4sd3_1 hold711 (.A(net1681),
    .X(net1217));
 sky130_fd_sc_hd__dlygate4sd3_1 hold712 (.A(net1651),
    .X(net1218));
 sky130_fd_sc_hd__dlygate4sd3_1 hold713 (.A(net1791),
    .X(net1219));
 sky130_fd_sc_hd__dlygate4sd3_1 hold714 (.A(\gpio_configure[22][2] ),
    .X(net1220));
 sky130_fd_sc_hd__dlygate4sd3_1 hold715 (.A(net1627),
    .X(net1221));
 sky130_fd_sc_hd__dlygate4sd3_1 hold716 (.A(\gpio_configure[3][7] ),
    .X(net1222));
 sky130_fd_sc_hd__dlygate4sd3_1 hold717 (.A(_3126_),
    .X(net1223));
 sky130_fd_sc_hd__dlygate4sd3_1 hold718 (.A(net1691),
    .X(net1224));
 sky130_fd_sc_hd__dlygate4sd3_1 hold719 (.A(net1785),
    .X(net1225));
 sky130_fd_sc_hd__dlygate4sd3_1 hold720 (.A(\gpio_configure[8][2] ),
    .X(net1226));
 sky130_fd_sc_hd__dlygate4sd3_1 hold721 (.A(_3171_),
    .X(net1227));
 sky130_fd_sc_hd__dlygate4sd3_1 hold722 (.A(net1718),
    .X(net1228));
 sky130_fd_sc_hd__dlygate4sd3_1 hold723 (.A(\gpio_configure[21][2] ),
    .X(net1229));
 sky130_fd_sc_hd__dlygate4sd3_1 hold724 (.A(net1629),
    .X(net1230));
 sky130_fd_sc_hd__dlygate4sd3_1 hold725 (.A(net1639),
    .X(net1231));
 sky130_fd_sc_hd__dlygate4sd3_1 hold726 (.A(_3109_),
    .X(net1232));
 sky130_fd_sc_hd__dlygate4sd3_1 hold727 (.A(net1720),
    .X(net1233));
 sky130_fd_sc_hd__dlygate4sd3_1 hold728 (.A(net1618),
    .X(net1234));
 sky130_fd_sc_hd__dlygate4sd3_1 hold729 (.A(_1680_),
    .X(net1235));
 sky130_fd_sc_hd__dlygate4sd3_1 hold730 (.A(\gpio_configure[19][6] ),
    .X(net1236));
 sky130_fd_sc_hd__dlygate4sd3_1 hold731 (.A(_3284_),
    .X(net1237));
 sky130_fd_sc_hd__dlygate4sd3_1 hold732 (.A(net1661),
    .X(net1238));
 sky130_fd_sc_hd__dlygate4sd3_1 hold733 (.A(\gpio_configure[13][6] ),
    .X(net1239));
 sky130_fd_sc_hd__dlygate4sd3_1 hold734 (.A(_3221_),
    .X(net1240));
 sky130_fd_sc_hd__dlygate4sd3_1 hold735 (.A(\gpio_configure[25][6] ),
    .X(net1241));
 sky130_fd_sc_hd__dlygate4sd3_1 hold736 (.A(_3340_),
    .X(net1242));
 sky130_fd_sc_hd__dlygate4sd3_1 hold737 (.A(net1697),
    .X(net1243));
 sky130_fd_sc_hd__dlygate4sd3_1 hold738 (.A(\gpio_configure[37][7] ),
    .X(net1244));
 sky130_fd_sc_hd__dlygate4sd3_1 hold739 (.A(_3454_),
    .X(net1245));
 sky130_fd_sc_hd__dlygate4sd3_1 hold740 (.A(\gpio_configure[27][6] ),
    .X(net1246));
 sky130_fd_sc_hd__dlygate4sd3_1 hold741 (.A(_3362_),
    .X(net1247));
 sky130_fd_sc_hd__dlygate4sd3_1 hold742 (.A(net1678),
    .X(net1248));
 sky130_fd_sc_hd__dlygate4sd3_1 hold743 (.A(\gpio_configure[0][2] ),
    .X(net1249));
 sky130_fd_sc_hd__dlygate4sd3_1 hold744 (.A(_3090_),
    .X(net1250));
 sky130_fd_sc_hd__dlygate4sd3_1 hold745 (.A(_3014_),
    .X(net1251));
 sky130_fd_sc_hd__dlygate4sd3_1 hold746 (.A(\gpio_configure[20][6] ),
    .X(net1252));
 sky130_fd_sc_hd__dlygate4sd3_1 hold747 (.A(_3293_),
    .X(net1253));
 sky130_fd_sc_hd__dlygate4sd3_1 hold748 (.A(_3041_),
    .X(net1254));
 sky130_fd_sc_hd__dlygate4sd3_1 hold749 (.A(net1745),
    .X(net1255));
 sky130_fd_sc_hd__dlygate4sd3_1 hold750 (.A(\gpio_configure[11][6] ),
    .X(net1256));
 sky130_fd_sc_hd__dlygate4sd3_1 hold751 (.A(_3203_),
    .X(net1257));
 sky130_fd_sc_hd__dlygate4sd3_1 hold752 (.A(_3045_),
    .X(net1258));
 sky130_fd_sc_hd__dlygate4sd3_1 hold753 (.A(\gpio_configure[9][10] ),
    .X(net1259));
 sky130_fd_sc_hd__dlygate4sd3_1 hold754 (.A(\gpio_configure[17][6] ),
    .X(net1260));
 sky130_fd_sc_hd__dlygate4sd3_1 hold755 (.A(_3263_),
    .X(net1261));
 sky130_fd_sc_hd__dlygate4sd3_1 hold756 (.A(\gpio_configure[21][6] ),
    .X(net1262));
 sky130_fd_sc_hd__dlygate4sd3_1 hold757 (.A(_3303_),
    .X(net1263));
 sky130_fd_sc_hd__dlygate4sd3_1 hold758 (.A(net1755),
    .X(net1264));
 sky130_fd_sc_hd__dlygate4sd3_1 hold759 (.A(\gpio_configure[15][6] ),
    .X(net1265));
 sky130_fd_sc_hd__dlygate4sd3_1 hold760 (.A(_3243_),
    .X(net1266));
 sky130_fd_sc_hd__dlygate4sd3_1 hold761 (.A(_1691_),
    .X(net1267));
 sky130_fd_sc_hd__dlygate4sd3_1 hold762 (.A(\gpio_configure[7][6] ),
    .X(net1268));
 sky130_fd_sc_hd__dlygate4sd3_1 hold763 (.A(_3165_),
    .X(net1269));
 sky130_fd_sc_hd__dlygate4sd3_1 hold764 (.A(net1733),
    .X(net1270));
 sky130_fd_sc_hd__dlygate4sd3_1 hold765 (.A(\gpio_configure[5][6] ),
    .X(net1271));
 sky130_fd_sc_hd__dlygate4sd3_1 hold766 (.A(_3144_),
    .X(net1272));
 sky130_fd_sc_hd__dlygate4sd3_1 hold767 (.A(_3044_),
    .X(net1273));
 sky130_fd_sc_hd__dlygate4sd3_1 hold768 (.A(net1637),
    .X(net1274));
 sky130_fd_sc_hd__dlygate4sd3_1 hold769 (.A(\gpio_configure[6][2] ),
    .X(net1275));
 sky130_fd_sc_hd__dlygate4sd3_1 hold770 (.A(_3149_),
    .X(net1276));
 sky130_fd_sc_hd__dlygate4sd3_1 hold771 (.A(net1623),
    .X(net1277));
 sky130_fd_sc_hd__dlygate4sd3_1 hold772 (.A(\gpio_configure[18][6] ),
    .X(net1278));
 sky130_fd_sc_hd__dlygate4sd3_1 hold773 (.A(_3272_),
    .X(net1279));
 sky130_fd_sc_hd__dlygate4sd3_1 hold774 (.A(\wbbd_addr[5] ),
    .X(net1280));
 sky130_fd_sc_hd__dlygate4sd3_1 hold775 (.A(_0838_),
    .X(net1281));
 sky130_fd_sc_hd__dlygate4sd3_1 hold776 (.A(_3008_),
    .X(net1282));
 sky130_fd_sc_hd__dlygate4sd3_1 hold777 (.A(net1690),
    .X(net1283));
 sky130_fd_sc_hd__dlygate4sd3_1 hold778 (.A(net1664),
    .X(net1284));
 sky130_fd_sc_hd__dlygate4sd3_1 hold779 (.A(\gpio_configure[2][2] ),
    .X(net1285));
 sky130_fd_sc_hd__dlygate4sd3_1 hold780 (.A(_3108_),
    .X(net1286));
 sky130_fd_sc_hd__dlygate4sd3_1 hold781 (.A(net1610),
    .X(net1287));
 sky130_fd_sc_hd__dlygate4sd3_1 hold782 (.A(net1609),
    .X(net1288));
 sky130_fd_sc_hd__dlygate4sd3_1 hold783 (.A(_3013_),
    .X(net1289));
 sky130_fd_sc_hd__dlygate4sd3_1 hold784 (.A(\gpio_configure[15][10] ),
    .X(net1290));
 sky130_fd_sc_hd__dlygate4sd3_1 hold785 (.A(\gpio_configure[3][6] ),
    .X(net1291));
 sky130_fd_sc_hd__dlygate4sd3_1 hold786 (.A(_3125_),
    .X(net1292));
 sky130_fd_sc_hd__dlygate4sd3_1 hold787 (.A(net1634),
    .X(net1293));
 sky130_fd_sc_hd__dlygate4sd3_1 hold788 (.A(\gpio_configure[13][10] ),
    .X(net1294));
 sky130_fd_sc_hd__dlygate4sd3_1 hold789 (.A(_3162_),
    .X(net1295));
 sky130_fd_sc_hd__dlygate4sd3_1 hold790 (.A(\gpio_configure[31][7] ),
    .X(net1296));
 sky130_fd_sc_hd__dlygate4sd3_1 hold791 (.A(_3399_),
    .X(net1297));
 sky130_fd_sc_hd__dlygate4sd3_1 hold792 (.A(_3007_),
    .X(net1298));
 sky130_fd_sc_hd__dlygate4sd3_1 hold793 (.A(net1611),
    .X(net1299));
 sky130_fd_sc_hd__dlygate4sd3_1 hold794 (.A(\gpio_configure[4][6] ),
    .X(net1300));
 sky130_fd_sc_hd__dlygate4sd3_1 hold795 (.A(_3134_),
    .X(net1301));
 sky130_fd_sc_hd__dlygate4sd3_1 hold796 (.A(net1628),
    .X(net1302));
 sky130_fd_sc_hd__dlygate4sd3_1 hold797 (.A(_1693_),
    .X(net1303));
 sky130_fd_sc_hd__dlygate4sd3_1 hold798 (.A(\gpio_configure[6][6] ),
    .X(net1304));
 sky130_fd_sc_hd__dlygate4sd3_1 hold799 (.A(_3153_),
    .X(net1305));
 sky130_fd_sc_hd__dlygate4sd3_1 hold800 (.A(\gpio_configure[1][2] ),
    .X(net1306));
 sky130_fd_sc_hd__dlygate4sd3_1 hold801 (.A(_3099_),
    .X(net1307));
 sky130_fd_sc_hd__dlygate4sd3_1 hold802 (.A(net1752),
    .X(net1308));
 sky130_fd_sc_hd__dlygate4sd3_1 hold803 (.A(net1706),
    .X(net1309));
 sky130_fd_sc_hd__dlygate4sd3_1 hold804 (.A(net1707),
    .X(net1310));
 sky130_fd_sc_hd__dlygate4sd3_1 hold805 (.A(\gpio_configure[1][5] ),
    .X(net1311));
 sky130_fd_sc_hd__dlygate4sd3_1 hold806 (.A(_3102_),
    .X(net1312));
 sky130_fd_sc_hd__dlygate4sd3_1 hold807 (.A(_3040_),
    .X(net1313));
 sky130_fd_sc_hd__dlygate4sd3_1 hold808 (.A(_3029_),
    .X(net1314));
 sky130_fd_sc_hd__dlygate4sd3_1 hold809 (.A(\gpio_configure[24][10] ),
    .X(net1315));
 sky130_fd_sc_hd__dlygate4sd3_1 hold810 (.A(_3004_),
    .X(net1316));
 sky130_fd_sc_hd__dlygate4sd3_1 hold811 (.A(\gpio_configure[22][10] ),
    .X(net1317));
 sky130_fd_sc_hd__dlygate4sd3_1 hold812 (.A(\gpio_configure[2][10] ),
    .X(net1318));
 sky130_fd_sc_hd__dlygate4sd3_1 hold813 (.A(_1980_),
    .X(net1319));
 sky130_fd_sc_hd__dlygate4sd3_1 hold814 (.A(\mgmt_gpio_data_buf[0] ),
    .X(net1320));
 sky130_fd_sc_hd__dlygate4sd3_1 hold815 (.A(_3078_),
    .X(net1321));
 sky130_fd_sc_hd__dlygate4sd3_1 hold816 (.A(\mgmt_gpio_data_buf[21] ),
    .X(net1322));
 sky130_fd_sc_hd__dlygate4sd3_1 hold817 (.A(_1709_),
    .X(net1323));
 sky130_fd_sc_hd__dlygate4sd3_1 hold818 (.A(_3075_),
    .X(net1324));
 sky130_fd_sc_hd__dlygate4sd3_1 hold819 (.A(_0448_),
    .X(net1325));
 sky130_fd_sc_hd__dlygate4sd3_1 hold820 (.A(net1693),
    .X(net1326));
 sky130_fd_sc_hd__dlygate4sd3_1 hold821 (.A(\mgmt_gpio_data_buf[22] ),
    .X(net1327));
 sky130_fd_sc_hd__dlygate4sd3_1 hold822 (.A(_1711_),
    .X(net1328));
 sky130_fd_sc_hd__dlygate4sd3_1 hold823 (.A(\gpio_configure[0][12] ),
    .X(net1329));
 sky130_fd_sc_hd__dlygate4sd3_1 hold824 (.A(\gpio_configure[10][6] ),
    .X(net1330));
 sky130_fd_sc_hd__dlygate4sd3_1 hold825 (.A(_3194_),
    .X(net1331));
 sky130_fd_sc_hd__dlygate4sd3_1 hold826 (.A(\gpio_configure[33][0] ),
    .X(net1332));
 sky130_fd_sc_hd__dlygate4sd3_1 hold827 (.A(\gpio_configure[0][0] ),
    .X(net1333));
 sky130_fd_sc_hd__dlygate4sd3_1 hold828 (.A(\mgmt_gpio_data_buf[16] ),
    .X(net1334));
 sky130_fd_sc_hd__dlygate4sd3_1 hold829 (.A(_1703_),
    .X(net1335));
 sky130_fd_sc_hd__dlygate4sd3_1 hold830 (.A(\gpio_configure[18][8] ),
    .X(net1336));
 sky130_fd_sc_hd__dlygate4sd3_1 hold831 (.A(net1710),
    .X(net1337));
 sky130_fd_sc_hd__dlygate4sd3_1 hold832 (.A(\gpio_configure[9][6] ),
    .X(net1338));
 sky130_fd_sc_hd__dlygate4sd3_1 hold833 (.A(_3184_),
    .X(net1339));
 sky130_fd_sc_hd__dlygate4sd3_1 hold834 (.A(\gpio_configure[12][6] ),
    .X(net1340));
 sky130_fd_sc_hd__dlygate4sd3_1 hold835 (.A(_3212_),
    .X(net1341));
 sky130_fd_sc_hd__dlygate4sd3_1 hold836 (.A(\gpio_configure[14][6] ),
    .X(net1342));
 sky130_fd_sc_hd__dlygate4sd3_1 hold837 (.A(_3234_),
    .X(net1343));
 sky130_fd_sc_hd__dlygate4sd3_1 hold838 (.A(\mgmt_gpio_data_buf[8] ),
    .X(net1344));
 sky130_fd_sc_hd__dlygate4sd3_1 hold839 (.A(_1716_),
    .X(net1345));
 sky130_fd_sc_hd__dlygate4sd3_1 hold840 (.A(\gpio_configure[8][0] ),
    .X(net1346));
 sky130_fd_sc_hd__dlygate4sd3_1 hold841 (.A(net1717),
    .X(net1347));
 sky130_fd_sc_hd__dlygate4sd3_1 hold842 (.A(\gpio_configure[36][0] ),
    .X(net1348));
 sky130_fd_sc_hd__dlygate4sd3_1 hold843 (.A(\gpio_configure[6][8] ),
    .X(net1349));
 sky130_fd_sc_hd__dlygate4sd3_1 hold844 (.A(_2028_),
    .X(net1350));
 sky130_fd_sc_hd__dlygate4sd3_1 hold845 (.A(net1756),
    .X(net1351));
 sky130_fd_sc_hd__dlygate4sd3_1 hold846 (.A(net1738),
    .X(net1352));
 sky130_fd_sc_hd__dlygate4sd3_1 hold847 (.A(net1772),
    .X(net1353));
 sky130_fd_sc_hd__dlygate4sd3_1 hold848 (.A(net1754),
    .X(net1354));
 sky130_fd_sc_hd__dlygate4sd3_1 hold849 (.A(net1602),
    .X(net1355));
 sky130_fd_sc_hd__dlygate4sd3_1 hold850 (.A(net1657),
    .X(net1356));
 sky130_fd_sc_hd__dlygate4sd3_1 hold851 (.A(net1674),
    .X(net1357));
 sky130_fd_sc_hd__dlygate4sd3_1 hold852 (.A(\gpio_configure[16][0] ),
    .X(net1358));
 sky130_fd_sc_hd__dlygate4sd3_1 hold853 (.A(\gpio_configure[11][0] ),
    .X(net1359));
 sky130_fd_sc_hd__dlygate4sd3_1 hold854 (.A(_3003_),
    .X(net1360));
 sky130_fd_sc_hd__dlygate4sd3_1 hold855 (.A(\gpio_configure[3][8] ),
    .X(net1361));
 sky130_fd_sc_hd__dlygate4sd3_1 hold856 (.A(_1995_),
    .X(net1362));
 sky130_fd_sc_hd__dlygate4sd3_1 hold857 (.A(\wbbd_addr[4] ),
    .X(net1363));
 sky130_fd_sc_hd__dlygate4sd3_1 hold858 (.A(_3115_),
    .X(net1364));
 sky130_fd_sc_hd__dlygate4sd3_1 hold859 (.A(\gpio_configure[37][0] ),
    .X(net1365));
 sky130_fd_sc_hd__dlygate4sd3_1 hold860 (.A(_1683_),
    .X(net1366));
 sky130_fd_sc_hd__dlygate4sd3_1 hold861 (.A(_3020_),
    .X(net1367));
 sky130_fd_sc_hd__dlygate4sd3_1 hold862 (.A(net1686),
    .X(net1368));
 sky130_fd_sc_hd__dlygate4sd3_1 hold863 (.A(_3006_),
    .X(net1369));
 sky130_fd_sc_hd__dlygate4sd3_1 hold864 (.A(_3037_),
    .X(net1370));
 sky130_fd_sc_hd__dlygate4sd3_1 hold865 (.A(net1680),
    .X(net1371));
 sky130_fd_sc_hd__dlygate4sd3_1 hold866 (.A(net1713),
    .X(net1372));
 sky130_fd_sc_hd__dlygate4sd3_1 hold867 (.A(net1708),
    .X(net1373));
 sky130_fd_sc_hd__dlygate4sd3_1 hold868 (.A(net1650),
    .X(net1374));
 sky130_fd_sc_hd__dlygate4sd3_1 hold869 (.A(net1644),
    .X(net1375));
 sky130_fd_sc_hd__dlygate4sd3_1 hold870 (.A(net1748),
    .X(net1376));
 sky130_fd_sc_hd__dlygate4sd3_1 hold871 (.A(\gpio_configure[4][0] ),
    .X(net1377));
 sky130_fd_sc_hd__dlygate4sd3_1 hold872 (.A(net1779),
    .X(net1378));
 sky130_fd_sc_hd__dlygate4sd3_1 hold873 (.A(\gpio_configure[32][0] ),
    .X(net1379));
 sky130_fd_sc_hd__dlygate4sd3_1 hold874 (.A(_3402_),
    .X(net1380));
 sky130_fd_sc_hd__dlygate4sd3_1 hold875 (.A(net1747),
    .X(net1381));
 sky130_fd_sc_hd__dlygate4sd3_1 hold876 (.A(\gpio_configure[15][0] ),
    .X(net1382));
 sky130_fd_sc_hd__dlygate4sd3_1 hold877 (.A(net1715),
    .X(net1383));
 sky130_fd_sc_hd__dlygate4sd3_1 hold878 (.A(\gpio_configure[24][0] ),
    .X(net1384));
 sky130_fd_sc_hd__dlygate4sd3_1 hold879 (.A(_3325_),
    .X(net1385));
 sky130_fd_sc_hd__dlygate4sd3_1 hold880 (.A(\gpio_configure[28][8] ),
    .X(net1386));
 sky130_fd_sc_hd__dlygate4sd3_1 hold881 (.A(net1736),
    .X(net1387));
 sky130_fd_sc_hd__dlygate4sd3_1 hold882 (.A(net1740),
    .X(net1388));
 sky130_fd_sc_hd__dlygate4sd3_1 hold883 (.A(net1622),
    .X(net1389));
 sky130_fd_sc_hd__dlygate4sd3_1 hold884 (.A(net1761),
    .X(net1390));
 sky130_fd_sc_hd__dlygate4sd3_1 hold885 (.A(_3012_),
    .X(net1391));
 sky130_fd_sc_hd__dlygate4sd3_1 hold886 (.A(_1969_),
    .X(net1392));
 sky130_fd_sc_hd__dlygate4sd3_1 hold887 (.A(\gpio_configure[25][0] ),
    .X(net1393));
 sky130_fd_sc_hd__dlygate4sd3_1 hold888 (.A(\gpio_configure[30][0] ),
    .X(net1394));
 sky130_fd_sc_hd__dlygate4sd3_1 hold889 (.A(\gpio_configure[21][0] ),
    .X(net1395));
 sky130_fd_sc_hd__dlygate4sd3_1 hold890 (.A(net1626),
    .X(net1396));
 sky130_fd_sc_hd__dlygate4sd3_1 hold891 (.A(net1684),
    .X(net1397));
 sky130_fd_sc_hd__dlygate4sd3_1 hold892 (.A(net1723),
    .X(net1398));
 sky130_fd_sc_hd__dlygate4sd3_1 hold893 (.A(\gpio_configure[6][0] ),
    .X(net1399));
 sky130_fd_sc_hd__dlygate4sd3_1 hold894 (.A(net1769),
    .X(net1400));
 sky130_fd_sc_hd__dlygate4sd3_1 hold895 (.A(net1615),
    .X(net1401));
 sky130_fd_sc_hd__dlygate4sd3_1 hold896 (.A(_1952_),
    .X(net1402));
 sky130_fd_sc_hd__dlygate4sd3_1 hold897 (.A(_0292_),
    .X(net1403));
 sky130_fd_sc_hd__dlygate4sd3_1 hold898 (.A(net1732),
    .X(net1404));
 sky130_fd_sc_hd__dlygate4sd3_1 hold899 (.A(net1757),
    .X(net1405));
 sky130_fd_sc_hd__dlygate4sd3_1 hold900 (.A(\gpio_configure[31][0] ),
    .X(net1406));
 sky130_fd_sc_hd__dlygate4sd3_1 hold901 (.A(net1652),
    .X(net1407));
 sky130_fd_sc_hd__dlygate4sd3_1 hold902 (.A(\gpio_configure[29][0] ),
    .X(net1408));
 sky130_fd_sc_hd__dlygate4sd3_1 hold903 (.A(net1702),
    .X(net1409));
 sky130_fd_sc_hd__dlygate4sd3_1 hold904 (.A(\gpio_configure[22][0] ),
    .X(net1410));
 sky130_fd_sc_hd__dlygate4sd3_1 hold905 (.A(\gpio_configure[13][0] ),
    .X(net1411));
 sky130_fd_sc_hd__dlygate4sd3_1 hold906 (.A(net1783),
    .X(net1412));
 sky130_fd_sc_hd__dlygate4sd3_1 hold907 (.A(_3039_),
    .X(net1413));
 sky130_fd_sc_hd__dlygate4sd3_1 hold908 (.A(\gpio_configure[1][0] ),
    .X(net1414));
 sky130_fd_sc_hd__dlygate4sd3_1 hold909 (.A(_3048_),
    .X(net1415));
 sky130_fd_sc_hd__dlygate4sd3_1 hold910 (.A(_0428_),
    .X(net1416));
 sky130_fd_sc_hd__dlygate4sd3_1 hold911 (.A(\gpio_configure[2][0] ),
    .X(net1417));
 sky130_fd_sc_hd__dlygate4sd3_1 hold912 (.A(\gpio_configure[5][0] ),
    .X(net1418));
 sky130_fd_sc_hd__dlygate4sd3_1 hold913 (.A(net1606),
    .X(net1419));
 sky130_fd_sc_hd__dlygate4sd3_1 hold914 (.A(\gpio_configure[14][0] ),
    .X(net1420));
 sky130_fd_sc_hd__dlygate4sd3_1 hold915 (.A(net1765),
    .X(net1421));
 sky130_fd_sc_hd__dlygate4sd3_1 hold916 (.A(net1729),
    .X(net1422));
 sky130_fd_sc_hd__dlygate4sd3_1 hold917 (.A(net1742),
    .X(net1423));
 sky130_fd_sc_hd__dlygate4sd3_1 hold918 (.A(net1642),
    .X(net1424));
 sky130_fd_sc_hd__dlygate4sd3_1 hold919 (.A(\gpio_configure[28][0] ),
    .X(net1425));
 sky130_fd_sc_hd__dlygate4sd3_1 hold920 (.A(\gpio_configure[7][0] ),
    .X(net1426));
 sky130_fd_sc_hd__dlygate4sd3_1 hold921 (.A(\gpio_configure[35][0] ),
    .X(net1427));
 sky130_fd_sc_hd__dlygate4sd3_1 hold922 (.A(\gpio_configure[10][0] ),
    .X(net1428));
 sky130_fd_sc_hd__dlygate4sd3_1 hold923 (.A(net1730),
    .X(net1429));
 sky130_fd_sc_hd__dlygate4sd3_1 hold924 (.A(\gpio_configure[26][0] ),
    .X(net1430));
 sky130_fd_sc_hd__dlygate4sd3_1 hold925 (.A(\gpio_configure[19][0] ),
    .X(net1431));
 sky130_fd_sc_hd__dlygate4sd3_1 hold926 (.A(\gpio_configure[9][0] ),
    .X(net1432));
 sky130_fd_sc_hd__dlygate4sd3_1 hold927 (.A(\gpio_configure[17][0] ),
    .X(net1433));
 sky130_fd_sc_hd__dlygate4sd3_1 hold928 (.A(\gpio_configure[18][0] ),
    .X(net1434));
 sky130_fd_sc_hd__dlygate4sd3_1 hold929 (.A(\gpio_configure[20][0] ),
    .X(net1435));
 sky130_fd_sc_hd__dlygate4sd3_1 hold930 (.A(net1607),
    .X(net1436));
 sky130_fd_sc_hd__dlygate4sd3_1 hold931 (.A(\gpio_configure[23][0] ),
    .X(net1437));
 sky130_fd_sc_hd__dlygate4sd3_1 hold932 (.A(net1683),
    .X(net1438));
 sky130_fd_sc_hd__dlygate4sd3_1 hold933 (.A(_3069_),
    .X(net1439));
 sky130_fd_sc_hd__dlygate4sd3_1 hold934 (.A(_0443_),
    .X(net1440));
 sky130_fd_sc_hd__dlygate4sd3_1 hold935 (.A(\gpio_configure[27][0] ),
    .X(net1441));
 sky130_fd_sc_hd__dlygate4sd3_1 hold936 (.A(\gpio_configure[34][0] ),
    .X(net1442));
 sky130_fd_sc_hd__dlygate4sd3_1 hold937 (.A(_1661_),
    .X(net1443));
 sky130_fd_sc_hd__dlygate4sd3_1 hold938 (.A(\gpio_configure[12][0] ),
    .X(net1444));
 sky130_fd_sc_hd__dlygate4sd3_1 hold939 (.A(net1656),
    .X(net1445));
 sky130_fd_sc_hd__dlygate4sd3_1 hold940 (.A(net1712),
    .X(net1446));
 sky130_fd_sc_hd__dlygate4sd3_1 hold941 (.A(net1703),
    .X(net1447));
 sky130_fd_sc_hd__dlygate4sd3_1 hold942 (.A(\wbbd_state[1] ),
    .X(net1448));
 sky130_fd_sc_hd__dlygate4sd3_1 hold943 (.A(\hkspi.ldata[0] ),
    .X(net1449));
 sky130_fd_sc_hd__dlygate4sd3_1 hold944 (.A(\hkspi.addr[7] ),
    .X(net1450));
 sky130_fd_sc_hd__dlygate4sd3_1 hold945 (.A(_0777_),
    .X(net1451));
 sky130_fd_sc_hd__dlygate4sd3_1 hold946 (.A(\serial_data_staging_2[0] ),
    .X(net1452));
 sky130_fd_sc_hd__dlygate4sd3_1 hold947 (.A(\serial_data_staging_1[1] ),
    .X(net1453));
 sky130_fd_sc_hd__dlygate4sd3_1 hold948 (.A(_0780_),
    .X(net1454));
 sky130_fd_sc_hd__dlygate4sd3_1 hold949 (.A(\hkspi.state[1] ),
    .X(net1455));
 sky130_fd_sc_hd__dlygate4sd3_1 hold950 (.A(_0005_),
    .X(net1456));
 sky130_fd_sc_hd__dlygate4sd3_1 hold951 (.A(\hkspi.state[4] ),
    .X(net1457));
 sky130_fd_sc_hd__dlygate4sd3_1 hold952 (.A(_0086_),
    .X(net1458));
 sky130_fd_sc_hd__dlygate4sd3_1 hold953 (.A(\serial_data_staging_1[0] ),
    .X(net1459));
 sky130_fd_sc_hd__dlygate4sd3_1 hold954 (.A(\serial_data_staging_2[4] ),
    .X(net1460));
 sky130_fd_sc_hd__dlygate4sd3_1 hold955 (.A(_0796_),
    .X(net1461));
 sky130_fd_sc_hd__dlygate4sd3_1 hold956 (.A(\hkspi.ldata[3] ),
    .X(net1462));
 sky130_fd_sc_hd__dlygate4sd3_1 hold957 (.A(_1223_),
    .X(net1463));
 sky130_fd_sc_hd__dlygate4sd3_1 hold958 (.A(\wbbd_state[4] ),
    .X(net1464));
 sky130_fd_sc_hd__dlygate4sd3_1 hold959 (.A(\serial_data_staging_2[8] ),
    .X(net1465));
 sky130_fd_sc_hd__dlygate4sd3_1 hold960 (.A(_0800_),
    .X(net1466));
 sky130_fd_sc_hd__dlygate4sd3_1 hold961 (.A(\hkspi.ldata[2] ),
    .X(net1467));
 sky130_fd_sc_hd__dlygate4sd3_1 hold962 (.A(_1287_),
    .X(net1468));
 sky130_fd_sc_hd__dlygate4sd3_1 hold963 (.A(\hkspi.ldata[6] ),
    .X(net1469));
 sky130_fd_sc_hd__dlygate4sd3_1 hold964 (.A(_1024_),
    .X(net1470));
 sky130_fd_sc_hd__dlygate4sd3_1 hold965 (.A(\hkspi.fixed[1] ),
    .X(net1471));
 sky130_fd_sc_hd__dlygate4sd3_1 hold966 (.A(_0082_),
    .X(net1472));
 sky130_fd_sc_hd__dlygate4sd3_1 hold967 (.A(\wbbd_state[3] ),
    .X(net1473));
 sky130_fd_sc_hd__dlygate4sd3_1 hold968 (.A(\serial_data_staging_2[2] ),
    .X(net1474));
 sky130_fd_sc_hd__dlygate4sd3_1 hold969 (.A(_0794_),
    .X(net1475));
 sky130_fd_sc_hd__dlygate4sd3_1 hold970 (.A(\serial_data_staging_2[11] ),
    .X(net1476));
 sky130_fd_sc_hd__dlygate4sd3_1 hold971 (.A(_0803_),
    .X(net1477));
 sky130_fd_sc_hd__dlygate4sd3_1 hold972 (.A(\hkspi.ldata[5] ),
    .X(net1478));
 sky130_fd_sc_hd__dlygate4sd3_1 hold973 (.A(_1064_),
    .X(net1479));
 sky130_fd_sc_hd__dlygate4sd3_1 hold974 (.A(\serial_data_staging_1[3] ),
    .X(net1480));
 sky130_fd_sc_hd__dlygate4sd3_1 hold975 (.A(_0782_),
    .X(net1481));
 sky130_fd_sc_hd__dlygate4sd3_1 hold976 (.A(\serial_data_staging_1[6] ),
    .X(net1482));
 sky130_fd_sc_hd__dlygate4sd3_1 hold977 (.A(_0785_),
    .X(net1483));
 sky130_fd_sc_hd__dlygate4sd3_1 hold978 (.A(\serial_data_staging_1[9] ),
    .X(net1484));
 sky130_fd_sc_hd__dlygate4sd3_1 hold979 (.A(_0788_),
    .X(net1485));
 sky130_fd_sc_hd__dlygate4sd3_1 hold980 (.A(\hkspi.ldata[1] ),
    .X(net1486));
 sky130_fd_sc_hd__dlygate4sd3_1 hold981 (.A(\wbbd_state[2] ),
    .X(net1487));
 sky130_fd_sc_hd__dlygate4sd3_1 hold982 (.A(\serial_data_staging_1[7] ),
    .X(net1488));
 sky130_fd_sc_hd__dlygate4sd3_1 hold983 (.A(\serial_data_staging_2[5] ),
    .X(net1489));
 sky130_fd_sc_hd__dlygate4sd3_1 hold984 (.A(\hkspi.SDO ),
    .X(net1490));
 sky130_fd_sc_hd__dlygate4sd3_1 hold985 (.A(\serial_data_staging_1[11] ),
    .X(net1491));
 sky130_fd_sc_hd__dlygate4sd3_1 hold986 (.A(_0790_),
    .X(net1492));
 sky130_fd_sc_hd__dlygate4sd3_1 hold987 (.A(\serial_data_staging_1[10] ),
    .X(net1493));
 sky130_fd_sc_hd__dlygate4sd3_1 hold988 (.A(_0791_),
    .X(net1494));
 sky130_fd_sc_hd__dlygate4sd3_1 hold989 (.A(\serial_data_staging_1[4] ),
    .X(net1495));
 sky130_fd_sc_hd__dlygate4sd3_1 hold990 (.A(\serial_data_staging_2[7] ),
    .X(net1496));
 sky130_fd_sc_hd__dlygate4sd3_1 hold991 (.A(_0799_),
    .X(net1497));
 sky130_fd_sc_hd__dlygate4sd3_1 hold992 (.A(\wbbd_state[6] ),
    .X(net1498));
 sky130_fd_sc_hd__dlygate4sd3_1 hold993 (.A(\pad_count_2[2] ),
    .X(net1499));
 sky130_fd_sc_hd__dlygate4sd3_1 hold994 (.A(\hkspi.pre_pass_thru_user ),
    .X(net1500));
 sky130_fd_sc_hd__dlygate4sd3_1 hold995 (.A(_0007_),
    .X(net1501));
 sky130_fd_sc_hd__dlygate4sd3_1 hold996 (.A(\wbbd_state[0] ),
    .X(net1502));
 sky130_fd_sc_hd__dlygate4sd3_1 hold997 (.A(\serial_data_staging_1[5] ),
    .X(net1503));
 sky130_fd_sc_hd__dlygate4sd3_1 hold998 (.A(_0804_),
    .X(net1504));
 sky130_fd_sc_hd__dlygate4sd3_1 hold999 (.A(\hkspi.pre_pass_thru_mgmt ),
    .X(net1505));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1000 (.A(\hkspi.fixed[0] ),
    .X(net1506));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1001 (.A(\serial_data_staging_2[9] ),
    .X(net1507));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1002 (.A(\serial_data_staging_2[1] ),
    .X(net1508));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1003 (.A(\hkspi.count[2] ),
    .X(net1509));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1004 (.A(serial_clock_pre),
    .X(net1510));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1005 (.A(\serial_data_staging_1[8] ),
    .X(net1511));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1006 (.A(\serial_data_staging_2[3] ),
    .X(net1512));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1007 (.A(\serial_data_staging_1[2] ),
    .X(net1513));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1008 (.A(\hkspi.state[2] ),
    .X(net1514));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1009 (.A(_0004_),
    .X(net1515));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1010 (.A(\pad_count_1[1] ),
    .X(net1516));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1011 (.A(\xfer_count[3] ),
    .X(net1517));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1012 (.A(\hkspi.writemode ),
    .X(net1518));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1013 (.A(\pad_count_2[1] ),
    .X(net1519));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1014 (.A(\serial_data_staging_2[6] ),
    .X(net1520));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1015 (.A(\wbbd_state[8] ),
    .X(net1521));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1016 (.A(_4309_),
    .X(net1522));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1017 (.A(_4311_),
    .X(net1523));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1018 (.A(\pad_count_2[4] ),
    .X(net1524));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1019 (.A(\xfer_state[3] ),
    .X(net1525));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1020 (.A(\serial_data_staging_2[10] ),
    .X(net1526));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1021 (.A(\pad_count_2[5] ),
    .X(net1527));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1022 (.A(\hkspi.count[1] ),
    .X(net1528));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1023 (.A(\pad_count_2[3] ),
    .X(net1529));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1024 (.A(\hkspi.rdstb ),
    .X(net1530));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1025 (.A(\xfer_count[1] ),
    .X(net1531));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1026 (.A(\wbbd_state[6] ),
    .X(net1532));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1027 (.A(\wbbd_data[6] ),
    .X(net1533));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1028 (.A(\hkspi.odata[6] ),
    .X(net1534));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1029 (.A(\hkspi.odata[1] ),
    .X(net1535));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1030 (.A(\hkspi.odata[4] ),
    .X(net1536));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1031 (.A(\wbbd_state[5] ),
    .X(net1537));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1032 (.A(\wbbd_state[7] ),
    .X(net1538));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1033 (.A(_1945_),
    .X(net1539));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1034 (.A(_0290_),
    .X(net1540));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1035 (.A(\wbbd_data[7] ),
    .X(net1541));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1036 (.A(_1677_),
    .X(net1542));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1037 (.A(net1705),
    .X(net1543));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1038 (.A(net1621),
    .X(net1544));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1039 (.A(net1667),
    .X(net1545));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1040 (.A(net1655),
    .X(net1546));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1041 (.A(net1692),
    .X(net1547));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1042 (.A(_1956_),
    .X(net1548));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1043 (.A(\gpio_configure[22][1] ),
    .X(net1549));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1044 (.A(\gpio_configure[26][1] ),
    .X(net1550));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1045 (.A(\gpio_configure[23][1] ),
    .X(net1551));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1046 (.A(\gpio_configure[30][1] ),
    .X(net1552));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1047 (.A(\wbbd_data[5] ),
    .X(net1553));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1048 (.A(_1671_),
    .X(net1554));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1049 (.A(\wbbd_state[5] ),
    .X(net1555));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1050 (.A(\hkspi.odata[5] ),
    .X(net1556));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1051 (.A(\wbbd_addr[2] ),
    .X(net1557));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1052 (.A(\wbbd_data[2] ),
    .X(net1558));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1053 (.A(\wbbd_data[0] ),
    .X(net1559));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1054 (.A(\hkspi.odata[6] ),
    .X(net1560));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1055 (.A(\hkspi.addr[3] ),
    .X(net1561));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1056 (.A(\hkspi.addr[0] ),
    .X(net1562));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1057 (.A(\wbbd_data[3] ),
    .X(net1563));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1058 (.A(\wbbd_data[5] ),
    .X(net1564));
 sky130_fd_sc_hd__buf_6 rebuffer3 (.A(clknet_0_wb_clk_i),
    .X(net509));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1059 (.A(_1918_),
    .X(net1565));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1060 (.A(_0277_),
    .X(net1566));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1061 (.A(_1916_),
    .X(net1567));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1062 (.A(_0276_),
    .X(net1568));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1063 (.A(_1914_),
    .X(net1569));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1064 (.A(_0275_),
    .X(net1570));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1065 (.A(_1926_),
    .X(net1571));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1066 (.A(_0281_),
    .X(net1572));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1067 (.A(_1954_),
    .X(net1573));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1068 (.A(_0293_),
    .X(net1574));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1069 (.A(_1941_),
    .X(net1575));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1070 (.A(_0288_),
    .X(net1576));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1071 (.A(_1943_),
    .X(net1577));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1072 (.A(_0289_),
    .X(net1578));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1073 (.A(_3032_),
    .X(net1579));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1074 (.A(_0415_),
    .X(net1580));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1075 (.A(_1933_),
    .X(net1581));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1076 (.A(_0284_),
    .X(net1582));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1077 (.A(_1924_),
    .X(net1583));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1078 (.A(_0280_),
    .X(net1584));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1079 (.A(_1922_),
    .X(net1585));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1080 (.A(_0279_),
    .X(net1586));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1081 (.A(_1920_),
    .X(net1587));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1082 (.A(_0278_),
    .X(net1588));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1083 (.A(_1928_),
    .X(net1589));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1084 (.A(_0282_),
    .X(net1590));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1085 (.A(_3328_),
    .X(net1591));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1086 (.A(_3250_),
    .X(net1592));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1087 (.A(_3309_),
    .X(net1593));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1088 (.A(_3348_),
    .X(net1594));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1089 (.A(_3318_),
    .X(net1595));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1090 (.A(_3395_),
    .X(net1596));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1091 (.A(_3386_),
    .X(net1597));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1092 (.A(\gpio_configure[32][12] ),
    .X(net1598));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1093 (.A(\gpio_configure[13][4] ),
    .X(net1599));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1094 (.A(_3219_),
    .X(net1600));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1095 (.A(\gpio_configure[26][5] ),
    .X(net1601));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1096 (.A(\gpio_configure[34][8] ),
    .X(net1602));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1097 (.A(\gpio_configure[24][4] ),
    .X(net1603));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1098 (.A(_3329_),
    .X(net1604));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1099 (.A(\gpio_configure[31][12] ),
    .X(net1605));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1100 (.A(\gpio_configure[37][8] ),
    .X(net1606));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1101 (.A(\gpio_configure[33][8] ),
    .X(net1607));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1102 (.A(\gpio_configure[9][11] ),
    .X(net1608));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1103 (.A(\gpio_configure[11][2] ),
    .X(net1609));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1104 (.A(\gpio_configure[9][2] ),
    .X(net1610));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1105 (.A(_3063_),
    .X(net1611));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1106 (.A(\gpio_configure[16][4] ),
    .X(net1612));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1107 (.A(_3251_),
    .X(net1613));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1108 (.A(\gpio_configure[32][11] ),
    .X(net1614));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1109 (.A(\gpio_configure[25][8] ),
    .X(net1615));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1110 (.A(\gpio_configure[5][12] ),
    .X(net1616));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1111 (.A(\gpio_configure[15][11] ),
    .X(net1617));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1112 (.A(\gpio_configure[34][9] ),
    .X(net1618));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1113 (.A(\gpio_configure[9][12] ),
    .X(net1619));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1114 (.A(_2054_),
    .X(net1620));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1115 (.A(_1939_),
    .X(net1621));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1116 (.A(\gpio_configure[9][8] ),
    .X(net1622));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1117 (.A(\gpio_configure[12][2] ),
    .X(net1623));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1118 (.A(\gpio_configure[8][4] ),
    .X(net1624));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1119 (.A(_3173_),
    .X(net1625));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1120 (.A(\gpio_configure[2][8] ),
    .X(net1626));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1121 (.A(\gpio_configure[24][2] ),
    .X(net1627));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1122 (.A(\gpio_configure[21][9] ),
    .X(net1628));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1123 (.A(\gpio_configure[29][2] ),
    .X(net1629));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1124 (.A(\gpio_configure[25][12] ),
    .X(net1630));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1125 (.A(\gpio_configure[25][11] ),
    .X(net1631));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1126 (.A(\gpio_configure[22][11] ),
    .X(net1632));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1127 (.A(\gpio_configure[32][9] ),
    .X(net1633));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1128 (.A(\gpio_configure[13][2] ),
    .X(net1634));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1129 (.A(_1937_),
    .X(net1635));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1130 (.A(\gpio_configure[14][9] ),
    .X(net1636));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1131 (.A(\gpio_configure[24][9] ),
    .X(net1637));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1132 (.A(\gpio_configure[31][4] ),
    .X(net1638));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1133 (.A(\gpio_configure[35][2] ),
    .X(net1639));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1134 (.A(\gpio_configure[29][9] ),
    .X(net1640));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1135 (.A(\gpio_configure[24][7] ),
    .X(net1641));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1136 (.A(\gpio_configure[32][8] ),
    .X(net1642));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1137 (.A(\gpio_configure[16][7] ),
    .X(net1643));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1138 (.A(\gpio_configure[22][8] ),
    .X(net1644));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1139 (.A(_1670_),
    .X(net1645));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1140 (.A(\gpio_configure[30][2] ),
    .X(net1646));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1141 (.A(\gpio_configure[12][4] ),
    .X(net1647));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1142 (.A(_3210_),
    .X(net1648));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1143 (.A(\gpio_configure[29][4] ),
    .X(net1649));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1144 (.A(_3064_),
    .X(net1650));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1145 (.A(\gpio_configure[24][11] ),
    .X(net1651));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1146 (.A(\gpio_configure[5][8] ),
    .X(net1652));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1147 (.A(\gpio_configure[36][9] ),
    .X(net1653));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1148 (.A(\gpio_configure[26][7] ),
    .X(net1654));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1149 (.A(_1935_),
    .X(net1655));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1150 (.A(\gpio_configure[15][8] ),
    .X(net1656));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1151 (.A(\gpio_configure[22][9] ),
    .X(net1657));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1152 (.A(\gpio_configure[13][12] ),
    .X(net1658));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1153 (.A(\gpio_configure[5][11] ),
    .X(net1659));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1154 (.A(\gpio_configure[8][9] ),
    .X(net1660));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1155 (.A(\gpio_configure[26][6] ),
    .X(net1661));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1156 (.A(\gpio_configure[21][11] ),
    .X(net1662));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1157 (.A(\gpio_configure[27][9] ),
    .X(net1663));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1158 (.A(\gpio_configure[10][2] ),
    .X(net1664));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1159 (.A(\gpio_configure[22][12] ),
    .X(net1665));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1160 (.A(_1870_),
    .X(net1666));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1161 (.A(_1960_),
    .X(net1667));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1162 (.A(\hkspi.odata[4] ),
    .X(net1668));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1163 (.A(_3301_),
    .X(net1669));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1164 (.A(\gpio_configure[8][11] ),
    .X(net1670));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1165 (.A(\gpio_configure[33][12] ),
    .X(net1671));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1166 (.A(\gpio_configure[23][4] ),
    .X(net1672));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1167 (.A(\gpio_configure[23][12] ),
    .X(net1673));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1168 (.A(\gpio_configure[2][11] ),
    .X(net1674));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1169 (.A(\gpio_configure[35][11] ),
    .X(net1675));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1170 (.A(_3053_),
    .X(net1676));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1171 (.A(\gpio_configure[33][11] ),
    .X(net1677));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1172 (.A(\gpio_configure[33][9] ),
    .X(net1678));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1173 (.A(\gpio_configure[15][4] ),
    .X(net1679));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1174 (.A(\gpio_configure[3][2] ),
    .X(net1680));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1175 (.A(\gpio_configure[23][2] ),
    .X(net1681));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1176 (.A(\gpio_configure[12][9] ),
    .X(net1682));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1177 (.A(\gpio_configure[13][8] ),
    .X(net1683));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1178 (.A(\gpio_configure[4][8] ),
    .X(net1684));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1179 (.A(_3052_),
    .X(net1685));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1180 (.A(\gpio_configure[36][8] ),
    .X(net1686));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1181 (.A(\gpio_configure[0][4] ),
    .X(net1687));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1182 (.A(\gpio_configure[10][9] ),
    .X(net1688));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1183 (.A(\gpio_configure[31][11] ),
    .X(net1689));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1184 (.A(\gpio_configure[22][6] ),
    .X(net1690));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1185 (.A(\gpio_configure[20][2] ),
    .X(net1691));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1186 (.A(_1962_),
    .X(net1692));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1187 (.A(\gpio_configure[26][8] ),
    .X(net1693));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1188 (.A(_1604_),
    .X(net1694));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1189 (.A(_0429_),
    .X(net1695));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1190 (.A(\gpio_configure[27][4] ),
    .X(net1696));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1191 (.A(\gpio_configure[31][2] ),
    .X(net1697));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1192 (.A(\gpio_configure[35][9] ),
    .X(net1698));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1193 (.A(\gpio_configure[37][10] ),
    .X(net1699));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1194 (.A(\gpio_configure[8][12] ),
    .X(net1700));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1195 (.A(\gpio_configure[14][4] ),
    .X(net1701));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1196 (.A(\gpio_configure[31][8] ),
    .X(net1702));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1197 (.A(\gpio_configure[21][8] ),
    .X(net1703));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1198 (.A(\gpio_configure[21][12] ),
    .X(net1704));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1199 (.A(_1966_),
    .X(net1705));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1200 (.A(_3067_),
    .X(net1706));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1201 (.A(\gpio_configure[15][12] ),
    .X(net1707));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1202 (.A(_3066_),
    .X(net1708));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1203 (.A(\gpio_configure[37][4] ),
    .X(net1709));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1204 (.A(\gpio_configure[30][8] ),
    .X(net1710));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1205 (.A(\gpio_configure[26][4] ),
    .X(net1711));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1206 (.A(\gpio_configure[0][8] ),
    .X(net1712));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1207 (.A(\gpio_configure[9][9] ),
    .X(net1713));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1208 (.A(\gpio_configure[23][5] ),
    .X(net1714));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1209 (.A(_1931_),
    .X(net1715));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1210 (.A(\gpio_configure[31][6] ),
    .X(net1716));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1211 (.A(\gpio_configure[21][7] ),
    .X(net1717));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1212 (.A(\gpio_configure[17][2] ),
    .X(net1718));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1213 (.A(_1958_),
    .X(net1719));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1214 (.A(\gpio_configure[23][6] ),
    .X(net1720));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1215 (.A(\gpio_configure[24][12] ),
    .X(net1721));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1216 (.A(\gpio_configure[37][9] ),
    .X(net1722));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1217 (.A(\gpio_configure[23][8] ),
    .X(net1723));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1218 (.A(\gpio_configure[29][12] ),
    .X(net1724));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1219 (.A(_3062_),
    .X(net1725));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1220 (.A(\gpio_configure[17][11] ),
    .X(net1726));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1221 (.A(_3218_),
    .X(net1727));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1222 (.A(\gpio_configure[30][6] ),
    .X(net1728));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1223 (.A(hkspi_disable),
    .X(net1729));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1224 (.A(\gpio_configure[17][8] ),
    .X(net1730));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1225 (.A(\gpio_configure[35][4] ),
    .X(net1731));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1226 (.A(\gpio_configure[8][8] ),
    .X(net1732));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1227 (.A(\gpio_configure[5][2] ),
    .X(net1733));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1228 (.A(\gpio_configure[19][9] ),
    .X(net1734));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1229 (.A(\gpio_configure[24][6] ),
    .X(net1735));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1230 (.A(\gpio_configure[10][8] ),
    .X(net1736));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1231 (.A(\gpio_configure[10][11] ),
    .X(net1737));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1232 (.A(\gpio_configure[14][8] ),
    .X(net1738));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1233 (.A(\gpio_configure[36][10] ),
    .X(net1739));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1234 (.A(\gpio_configure[27][8] ),
    .X(net1740));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1235 (.A(\gpio_configure[17][9] ),
    .X(net1741));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1236 (.A(\gpio_configure[1][8] ),
    .X(net1742));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1237 (.A(\gpio_configure[23][9] ),
    .X(net1743));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1238 (.A(\gpio_configure[15][2] ),
    .X(net1744));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1239 (.A(\gpio_configure[15][9] ),
    .X(net1745));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1240 (.A(_3229_),
    .X(net1746));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1241 (.A(_3031_),
    .X(net1747));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1242 (.A(\gpio_configure[29][8] ),
    .X(net1748));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1243 (.A(\hkspi.addr[3] ),
    .X(net1749));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1244 (.A(_1608_),
    .X(net1750));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1245 (.A(\gpio_configure[30][9] ),
    .X(net1751));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1246 (.A(_3036_),
    .X(net1752));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1247 (.A(\gpio_configure[16][6] ),
    .X(net1753));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1248 (.A(\gpio_configure[14][7] ),
    .X(net1754));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1249 (.A(_3017_),
    .X(net1755));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1250 (.A(\gpio_configure[35][8] ),
    .X(net1756));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1251 (.A(\gpio_configure[12][8] ),
    .X(net1757));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1252 (.A(_3140_),
    .X(net1758));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1253 (.A(\gpio_configure[5][9] ),
    .X(net1759));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1254 (.A(_3450_),
    .X(net1760));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1255 (.A(\gpio_configure[7][8] ),
    .X(net1761));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1256 (.A(\gpio_configure[26][11] ),
    .X(net1762));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1257 (.A(\gpio_configure[11][9] ),
    .X(net1763));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1258 (.A(_3034_),
    .X(net1764));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1259 (.A(\gpio_configure[24][8] ),
    .X(net1765));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1260 (.A(\gpio_configure[10][12] ),
    .X(net1766));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1261 (.A(\gpio_configure[25][9] ),
    .X(net1767));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1262 (.A(\gpio_configure[31][9] ),
    .X(net1768));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1263 (.A(\gpio_configure[16][8] ),
    .X(net1769));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1264 (.A(\gpio_configure[11][11] ),
    .X(net1770));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1265 (.A(\gpio_configure[27][11] ),
    .X(net1771));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1266 (.A(\gpio_configure[19][8] ),
    .X(net1772));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1267 (.A(\gpio_configure[30][4] ),
    .X(net1773));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1268 (.A(\gpio_configure[19][11] ),
    .X(net1774));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1269 (.A(\gpio_configure[17][12] ),
    .X(net1775));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1270 (.A(\gpio_configure[12][11] ),
    .X(net1776));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1271 (.A(\gpio_configure[13][11] ),
    .X(net1777));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1272 (.A(_3056_),
    .X(net1778));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1273 (.A(\gpio_configure[20][8] ),
    .X(net1779));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1274 (.A(_3209_),
    .X(net1780));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1275 (.A(_3033_),
    .X(net1781));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1276 (.A(\gpio_configure[29][11] ),
    .X(net1782));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1277 (.A(\gpio_configure[11][8] ),
    .X(net1783));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1278 (.A(\gpio_configure[13][9] ),
    .X(net1784));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1279 (.A(\gpio_configure[18][2] ),
    .X(net1785));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1280 (.A(\gpio_configure[16][2] ),
    .X(net1786));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1281 (.A(\gpio_configure[20][9] ),
    .X(net1787));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1282 (.A(_3200_),
    .X(net1788));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1283 (.A(\gpio_configure[14][11] ),
    .X(net1789));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1284 (.A(_3091_),
    .X(net1790));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1285 (.A(\gpio_configure[19][2] ),
    .X(net1791));
 sky130_fd_sc_hd__diode_2 ANTENNA_1 (.DIODE(_0276_));
 sky130_fd_sc_hd__diode_2 ANTENNA_2 (.DIODE(_0284_));
 sky130_fd_sc_hd__diode_2 ANTENNA_3 (.DIODE(_0291_));
 sky130_fd_sc_hd__diode_2 ANTENNA_4 (.DIODE(_0291_));
 sky130_fd_sc_hd__diode_2 ANTENNA_5 (.DIODE(_0304_));
 sky130_fd_sc_hd__diode_2 ANTENNA_6 (.DIODE(_0348_));
 sky130_fd_sc_hd__diode_2 ANTENNA_7 (.DIODE(_0350_));
 sky130_fd_sc_hd__diode_2 ANTENNA_8 (.DIODE(_0402_));
 sky130_fd_sc_hd__diode_2 ANTENNA_9 (.DIODE(_0414_));
 sky130_fd_sc_hd__diode_2 ANTENNA_10 (.DIODE(_0415_));
 sky130_fd_sc_hd__diode_2 ANTENNA_11 (.DIODE(_0417_));
 sky130_fd_sc_hd__diode_2 ANTENNA_12 (.DIODE(_0612_));
 sky130_fd_sc_hd__diode_2 ANTENNA_13 (.DIODE(_0776_));
 sky130_fd_sc_hd__diode_2 ANTENNA_14 (.DIODE(_0890_));
 sky130_fd_sc_hd__diode_2 ANTENNA_15 (.DIODE(_0890_));
 sky130_fd_sc_hd__diode_2 ANTENNA_16 (.DIODE(_0890_));
 sky130_fd_sc_hd__diode_2 ANTENNA_17 (.DIODE(_0898_));
 sky130_fd_sc_hd__diode_2 ANTENNA_18 (.DIODE(_0898_));
 sky130_fd_sc_hd__diode_2 ANTENNA_19 (.DIODE(_0909_));
 sky130_fd_sc_hd__diode_2 ANTENNA_20 (.DIODE(_0916_));
 sky130_fd_sc_hd__diode_2 ANTENNA_21 (.DIODE(_0935_));
 sky130_fd_sc_hd__diode_2 ANTENNA_22 (.DIODE(_0935_));
 sky130_fd_sc_hd__diode_2 ANTENNA_23 (.DIODE(_0935_));
 sky130_fd_sc_hd__diode_2 ANTENNA_24 (.DIODE(_1005_));
 sky130_fd_sc_hd__diode_2 ANTENNA_25 (.DIODE(_1015_));
 sky130_fd_sc_hd__diode_2 ANTENNA_26 (.DIODE(_1039_));
 sky130_fd_sc_hd__diode_2 ANTENNA_27 (.DIODE(_1039_));
 sky130_fd_sc_hd__diode_2 ANTENNA_28 (.DIODE(_1041_));
 sky130_fd_sc_hd__diode_2 ANTENNA_29 (.DIODE(_1041_));
 sky130_fd_sc_hd__diode_2 ANTENNA_30 (.DIODE(_1048_));
 sky130_fd_sc_hd__diode_2 ANTENNA_31 (.DIODE(_1053_));
 sky130_fd_sc_hd__diode_2 ANTENNA_32 (.DIODE(_1065_));
 sky130_fd_sc_hd__diode_2 ANTENNA_33 (.DIODE(_1088_));
 sky130_fd_sc_hd__diode_2 ANTENNA_34 (.DIODE(_1112_));
 sky130_fd_sc_hd__diode_2 ANTENNA_35 (.DIODE(_1121_));
 sky130_fd_sc_hd__diode_2 ANTENNA_36 (.DIODE(_1121_));
 sky130_fd_sc_hd__diode_2 ANTENNA_37 (.DIODE(_1126_));
 sky130_fd_sc_hd__diode_2 ANTENNA_38 (.DIODE(_1146_));
 sky130_fd_sc_hd__diode_2 ANTENNA_39 (.DIODE(_1151_));
 sky130_fd_sc_hd__diode_2 ANTENNA_40 (.DIODE(_1154_));
 sky130_fd_sc_hd__diode_2 ANTENNA_41 (.DIODE(_1154_));
 sky130_fd_sc_hd__diode_2 ANTENNA_42 (.DIODE(_1170_));
 sky130_fd_sc_hd__diode_2 ANTENNA_43 (.DIODE(_1207_));
 sky130_fd_sc_hd__diode_2 ANTENNA_44 (.DIODE(_1226_));
 sky130_fd_sc_hd__diode_2 ANTENNA_45 (.DIODE(_1226_));
 sky130_fd_sc_hd__diode_2 ANTENNA_46 (.DIODE(_1233_));
 sky130_fd_sc_hd__diode_2 ANTENNA_47 (.DIODE(_1252_));
 sky130_fd_sc_hd__diode_2 ANTENNA_48 (.DIODE(_1275_));
 sky130_fd_sc_hd__diode_2 ANTENNA_49 (.DIODE(_1283_));
 sky130_fd_sc_hd__diode_2 ANTENNA_50 (.DIODE(_1315_));
 sky130_fd_sc_hd__diode_2 ANTENNA_51 (.DIODE(_1331_));
 sky130_fd_sc_hd__diode_2 ANTENNA_52 (.DIODE(_1344_));
 sky130_fd_sc_hd__diode_2 ANTENNA_53 (.DIODE(_1352_));
 sky130_fd_sc_hd__diode_2 ANTENNA_54 (.DIODE(_1352_));
 sky130_fd_sc_hd__diode_2 ANTENNA_55 (.DIODE(_1399_));
 sky130_fd_sc_hd__diode_2 ANTENNA_56 (.DIODE(_1399_));
 sky130_fd_sc_hd__diode_2 ANTENNA_57 (.DIODE(_1399_));
 sky130_fd_sc_hd__diode_2 ANTENNA_58 (.DIODE(_1399_));
 sky130_fd_sc_hd__diode_2 ANTENNA_59 (.DIODE(_1399_));
 sky130_fd_sc_hd__diode_2 ANTENNA_60 (.DIODE(_1413_));
 sky130_fd_sc_hd__diode_2 ANTENNA_61 (.DIODE(_1466_));
 sky130_fd_sc_hd__diode_2 ANTENNA_62 (.DIODE(_1466_));
 sky130_fd_sc_hd__diode_2 ANTENNA_63 (.DIODE(_1466_));
 sky130_fd_sc_hd__diode_2 ANTENNA_64 (.DIODE(_1466_));
 sky130_fd_sc_hd__diode_2 ANTENNA_65 (.DIODE(_1466_));
 sky130_fd_sc_hd__diode_2 ANTENNA_66 (.DIODE(_1487_));
 sky130_fd_sc_hd__diode_2 ANTENNA_67 (.DIODE(_1564_));
 sky130_fd_sc_hd__diode_2 ANTENNA_68 (.DIODE(_1565_));
 sky130_fd_sc_hd__diode_2 ANTENNA_69 (.DIODE(_1567_));
 sky130_fd_sc_hd__diode_2 ANTENNA_70 (.DIODE(_1578_));
 sky130_fd_sc_hd__diode_2 ANTENNA_71 (.DIODE(_1582_));
 sky130_fd_sc_hd__diode_2 ANTENNA_72 (.DIODE(_1600_));
 sky130_fd_sc_hd__diode_2 ANTENNA_73 (.DIODE(_1600_));
 sky130_fd_sc_hd__diode_2 ANTENNA_74 (.DIODE(_1600_));
 sky130_fd_sc_hd__diode_2 ANTENNA_75 (.DIODE(_1600_));
 sky130_fd_sc_hd__diode_2 ANTENNA_76 (.DIODE(_1601_));
 sky130_fd_sc_hd__diode_2 ANTENNA_77 (.DIODE(_1607_));
 sky130_fd_sc_hd__diode_2 ANTENNA_78 (.DIODE(_1615_));
 sky130_fd_sc_hd__diode_2 ANTENNA_79 (.DIODE(_1615_));
 sky130_fd_sc_hd__diode_2 ANTENNA_80 (.DIODE(_1615_));
 sky130_fd_sc_hd__diode_2 ANTENNA_81 (.DIODE(_1615_));
 sky130_fd_sc_hd__diode_2 ANTENNA_82 (.DIODE(_1658_));
 sky130_fd_sc_hd__diode_2 ANTENNA_83 (.DIODE(_1662_));
 sky130_fd_sc_hd__diode_2 ANTENNA_84 (.DIODE(_1664_));
 sky130_fd_sc_hd__diode_2 ANTENNA_85 (.DIODE(_1668_));
 sky130_fd_sc_hd__diode_2 ANTENNA_86 (.DIODE(_1708_));
 sky130_fd_sc_hd__diode_2 ANTENNA_87 (.DIODE(_1708_));
 sky130_fd_sc_hd__diode_2 ANTENNA_88 (.DIODE(_1708_));
 sky130_fd_sc_hd__diode_2 ANTENNA_89 (.DIODE(_1710_));
 sky130_fd_sc_hd__diode_2 ANTENNA_90 (.DIODE(_1710_));
 sky130_fd_sc_hd__diode_2 ANTENNA_91 (.DIODE(_1731_));
 sky130_fd_sc_hd__diode_2 ANTENNA_92 (.DIODE(_1731_));
 sky130_fd_sc_hd__diode_2 ANTENNA_93 (.DIODE(_1801_));
 sky130_fd_sc_hd__diode_2 ANTENNA_94 (.DIODE(_1801_));
 sky130_fd_sc_hd__diode_2 ANTENNA_95 (.DIODE(_1801_));
 sky130_fd_sc_hd__diode_2 ANTENNA_96 (.DIODE(_1801_));
 sky130_fd_sc_hd__diode_2 ANTENNA_97 (.DIODE(_1838_));
 sky130_fd_sc_hd__diode_2 ANTENNA_98 (.DIODE(_1905_));
 sky130_fd_sc_hd__diode_2 ANTENNA_99 (.DIODE(_1905_));
 sky130_fd_sc_hd__diode_2 ANTENNA_100 (.DIODE(_1905_));
 sky130_fd_sc_hd__diode_2 ANTENNA_101 (.DIODE(_1905_));
 sky130_fd_sc_hd__diode_2 ANTENNA_102 (.DIODE(_1913_));
 sky130_fd_sc_hd__diode_2 ANTENNA_103 (.DIODE(_1996_));
 sky130_fd_sc_hd__diode_2 ANTENNA_104 (.DIODE(_1996_));
 sky130_fd_sc_hd__diode_2 ANTENNA_105 (.DIODE(_2030_));
 sky130_fd_sc_hd__diode_2 ANTENNA_106 (.DIODE(_2030_));
 sky130_fd_sc_hd__diode_2 ANTENNA_107 (.DIODE(_2030_));
 sky130_fd_sc_hd__diode_2 ANTENNA_108 (.DIODE(_2030_));
 sky130_fd_sc_hd__diode_2 ANTENNA_109 (.DIODE(_2032_));
 sky130_fd_sc_hd__diode_2 ANTENNA_110 (.DIODE(_2032_));
 sky130_fd_sc_hd__diode_2 ANTENNA_111 (.DIODE(_2032_));
 sky130_fd_sc_hd__diode_2 ANTENNA_112 (.DIODE(_2032_));
 sky130_fd_sc_hd__diode_2 ANTENNA_113 (.DIODE(_2034_));
 sky130_fd_sc_hd__diode_2 ANTENNA_114 (.DIODE(_2034_));
 sky130_fd_sc_hd__diode_2 ANTENNA_115 (.DIODE(_2034_));
 sky130_fd_sc_hd__diode_2 ANTENNA_116 (.DIODE(_2034_));
 sky130_fd_sc_hd__diode_2 ANTENNA_117 (.DIODE(_2051_));
 sky130_fd_sc_hd__diode_2 ANTENNA_118 (.DIODE(_2100_));
 sky130_fd_sc_hd__diode_2 ANTENNA_119 (.DIODE(_2171_));
 sky130_fd_sc_hd__diode_2 ANTENNA_120 (.DIODE(_2174_));
 sky130_fd_sc_hd__diode_2 ANTENNA_121 (.DIODE(_2193_));
 sky130_fd_sc_hd__diode_2 ANTENNA_122 (.DIODE(_2653_));
 sky130_fd_sc_hd__diode_2 ANTENNA_123 (.DIODE(_3070_));
 sky130_fd_sc_hd__diode_2 ANTENNA_124 (.DIODE(_3117_));
 sky130_fd_sc_hd__diode_2 ANTENNA_125 (.DIODE(_3117_));
 sky130_fd_sc_hd__diode_2 ANTENNA_126 (.DIODE(_3136_));
 sky130_fd_sc_hd__diode_2 ANTENNA_127 (.DIODE(_3154_));
 sky130_fd_sc_hd__diode_2 ANTENNA_128 (.DIODE(_3154_));
 sky130_fd_sc_hd__diode_2 ANTENNA_129 (.DIODE(_3156_));
 sky130_fd_sc_hd__diode_2 ANTENNA_130 (.DIODE(_3275_));
 sky130_fd_sc_hd__diode_2 ANTENNA_131 (.DIODE(_3275_));
 sky130_fd_sc_hd__diode_2 ANTENNA_132 (.DIODE(_3345_));
 sky130_fd_sc_hd__diode_2 ANTENNA_133 (.DIODE(_3345_));
 sky130_fd_sc_hd__diode_2 ANTENNA_134 (.DIODE(_3401_));
 sky130_fd_sc_hd__diode_2 ANTENNA_135 (.DIODE(_3419_));
 sky130_fd_sc_hd__diode_2 ANTENNA_136 (.DIODE(_3437_));
 sky130_fd_sc_hd__diode_2 ANTENNA_137 (.DIODE(_3469_));
 sky130_fd_sc_hd__diode_2 ANTENNA_138 (.DIODE(_3484_));
 sky130_fd_sc_hd__diode_2 ANTENNA_139 (.DIODE(_3500_));
 sky130_fd_sc_hd__diode_2 ANTENNA_140 (.DIODE(_3500_));
 sky130_fd_sc_hd__diode_2 ANTENNA_141 (.DIODE(_3500_));
 sky130_fd_sc_hd__diode_2 ANTENNA_142 (.DIODE(_3500_));
 sky130_fd_sc_hd__diode_2 ANTENNA_143 (.DIODE(_3509_));
 sky130_fd_sc_hd__diode_2 ANTENNA_144 (.DIODE(_3511_));
 sky130_fd_sc_hd__diode_2 ANTENNA_145 (.DIODE(_3511_));
 sky130_fd_sc_hd__diode_2 ANTENNA_146 (.DIODE(_3511_));
 sky130_fd_sc_hd__diode_2 ANTENNA_147 (.DIODE(_3511_));
 sky130_fd_sc_hd__diode_2 ANTENNA_148 (.DIODE(_3511_));
 sky130_fd_sc_hd__diode_2 ANTENNA_149 (.DIODE(_3515_));
 sky130_fd_sc_hd__diode_2 ANTENNA_150 (.DIODE(_3515_));
 sky130_fd_sc_hd__diode_2 ANTENNA_151 (.DIODE(_3517_));
 sky130_fd_sc_hd__diode_2 ANTENNA_152 (.DIODE(_3526_));
 sky130_fd_sc_hd__diode_2 ANTENNA_153 (.DIODE(_3528_));
 sky130_fd_sc_hd__diode_2 ANTENNA_154 (.DIODE(_3528_));
 sky130_fd_sc_hd__diode_2 ANTENNA_155 (.DIODE(_3528_));
 sky130_fd_sc_hd__diode_2 ANTENNA_156 (.DIODE(_3535_));
 sky130_fd_sc_hd__diode_2 ANTENNA_157 (.DIODE(_3535_));
 sky130_fd_sc_hd__diode_2 ANTENNA_158 (.DIODE(_3535_));
 sky130_fd_sc_hd__diode_2 ANTENNA_159 (.DIODE(_3535_));
 sky130_fd_sc_hd__diode_2 ANTENNA_160 (.DIODE(_3536_));
 sky130_fd_sc_hd__diode_2 ANTENNA_161 (.DIODE(_3537_));
 sky130_fd_sc_hd__diode_2 ANTENNA_162 (.DIODE(_3537_));
 sky130_fd_sc_hd__diode_2 ANTENNA_163 (.DIODE(_3537_));
 sky130_fd_sc_hd__diode_2 ANTENNA_164 (.DIODE(_3537_));
 sky130_fd_sc_hd__diode_2 ANTENNA_165 (.DIODE(_3544_));
 sky130_fd_sc_hd__diode_2 ANTENNA_166 (.DIODE(_3544_));
 sky130_fd_sc_hd__diode_2 ANTENNA_167 (.DIODE(_3544_));
 sky130_fd_sc_hd__diode_2 ANTENNA_168 (.DIODE(_3544_));
 sky130_fd_sc_hd__diode_2 ANTENNA_169 (.DIODE(_3548_));
 sky130_fd_sc_hd__diode_2 ANTENNA_170 (.DIODE(_3548_));
 sky130_fd_sc_hd__diode_2 ANTENNA_171 (.DIODE(_3548_));
 sky130_fd_sc_hd__diode_2 ANTENNA_172 (.DIODE(_3550_));
 sky130_fd_sc_hd__diode_2 ANTENNA_173 (.DIODE(_3550_));
 sky130_fd_sc_hd__diode_2 ANTENNA_174 (.DIODE(_3555_));
 sky130_fd_sc_hd__diode_2 ANTENNA_175 (.DIODE(_3557_));
 sky130_fd_sc_hd__diode_2 ANTENNA_176 (.DIODE(_3557_));
 sky130_fd_sc_hd__diode_2 ANTENNA_177 (.DIODE(_3559_));
 sky130_fd_sc_hd__diode_2 ANTENNA_178 (.DIODE(_3561_));
 sky130_fd_sc_hd__diode_2 ANTENNA_179 (.DIODE(_3561_));
 sky130_fd_sc_hd__diode_2 ANTENNA_180 (.DIODE(_3561_));
 sky130_fd_sc_hd__diode_2 ANTENNA_181 (.DIODE(_3565_));
 sky130_fd_sc_hd__diode_2 ANTENNA_182 (.DIODE(_3567_));
 sky130_fd_sc_hd__diode_2 ANTENNA_183 (.DIODE(_3569_));
 sky130_fd_sc_hd__diode_2 ANTENNA_184 (.DIODE(_3578_));
 sky130_fd_sc_hd__diode_2 ANTENNA_185 (.DIODE(_3578_));
 sky130_fd_sc_hd__diode_2 ANTENNA_186 (.DIODE(_3581_));
 sky130_fd_sc_hd__diode_2 ANTENNA_187 (.DIODE(_3581_));
 sky130_fd_sc_hd__diode_2 ANTENNA_188 (.DIODE(_3585_));
 sky130_fd_sc_hd__diode_2 ANTENNA_189 (.DIODE(_3585_));
 sky130_fd_sc_hd__diode_2 ANTENNA_190 (.DIODE(_3585_));
 sky130_fd_sc_hd__diode_2 ANTENNA_191 (.DIODE(_3585_));
 sky130_fd_sc_hd__diode_2 ANTENNA_192 (.DIODE(_3585_));
 sky130_fd_sc_hd__diode_2 ANTENNA_193 (.DIODE(_3589_));
 sky130_fd_sc_hd__diode_2 ANTENNA_194 (.DIODE(_3589_));
 sky130_fd_sc_hd__diode_2 ANTENNA_195 (.DIODE(_3589_));
 sky130_fd_sc_hd__diode_2 ANTENNA_196 (.DIODE(_3589_));
 sky130_fd_sc_hd__diode_2 ANTENNA_197 (.DIODE(_3589_));
 sky130_fd_sc_hd__diode_2 ANTENNA_198 (.DIODE(_3589_));
 sky130_fd_sc_hd__diode_2 ANTENNA_199 (.DIODE(_3589_));
 sky130_fd_sc_hd__diode_2 ANTENNA_200 (.DIODE(_3621_));
 sky130_fd_sc_hd__diode_2 ANTENNA_201 (.DIODE(_3689_));
 sky130_fd_sc_hd__diode_2 ANTENNA_202 (.DIODE(_3879_));
 sky130_fd_sc_hd__diode_2 ANTENNA_203 (.DIODE(_3884_));
 sky130_fd_sc_hd__diode_2 ANTENNA_204 (.DIODE(_3884_));
 sky130_fd_sc_hd__diode_2 ANTENNA_205 (.DIODE(_3884_));
 sky130_fd_sc_hd__diode_2 ANTENNA_206 (.DIODE(_3885_));
 sky130_fd_sc_hd__diode_2 ANTENNA_207 (.DIODE(_3887_));
 sky130_fd_sc_hd__diode_2 ANTENNA_208 (.DIODE(_3900_));
 sky130_fd_sc_hd__diode_2 ANTENNA_209 (.DIODE(_3908_));
 sky130_fd_sc_hd__diode_2 ANTENNA_210 (.DIODE(_3920_));
 sky130_fd_sc_hd__diode_2 ANTENNA_211 (.DIODE(_3920_));
 sky130_fd_sc_hd__diode_2 ANTENNA_212 (.DIODE(_3920_));
 sky130_fd_sc_hd__diode_2 ANTENNA_213 (.DIODE(_3921_));
 sky130_fd_sc_hd__diode_2 ANTENNA_214 (.DIODE(_3941_));
 sky130_fd_sc_hd__diode_2 ANTENNA_215 (.DIODE(_3963_));
 sky130_fd_sc_hd__diode_2 ANTENNA_216 (.DIODE(_3964_));
 sky130_fd_sc_hd__diode_2 ANTENNA_217 (.DIODE(_3964_));
 sky130_fd_sc_hd__diode_2 ANTENNA_218 (.DIODE(_3965_));
 sky130_fd_sc_hd__diode_2 ANTENNA_219 (.DIODE(_3974_));
 sky130_fd_sc_hd__diode_2 ANTENNA_220 (.DIODE(clk1_output_dest));
 sky130_fd_sc_hd__diode_2 ANTENNA_221 (.DIODE(\gpio_configure[0][3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_222 (.DIODE(\gpio_configure[14][8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_223 (.DIODE(\gpio_configure[16][6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_224 (.DIODE(\gpio_configure[1][9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_225 (.DIODE(\gpio_configure[1][9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_226 (.DIODE(\gpio_configure[22][3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_227 (.DIODE(\gpio_configure[23][9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_228 (.DIODE(\gpio_configure[26][2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_229 (.DIODE(\gpio_configure[30][0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_230 (.DIODE(\gpio_configure[31][1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_231 (.DIODE(\gpio_configure[31][1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_232 (.DIODE(\gpio_configure[35][3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_233 (.DIODE(\gpio_configure[35][3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_234 (.DIODE(\gpio_configure[35][8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_235 (.DIODE(\gpio_configure[3][4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_236 (.DIODE(\gpio_configure[3][4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_237 (.DIODE(\gpio_configure[5][9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_238 (.DIODE(\gpio_configure[7][0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_239 (.DIODE(\hkspi.pass_thru_user_delay ));
 sky130_fd_sc_hd__diode_2 ANTENNA_240 (.DIODE(hkspi_disable));
 sky130_fd_sc_hd__diode_2 ANTENNA_241 (.DIODE(\mgmt_gpio_data[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_242 (.DIODE(user_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA_243 (.DIODE(user_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA_244 (.DIODE(wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_245 (.DIODE(wb_dat_i[21]));
 sky130_fd_sc_hd__diode_2 ANTENNA_246 (.DIODE(wb_dat_i[22]));
 sky130_fd_sc_hd__diode_2 ANTENNA_247 (.DIODE(wb_dat_i[23]));
 sky130_fd_sc_hd__diode_2 ANTENNA_248 (.DIODE(wb_dat_i[25]));
 sky130_fd_sc_hd__diode_2 ANTENNA_249 (.DIODE(wb_dat_i[27]));
 sky130_fd_sc_hd__diode_2 ANTENNA_250 (.DIODE(wb_sel_i[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA_251 (.DIODE(wb_sel_i[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA_252 (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA_253 (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA_254 (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA_255 (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA_256 (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA_257 (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA_258 (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA_259 (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA_260 (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA_261 (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA_262 (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA_263 (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA_264 (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA_265 (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA_266 (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA_267 (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA_268 (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA_269 (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA_270 (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA_271 (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA_272 (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA_273 (.DIODE(net58));
 sky130_fd_sc_hd__diode_2 ANTENNA_274 (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA_275 (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA_276 (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA_277 (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA_278 (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA_279 (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA_280 (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA_281 (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA_282 (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA_283 (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA_284 (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA_285 (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA_286 (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA_287 (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA_288 (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA_289 (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA_290 (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA_291 (.DIODE(net267));
 sky130_fd_sc_hd__diode_2 ANTENNA_292 (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA_293 (.DIODE(net272));
 sky130_fd_sc_hd__diode_2 ANTENNA_294 (.DIODE(net308));
 sky130_fd_sc_hd__diode_2 ANTENNA_295 (.DIODE(net359));
 sky130_fd_sc_hd__diode_2 ANTENNA_296 (.DIODE(net361));
 sky130_fd_sc_hd__diode_2 ANTENNA_297 (.DIODE(net372));
 sky130_fd_sc_hd__diode_2 ANTENNA_298 (.DIODE(net372));
 sky130_fd_sc_hd__diode_2 ANTENNA_299 (.DIODE(net372));
 sky130_fd_sc_hd__diode_2 ANTENNA_300 (.DIODE(net372));
 sky130_fd_sc_hd__diode_2 ANTENNA_301 (.DIODE(net374));
 sky130_fd_sc_hd__diode_2 ANTENNA_302 (.DIODE(net374));
 sky130_fd_sc_hd__diode_2 ANTENNA_303 (.DIODE(net374));
 sky130_fd_sc_hd__diode_2 ANTENNA_304 (.DIODE(net377));
 sky130_fd_sc_hd__diode_2 ANTENNA_305 (.DIODE(net385));
 sky130_fd_sc_hd__diode_2 ANTENNA_306 (.DIODE(net387));
 sky130_fd_sc_hd__diode_2 ANTENNA_307 (.DIODE(net388));
 sky130_fd_sc_hd__diode_2 ANTENNA_308 (.DIODE(net390));
 sky130_fd_sc_hd__diode_2 ANTENNA_309 (.DIODE(net498));
 sky130_fd_sc_hd__diode_2 ANTENNA_310 (.DIODE(net504));
 sky130_fd_sc_hd__diode_2 ANTENNA_311 (.DIODE(net504));
 sky130_fd_sc_hd__diode_2 ANTENNA_312 (.DIODE(clknet_3_2_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_313 (.DIODE(net511));
 sky130_fd_sc_hd__diode_2 ANTENNA_314 (.DIODE(net521));
 sky130_fd_sc_hd__diode_2 ANTENNA_315 (.DIODE(net552));
 sky130_fd_sc_hd__diode_2 ANTENNA_316 (.DIODE(net939));
 sky130_fd_sc_hd__diode_2 ANTENNA_317 (.DIODE(net1581));
 sky130_fd_sc_hd__diode_2 ANTENNA_318 (.DIODE(net1586));
 sky130_fd_sc_hd__diode_2 ANTENNA_319 (.DIODE(_0099_));
 sky130_fd_sc_hd__diode_2 ANTENNA_320 (.DIODE(_0430_));
 sky130_fd_sc_hd__diode_2 ANTENNA_321 (.DIODE(_0435_));
 sky130_fd_sc_hd__diode_2 ANTENNA_322 (.DIODE(_0628_));
 sky130_fd_sc_hd__diode_2 ANTENNA_323 (.DIODE(_0644_));
 sky130_fd_sc_hd__diode_2 ANTENNA_324 (.DIODE(_0700_));
 sky130_fd_sc_hd__diode_2 ANTENNA_325 (.DIODE(_1005_));
 sky130_fd_sc_hd__diode_2 ANTENNA_326 (.DIODE(_1022_));
 sky130_fd_sc_hd__diode_2 ANTENNA_327 (.DIODE(_1347_));
 sky130_fd_sc_hd__diode_2 ANTENNA_328 (.DIODE(_1466_));
 sky130_fd_sc_hd__diode_2 ANTENNA_329 (.DIODE(_1466_));
 sky130_fd_sc_hd__diode_2 ANTENNA_330 (.DIODE(_1557_));
 sky130_fd_sc_hd__diode_2 ANTENNA_331 (.DIODE(_1575_));
 sky130_fd_sc_hd__diode_2 ANTENNA_332 (.DIODE(_1598_));
 sky130_fd_sc_hd__diode_2 ANTENNA_333 (.DIODE(_1598_));
 sky130_fd_sc_hd__diode_2 ANTENNA_334 (.DIODE(_1607_));
 sky130_fd_sc_hd__diode_2 ANTENNA_335 (.DIODE(_1618_));
 sky130_fd_sc_hd__diode_2 ANTENNA_336 (.DIODE(_1658_));
 sky130_fd_sc_hd__diode_2 ANTENNA_337 (.DIODE(_1658_));
 sky130_fd_sc_hd__diode_2 ANTENNA_338 (.DIODE(_1672_));
 sky130_fd_sc_hd__diode_2 ANTENNA_339 (.DIODE(_1710_));
 sky130_fd_sc_hd__diode_2 ANTENNA_340 (.DIODE(_1712_));
 sky130_fd_sc_hd__diode_2 ANTENNA_341 (.DIODE(_1731_));
 sky130_fd_sc_hd__diode_2 ANTENNA_342 (.DIODE(_1993_));
 sky130_fd_sc_hd__diode_2 ANTENNA_343 (.DIODE(_2011_));
 sky130_fd_sc_hd__diode_2 ANTENNA_344 (.DIODE(_2032_));
 sky130_fd_sc_hd__diode_2 ANTENNA_345 (.DIODE(_2032_));
 sky130_fd_sc_hd__diode_2 ANTENNA_346 (.DIODE(_3070_));
 sky130_fd_sc_hd__diode_2 ANTENNA_347 (.DIODE(_3070_));
 sky130_fd_sc_hd__diode_2 ANTENNA_348 (.DIODE(_3117_));
 sky130_fd_sc_hd__diode_2 ANTENNA_349 (.DIODE(_3117_));
 sky130_fd_sc_hd__diode_2 ANTENNA_350 (.DIODE(_3127_));
 sky130_fd_sc_hd__diode_2 ANTENNA_351 (.DIODE(_3156_));
 sky130_fd_sc_hd__diode_2 ANTENNA_352 (.DIODE(_3156_));
 sky130_fd_sc_hd__diode_2 ANTENNA_353 (.DIODE(_3158_));
 sky130_fd_sc_hd__diode_2 ANTENNA_354 (.DIODE(_3246_));
 sky130_fd_sc_hd__diode_2 ANTENNA_355 (.DIODE(_3410_));
 sky130_fd_sc_hd__diode_2 ANTENNA_356 (.DIODE(_3521_));
 sky130_fd_sc_hd__diode_2 ANTENNA_357 (.DIODE(_3538_));
 sky130_fd_sc_hd__diode_2 ANTENNA_358 (.DIODE(_3540_));
 sky130_fd_sc_hd__diode_2 ANTENNA_359 (.DIODE(_3544_));
 sky130_fd_sc_hd__diode_2 ANTENNA_360 (.DIODE(_3557_));
 sky130_fd_sc_hd__diode_2 ANTENNA_361 (.DIODE(_3587_));
 sky130_fd_sc_hd__diode_2 ANTENNA_362 (.DIODE(_3591_));
 sky130_fd_sc_hd__diode_2 ANTENNA_363 (.DIODE(_3921_));
 sky130_fd_sc_hd__diode_2 ANTENNA_364 (.DIODE(_3954_));
 sky130_fd_sc_hd__diode_2 ANTENNA_365 (.DIODE(_3959_));
 sky130_fd_sc_hd__diode_2 ANTENNA_366 (.DIODE(\gpio_configure[19][4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_367 (.DIODE(\gpio_configure[29][12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_368 (.DIODE(\gpio_configure[5][10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_369 (.DIODE(\gpio_configure[7][5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_370 (.DIODE(\hkspi.pass_thru_user ));
 sky130_fd_sc_hd__diode_2 ANTENNA_371 (.DIODE(irq_1_inputsrc));
 sky130_fd_sc_hd__diode_2 ANTENNA_372 (.DIODE(wb_dat_i[24]));
 sky130_fd_sc_hd__diode_2 ANTENNA_373 (.DIODE(wb_dat_i[26]));
 sky130_fd_sc_hd__diode_2 ANTENNA_374 (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA_375 (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA_376 (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA_377 (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA_378 (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA_379 (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA_380 (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA_381 (.DIODE(net307));
 sky130_fd_sc_hd__diode_2 ANTENNA_382 (.DIODE(net316));
 sky130_fd_sc_hd__diode_2 ANTENNA_383 (.DIODE(net390));
 sky130_fd_sc_hd__diode_2 ANTENNA_384 (.DIODE(net457));
 sky130_fd_sc_hd__diode_2 ANTENNA_385 (.DIODE(net457));
 sky130_fd_sc_hd__diode_2 ANTENNA_386 (.DIODE(net457));
 sky130_fd_sc_hd__diode_2 ANTENNA_387 (.DIODE(net533));
 sky130_fd_sc_hd__diode_2 ANTENNA_388 (.DIODE(net552));
 sky130_fd_sc_hd__diode_2 ANTENNA_389 (.DIODE(net1590));
 sky130_fd_sc_hd__diode_2 ANTENNA_390 (.DIODE(_0763_));
 sky130_fd_sc_hd__diode_2 ANTENNA_391 (.DIODE(_0973_));
 sky130_fd_sc_hd__diode_2 ANTENNA_392 (.DIODE(_1710_));
 sky130_fd_sc_hd__diode_2 ANTENNA_393 (.DIODE(_1712_));
 sky130_fd_sc_hd__diode_2 ANTENNA_394 (.DIODE(_1996_));
 sky130_fd_sc_hd__diode_2 ANTENNA_395 (.DIODE(_1996_));
 sky130_fd_sc_hd__diode_2 ANTENNA_396 (.DIODE(_1996_));
 sky130_fd_sc_hd__diode_2 ANTENNA_397 (.DIODE(_2032_));
 sky130_fd_sc_hd__diode_2 ANTENNA_398 (.DIODE(_2034_));
 sky130_fd_sc_hd__diode_2 ANTENNA_399 (.DIODE(_3068_));
 sky130_fd_sc_hd__diode_2 ANTENNA_400 (.DIODE(_3156_));
 sky130_fd_sc_hd__diode_2 ANTENNA_401 (.DIODE(_3475_));
 sky130_fd_sc_hd__diode_2 ANTENNA_402 (.DIODE(_3538_));
 sky130_fd_sc_hd__diode_2 ANTENNA_403 (.DIODE(\hkspi.pass_thru_user ));
 sky130_fd_sc_hd__diode_2 ANTENNA_404 (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA_405 (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA_406 (.DIODE(net533));
 sky130_fd_sc_hd__decap_6 FILLER_0_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_511 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_547 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_566 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_573 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_622 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_683 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_775 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_12 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_16 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_20 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_34 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_90 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_242 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_267 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_423 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_491 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_500 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_534 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_566 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_578 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_591 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_622 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_626 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_650 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_683 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_711 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_715 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_759 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_34 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_99 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_332 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_396 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_448 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_500 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_557 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_587 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_604 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_616 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_623 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_655 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_663 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_738 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_775 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_12 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_20 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_25 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_34 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_90 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_179 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_254 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_480 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_500 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_580 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_644 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_682 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_686 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_739 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_747 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_754 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_758 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_44 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_52 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_67 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_78 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_164 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_339 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_384 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_452 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_482 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_522 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_552 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_564 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_572 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_622 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_634 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_651 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_680 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_686 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_724 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_736 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_32 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_86 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_123 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_240 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_415 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_432 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_543 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_574 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_581 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_594 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_628 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_636 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_659 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_691 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_702 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_706 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_715 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_763 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_775 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_49 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_58 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_151 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_227 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_298 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_320 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_340 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_451 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_466 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_491 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_508 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_522 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_543 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_584 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_619 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_632 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_662 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_691 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_25 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_36 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_136 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_189 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_196 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_420 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_432 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_515 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_540 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_558 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_642 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_651 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_664 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_678 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_703 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_739 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_747 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_768 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_775 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_14 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_52 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_102 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_290 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_319 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_384 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_418 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_452 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_492 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_514 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_547 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_551 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_558 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_562 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_599 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_611 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_619 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_642 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_698 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_715 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_728 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_767 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_75 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_198 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_354 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_366 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_422 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_454 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_460 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_482 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_515 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_528 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_534 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_586 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_639 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_651 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_659 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_684 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_726 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_775 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_10 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_17 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_62 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_66 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_104 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_114 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_226 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_276 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_338 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_386 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_443 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_519 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_547 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_555 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_611 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_642 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_656 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_676 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_711 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_747 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_25 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_31 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_40 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_70 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_87 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_127 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_232 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_436 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_484 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_525 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_576 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_621 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_631 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_647 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_659 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_680 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_750 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_772 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_34 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_102 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_114 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_163 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_170 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_217 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_238 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_272 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_284 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_395 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_410 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_448 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_463 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_473 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_483 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_530 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_560 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_594 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_670 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_674 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_711 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_735 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_767 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_775 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_14 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_74 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_86 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_176 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_311 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_415 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_492 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_525 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_584 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_615 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_623 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_662 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_669 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_690 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_703 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_715 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_748 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_46 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_89 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_170 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_224 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_282 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_360 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_384 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_435 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_484 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_522 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_530 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_611 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_623 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_653 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_711 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_724 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_730 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_766 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_775 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_31 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_42 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_64 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_143 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_198 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_296 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_386 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_420 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_478 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_491 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_527 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_543 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_574 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_639 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_651 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_690 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_751 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_763 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_60 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_96 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_104 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_215 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_272 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_284 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_292 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_327 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_340 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_397 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_442 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_460 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_499 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_506 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_518 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_553 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_584 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_618 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_630 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_640 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_654 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_666 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_687 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_711 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_735 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_743 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_767 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_32 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_70 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_88 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_135 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_235 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_267 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_296 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_359 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_479 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_535 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_570 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_594 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_606 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_622 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_626 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_650 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_662 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_704 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_104 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_179 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_282 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_331 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_360 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_371 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_500 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_551 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_570 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_596 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_609 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_663 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_767 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_68 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_135 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_142 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_242 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_246 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_355 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_368 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_503 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_528 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_532 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_554 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_592 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_604 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_625 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_650 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_658 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_684 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_711 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_740 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_752 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_758 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_13 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_96 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_168 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_212 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_436 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_556 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_564 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_594 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_598 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_620 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_626 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_653 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_687 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_711 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_731 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_763 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_775 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_179 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_398 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_459 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_491 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_510 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_518 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_547 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_639 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_652 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_660 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_695 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_707 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_713 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_764 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_17 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_56 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_98 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_224 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_228 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_232 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_395 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_458 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_515 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_530 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_603 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_615 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_655 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_667 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_675 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_724 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_734 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_19 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_86 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_117 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_144 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_160 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_200 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_255 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_411 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_423 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_442 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_502 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_534 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_570 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_580 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_590 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_627 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_683 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_714 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_751 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_761 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_771 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_17 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_44 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_186 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_228 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_275 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_282 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_341 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_392 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_437 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_487 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_507 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_516 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_555 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_566 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_612 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_624 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_670 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_711 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_731 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_738 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_767 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_775 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_16 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_28 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_39 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_50 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_149 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_199 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_355 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_408 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_420 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_510 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_536 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_582 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_592 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_604 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_608 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_641 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_696 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_708 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_714 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_734 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_762 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_766 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_48 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_56 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_155 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_202 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_263 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_329 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_445 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_504 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_555 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_602 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_612 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_643 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_674 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_727 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_733 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_767 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_774 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_30 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_77 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_260 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_367 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_380 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_465 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_492 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_542 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_571 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_581 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_622 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_646 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_670 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_700 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_747 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_772 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_61 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_104 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_152 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_170 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_179 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_188 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_212 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_224 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_230 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_259 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_275 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_340 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_379 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_442 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_454 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_475 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_528 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_543 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_556 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_562 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_570 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_586 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_598 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_650 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_670 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_682 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_698 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_705 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_775 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_18 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_22 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_31 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_180 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_208 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_256 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_295 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_302 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_415 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_460 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_478 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_528 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_558 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_574 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_640 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_671 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_17 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_40 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_58 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_115 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_130 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_272 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_326 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_343 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_358 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_382 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_554 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_586 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_610 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_642 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_651 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_678 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_682 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_724 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_728 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_738 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_762 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_766 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_775 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_16 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_63 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_80 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_123 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_130 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_147 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_179 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_191 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_263 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_467 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_478 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_516 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_528 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_534 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_579 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_602 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_639 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_651 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_659 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_679 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_754 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_758 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_775 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_10 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_26 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_56 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_73 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_78 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_151 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_171 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_206 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_218 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_226 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_286 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_340 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_356 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_379 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_513 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_547 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_586 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_606 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_640 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_698 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_715 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_743 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_763 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_775 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_10 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_31 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_79 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_196 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_235 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_247 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_303 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_366 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_436 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_519 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_591 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_596 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_600 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_610 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_624 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_632 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_641 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_671 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_775 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_13 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_47 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_60 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_74 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_105 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_180 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_282 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_394 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_491 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_543 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_555 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_563 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_567 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_600 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_608 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_612 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_619 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_658 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_711 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_715 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_724 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_736 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_767 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_774 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_13 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_84 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_301 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_313 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_333 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_343 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_479 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_503 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_532 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_582 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_594 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_598 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_614 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_644 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_656 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_684 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_688 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_695 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_37 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_58 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_67 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_94 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_151 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_159 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_171 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_262 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_344 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_396 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_507 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_555 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_566 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_596 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_608 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_662 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_687 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_726 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_730 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_13 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_17 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_25 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_30 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_78 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_123 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_148 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_190 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_231 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_311 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_344 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_368 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_431 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_519 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_535 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_556 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_572 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_578 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_590 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_614 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_628 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_632 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_636 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_670 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_17 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_25 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_44 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_56 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_64 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_107 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_218 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_226 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_323 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_336 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_430 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_442 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_512 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_566 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_586 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_595 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_603 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_615 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_622 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_668 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_674 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_687 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_724 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_736 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_767 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_10 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_88 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_189 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_200 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_368 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_459 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_471 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_542 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_573 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_593 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_648 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_668 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_679 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_703 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_775 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_60 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_72 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_130 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_151 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_288 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_300 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_331 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_500 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_543 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_555 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_567 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_611 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_620 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_711 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_715 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_739 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_768 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_775 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_30 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_37 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_88 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_108 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_119 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_140 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_305 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_352 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_370 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_380 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_407 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_502 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_519 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_543 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_571 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_575 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_583 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_698 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_710 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_734 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_738 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_747 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_771 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_50 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_154 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_190 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_226 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_326 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_347 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_441 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_506 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_510 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_520 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_537 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_612 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_616 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_620 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_654 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_658 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_662 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_675 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_682 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_686 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_762 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_14 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_22 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_63 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_77 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_134 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_155 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_162 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_198 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_220 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_243 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_252 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_308 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_388 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_424 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_428 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_503 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_517 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_535 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_538 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_642 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_670 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_690 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_754 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_767 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_16 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_37 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_99 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_103 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_115 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_172 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_282 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_326 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_448 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_501 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_555 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_564 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_580 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_619 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_656 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_660 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_680 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_699 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_716 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_723 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_738 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_768 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_43 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_48 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_68 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_75 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_148 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_179 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_191 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_261 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_305 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_366 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_455 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_469 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_491 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_528 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_558 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_569 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_578 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_586 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_678 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_682 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_704 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_739 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_747 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_768 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_48 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_58 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_66 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_95 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_107 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_152 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_291 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_458 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_550 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_604 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_614 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_658 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_665 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_723 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_8 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_30 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_90 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_179 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_305 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_323 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_386 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_407 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_427 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_460 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_484 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_496 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_523 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_535 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_573 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_591 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_600 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_640 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_652 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_684 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_704 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_715 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_739 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_746 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_772 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_38 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_47 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_58 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_112 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_378 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_402 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_414 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_603 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_615 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_631 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_667 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_680 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_684 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_768 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_775 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_13 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_37 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_179 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_189 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_411 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_422 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_503 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_519 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_535 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_547 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_571 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_583 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_606 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_622 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_641 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_696 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_775 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_17 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_46 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_58 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_106 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_163 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_170 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_176 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_248 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_268 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_288 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_379 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_431 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_435 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_474 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_494 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_506 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_514 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_544 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_612 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_624 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_650 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_658 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_682 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_712 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_720 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_768 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_36 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_64 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_71 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_98 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_110 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_179 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_191 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_245 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_470 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_529 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_549 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_554 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_626 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_632 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_642 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_648 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_670 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_687 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_697 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_707 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_751 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_767 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_46 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_211 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_264 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_605 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_650 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_658 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_662 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_674 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_684 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_708 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_767 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_46 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_78 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_298 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_310 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_407 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_484 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_529 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_585 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_635 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_647 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_685 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_711 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_749 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_773 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_108 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_160 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_172 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_217 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_224 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_232 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_319 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_323 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_392 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_431 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_613 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_638 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_708 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_714 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_721 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_731 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_743 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_9 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_32 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_79 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_91 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_143 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_196 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_208 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_303 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_368 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_478 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_573 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_591 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_629 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_650 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_683 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_695 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_702 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_714 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_727 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_746 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_770 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_776 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_96 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_206 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_288 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_401 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_452 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_543 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_555 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_585 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_627 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_655 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_667 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_719 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_728 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_734 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_768 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_775 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_28 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_143 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_176 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_186 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_198 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_458 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_594 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_627 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_639 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_651 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_727 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_742 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_746 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_767 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_775 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_56 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_104 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_116 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_434 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_458 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_622 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_767 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_774 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_135 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_179 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_191 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_709 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_726 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_758 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_771 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_36 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_116 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_157 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_206 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_374 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_402 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_654 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_658 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_682 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_694 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_767 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_25 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_88 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_231 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_240 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_252 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_260 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_268 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_316 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_408 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_420 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_471 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_515 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_539 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_595 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_615 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_631 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_655 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_664 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_688 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_700 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_712 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_722 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_754 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_766 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_775 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_22 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_67 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_98 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_157 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_224 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_339 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_441 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_450 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_507 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_514 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_526 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_544 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_568 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_643 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_651 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_654 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_664 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_676 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_688 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_721 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_767 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_13 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_22 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_48 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_61 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_148 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_200 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_541 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_579 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_592 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_633 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_642 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_654 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_693 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_705 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_726 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_747 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_771 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_48 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_80 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_158 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_170 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_208 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_336 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_375 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_398 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_485 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_657 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_697 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_710 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_718 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_738 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_775 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_30 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_124 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_142 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_179 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_258 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_709 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_726 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_748 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_772 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_776 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_39 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_95 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_116 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_163 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_207 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_219 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_315 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_336 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_431 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_443 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_546 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_568 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_609 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_620 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_626 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_665 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_679 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_728 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_739 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_743 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_768 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_136 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_260 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_422 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_462 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_466 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_529 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_575 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_583 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_596 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_608 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_715 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_40 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_44 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_102 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_127 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_134 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_154 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_275 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_443 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_550 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_597 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_609 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_621 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_641 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_656 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_668 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_680 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_692 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_762 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_766 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_775 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_34 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_75 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_132 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_238 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_247 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_267 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_292 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_324 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_525 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_693 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_704 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_726 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_743 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_766 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_90 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_107 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_115 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_207 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_219 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_322 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_375 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_512 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_549 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_613 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_625 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_636 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_659 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_706 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_718 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_732 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_743 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_754 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_761 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_770 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_776 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_68 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_80 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_198 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_302 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_318 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_411 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_422 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_430 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_456 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_480 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_529 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_588 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_612 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_629 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_642 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_650 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_682 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_693 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_705 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_743 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_767 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_152 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_263 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_275 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_318 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_322 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_458 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_632 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_699 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_716 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_720 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_726 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_734 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_44 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_79 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_86 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_92 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_146 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_193 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_239 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_397 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_411 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_420 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_431 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_470 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_502 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_511 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_532 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_582 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_629 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_660 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_697 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_709 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_720 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_735 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_744 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_750 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_771 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_13 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_40 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_96 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_157 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_269 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_499 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_723 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_732 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_767 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_16 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_30 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_37 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_87 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_118 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_199 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_299 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_311 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_319 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_347 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_357 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_454 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_515 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_539 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_559 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_572 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_596 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_608 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_629 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_654 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_666 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_775 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_10 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_22 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_42 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_70 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_340 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_560 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_572 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_667 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_687 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_711 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_767 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_67 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_79 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_140 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_144 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_180 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_208 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_232 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_467 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_633 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_641 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_692 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_705 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_64 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_72 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_202 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_214 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_226 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_487 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_499 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_555 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_567 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_607 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_699 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_715 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_730 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_767 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_774 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_14 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_30 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_90 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_148 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_432 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_442 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_483 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_529 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_541 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_581 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_592 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_598 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_627 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_639 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_651 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_727 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_743 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_767 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_775 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_159 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_318 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_330 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_346 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_379 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_598 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_606 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_618 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_630 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_662 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_767 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_32 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_63 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_72 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_140 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_368 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_374 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_480 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_548 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_596 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_626 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_638 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_648 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_683 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_687 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_699 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_711 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_722 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_767 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_34 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_42 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_82 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_151 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_163 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_207 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_398 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_487 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_555 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_559 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_599 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_611 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_623 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_643 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_658 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_682 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_694 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_723 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_735 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_775 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_160 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_274 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_310 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_413 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_422 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_582 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_593 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_641 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_653 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_664 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_752 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_764 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_96 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_116 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_172 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_206 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_339 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_487 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_499 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_620 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_632 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_669 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_681 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_692 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_707 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_716 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_722 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_726 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_753 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_775 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_75 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_200 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_347 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_359 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_371 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_458 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_693 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_703 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_715 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_51 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_112 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_136 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_163 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_203 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_213 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_270 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_282 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_320 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_398 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_458 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_564 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_576 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_595 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_608 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_620 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_654 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_665 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_677 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_733 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_744 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_768 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_775 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_10 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_14 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_74 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_86 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_150 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_179 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_214 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_301 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_323 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_330 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_366 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_462 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_581 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_591 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_685 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_697 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_705 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_735 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_40 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_112 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_318 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_327 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_339 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_531 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_550 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_667 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_677 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_737 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_743 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_752 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_21 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_28 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_98 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_102 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_109 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_119 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_143 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_155 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_312 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_418 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_476 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_542 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_588 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_592 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_627 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_636 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_648 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_660 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_714 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_740 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_744 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_90 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_152 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_208 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_244 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_347 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_612 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_631 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_655 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_667 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_679 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_718 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_767 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_20 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_25 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_92 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_295 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_347 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_420 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_496 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_519 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_540 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_685 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_705 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_151 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_207 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_219 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_378 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_394 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_460 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_488 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_500 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_506 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_543 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_555 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_567 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_657 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_677 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_749 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_754 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_761 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_770 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_776 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_10 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_36 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_70 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_311 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_346 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_368 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_469 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_540 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_552 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_579 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_598 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_610 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_627 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_639 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_651 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_727 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_735 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_745 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_775 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_12 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_49 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_103 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_152 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_164 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_176 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_184 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_319 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_495 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_504 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_516 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_543 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_548 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_560 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_627 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_655 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_675 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_689 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_712 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_716 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_728 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_732 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_767 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_235 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_239 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_347 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_415 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_485 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_502 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_534 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_628 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_652 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_664 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_685 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_726 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_775 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_18 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_35 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_51 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_107 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_136 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_297 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_302 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_319 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_326 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_376 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_492 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_504 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_508 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_611 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_638 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_699 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_715 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_735 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_753 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_763 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_21 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_71 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_90 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_136 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_160 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_200 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_357 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_468 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_476 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_577 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_586 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_592 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_631 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_685 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_708 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_720 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_735 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_749 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_760 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_764 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_34 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_82 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_172 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_184 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_215 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_227 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_272 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_322 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_346 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_375 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_553 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_565 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_611 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_618 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_654 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_658 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_670 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_674 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_682 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_711 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_723 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_731 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_743 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_768 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_21 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_133 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_180 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_241 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_415 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_469 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_478 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_510 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_522 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_534 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_543 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_547 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_573 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_598 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_610 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_626 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_652 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_656 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_666 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_692 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_704 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_716 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_742 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_754 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_766 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_774 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_18 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_63 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_327 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_339 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_507 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_542 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_554 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_566 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_572 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_606 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_616 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_36 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_162 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_182 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_202 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_258 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_416 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_515 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_528 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_546 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_697 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_715 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_722 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_756 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_763 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_46 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_58 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_132 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_158 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_170 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_176 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_336 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_342 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_379 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_395 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_435 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_514 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_526 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_562 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_566 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_576 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_657 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_675 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_709 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_728 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_733 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_753 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_774 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_38 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_180 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_200 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_243 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_252 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_260 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_403 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_476 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_615 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_627 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_639 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_651 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_671 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_683 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_703 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_710 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_722 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_749 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_46 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_58 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_64 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_219 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_414 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_432 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_530 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_557 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_567 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_625 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_642 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_661 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_711 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_723 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_735 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_755 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_763 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_36 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_52 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_84 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_108 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_122 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_142 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_212 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_267 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_346 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_354 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_364 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_411 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_420 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_583 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_595 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_615 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_632 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_644 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_693 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_702 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_735 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_738 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_749 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_34 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_60 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_68 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_102 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_114 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_190 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_475 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_600 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_611 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_623 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_655 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_667 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_679 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_762 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_773 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_19 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_76 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_118 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_142 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_146 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_191 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_291 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_303 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_429 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_466 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_46 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_58 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_90 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_163 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_230 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_327 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_339 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_392 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_437 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_463 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_602 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_606 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_624 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_636 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_669 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_680 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_775 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_26 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_82 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_94 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_102 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_179 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_261 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_308 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_368 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_415 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_424 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_482 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_502 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_515 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_583 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_595 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_694 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_706 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_718 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_746 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_48 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_56 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_80 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_94 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_104 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_116 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_168 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_207 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_219 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_290 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_374 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_398 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_490 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_514 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_568 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_724 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_736 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_748 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_753 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_770 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_32 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_36 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_78 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_129 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_136 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_148 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_346 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_350 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_455 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_465 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_559 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_572 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_576 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_588 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_612 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_639 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_649 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_685 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_705 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_747 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_752 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_760 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_766 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_62 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_82 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_99 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_132 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_152 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_210 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_219 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_656 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_660 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_672 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_684 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_712 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_762 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_774 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_18 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_25 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_32 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_42 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_110 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_135 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_154 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_212 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_243 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_247 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_259 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_292 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_296 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_312 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_626 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_646 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_655 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_687 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_63 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_104 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_150 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_159 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_219 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_378 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_402 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_439 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_448 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_504 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_528 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_547 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_669 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_713 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_773 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_12 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_36 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_80 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_95 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_243 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_255 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_291 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_303 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_347 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_367 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_473 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_485 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_535 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_577 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_727 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_96 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_150 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_157 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_203 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_215 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_227 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_340 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_543 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_555 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_573 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_730 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_21 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_34 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_75 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_87 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_180 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_214 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_236 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_240 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_295 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_310 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_347 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_399 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_406 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_523 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_532 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_592 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_604 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_691 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_727 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_760 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_772 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_104 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_116 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_158 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_248 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_259 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_286 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_555 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_570 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_582 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_603 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_607 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_620 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_632 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_669 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_721 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_733 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_34 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_75 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_118 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_185 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_235 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_247 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_291 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_303 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_487 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_496 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_542 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_559 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_572 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_588 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_612 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_630 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_650 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_670 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_681 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_690 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_705 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_62 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_92 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_102 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_114 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_267 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_339 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_441 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_459 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_555 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_664 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_676 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_688 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_767 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_28 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_44 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_48 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_79 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_95 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_180 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_188 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_196 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_211 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_424 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_513 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_524 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_540 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_574 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_583 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_595 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_49 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_92 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_112 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_202 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_228 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_263 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_267 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_322 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_376 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_394 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_549 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_608 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_620 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_632 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_665 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_674 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_767 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_34 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_46 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_79 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_120 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_127 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_145 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_176 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_200 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_348 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_384 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_420 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_458 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_466 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_517 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_591 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_637 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_651 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_671 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_693 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_705 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_749 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_755 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_764 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_46 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_56 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_101 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_114 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_152 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_224 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_282 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_450 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_488 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_510 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_540 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_544 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_568 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_620 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_632 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_669 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_681 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_698 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_716 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_747 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_754 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_763 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_72 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_134 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_186 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_198 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_221 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_231 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_252 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_291 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_347 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_364 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_413 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_480 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_581 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_628 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_652 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_664 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_727 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_748 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_773 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_126 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_156 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_168 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_210 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_218 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_226 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_296 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_401 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_434 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_458 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_485 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_507 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_569 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_711 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_738 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_28 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_62 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_86 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_90 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_133 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_151 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_196 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_208 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_216 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_301 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_315 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_370 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_515 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_539 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_598 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_610 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_641 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_653 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_664 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_703 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_725 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_738 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_75 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_170 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_203 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_207 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_227 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_264 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_276 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_443 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_564 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_576 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_661 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_669 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_725 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_768 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_92 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_100 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_119 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_143 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_182 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_191 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_129_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_302 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_311 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_346 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_431 ();
 sky130_fd_sc_hd__decap_3 FILLER_129_439 ();
 sky130_fd_sc_hd__decap_3 FILLER_129_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_472 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_484 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_525 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_534 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_542 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_558 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_577 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_588 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_612 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_638 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_650 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_722 ();
 sky130_fd_sc_hd__decap_3 FILLER_129_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_46 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_58 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_71 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_102 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_112 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_120 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_208 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_232 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_275 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_288 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_437 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_488 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_711 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_724 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_730 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_762 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_770 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_131_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_90 ();
 sky130_fd_sc_hd__decap_3 FILLER_131_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_110 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_129 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_131_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_210 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_252 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_302 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_413 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_423 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_131_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_471 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_131_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_590 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_651 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_131_693 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_705 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_747 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_62 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_134 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_170 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_190 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_213 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_347 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_375 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_387 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_443 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_484 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_504 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_516 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_543 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_555 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_575 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_585 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_600 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_612 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_623 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_657 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_712 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_724 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_736 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_753 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_770 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_21 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_122 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_134 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_146 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_183 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_187 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_254 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_359 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_413 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_583 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_595 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_637 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_648 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_660 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_704 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_716 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_738 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_747 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_759 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_763 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_767 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_33 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_42 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_66 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_105 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_224 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_236 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_282 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_331 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_431 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_563 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_575 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_620 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_632 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_657 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_668 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_713 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_764 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_771 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_21 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_28 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_43 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_64 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_88 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_127 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_174 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_206 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_238 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_256 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_291 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_466 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_472 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_484 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_492 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_633 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_646 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_693 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_724 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_744 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_771 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_64 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_103 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_150 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_262 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_320 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_398 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_430 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_492 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_514 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_669 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_733 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_28 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_63 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_75 ();
 sky130_fd_sc_hd__decap_3 FILLER_137_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_122 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_134 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_150 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_137_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_254 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_314 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_348 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_516 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_528 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_547 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_558 ();
 sky130_fd_sc_hd__decap_3 FILLER_137_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_590 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_628 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_652 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_664 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_711 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_750 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_34 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_42 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_64 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_134 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_159 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_171 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_179 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_227 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_288 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_375 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_494 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_531 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_543 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_555 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_600 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_611 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_623 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_654 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_666 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_678 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_722 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_732 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_742 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_767 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_34 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_75 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_92 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_100 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_140 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_151 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_162 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_182 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_245 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_252 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_384 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_526 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_538 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_554 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_653 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_695 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_726 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_738 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_742 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_43 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_140_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_140_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_172 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_184 ();
 sky130_fd_sc_hd__decap_3 FILLER_140_193 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_203 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_227 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_286 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_510 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_530 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_539 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_547 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_566 ();
 sky130_fd_sc_hd__decap_3 FILLER_140_574 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_625 ();
 sky130_fd_sc_hd__decap_3 FILLER_140_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_665 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_140_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_710 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_716 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_735 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_750 ();
 sky130_fd_sc_hd__decap_3 FILLER_140_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_763 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_141_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_63 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_70 ();
 sky130_fd_sc_hd__decap_3 FILLER_141_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_92 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_120 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_127 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_164 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_199 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_211 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_141_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_141_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_368 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_591 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_726 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_743 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_768 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_66 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_116 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_158 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_170 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_208 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_244 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_327 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_339 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_398 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_443 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_455 ();
 sky130_fd_sc_hd__decap_3 FILLER_142_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_486 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_510 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_530 ();
 sky130_fd_sc_hd__decap_3 FILLER_142_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_538 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_548 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_560 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_602 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_626 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_638 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_660 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_672 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_696 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_142_721 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_730 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_755 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_21 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_34 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_73 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_88 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_92 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_135 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_196 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_255 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_308 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_467 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_479 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_491 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_500 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_516 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_540 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_571 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_583 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_591 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_628 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_632 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_644 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_668 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_697 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_715 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_726 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_736 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_746 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_752 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_44 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_56 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_74 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_92 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_170 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_214 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_236 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_319 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_331 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_501 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_531 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_539 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_543 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_555 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_567 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_582 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_609 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_642 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_651 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_659 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_699 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_714 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_721 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_728 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_734 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_740 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_763 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_775 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_182 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_243 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_292 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_300 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_355 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_364 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_484 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_496 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_536 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_548 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_582 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_639 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_647 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_710 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_720 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_738 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_749 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_34 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_62 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_95 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_208 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_236 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_346 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_432 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_488 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_520 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_556 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_582 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_608 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_621 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_146_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_727 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_731 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_747 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_767 ();
 sky130_fd_sc_hd__decap_3 FILLER_146_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_63 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_75 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_87 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_98 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_123 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_130 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_186 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_292 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_326 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_347 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_415 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_500 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_535 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_584 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_614 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_628 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_632 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_671 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_679 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_689 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_714 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_724 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_46 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_58 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_104 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_122 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_172 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_204 ();
 sky130_fd_sc_hd__decap_3 FILLER_148_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_148_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_375 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_148_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_490 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_566 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_578 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_586 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_618 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_630 ();
 sky130_fd_sc_hd__decap_3 FILLER_148_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_665 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_680 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_696 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_710 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_717 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_767 ();
 sky130_fd_sc_hd__decap_3 FILLER_148_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_34 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_140 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_151 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_185 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_196 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_211 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_218 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_149_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_243 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_252 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_409 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_465 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_473 ();
 sky130_fd_sc_hd__decap_3 FILLER_149_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_524 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_558 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_584 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_642 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_654 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_670 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_691 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_707 ();
 sky130_fd_sc_hd__decap_3 FILLER_149_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_738 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_150_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_56 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_150_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_273 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_296 ();
 sky130_fd_sc_hd__decap_3 FILLER_150_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_338 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_150_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_428 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_452 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_512 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_531 ();
 sky130_fd_sc_hd__decap_3 FILLER_150_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_600 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_620 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_664 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_670 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_674 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_687 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_698 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_708 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_715 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_722 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_767 ();
 sky130_fd_sc_hd__decap_3 FILLER_150_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_63 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_75 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_120 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_156 ();
 sky130_fd_sc_hd__decap_3 FILLER_151_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_184 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_196 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_256 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_290 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_310 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_359 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_372 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_510 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_536 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_151_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_583 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_635 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_642 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_670 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_688 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_695 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_702 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_58 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_217 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_326 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_330 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_416 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_435 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_500 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_504 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_508 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_543 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_555 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_564 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_575 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_599 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_608 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_654 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_663 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_670 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_698 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_768 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_88 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_303 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_360 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_424 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_581 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_594 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_600 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_622 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_637 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_670 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_682 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_702 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_759 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_768 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_46 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_58 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_130 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_171 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_259 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_346 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_495 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_504 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_600 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_604 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_626 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_650 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_662 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_666 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_670 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_674 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_678 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_687 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_738 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_155_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_92 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_104 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_142 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_151 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_155_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_155_301 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_356 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_375 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_384 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_155_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_155_445 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_476 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_586 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_590 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_640 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_647 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_664 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_688 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_692 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_739 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_747 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_768 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_39 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_63 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_115 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_158 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_168 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_183 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_190 ();
 sky130_fd_sc_hd__decap_3 FILLER_156_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_228 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_239 ();
 sky130_fd_sc_hd__decap_3 FILLER_156_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_339 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_375 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_387 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_466 ();
 sky130_fd_sc_hd__decap_3 FILLER_156_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_515 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_552 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_562 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_643 ();
 sky130_fd_sc_hd__decap_3 FILLER_156_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_651 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_676 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_156_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_768 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_21 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_34 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_50 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_70 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_82 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_91 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_124 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_135 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_143 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_183 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_198 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_206 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_247 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_292 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_423 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_510 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_514 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_536 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_548 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_556 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_573 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_634 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_638 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_648 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_696 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_715 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_110 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_119 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_148 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_173 ();
 sky130_fd_sc_hd__decap_3 FILLER_158_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_226 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_158_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_376 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_396 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_443 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_500 ();
 sky130_fd_sc_hd__decap_3 FILLER_158_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_524 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_564 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_604 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_665 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_158_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_711 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_715 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_736 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_768 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_34 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_70 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_164 ();
 sky130_fd_sc_hd__decap_3 FILLER_159_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_203 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_303 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_359 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_375 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_384 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_424 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_159_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_159_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_556 ();
 sky130_fd_sc_hd__decap_3 FILLER_159_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_590 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_594 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_604 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_683 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_703 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_739 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_747 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_34 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_49 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_58 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_203 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_213 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_258 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_276 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_283 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_329 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_340 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_371 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_392 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_436 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_448 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_499 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_506 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_519 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_526 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_547 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_578 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_663 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_698 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_706 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_730 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_738 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_762 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_64 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_88 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_189 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_161_202 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_236 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_257 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_478 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_490 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_516 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_558 ();
 sky130_fd_sc_hd__decap_3 FILLER_161_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_574 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_581 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_594 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_641 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_653 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_688 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_698 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_702 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_739 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_747 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_771 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_162_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_75 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_116 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_172 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_162_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_228 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_375 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_387 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_407 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_445 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_528 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_539 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_543 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_563 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_570 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_606 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_610 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_666 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_678 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_711 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_718 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_724 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_734 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_747 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_768 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_28 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_75 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_134 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_148 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_179 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_186 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_198 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_270 ();
 sky130_fd_sc_hd__decap_3 FILLER_163_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_163_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_354 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_420 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_469 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_558 ();
 sky130_fd_sc_hd__decap_3 FILLER_163_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_578 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_590 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_598 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_639 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_646 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_703 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_39 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_49 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_60 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_78 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_122 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_168 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_192 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_203 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_207 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_260 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_295 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_320 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_338 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_402 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_414 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_563 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_586 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_622 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_634 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_642 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_651 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_660 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_687 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_723 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_747 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_767 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_86 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_130 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_142 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_160 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_198 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_165_245 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_254 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_165_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_368 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_403 ();
 sky130_fd_sc_hd__decap_3 FILLER_165_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_479 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_491 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_547 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_566 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_588 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_614 ();
 sky130_fd_sc_hd__decap_3 FILLER_165_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_628 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_632 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_637 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_644 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_658 ();
 sky130_fd_sc_hd__decap_3 FILLER_165_669 ();
 sky130_fd_sc_hd__decap_3 FILLER_165_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_684 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_696 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_726 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_735 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_745 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_49 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_72 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_204 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_216 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_228 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_236 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_268 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_283 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_296 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_324 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_336 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_450 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_472 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_491 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_503 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_555 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_566 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_576 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_596 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_609 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_642 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_684 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_731 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_768 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_28 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_176 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_200 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_242 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_308 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_167_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_167_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_479 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_500 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_519 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_532 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_546 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_559 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_575 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_582 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_684 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_688 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_775 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_14 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_18 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_24 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_64 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_76 ();
 sky130_fd_sc_hd__decap_3 FILLER_168_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_116 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_238 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_282 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_339 ();
 sky130_fd_sc_hd__decap_3 FILLER_168_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_376 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_394 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_652 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_677 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_683 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_712 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_767 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_79 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_103 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_124 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_143 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_152 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_367 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_407 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_436 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_500 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_525 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_550 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_603 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_639 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_646 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_683 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_698 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_710 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_763 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_775 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_48 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_61 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_228 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_236 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_282 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_336 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_383 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_438 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_448 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_506 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_555 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_626 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_655 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_662 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_676 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_690 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_723 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_731 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_768 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_775 ();
 sky130_fd_sc_hd__decap_3 FILLER_171_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_21 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_26 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_104 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_142 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_171_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_242 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_303 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_320 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_348 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_366 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_171_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_459 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_550 ();
 sky130_fd_sc_hd__decap_3 FILLER_171_557 ();
 sky130_fd_sc_hd__decap_3 FILLER_171_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_595 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_622 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_650 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_695 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_764 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_768 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_46 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_52 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_127 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_134 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_171 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_179 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_215 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_227 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_266 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_172_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_396 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_444 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_499 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_611 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_623 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_636 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_683 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_687 ();
 sky130_fd_sc_hd__decap_3 FILLER_172_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_9 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_16 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_75 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_119 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_142 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_174 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_198 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_208 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_230 ();
 sky130_fd_sc_hd__decap_3 FILLER_173_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_247 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_173_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_287 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_409 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_429 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_454 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_479 ();
 sky130_fd_sc_hd__decap_3 FILLER_173_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_527 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_649 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_655 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_671 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_173_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_740 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_116 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_128 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_155 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_248 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_267 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_351 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_372 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_400 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_514 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_594 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_600 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_610 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_618 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_665 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_669 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_680 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_712 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_723 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_738 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_742 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_767 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_21 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_32 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_40 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_101 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_186 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_198 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_242 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_175_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_304 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_386 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_422 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_446 ();
 sky130_fd_sc_hd__decap_3 FILLER_175_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_510 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_542 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_579 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_634 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_646 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_656 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_678 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_682 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_703 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_716 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_763 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_775 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_56 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_71 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_102 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_127 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_264 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_176_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_463 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_470 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_486 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_507 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_572 ();
 sky130_fd_sc_hd__decap_3 FILLER_176_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_596 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_623 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_663 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_672 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_684 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_698 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_716 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_176_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_767 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_771 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_44 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_64 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_88 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_140 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_303 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_311 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_574 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_695 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_702 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_754 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_766 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_775 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_38 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_46 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_82 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_178_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_182 ();
 sky130_fd_sc_hd__decap_3 FILLER_178_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_204 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_216 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_242 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_282 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_339 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_348 ();
 sky130_fd_sc_hd__decap_3 FILLER_178_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_385 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_458 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_552 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_595 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_622 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_628 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_659 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_680 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_706 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_710 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_720 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_732 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_762 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_766 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_179_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_37 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_64 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_87 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_179_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_132 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_152 ();
 sky130_fd_sc_hd__decap_3 FILLER_179_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_198 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_255 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_310 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_368 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_414 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_424 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_435 ();
 sky130_fd_sc_hd__decap_3 FILLER_179_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_459 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_479 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_559 ();
 sky130_fd_sc_hd__decap_3 FILLER_179_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_570 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_625 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_652 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_684 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_704 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_739 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_751 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_772 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_13 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_17 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_180_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_180_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_48 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_58 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_82 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_99 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_320 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_397 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_444 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_452 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_458 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_586 ();
 sky130_fd_sc_hd__decap_3 FILLER_180_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_659 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_680 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_712 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_724 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_730 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_739 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_775 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_10 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_18 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_181_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_238 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_367 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_594 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_636 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_640 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_662 ();
 sky130_fd_sc_hd__decap_3 FILLER_181_669 ();
 sky130_fd_sc_hd__decap_3 FILLER_181_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_696 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_700 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_739 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_743 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_764 ();
 sky130_fd_sc_hd__decap_3 FILLER_181_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_36 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_64 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_116 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_168 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_216 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_228 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_272 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_320 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_394 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_451 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_464 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_572 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_600 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_627 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_670 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_674 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_678 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_725 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_737 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_754 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_768 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_30 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_76 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_86 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_100 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_134 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_144 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_206 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_252 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_297 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_388 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_399 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_423 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_484 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_508 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_537 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_571 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_598 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_614 ();
 sky130_fd_sc_hd__decap_3 FILLER_183_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_641 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_654 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_666 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_697 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_775 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_39 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_49 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_90 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_102 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_107 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_172 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_184_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_208 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_242 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_282 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_338 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_474 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_494 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_506 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_514 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_614 ();
 sky130_fd_sc_hd__decap_3 FILLER_184_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_667 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_679 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_698 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_714 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_738 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_750 ();
 sky130_fd_sc_hd__decap_3 FILLER_184_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_768 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_775 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_31 ();
 sky130_fd_sc_hd__decap_8 FILLER_185_40 ();
 sky130_fd_sc_hd__decap_3 FILLER_185_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_62 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_76 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_86 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_95 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_134 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_185_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_185_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_247 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_252 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_294 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_359 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_376 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_185_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_185_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_459 ();
 sky130_fd_sc_hd__decap_8 FILLER_185_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_515 ();
 sky130_fd_sc_hd__decap_8 FILLER_185_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_535 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_583 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_639 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_651 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_695 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_767 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_26 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_39 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_59 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_96 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_106 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_210 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_219 ();
 sky130_fd_sc_hd__decap_3 FILLER_186_227 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_325 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_374 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_458 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_470 ();
 sky130_fd_sc_hd__decap_3 FILLER_186_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_558 ();
 sky130_fd_sc_hd__decap_3 FILLER_186_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_611 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_667 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_679 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_711 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_723 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_754 ();
 sky130_fd_sc_hd__decap_3 FILLER_186_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_768 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_44 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_78 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_120 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_131 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_142 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_150 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_189 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_200 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_245 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_308 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_436 ();
 sky130_fd_sc_hd__decap_3 FILLER_187_445 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_502 ();
 sky130_fd_sc_hd__decap_3 FILLER_187_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_581 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_594 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_695 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_739 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_743 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_764 ();
 sky130_fd_sc_hd__decap_3 FILLER_187_774 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_10 ();
 sky130_fd_sc_hd__decap_8 FILLER_188_14 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_46 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_59 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_66 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_78 ();
 sky130_fd_sc_hd__decap_3 FILLER_188_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_103 ();
 sky130_fd_sc_hd__decap_8 FILLER_188_114 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_152 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_161 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_173 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_188_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_188_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_188_244 ();
 sky130_fd_sc_hd__decap_3 FILLER_188_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_319 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_329 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_188_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_375 ();
 sky130_fd_sc_hd__decap_3 FILLER_188_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_395 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_410 ();
 sky130_fd_sc_hd__decap_3 FILLER_188_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_432 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_502 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_556 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_568 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_574 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_611 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_626 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_667 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_679 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_723 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_189_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_189_23 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_74 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_189_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_198 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_189_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_189_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_310 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_366 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_415 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_428 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_189_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_478 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_540 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_559 ();
 sky130_fd_sc_hd__decap_3 FILLER_189_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_584 ();
 sky130_fd_sc_hd__decap_8 FILLER_189_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_679 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_693 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_189_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_775 ();
 sky130_fd_sc_hd__decap_8 FILLER_190_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_190_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_17 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_26 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_52 ();
 sky130_fd_sc_hd__decap_8 FILLER_190_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_190_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_190_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_190_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_170 ();
 sky130_fd_sc_hd__decap_8 FILLER_190_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_190_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_331 ();
 sky130_fd_sc_hd__decap_8 FILLER_190_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_190_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_392 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_190_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_564 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_584 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_190_641 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_651 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_724 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_728 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_13 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_42 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_50 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_98 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_123 ();
 sky130_fd_sc_hd__decap_8 FILLER_191_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_143 ();
 sky130_fd_sc_hd__decap_8 FILLER_191_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_252 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_301 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_313 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_354 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_358 ();
 sky130_fd_sc_hd__decap_8 FILLER_191_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_378 ();
 sky130_fd_sc_hd__decap_3 FILLER_191_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_191_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_502 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_532 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_584 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_615 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_670 ();
 sky130_fd_sc_hd__decap_8 FILLER_191_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_702 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_712 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_726 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_735 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_752 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_758 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_775 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_12 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_20 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_48 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_59 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_94 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_112 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_164 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_226 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_340 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_192_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_386 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_441 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_463 ();
 sky130_fd_sc_hd__decap_3 FILLER_192_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_483 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_549 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_566 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_719 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_746 ();
 sky130_fd_sc_hd__decap_3 FILLER_192_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_775 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_71 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_82 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_110 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_193_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_267 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_193_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_319 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_330 ();
 sky130_fd_sc_hd__decap_3 FILLER_193_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_193_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_558 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_747 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_775 ();
endmodule
