VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO caravan_signal_routing
  CLASS BLOCK ;
  FOREIGN caravan_signal_routing ;
  ORIGIN -98.815 -4489.235 ;
  SIZE 3390.220 BY 600.000 ;
  OBS
      LAYER met3 ;
        RECT 198.820 4489.235 3389.030 4989.230 ;
        POLYGON 322.540 4214.800 322.540 4212.290 320.030 4212.290 ;
        RECT 322.540 4212.290 326.540 4214.800 ;
        RECT 199.500 4190.800 326.540 4212.290 ;
        RECT 199.500 4188.390 320.760 4190.800 ;
        POLYGON 320.760 4190.800 323.170 4190.800 320.760 4188.390 ;
        RECT 3246.540 4166.505 3250.540 4170.400 ;
        POLYGON 322.540 4164.800 322.540 4162.395 320.135 4162.395 ;
        RECT 322.540 4162.395 326.540 4164.800 ;
        RECT 199.500 4140.800 326.540 4162.395 ;
        RECT 3246.540 4146.400 3388.160 4166.505 ;
        RECT 3249.290 4142.605 3388.160 4146.400 ;
        RECT 249.460 4140.795 323.170 4140.800 ;
        RECT 199.500 4138.495 320.870 4140.795 ;
        POLYGON 320.870 4140.795 323.170 4140.795 320.870 4138.495 ;
        RECT 3246.540 4116.610 3250.540 4120.400 ;
        RECT 3246.540 4096.400 3388.160 4116.610 ;
        RECT 3249.290 4092.710 3388.160 4096.400 ;
        RECT 3246.540 2593.505 3250.540 2593.740 ;
        RECT 3246.540 2569.740 3388.160 2593.505 ;
        RECT 3250.290 2569.605 3335.580 2569.740 ;
        RECT 3246.540 2543.610 3250.540 2543.740 ;
        RECT 3246.540 2519.740 3388.160 2543.610 ;
        RECT 3250.330 2519.710 3335.620 2519.740 ;
        POLYGON 322.540 2492.030 322.540 2489.290 319.800 2489.290 ;
        RECT 322.540 2489.290 326.540 2492.030 ;
        RECT 199.500 2468.030 326.540 2489.290 ;
        RECT 199.500 2465.390 320.060 2468.030 ;
        POLYGON 320.060 2468.030 322.700 2468.030 320.060 2465.390 ;
        POLYGON 322.540 2442.025 322.540 2439.395 319.910 2439.395 ;
        RECT 322.540 2439.395 326.540 2442.030 ;
        RECT 199.500 2418.030 326.540 2439.395 ;
        RECT 199.500 2415.495 320.205 2418.030 ;
        POLYGON 320.205 2418.030 322.740 2418.030 320.205 2415.495 ;
        RECT 3246.540 2373.500 3250.540 2374.740 ;
        RECT 3246.540 2350.740 3380.890 2373.500 ;
        RECT 3250.210 2349.500 3380.890 2350.740 ;
        RECT 3246.540 2323.245 3250.540 2324.740 ;
        RECT 3246.540 2300.740 3380.890 2323.245 ;
        RECT 3250.210 2299.300 3380.890 2300.740 ;
        POLYGON 322.540 2282.030 322.540 2278.700 319.210 2278.700 ;
        RECT 322.540 2278.700 326.540 2282.030 ;
        RECT 207.000 2258.030 326.540 2278.700 ;
        RECT 207.000 2254.755 319.635 2258.030 ;
        POLYGON 319.635 2258.030 322.910 2258.030 319.635 2254.755 ;
        POLYGON 322.540 2232.030 322.540 2228.500 319.010 2228.500 ;
        RECT 322.540 2228.500 326.540 2232.030 ;
        RECT 207.000 2208.030 326.540 2228.500 ;
        RECT 207.000 2204.500 319.290 2208.030 ;
        POLYGON 319.290 2208.030 322.820 2208.030 319.290 2204.500 ;
        RECT 3250.340 2151.740 3388.380 2152.505 ;
        RECT 3246.540 2128.605 3388.380 2151.740 ;
        RECT 3246.540 2127.810 3385.120 2128.605 ;
        RECT 3246.540 2127.740 3250.540 2127.810 ;
        RECT 3250.290 2101.740 3388.380 2102.610 ;
        RECT 3246.540 2078.710 3388.380 2101.740 ;
        RECT 3246.540 2077.740 3250.540 2078.710 ;
      LAYER met4 ;
        RECT 1105.000 4913.590 2046.000 4980.100 ;
      LAYER met5 ;
        RECT 1105.000 4913.590 2046.000 4980.100 ;
  END
END caravan_signal_routing
END LIBRARY

