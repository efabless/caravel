* NGSPICE file created from housekeeping.ext - technology: sky130A

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_2 abstract view
.subckt sky130_fd_sc_hd__dfstp_2 CLK D SET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_4 abstract view
.subckt sky130_fd_sc_hd__dfrtp_4 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_1 abstract view
.subckt sky130_fd_sc_hd__dfrtp_1 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_4 abstract view
.subckt sky130_fd_sc_hd__or3b_4 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_1 abstract view
.subckt sky130_fd_sc_hd__o32a_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd3_1 abstract view
.subckt sky130_fd_sc_hd__dlygate4sd3_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_1 abstract view
.subckt sky130_fd_sc_hd__nand3b_1 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_2 abstract view
.subckt sky130_fd_sc_hd__o21a_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_1 abstract view
.subckt sky130_fd_sc_hd__o41a_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_2 abstract view
.subckt sky130_fd_sc_hd__dfrtp_2 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_4 abstract view
.subckt sky130_fd_sc_hd__and3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_12 abstract view
.subckt sky130_fd_sc_hd__buf_12 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_1 abstract view
.subckt sky130_fd_sc_hd__dfstp_1 CLK D SET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_2 abstract view
.subckt sky130_fd_sc_hd__a22o_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_8 abstract view
.subckt sky130_fd_sc_hd__nor2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_4 abstract view
.subckt sky130_fd_sc_hd__or4b_4 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_1 abstract view
.subckt sky130_fd_sc_hd__o311a_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4b_1 abstract view
.subckt sky130_fd_sc_hd__nor4b_1 A B C D_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_4 abstract view
.subckt sky130_fd_sc_hd__o221ai_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_1 abstract view
.subckt sky130_fd_sc_hd__o31ai_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_4 abstract view
.subckt sky130_fd_sc_hd__or2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_4 abstract view
.subckt sky130_fd_sc_hd__dfstp_4 CLK D SET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_1 abstract view
.subckt sky130_fd_sc_hd__a2111o_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_1 abstract view
.subckt sky130_fd_sc_hd__and4b_1 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_2 abstract view
.subckt sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_4 abstract view
.subckt sky130_fd_sc_hd__nand2b_4 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_4 abstract view
.subckt sky130_fd_sc_hd__and2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_1 abstract view
.subckt sky130_fd_sc_hd__a41o_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_8 abstract view
.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_1 abstract view
.subckt sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_4 abstract view
.subckt sky130_fd_sc_hd__nor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_1 abstract view
.subckt sky130_fd_sc_hd__and4bb_1 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_8 abstract view
.subckt sky130_fd_sc_hd__nand2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_2 abstract view
.subckt sky130_fd_sc_hd__and2b_2 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_2 abstract view
.subckt sky130_fd_sc_hd__or3b_2 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_4 abstract view
.subckt sky130_fd_sc_hd__and3b_4 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_1 abstract view
.subckt sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_1 abstract view
.subckt sky130_fd_sc_hd__nor4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_1 abstract view
.subckt sky130_fd_sc_hd__nand4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_2 abstract view
.subckt sky130_fd_sc_hd__a221o_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_2 abstract view
.subckt sky130_fd_sc_hd__clkinv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_1 abstract view
.subckt sky130_fd_sc_hd__o2111a_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_1 abstract view
.subckt sky130_fd_sc_hd__a221oi_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_2 abstract view
.subckt sky130_fd_sc_hd__a2111o_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_2 abstract view
.subckt sky130_fd_sc_hd__and4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_1 abstract view
.subckt sky130_fd_sc_hd__o211ai_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_1 abstract view
.subckt sky130_fd_sc_hd__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_4 abstract view
.subckt sky130_fd_sc_hd__o221a_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_2 abstract view
.subckt sky130_fd_sc_hd__nor4_2 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_1 abstract view
.subckt sky130_fd_sc_hd__a211oi_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_4 abstract view
.subckt sky130_fd_sc_hd__a2111o_4 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_4 abstract view
.subckt sky130_fd_sc_hd__mux2_4 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_1 abstract view
.subckt sky130_fd_sc_hd__or4bb_1 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_4 abstract view
.subckt sky130_fd_sc_hd__a221oi_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_4 abstract view
.subckt sky130_fd_sc_hd__and2b_4 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_4 abstract view
.subckt sky130_fd_sc_hd__nand3b_4 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_1 abstract view
.subckt sky130_fd_sc_hd__nand2b_1 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtn_1 abstract view
.subckt sky130_fd_sc_hd__dfrtn_1 CLK_N D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_4 abstract view
.subckt sky130_fd_sc_hd__a221o_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_2 abstract view
.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_2 abstract view
.subckt sky130_fd_sc_hd__o211a_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_4 abstract view
.subckt sky130_fd_sc_hd__and4b_4 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_2 abstract view
.subckt sky130_fd_sc_hd__mux2_2 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_2 abstract view
.subckt sky130_fd_sc_hd__or4b_2 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_2 abstract view
.subckt sky130_fd_sc_hd__nor3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_2 abstract view
.subckt sky130_fd_sc_hd__a211o_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_2 abstract view
.subckt sky130_fd_sc_hd__o221a_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_2 abstract view
.subckt sky130_fd_sc_hd__and3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_4 abstract view
.subckt sky130_fd_sc_hd__a21oi_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_4 abstract view
.subckt sky130_fd_sc_hd__o21ai_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_4 abstract view
.subckt sky130_fd_sc_hd__a41o_4 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4b_1 abstract view
.subckt sky130_fd_sc_hd__nand4b_1 A_N B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_1 abstract view
.subckt sky130_fd_sc_hd__o221ai_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_4 abstract view
.subckt sky130_fd_sc_hd__or4bb_4 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_1 abstract view
.subckt sky130_fd_sc_hd__a22oi_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_8 abstract view
.subckt sky130_fd_sc_hd__mux2_8 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_4 abstract view
.subckt sky130_fd_sc_hd__xnor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_4 abstract view
.subckt sky130_fd_sc_hd__o211ai_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_4 abstract view
.subckt sky130_fd_sc_hd__nor3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_2 abstract view
.subckt sky130_fd_sc_hd__nand3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_2 abstract view
.subckt sky130_fd_sc_hd__and3b_2 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_4 abstract view
.subckt sky130_fd_sc_hd__nor3b_4 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_6 abstract view
.subckt sky130_fd_sc_hd__inv_6 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_4 abstract view
.subckt sky130_fd_sc_hd__nand3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

.subckt housekeeping VGND VPWR debug_in debug_mode debug_oeb debug_out irq[0] irq[1]
+ irq[2] mask_rev_in[0] mask_rev_in[10] mask_rev_in[11] mask_rev_in[12] mask_rev_in[13]
+ mask_rev_in[14] mask_rev_in[15] mask_rev_in[16] mask_rev_in[17] mask_rev_in[18]
+ mask_rev_in[19] mask_rev_in[1] mask_rev_in[20] mask_rev_in[21] mask_rev_in[22] mask_rev_in[23]
+ mask_rev_in[24] mask_rev_in[25] mask_rev_in[26] mask_rev_in[27] mask_rev_in[28]
+ mask_rev_in[29] mask_rev_in[2] mask_rev_in[30] mask_rev_in[31] mask_rev_in[3] mask_rev_in[4]
+ mask_rev_in[5] mask_rev_in[6] mask_rev_in[7] mask_rev_in[8] mask_rev_in[9] mgmt_gpio_in[0]
+ mgmt_gpio_in[10] mgmt_gpio_in[11] mgmt_gpio_in[12] mgmt_gpio_in[13] mgmt_gpio_in[14]
+ mgmt_gpio_in[15] mgmt_gpio_in[16] mgmt_gpio_in[17] mgmt_gpio_in[18] mgmt_gpio_in[19]
+ mgmt_gpio_in[1] mgmt_gpio_in[20] mgmt_gpio_in[21] mgmt_gpio_in[22] mgmt_gpio_in[23]
+ mgmt_gpio_in[24] mgmt_gpio_in[25] mgmt_gpio_in[26] mgmt_gpio_in[27] mgmt_gpio_in[28]
+ mgmt_gpio_in[29] mgmt_gpio_in[2] mgmt_gpio_in[30] mgmt_gpio_in[31] mgmt_gpio_in[32]
+ mgmt_gpio_in[33] mgmt_gpio_in[34] mgmt_gpio_in[35] mgmt_gpio_in[36] mgmt_gpio_in[37]
+ mgmt_gpio_in[3] mgmt_gpio_in[4] mgmt_gpio_in[5] mgmt_gpio_in[6] mgmt_gpio_in[7]
+ mgmt_gpio_in[8] mgmt_gpio_in[9] mgmt_gpio_oeb[0] mgmt_gpio_oeb[10] mgmt_gpio_oeb[11]
+ mgmt_gpio_oeb[12] mgmt_gpio_oeb[13] mgmt_gpio_oeb[14] mgmt_gpio_oeb[15] mgmt_gpio_oeb[16]
+ mgmt_gpio_oeb[17] mgmt_gpio_oeb[18] mgmt_gpio_oeb[19] mgmt_gpio_oeb[1] mgmt_gpio_oeb[20]
+ mgmt_gpio_oeb[21] mgmt_gpio_oeb[22] mgmt_gpio_oeb[23] mgmt_gpio_oeb[24] mgmt_gpio_oeb[25]
+ mgmt_gpio_oeb[26] mgmt_gpio_oeb[27] mgmt_gpio_oeb[28] mgmt_gpio_oeb[29] mgmt_gpio_oeb[2]
+ mgmt_gpio_oeb[30] mgmt_gpio_oeb[31] mgmt_gpio_oeb[32] mgmt_gpio_oeb[33] mgmt_gpio_oeb[34]
+ mgmt_gpio_oeb[35] mgmt_gpio_oeb[36] mgmt_gpio_oeb[37] mgmt_gpio_oeb[3] mgmt_gpio_oeb[4]
+ mgmt_gpio_oeb[5] mgmt_gpio_oeb[6] mgmt_gpio_oeb[7] mgmt_gpio_oeb[8] mgmt_gpio_oeb[9]
+ mgmt_gpio_out[0] mgmt_gpio_out[10] mgmt_gpio_out[11] mgmt_gpio_out[12] mgmt_gpio_out[13]
+ mgmt_gpio_out[14] mgmt_gpio_out[15] mgmt_gpio_out[16] mgmt_gpio_out[17] mgmt_gpio_out[18]
+ mgmt_gpio_out[19] mgmt_gpio_out[1] mgmt_gpio_out[20] mgmt_gpio_out[21] mgmt_gpio_out[22]
+ mgmt_gpio_out[23] mgmt_gpio_out[24] mgmt_gpio_out[25] mgmt_gpio_out[26] mgmt_gpio_out[27]
+ mgmt_gpio_out[28] mgmt_gpio_out[29] mgmt_gpio_out[2] mgmt_gpio_out[30] mgmt_gpio_out[31]
+ mgmt_gpio_out[32] mgmt_gpio_out[33] mgmt_gpio_out[34] mgmt_gpio_out[35] mgmt_gpio_out[36]
+ mgmt_gpio_out[37] mgmt_gpio_out[3] mgmt_gpio_out[4] mgmt_gpio_out[5] mgmt_gpio_out[6]
+ mgmt_gpio_out[7] mgmt_gpio_out[8] mgmt_gpio_out[9] pad_flash_clk pad_flash_clk_oeb
+ pad_flash_csb pad_flash_csb_oeb pad_flash_io0_di pad_flash_io0_do pad_flash_io0_ieb
+ pad_flash_io0_oeb pad_flash_io1_di pad_flash_io1_do pad_flash_io1_ieb pad_flash_io1_oeb
+ pll90_sel[0] pll90_sel[1] pll90_sel[2] pll_bypass pll_dco_ena pll_div[0] pll_div[1]
+ pll_div[2] pll_div[3] pll_div[4] pll_ena pll_sel[0] pll_sel[1] pll_sel[2] pll_trim[0]
+ pll_trim[10] pll_trim[11] pll_trim[12] pll_trim[13] pll_trim[14] pll_trim[15] pll_trim[16]
+ pll_trim[17] pll_trim[18] pll_trim[19] pll_trim[1] pll_trim[20] pll_trim[21] pll_trim[22]
+ pll_trim[23] pll_trim[24] pll_trim[25] pll_trim[2] pll_trim[3] pll_trim[4] pll_trim[5]
+ pll_trim[6] pll_trim[7] pll_trim[8] pll_trim[9] porb pwr_ctrl_out[0] pwr_ctrl_out[1]
+ pwr_ctrl_out[2] pwr_ctrl_out[3] qspi_enabled reset ser_rx ser_tx serial_clock serial_data_1
+ serial_data_2 serial_load serial_resetn spi_csb spi_enabled spi_sck spi_sdi spi_sdo
+ spi_sdoenb spimemio_flash_clk spimemio_flash_csb spimemio_flash_io0_di spimemio_flash_io0_do
+ spimemio_flash_io0_oeb spimemio_flash_io1_di spimemio_flash_io1_do spimemio_flash_io1_oeb
+ spimemio_flash_io2_di spimemio_flash_io2_do spimemio_flash_io2_oeb spimemio_flash_io3_di
+ spimemio_flash_io3_do spimemio_flash_io3_oeb trap uart_enabled user_clock usr1_vcc_pwrgood
+ usr1_vdd_pwrgood usr2_vcc_pwrgood usr2_vdd_pwrgood wb_ack_o wb_adr_i[0] wb_adr_i[10]
+ wb_adr_i[11] wb_adr_i[12] wb_adr_i[13] wb_adr_i[14] wb_adr_i[15] wb_adr_i[16] wb_adr_i[17]
+ wb_adr_i[18] wb_adr_i[19] wb_adr_i[1] wb_adr_i[20] wb_adr_i[21] wb_adr_i[22] wb_adr_i[23]
+ wb_adr_i[24] wb_adr_i[25] wb_adr_i[26] wb_adr_i[27] wb_adr_i[28] wb_adr_i[29] wb_adr_i[2]
+ wb_adr_i[30] wb_adr_i[31] wb_adr_i[3] wb_adr_i[4] wb_adr_i[5] wb_adr_i[6] wb_adr_i[7]
+ wb_adr_i[8] wb_adr_i[9] wb_clk_i wb_cyc_i wb_dat_i[0] wb_dat_i[10] wb_dat_i[11]
+ wb_dat_i[12] wb_dat_i[13] wb_dat_i[14] wb_dat_i[15] wb_dat_i[16] wb_dat_i[17] wb_dat_i[18]
+ wb_dat_i[19] wb_dat_i[1] wb_dat_i[20] wb_dat_i[21] wb_dat_i[22] wb_dat_i[23] wb_dat_i[24]
+ wb_dat_i[25] wb_dat_i[26] wb_dat_i[27] wb_dat_i[28] wb_dat_i[29] wb_dat_i[2] wb_dat_i[30]
+ wb_dat_i[31] wb_dat_i[3] wb_dat_i[4] wb_dat_i[5] wb_dat_i[6] wb_dat_i[7] wb_dat_i[8]
+ wb_dat_i[9] wb_dat_o[0] wb_dat_o[10] wb_dat_o[11] wb_dat_o[12] wb_dat_o[13] wb_dat_o[14]
+ wb_dat_o[15] wb_dat_o[16] wb_dat_o[17] wb_dat_o[18] wb_dat_o[19] wb_dat_o[1] wb_dat_o[20]
+ wb_dat_o[21] wb_dat_o[22] wb_dat_o[23] wb_dat_o[24] wb_dat_o[25] wb_dat_o[26] wb_dat_o[27]
+ wb_dat_o[28] wb_dat_o[29] wb_dat_o[2] wb_dat_o[30] wb_dat_o[31] wb_dat_o[3] wb_dat_o[4]
+ wb_dat_o[5] wb_dat_o[6] wb_dat_o[7] wb_dat_o[8] wb_dat_o[9] wb_rstn_i wb_sel_i[0]
+ wb_sel_i[1] wb_sel_i[2] wb_sel_i[3] wb_stb_i wb_we_i
XFILLER_67_520 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6914_ _7010_/CLK _6914_/D fanout498/X VGND VGND VPWR VPWR _6914_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_35_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6845_ _7069_/CLK _6845_/D fanout516/X VGND VGND VPWR VPWR _6845_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_52_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6776_ _6881_/CLK _6776_/D fanout523/X VGND VGND VPWR VPWR _7195_/A sky130_fd_sc_hd__dfrtp_1
X_3988_ hold499/X _5491_/A1 _3992_/S VGND VGND VPWR VPWR _3988_/X sky130_fd_sc_hd__mux2_1
XFILLER_50_486 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_330 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5727_ _7005_/Q _5912_/A2 _5618_/X _6877_/Q VGND VGND VPWR VPWR _5727_/X sky130_fd_sc_hd__a22o_1
XFILLER_136_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5658_ _6802_/Q _5639_/X _5642_/X _6978_/Q _5641_/Y VGND VGND VPWR VPWR _5658_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_163_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4609_ _4614_/A _4609_/B _4613_/C VGND VGND VPWR VPWR _4701_/A sky130_fd_sc_hd__or3b_4
XFILLER_191_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_190_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5589_ _5609_/B _5981_/A _5977_/A _5565_/X _7098_/Q VGND VGND VPWR VPWR _7098_/D
+ sky130_fd_sc_hd__o32a_1
XFILLER_151_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold340 _5229_/X VGND VGND VPWR VPWR _6804_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_117_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_190_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold351 _6909_/Q VGND VGND VPWR VPWR hold351/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold362 _5364_/X VGND VGND VPWR VPWR _6924_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold373 _6504_/Q VGND VGND VPWR VPWR hold373/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_117_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold384 _5175_/X VGND VGND VPWR VPWR _6759_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold395 hold395/A VGND VGND VPWR VPWR hold395/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_132_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_520 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1040 _6819_/Q VGND VGND VPWR VPWR _5246_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_133_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1051 _5480_/X VGND VGND VPWR VPWR _7027_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1062 _6986_/Q VGND VGND VPWR VPWR _5434_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_58_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1073 _7002_/Q VGND VGND VPWR VPWR _5452_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1084 _5470_/X VGND VGND VPWR VPWR _7018_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_172_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_202 _5918_/A2 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1095 _7022_/Q VGND VGND VPWR VPWR _5474_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_213 _5460_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_464 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_260 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_403 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_190_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4960_ _4959_/C _4960_/B _4960_/C VGND VGND VPWR VPWR _4960_/Y sky130_fd_sc_hd__nand3b_1
X_3911_ _6487_/Q _3910_/Y _3749_/S VGND VGND VPWR VPWR _7157_/D sky130_fd_sc_hd__o21a_2
XFILLER_32_431 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4891_ _4885_/A _4737_/B _4430_/C _4885_/B _4740_/X VGND VGND VPWR VPWR _5073_/A
+ sky130_fd_sc_hd__o41a_1
XFILLER_177_403 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6630_ _6630_/CLK _6630_/D fanout496/X VGND VGND VPWR VPWR _6630_/Q sky130_fd_sc_hd__dfrtp_4
X_3842_ hold56/A _3842_/B VGND VGND VPWR VPWR _3843_/B sky130_fd_sc_hd__nand2_1
XFILLER_177_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6561_ _6630_/CLK _6561_/D _6401_/A VGND VGND VPWR VPWR _6561_/Q sky130_fd_sc_hd__dfrtp_2
X_3773_ _6962_/Q _5406_/A _3374_/Y _6850_/Q VGND VGND VPWR VPWR _3773_/X sky130_fd_sc_hd__a22o_1
XFILLER_192_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_660 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5512_ _5512_/A0 _5530_/A1 _5519_/S VGND VGND VPWR VPWR _5512_/X sky130_fd_sc_hd__mux2_1
XFILLER_145_311 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6492_ _6527_/CLK _6492_/D fanout524/X VGND VGND VPWR VPWR _7183_/A sky130_fd_sc_hd__dfrtp_1
XFILLER_118_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5443_ _5443_/A0 _5488_/A1 _5450_/S VGND VGND VPWR VPWR _5443_/X sky130_fd_sc_hd__mux2_1
XFILLER_172_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5374_ hold709/X _5542_/A1 hold42/X VGND VGND VPWR VPWR _5374_/X sky130_fd_sc_hd__mux2_1
X_7113_ _7123_/CLK _7113_/D fanout502/X VGND VGND VPWR VPWR _7113_/Q sky130_fd_sc_hd__dfrtp_1
X_4325_ hold555/X _5491_/A1 _4326_/S VGND VGND VPWR VPWR _4325_/X sky130_fd_sc_hd__mux2_1
XFILLER_87_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7044_ _7046_/CLK _7044_/D fanout503/X VGND VGND VPWR VPWR _7044_/Q sky130_fd_sc_hd__dfrtp_1
X_4256_ _4256_/A0 _6353_/A1 _4260_/S VGND VGND VPWR VPWR _4256_/X sky130_fd_sc_hd__mux2_1
XFILLER_74_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3207_ _6901_/Q VGND VGND VPWR VPWR _3207_/Y sky130_fd_sc_hd__inv_2
XFILLER_28_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4187_ _3471_/X _4187_/A1 _4189_/S VGND VGND VPWR VPWR _6596_/D sky130_fd_sc_hd__mux2_1
XFILLER_27_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6828_ _7041_/CLK _6828_/D fanout518/X VGND VGND VPWR VPWR _6828_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_10_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6759_ _6976_/CLK _6759_/D fanout497/X VGND VGND VPWR VPWR _6759_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_11_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_163_130 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_164_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold170 _4006_/X VGND VGND VPWR VPWR _6453_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold181 _4116_/X VGND VGND VPWR VPWR _6535_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_105_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold192 _3981_/X VGND VGND VPWR VPWR _6431_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_120_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_263 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_160_52 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_515 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_458 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4110_ hold221/X _5476_/A1 _4111_/S VGND VGND VPWR VPWR _4110_/X sky130_fd_sc_hd__mux2_1
X_5090_ _5090_/A _5090_/B VGND VGND VPWR VPWR _5091_/A sky130_fd_sc_hd__nand2_1
XFILLER_68_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4041_ hold753/X _5505_/A1 _4043_/S VGND VGND VPWR VPWR _4041_/X sky130_fd_sc_hd__mux2_1
XFILLER_64_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5992_ _7026_/Q _6291_/A2 _5980_/Y _7018_/Q _5991_/X VGND VGND VPWR VPWR _5992_/X
+ sky130_fd_sc_hd__a221o_1
X_4943_ _4943_/A _4943_/B _4943_/C VGND VGND VPWR VPWR _5026_/B sky130_fd_sc_hd__and3_4
XFILLER_178_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4874_ _4748_/B _4973_/A _4745_/B _4901_/B VGND VGND VPWR VPWR _4877_/B sky130_fd_sc_hd__o22a_1
XFILLER_177_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_178_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_177_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6613_ _6632_/CLK _6613_/D _3264_/A VGND VGND VPWR VPWR _6613_/Q sky130_fd_sc_hd__dfrtp_1
X_3825_ _6415_/Q _3825_/B VGND VGND VPWR VPWR _3826_/B sky130_fd_sc_hd__and2b_1
XFILLER_165_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6544_ _6630_/CLK _6544_/D fanout495/X VGND VGND VPWR VPWR _6544_/Q sky130_fd_sc_hd__dfstp_2
X_3756_ _6418_/Q _3958_/A _4255_/A _6660_/Q VGND VGND VPWR VPWR _3756_/X sky130_fd_sc_hd__a22o_1
XFILLER_192_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_3_5_0_csclk clkbuf_3_5_0_csclk/A VGND VGND VPWR VPWR clkbuf_3_5_0_csclk/X
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_118_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6475_ _6707_/CLK _6475_/D fanout486/X VGND VGND VPWR VPWR _6475_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_145_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3687_ _6711_/Q _4315_/A _4309_/A _6706_/Q VGND VGND VPWR VPWR _3687_/X sky130_fd_sc_hd__a22o_1
XFILLER_118_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5426_ _5426_/A0 _5495_/A1 _5432_/S VGND VGND VPWR VPWR _5426_/X sky130_fd_sc_hd__mux2_1
XFILLER_145_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_160_122 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput220 _7183_/X VGND VGND VPWR VPWR mgmt_gpio_out[18] sky130_fd_sc_hd__buf_12
Xoutput231 _7193_/X VGND VGND VPWR VPWR mgmt_gpio_out[28] sky130_fd_sc_hd__buf_12
Xoutput242 _7175_/X VGND VGND VPWR VPWR mgmt_gpio_out[3] sky130_fd_sc_hd__buf_12
Xoutput253 _3942_/Y VGND VGND VPWR VPWR pad_flash_io0_oeb sky130_fd_sc_hd__buf_12
Xoutput264 _6739_/Q VGND VGND VPWR VPWR pll_div[2] sky130_fd_sc_hd__buf_12
XFILLER_102_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5357_ _5357_/A0 _5465_/A1 _5360_/S VGND VGND VPWR VPWR _5357_/X sky130_fd_sc_hd__mux2_1
Xoutput275 _6431_/Q VGND VGND VPWR VPWR pll_trim[13] sky130_fd_sc_hd__buf_12
XFILLER_160_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput286 _6425_/Q VGND VGND VPWR VPWR pll_trim[23] sky130_fd_sc_hd__buf_12
Xoutput297 _6751_/Q VGND VGND VPWR VPWR pwr_ctrl_out[0] sky130_fd_sc_hd__buf_12
XFILLER_58_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4308_ hold391/X _5534_/A1 _4308_/S VGND VGND VPWR VPWR _4308_/X sky130_fd_sc_hd__mux2_1
XFILLER_102_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5288_ hold660/X _5537_/A1 _5288_/S VGND VGND VPWR VPWR _5288_/X sky130_fd_sc_hd__mux2_1
XFILLER_141_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7027_ _7027_/CLK _7027_/D fanout499/X VGND VGND VPWR VPWR _7027_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_59_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4239_ hold951/X _6354_/A1 _4242_/S VGND VGND VPWR VPWR _4239_/X sky130_fd_sc_hd__mux2_1
XFILLER_75_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_168_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_183_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire347 _3777_/Y VGND VGND VPWR VPWR wire347/X sky130_fd_sc_hd__clkbuf_1
XFILLER_109_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_137_642 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire358 _4642_/Y VGND VGND VPWR VPWR _5058_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_139_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_183_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_347 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7103__531 VGND VGND VPWR VPWR _7103_/D _7103__531/LO sky130_fd_sc_hd__conb_1
XFILLER_120_553 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout480 _6401_/B VGND VGND VPWR VPWR _6399_/B sky130_fd_sc_hd__buf_4
XFILLER_120_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_171_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout491 fanout492/X VGND VGND VPWR VPWR _6399_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_46_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_44 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_715 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_174_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3610_ _6933_/Q hold41/A _4309_/A _6708_/Q VGND VGND VPWR VPWR _3610_/X sky130_fd_sc_hd__a22o_2
X_4590_ _4590_/A _4632_/B VGND VGND VPWR VPWR _4985_/A sky130_fd_sc_hd__or2_1
X_3541_ _3563_/A hold53/A VGND VGND VPWR VPWR _6352_/A sky130_fd_sc_hd__nor2_8
Xhold906 _5463_/X VGND VGND VPWR VPWR _7012_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold917 _6859_/Q VGND VGND VPWR VPWR hold917/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_128_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold928 _5453_/X VGND VGND VPWR VPWR _7003_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_50_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold939 _6851_/Q VGND VGND VPWR VPWR hold939/X sky130_fd_sc_hd__dlygate4sd3_1
X_6260_ _6688_/Q _5942_/X _5979_/X _6453_/Q _6259_/X VGND VGND VPWR VPWR _6268_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_142_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3472_ _6731_/Q _3471_/X _3685_/S VGND VGND VPWR VPWR _3472_/X sky130_fd_sc_hd__mux2_1
XFILLER_143_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5211_ hold365/X _5532_/A1 _5216_/S VGND VGND VPWR VPWR _5211_/X sky130_fd_sc_hd__mux2_1
X_6191_ _6685_/Q _5942_/X _5972_/B _6690_/Q _6184_/X VGND VGND VPWR VPWR _6201_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_97_710 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5142_ _5142_/A _6352_/B VGND VGND VPWR VPWR _5144_/S sky130_fd_sc_hd__and2_1
XFILLER_123_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_404 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5073_ _5073_/A _5073_/B _5073_/C VGND VGND VPWR VPWR _5136_/C sky130_fd_sc_hd__and3_1
XFILLER_111_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4024_ hold513/X _5491_/A1 _4025_/S VGND VGND VPWR VPWR _4024_/X sky130_fd_sc_hd__mux2_1
XFILLER_49_191 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5975_ _5975_/A _5975_/B _5975_/C _5969_/Y VGND VGND VPWR VPWR _5975_/X sky130_fd_sc_hd__or4b_4
XFILLER_52_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4926_ _4721_/B _5026_/A _4788_/A _4612_/X _4818_/A VGND VGND VPWR VPWR _5108_/B
+ sky130_fd_sc_hd__o311a_1
XFILLER_52_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4857_ _4789_/B _4962_/C _4630_/B _4717_/B _4856_/X VGND VGND VPWR VPWR _4857_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_20_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_166_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3808_ _6858_/Q _5289_/A _4291_/A _6690_/Q _3807_/X VGND VGND VPWR VPWR _3814_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_165_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4788_ _4788_/A _4788_/B VGND VGND VPWR VPWR _4812_/B sky130_fd_sc_hd__or2_1
XFILLER_118_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6527_ _6527_/CLK _6527_/D fanout524/X VGND VGND VPWR VPWR _6527_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_4_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3739_ _6795_/Q _5217_/A _3629_/Y _6766_/Q VGND VGND VPWR VPWR _3739_/X sky130_fd_sc_hd__a22o_1
XFILLER_193_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_180_239 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6458_ _6565_/CLK _6458_/D fanout495/X VGND VGND VPWR VPWR _6458_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_134_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5409_ hold281/X _5541_/A1 _5414_/S VGND VGND VPWR VPWR _5409_/X sky130_fd_sc_hd__mux2_1
XFILLER_133_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6389_ _6399_/A _6399_/B VGND VGND VPWR VPWR _6389_/X sky130_fd_sc_hd__and2_1
XFILLER_102_520 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_264 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_43 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_188_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_188_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_184_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_51 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_404 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_275 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_94_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_651 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5760_ _6847_/Q _5922_/B1 _5651_/X _6799_/Q _5759_/X VGND VGND VPWR VPWR _5760_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_98_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4711_ _4711_/A _4711_/B _4710_/X VGND VGND VPWR VPWR _4711_/X sky130_fd_sc_hd__or3b_1
XTAP_1290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5691_ _5691_/A1 _6305_/A2 _5689_/X _5690_/X VGND VGND VPWR VPWR _7107_/D sky130_fd_sc_hd__o22a_1
XFILLER_187_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4642_ _5026_/A _4788_/A _4924_/B _4634_/B VGND VGND VPWR VPWR _4642_/Y sky130_fd_sc_hd__nor4b_1
XFILLER_147_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_163_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4573_ _4573_/A _4947_/B _4947_/C VGND VGND VPWR VPWR _4574_/B sky130_fd_sc_hd__and3_1
Xmax_cap400 _5648_/X VGND VGND VPWR VPWR _5925_/B1 sky130_fd_sc_hd__buf_12
Xmax_cap411 _5629_/X VGND VGND VPWR VPWR _5929_/B1 sky130_fd_sc_hd__buf_12
Xhold703 _6445_/Q VGND VGND VPWR VPWR hold703/X sky130_fd_sc_hd__dlygate4sd3_1
X_6312_ _3625_/X _6312_/A1 _6316_/S VGND VGND VPWR VPWR _7136_/D sky130_fd_sc_hd__mux2_1
Xhold714 _5542_/X VGND VGND VPWR VPWR _7082_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3524_ _6608_/Q _4196_/A _4145_/A _6564_/Q VGND VGND VPWR VPWR _3524_/X sky130_fd_sc_hd__a22o_1
XFILLER_116_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold725 _6951_/Q VGND VGND VPWR VPWR hold725/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold736 _5356_/X VGND VGND VPWR VPWR _6917_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_171_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold747 _6863_/Q VGND VGND VPWR VPWR hold747/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold758 _5313_/X VGND VGND VPWR VPWR _6879_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6243_ _6627_/Q _5973_/A _5971_/B _6611_/Q _6242_/X VGND VGND VPWR VPWR _6251_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_170_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold769 hold769/A VGND VGND VPWR VPWR hold769/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3455_ _6999_/Q _5442_/A _5289_/A _6863_/Q _3436_/X VGND VGND VPWR VPWR _3460_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_170_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6174_ _7078_/Q _6289_/A2 _5975_/A _6857_/Q VGND VGND VPWR VPWR _6174_/X sky130_fd_sc_hd__a22o_1
X_3386_ _3719_/A _3525_/A VGND VGND VPWR VPWR _5289_/A sky130_fd_sc_hd__nor2_8
XFILLER_85_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5125_ _4828_/A _5025_/Y _5027_/Y _4537_/B _5035_/C VGND VGND VPWR VPWR _5134_/B
+ sky130_fd_sc_hd__o221ai_4
Xhold1403 _6591_/Q VGND VGND VPWR VPWR _4182_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_111_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1414 _7136_/Q VGND VGND VPWR VPWR _6312_/A1 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1425 _6597_/Q VGND VGND VPWR VPWR _4188_/A1 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1436 _6728_/Q VGND VGND VPWR VPWR _3749_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_85_746 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1447 _6639_/Q VGND VGND VPWR VPWR _3873_/B1 sky130_fd_sc_hd__dlygate4sd3_1
X_5056_ _4692_/C _4691_/C _4965_/C _4978_/X VGND VGND VPWR VPWR _5118_/B sky130_fd_sc_hd__o31ai_1
Xhold1458 _6636_/Q VGND VGND VPWR VPWR _6641_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_38_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1469 hold92/A VGND VGND VPWR VPWR _6328_/A1 sky130_fd_sc_hd__dlygate4sd3_1
X_4007_ _4007_/A0 _4236_/A1 _4007_/S VGND VGND VPWR VPWR _4007_/X sky130_fd_sc_hd__mux2_1
XTAP_2908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_0_1_wb_clk_i clkbuf_1_0_1_wb_clk_i/A VGND VGND VPWR VPWR clkbuf_2_1_0_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_80_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5958_ _7099_/Q _7101_/Q _7102_/Q _7100_/Q VGND VGND VPWR VPWR _5965_/B sky130_fd_sc_hd__or4b_4
XFILLER_52_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4909_ _5008_/D _5135_/B _5016_/B VGND VGND VPWR VPWR _4913_/B sky130_fd_sc_hd__and3_1
X_5889_ _5889_/A1 _6305_/A2 _5887_/X _5888_/X VGND VGND VPWR VPWR _7116_/D sky130_fd_sc_hd__o22a_1
XFILLER_139_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_269 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_166_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_2_2_0_csclk clkbuf_2_3_0_csclk/A VGND VGND VPWR VPWR clkbuf_3_5_0_csclk/A
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_106_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_136_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold30 hold30/A VGND VGND VPWR VPWR hold30/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold41 hold41/A VGND VGND VPWR VPWR hold41/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_130_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold52 hold52/A VGND VGND VPWR VPWR hold52/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold63 hold63/A VGND VGND VPWR VPWR hold63/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold74 hold74/A VGND VGND VPWR VPWR hold74/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_152_64 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold85 hold85/A VGND VGND VPWR VPWR hold85/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold96 hold96/A VGND VGND VPWR VPWR hold96/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_91_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_40 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_334 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_188_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_188_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_176_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_145_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_375 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_5 _5208_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_153_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_112_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3240_ _3240_/A _3819_/B VGND VGND VPWR VPWR _3256_/S sky130_fd_sc_hd__or2_4
XFILLER_140_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3171_ _6813_/Q VGND VGND VPWR VPWR _3171_/Y sky130_fd_sc_hd__inv_2
XFILLER_79_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_212 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6930_ _6988_/CLK _6930_/D fanout513/X VGND VGND VPWR VPWR _6930_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_19_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_248 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6861_ _7017_/CLK _6861_/D fanout515/X VGND VGND VPWR VPWR _6861_/Q sky130_fd_sc_hd__dfrtp_4
Xclkbuf_leaf_6_csclk clkbuf_3_1_0_csclk/X VGND VGND VPWR VPWR _6630_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_62_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_179_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5812_ _6977_/Q _5644_/X _5806_/X _5807_/X _5811_/X VGND VGND VPWR VPWR _5812_/X
+ sky130_fd_sc_hd__a2111o_1
X_6792_ _7072_/CLK _6792_/D fanout507/X VGND VGND VPWR VPWR _6792_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_50_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5743_ _6838_/Q _5928_/A2 _5929_/B1 _7022_/Q _5742_/X VGND VGND VPWR VPWR _5743_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_148_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_148_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5674_ _7019_/Q _5629_/X _5631_/X _6859_/Q _5673_/X VGND VGND VPWR VPWR _5674_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_30_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_163_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4625_ input99/X _4409_/B _4707_/C _4888_/A VGND VGND VPWR VPWR _4778_/C sky130_fd_sc_hd__a31o_1
XFILLER_190_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold500 _3988_/X VGND VGND VPWR VPWR _6437_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_163_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold511 _6845_/Q VGND VGND VPWR VPWR hold511/X sky130_fd_sc_hd__dlygate4sd3_1
X_4556_ _4556_/A _4962_/C VGND VGND VPWR VPWR _4942_/B sky130_fd_sc_hd__or2_1
Xhold522 _4004_/X VGND VGND VPWR VPWR _6451_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold533 _6985_/Q VGND VGND VPWR VPWR hold533/X sky130_fd_sc_hd__dlygate4sd3_1
X_3507_ _3553_/A _3628_/B VGND VGND VPWR VPWR _4273_/A sky130_fd_sc_hd__nor2_8
Xhold544 _4171_/X VGND VGND VPWR VPWR _6582_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold555 _6718_/Q VGND VGND VPWR VPWR hold555/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_190_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold566 _4010_/X VGND VGND VPWR VPWR _6456_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4487_ _4490_/B _4561_/B VGND VGND VPWR VPWR _4588_/B sky130_fd_sc_hd__or2_4
Xhold577 _6471_/Q VGND VGND VPWR VPWR hold577/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold588 _3959_/X VGND VGND VPWR VPWR hold588/X sky130_fd_sc_hd__dlygate4sd3_1
X_6226_ _6610_/Q _5971_/B _6223_/X _6225_/X VGND VGND VPWR VPWR _6227_/C sky130_fd_sc_hd__a211o_1
Xhold599 _4289_/X VGND VGND VPWR VPWR _6688_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3438_ _5183_/A _3628_/B VGND VGND VPWR VPWR _5151_/A sky130_fd_sc_hd__nor2_8
XFILLER_131_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6157_ _7025_/Q _6290_/B1 _5981_/X _6937_/Q _6156_/X VGND VGND VPWR VPWR _6157_/X
+ sky130_fd_sc_hd__a221o_1
XTAP_871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1200 _5353_/X VGND VGND VPWR VPWR _6914_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3369_ _6441_/Q _3984_/A _5325_/A _6897_/Q _3365_/X VGND VGND VPWR VPWR _3369_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_112_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1211 _6426_/Q VGND VGND VPWR VPWR _3976_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1222 _4286_/X VGND VGND VPWR VPWR _6685_/D sky130_fd_sc_hd__dlygate4sd3_1
X_5108_ _5108_/A _5108_/B _5108_/C VGND VGND VPWR VPWR _5108_/Y sky130_fd_sc_hd__nand3_1
Xhold1233 _6670_/Q VGND VGND VPWR VPWR _4268_/A0 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1244 _5512_/X VGND VGND VPWR VPWR _7055_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6088_ _6990_/Q _6286_/B1 _5971_/A _6870_/Q VGND VGND VPWR VPWR _6088_/X sky130_fd_sc_hd__a22o_1
Xhold1255 _7151_/Q VGND VGND VPWR VPWR _6353_/A0 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1266 _5344_/X VGND VGND VPWR VPWR _6906_/D sky130_fd_sc_hd__dlygate4sd3_1
X_5039_ _5038_/X _5087_/C _5087_/B _5087_/A VGND VGND VPWR VPWR _5039_/X sky130_fd_sc_hd__and4b_1
XTAP_2705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1277 _6830_/Q VGND VGND VPWR VPWR _5258_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_73_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1288 _5222_/X VGND VGND VPWR VPWR _6798_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1299 _6522_/Q VGND VGND VPWR VPWR _4101_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_21 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_193_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_162_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_163_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput120 wb_adr_i[29] VGND VGND VPWR VPWR _3895_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_88_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput131 wb_cyc_i VGND VGND VPWR VPWR _3894_/C sky130_fd_sc_hd__clkbuf_1
Xinput142 wb_dat_i[19] VGND VGND VPWR VPWR _6333_/A2 sky130_fd_sc_hd__clkbuf_1
XFILLER_76_543 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput153 wb_dat_i[29] VGND VGND VPWR VPWR _6338_/A2 sky130_fd_sc_hd__clkbuf_1
Xinput164 wb_rstn_i VGND VGND VPWR VPWR input164/X sky130_fd_sc_hd__clkbuf_4
XFILLER_29_481 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_546 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4410_ _4513_/A _4943_/A VGND VGND VPWR VPWR _4410_/X sky130_fd_sc_hd__or2_1
XFILLER_145_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5390_ _5390_/A0 _5495_/A1 _5396_/S VGND VGND VPWR VPWR _5390_/X sky130_fd_sc_hd__mux2_1
XFILLER_172_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_132_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4341_ _4613_/C _4614_/A VGND VGND VPWR VPWR _4592_/A sky130_fd_sc_hd__and2_2
XFILLER_125_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_423 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_592 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_294 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7060_ _7060_/CLK _7060_/D fanout521/X VGND VGND VPWR VPWR _7060_/Q sky130_fd_sc_hd__dfrtp_1
X_4272_ hold551/X _6357_/A1 _4272_/S VGND VGND VPWR VPWR _4272_/X sky130_fd_sc_hd__mux2_1
XFILLER_86_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_141_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6011_ _6963_/Q _5955_/X _5975_/C _7048_/Q VGND VGND VPWR VPWR _6011_/X sky130_fd_sc_hd__a22o_1
X_3223_ _6920_/Q VGND VGND VPWR VPWR _3223_/Y sky130_fd_sc_hd__inv_2
XFILLER_140_286 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_532 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6913_ _6969_/CLK _6913_/D fanout506/X VGND VGND VPWR VPWR _6913_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_35_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6844_ _7041_/CLK _6844_/D fanout520/X VGND VGND VPWR VPWR _6844_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_50_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3987_ hold795/X _6355_/A1 _3992_/S VGND VGND VPWR VPWR _3987_/X sky130_fd_sc_hd__mux2_1
X_6775_ _6881_/CLK _6775_/D fanout523/X VGND VGND VPWR VPWR _7194_/A sky130_fd_sc_hd__dfrtp_1
XFILLER_167_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_498 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5726_ _6901_/Q _5623_/X _5637_/X _6853_/Q _5725_/X VGND VGND VPWR VPWR _5726_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_148_342 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_176_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5657_ _6954_/Q _5630_/X _5653_/X _5654_/X _5656_/X VGND VGND VPWR VPWR _5657_/X
+ sky130_fd_sc_hd__a2111o_1
XFILLER_163_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4608_ _4973_/A _4972_/A _4748_/B VGND VGND VPWR VPWR _4662_/A sky130_fd_sc_hd__a21o_1
XFILLER_163_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5588_ _7098_/Q _7097_/Q VGND VGND VPWR VPWR _5980_/A sky130_fd_sc_hd__nand2b_4
XFILLER_151_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold330 _5301_/X VGND VGND VPWR VPWR _6868_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold341 _6692_/Q VGND VGND VPWR VPWR hold341/X sky130_fd_sc_hd__dlygate4sd3_1
X_4539_ _4575_/A _4629_/B VGND VGND VPWR VPWR _4649_/A sky130_fd_sc_hd__or2_4
Xhold352 _5347_/X VGND VGND VPWR VPWR _6909_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_190_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold363 _6534_/Q VGND VGND VPWR VPWR hold363/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold374 _4076_/X VGND VGND VPWR VPWR _6504_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold385 _6649_/Q VGND VGND VPWR VPWR hold385/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_117_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_132_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold396 _5205_/X VGND VGND VPWR VPWR _6783_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6209_ _6600_/Q _5939_/X _5977_/X _6666_/Q VGND VGND VPWR VPWR _6209_/X sky130_fd_sc_hd__a22o_1
XFILLER_104_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_131_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7189_ _7189_/A VGND VGND VPWR VPWR _7189_/X sky130_fd_sc_hd__clkbuf_2
XTAP_690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1030 _6752_/Q VGND VGND VPWR VPWR _5165_/A0 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1041 _5246_/X VGND VGND VPWR VPWR _6819_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_46_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1052 _6954_/Q VGND VGND VPWR VPWR _5398_/A0 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1063 _5434_/X VGND VGND VPWR VPWR _6986_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1074 _5452_/X VGND VGND VPWR VPWR _7002_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1085 _6850_/Q VGND VGND VPWR VPWR _5281_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_203 _5912_/A2 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1096 _5474_/X VGND VGND VPWR VPWR _7022_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_214 _3384_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3221__1 net499_2/A VGND VGND VPWR VPWR _7157_/CLK sky130_fd_sc_hd__inv_2
XTAP_2546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_165_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_166_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_71_csclk clkbuf_3_1_0_csclk/X VGND VGND VPWR VPWR _6696_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_190_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3910_ _6486_/Q _6489_/Q VGND VGND VPWR VPWR _3910_/Y sky130_fd_sc_hd__nor2_1
XFILLER_32_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4890_ _4549_/B _4495_/X _4597_/Y _4901_/B _4889_/X VGND VGND VPWR VPWR _5135_/B
+ sky130_fd_sc_hd__o221a_1
XFILLER_32_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3841_ _3857_/S _3841_/B hold29/A VGND VGND VPWR VPWR _3843_/A sky130_fd_sc_hd__or3b_1
XFILLER_80_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3772_ _6978_/Q _5424_/A _5145_/A _6737_/Q _3771_/X VGND VGND VPWR VPWR _3777_/B
+ sky130_fd_sc_hd__a221o_1
X_6560_ _6630_/CLK _6560_/D fanout495/X VGND VGND VPWR VPWR _6560_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_158_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5511_ _5511_/A _5511_/B VGND VGND VPWR VPWR _5519_/S sky130_fd_sc_hd__and2_4
X_6491_ _6527_/CLK _6491_/D fanout524/X VGND VGND VPWR VPWR _7182_/A sky130_fd_sc_hd__dfrtp_1
XFILLER_145_323 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5442_ _5442_/A _5529_/B VGND VGND VPWR VPWR _5450_/S sky130_fd_sc_hd__and2_4
XFILLER_173_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5373_ hold433/X _5541_/A1 hold42/X VGND VGND VPWR VPWR _5373_/X sky130_fd_sc_hd__mux2_1
XFILLER_172_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_24_csclk clkbuf_3_6_0_csclk/X VGND VGND VPWR VPWR _6965_/CLK sky130_fd_sc_hd__clkbuf_16
X_7112_ _7124_/CLK _7112_/D fanout502/X VGND VGND VPWR VPWR _7112_/Q sky130_fd_sc_hd__dfrtp_1
X_4324_ hold616/X _5505_/A1 _4326_/S VGND VGND VPWR VPWR _4324_/X sky130_fd_sc_hd__mux2_1
XFILLER_114_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7043_ _7043_/CLK _7043_/D fanout513/X VGND VGND VPWR VPWR _7043_/Q sky130_fd_sc_hd__dfrtp_2
X_4255_ _4255_/A _6352_/B VGND VGND VPWR VPWR _4260_/S sky130_fd_sc_hd__and2_4
XFILLER_86_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3206_ _6909_/Q VGND VGND VPWR VPWR _3206_/Y sky130_fd_sc_hd__inv_2
X_4186_ _4186_/A0 _4186_/A1 _4189_/S VGND VGND VPWR VPWR _6595_/D sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_39_csclk clkbuf_3_7_0_csclk/X VGND VGND VPWR VPWR _6961_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_55_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_3_1_0_csclk clkbuf_3_1_0_csclk/A VGND VGND VPWR VPWR clkbuf_3_1_0_csclk/X
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_103_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_546 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6827_ _7046_/CLK _6827_/D fanout500/X VGND VGND VPWR VPWR _6827_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_50_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6758_ _6976_/CLK _6758_/D fanout501/X VGND VGND VPWR VPWR _6758_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_149_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_11 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5709_ _6444_/Q _5917_/B1 _5692_/X _5708_/X VGND VGND VPWR VPWR _5709_/X sky130_fd_sc_hd__a211o_1
XFILLER_176_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6689_ _6689_/CLK _6689_/D fanout510/X VGND VGND VPWR VPWR _6689_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_164_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_163_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_151_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_163_175 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold160 _5358_/X VGND VGND VPWR VPWR _6919_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_105_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold171 _6693_/Q VGND VGND VPWR VPWR hold171/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold182 _6955_/Q VGND VGND VPWR VPWR hold182/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_78_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold193 _6813_/Q VGND VGND VPWR VPWR hold193/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_120_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_262 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_169_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_139_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_186_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_170_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_108_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4040_ _4040_/A0 _5189_/A1 _4043_/S VGND VGND VPWR VPWR _4040_/X sky130_fd_sc_hd__mux2_1
XFILLER_77_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_267 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5991_ _6794_/Q _5948_/X _5963_/X _6826_/Q VGND VGND VPWR VPWR _5991_/X sky130_fd_sc_hd__a22o_1
X_4942_ _4531_/X _4942_/B _4942_/C VGND VGND VPWR VPWR _5087_/C sky130_fd_sc_hd__and3b_1
XFILLER_17_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_178_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4873_ _4973_/A _4972_/A _4745_/B _4872_/X _4855_/X VGND VGND VPWR VPWR _4877_/A
+ sky130_fd_sc_hd__a41o_1
XFILLER_178_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6612_ _7155_/CLK hold47/X _6370_/A VGND VGND VPWR VPWR _6612_/Q sky130_fd_sc_hd__dfrtp_4
X_3824_ _3824_/A _3824_/B VGND VGND VPWR VPWR _6416_/D sky130_fd_sc_hd__nor2_1
XFILLER_193_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6543_ _6697_/CLK _6543_/D fanout485/X VGND VGND VPWR VPWR _6543_/Q sky130_fd_sc_hd__dfstp_2
X_3755_ _6550_/Q _4133_/A _5187_/A _6768_/Q VGND VGND VPWR VPWR _3755_/X sky130_fd_sc_hd__a22o_1
XFILLER_118_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3686_ _3685_/X _3686_/A1 _3749_/S VGND VGND VPWR VPWR _6729_/D sky130_fd_sc_hd__mux2_1
X_6474_ _6699_/CLK _6474_/D fanout509/X VGND VGND VPWR VPWR _6474_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_118_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_146_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5425_ _5425_/A0 _5488_/A1 _5432_/S VGND VGND VPWR VPWR _5425_/X sky130_fd_sc_hd__mux2_1
Xoutput210 _3214_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[7] sky130_fd_sc_hd__buf_12
XFILLER_161_635 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput221 _7184_/X VGND VGND VPWR VPWR mgmt_gpio_out[19] sky130_fd_sc_hd__buf_12
XFILLER_133_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput232 _7194_/X VGND VGND VPWR VPWR mgmt_gpio_out[29] sky130_fd_sc_hd__buf_12
Xoutput243 _7176_/X VGND VGND VPWR VPWR mgmt_gpio_out[4] sky130_fd_sc_hd__buf_12
Xoutput254 _7198_/X VGND VGND VPWR VPWR pad_flash_io1_do sky130_fd_sc_hd__buf_12
X_5356_ hold735/X _5542_/A1 _5360_/S VGND VGND VPWR VPWR _5356_/X sky130_fd_sc_hd__mux2_1
Xoutput265 _6740_/Q VGND VGND VPWR VPWR pll_div[3] sky130_fd_sc_hd__buf_12
Xoutput276 _6432_/Q VGND VGND VPWR VPWR pll_trim[14] sky130_fd_sc_hd__buf_12
XFILLER_58_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput287 _6748_/Q VGND VGND VPWR VPWR pll_trim[24] sky130_fd_sc_hd__buf_12
X_4307_ hold495/X _5491_/A1 _4308_/S VGND VGND VPWR VPWR _4307_/X sky130_fd_sc_hd__mux2_1
Xoutput298 _6752_/Q VGND VGND VPWR VPWR pwr_ctrl_out[1] sky130_fd_sc_hd__buf_12
X_5287_ hold132/X _5476_/A1 _5288_/S VGND VGND VPWR VPWR _5287_/X sky130_fd_sc_hd__mux2_1
XFILLER_87_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7026_ _7027_/CLK _7026_/D fanout499/X VGND VGND VPWR VPWR _7026_/Q sky130_fd_sc_hd__dfstp_1
X_4238_ _4238_/A0 _6353_/A1 _4242_/S VGND VGND VPWR VPWR _4238_/X sky130_fd_sc_hd__mux2_1
XFILLER_74_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4169_ hold835/X _5505_/A1 _4171_/S VGND VGND VPWR VPWR _4169_/X sky130_fd_sc_hd__mux2_1
XFILLER_83_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_652 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_708 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_183_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_139_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire348 _3666_/Y VGND VGND VPWR VPWR wire348/X sky130_fd_sc_hd__clkbuf_2
XFILLER_128_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_654 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_602 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_191_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_152_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_93_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout470 hold6/X VGND VGND VPWR VPWR _5529_/B sky130_fd_sc_hd__buf_8
XFILLER_48_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout481 _6396_/B VGND VGND VPWR VPWR _6401_/B sky130_fd_sc_hd__buf_4
XFILLER_93_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout492 fanout496/X VGND VGND VPWR VPWR fanout492/X sky130_fd_sc_hd__buf_8
XFILLER_93_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_175_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_187_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3540_ _6974_/Q _5415_/A _5487_/A _7038_/Q _3539_/X VGND VGND VPWR VPWR _3548_/A
+ sky130_fd_sc_hd__a221o_1
Xhold907 _6613_/Q VGND VGND VPWR VPWR hold907/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold918 _5291_/X VGND VGND VPWR VPWR _6859_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_127_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold929 _6738_/Q VGND VGND VPWR VPWR hold929/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_115_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3471_ _3471_/A _3471_/B _3471_/C _3470_/Y VGND VGND VPWR VPWR _3471_/X sky130_fd_sc_hd__or4b_4
XFILLER_170_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5210_ _5210_/A0 _5495_/A1 _5216_/S VGND VGND VPWR VPWR _5210_/X sky130_fd_sc_hd__mux2_1
XFILLER_170_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6190_ _6455_/Q _6291_/A2 _6182_/X _6187_/X _6189_/X VGND VGND VPWR VPWR _6202_/B
+ sky130_fd_sc_hd__a2111o_1
XFILLER_97_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5141_ _5112_/X _5131_/X _5139_/X _5140_/X VGND VGND VPWR VPWR _6726_/D sky130_fd_sc_hd__a211o_1
XFILLER_130_329 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_435 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5072_ _4676_/B _4683_/B _4506_/A _4506_/B VGND VGND VPWR VPWR _5073_/C sky130_fd_sc_hd__o211a_1
XFILLER_84_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4023_ hold777/X _6355_/A1 _4025_/S VGND VGND VPWR VPWR _4023_/X sky130_fd_sc_hd__mux2_1
XFILLER_65_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5974_ _5981_/B _5974_/B _5974_/C _5973_/Y VGND VGND VPWR VPWR _5975_/B sky130_fd_sc_hd__or4b_1
X_4925_ _4701_/A _4861_/B _4816_/A _4585_/X VGND VGND VPWR VPWR _5064_/B sky130_fd_sc_hd__o211a_1
XFILLER_80_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4856_ _4620_/B _4715_/B _4855_/X _4597_/Y VGND VGND VPWR VPWR _4856_/X sky130_fd_sc_hd__o22a_1
XFILLER_166_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_178_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3807_ _6465_/Q _4020_/A _5163_/A _6751_/Q VGND VGND VPWR VPWR _3807_/X sky130_fd_sc_hd__a22o_1
XFILLER_119_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4787_ _5043_/B _4615_/B _4786_/Y _4921_/A VGND VGND VPWR VPWR _4788_/B sky130_fd_sc_hd__o22a_1
XFILLER_118_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6526_ _6887_/CLK _6526_/D fanout524/X VGND VGND VPWR VPWR _6526_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_193_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3738_ _6899_/Q _5334_/A _5520_/A _7064_/Q _3737_/X VGND VGND VPWR VPWR _3745_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_146_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_146_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6457_ _7038_/CLK _6457_/D fanout490/X VGND VGND VPWR VPWR _6457_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_161_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3669_ input45/X _3343_/Y _4112_/B _3247_/A _3668_/X VGND VGND VPWR VPWR _3674_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_118_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5408_ hold889/X _5531_/A1 _5414_/S VGND VGND VPWR VPWR _5408_/X sky130_fd_sc_hd__mux2_1
XFILLER_192_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6388_ _6399_/A _6399_/B VGND VGND VPWR VPWR _6388_/X sky130_fd_sc_hd__and2_1
XFILLER_121_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5339_ _5339_/A0 hold23/X _5342_/S VGND VGND VPWR VPWR hold24/A sky130_fd_sc_hd__mux2_1
XFILLER_0_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_565 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7009_ _7033_/CLK _7009_/D fanout506/X VGND VGND VPWR VPWR _7009_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_75_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_655 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_156_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_96 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_432 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_180_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_112_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4710_ _5043_/A _4965_/A _4701_/A _4678_/A VGND VGND VPWR VPWR _4710_/X sky130_fd_sc_hd__a211o_1
XTAP_1291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5690_ _5690_/A1 _5612_/A _5612_/B VGND VGND VPWR VPWR _5690_/X sky130_fd_sc_hd__o21a_1
XFILLER_148_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_187_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4641_ _4596_/B _4575_/B _4615_/B _4640_/X VGND VGND VPWR VPWR _4641_/X sky130_fd_sc_hd__o31a_1
XFILLER_147_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4572_ _4573_/A _4947_/B VGND VGND VPWR VPWR _5021_/B sky130_fd_sc_hd__nand2_2
XFILLER_162_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmax_cap401 _5647_/X VGND VGND VPWR VPWR _5912_/B1 sky130_fd_sc_hd__buf_12
Xmax_cap412 _5628_/X VGND VGND VPWR VPWR _5922_/A2 sky130_fd_sc_hd__buf_12
X_6311_ _3684_/X _6311_/A1 _6316_/S VGND VGND VPWR VPWR _7135_/D sky130_fd_sc_hd__mux2_1
Xhold704 _3997_/X VGND VGND VPWR VPWR _6445_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3523_ _3523_/A _3538_/B VGND VGND VPWR VPWR _4145_/A sky130_fd_sc_hd__nor2_4
Xhold715 _6973_/Q VGND VGND VPWR VPWR hold715/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_155_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold726 _5394_/X VGND VGND VPWR VPWR _6951_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold737 _6855_/Q VGND VGND VPWR VPWR hold737/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_668 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold748 _5295_/X VGND VGND VPWR VPWR _6863_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3454_ _3454_/A _3454_/B VGND VGND VPWR VPWR _3461_/C sky130_fd_sc_hd__or2_2
X_6242_ _6580_/Q _5946_/X _5959_/Y _6616_/Q VGND VGND VPWR VPWR _6242_/X sky130_fd_sc_hd__a22o_1
Xhold759 _7192_/A VGND VGND VPWR VPWR hold759/X sky130_fd_sc_hd__dlygate4sd3_1
X_6173_ _6449_/Q _5601_/Y _6285_/B1 _7017_/Q VGND VGND VPWR VPWR _6173_/X sky130_fd_sc_hd__a22o_1
X_3385_ _6953_/Q _5388_/A _3384_/Y input28/X VGND VGND VPWR VPWR _3385_/X sky130_fd_sc_hd__a22o_1
XFILLER_97_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5124_ _5124_/A _5124_/B _5123_/X VGND VGND VPWR VPWR _5126_/A sky130_fd_sc_hd__or3b_1
XFILLER_57_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1404 _6586_/Q VGND VGND VPWR VPWR _4176_/A1 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1415 _6583_/Q VGND VGND VPWR VPWR _4173_/A1 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1426 _6588_/Q VGND VGND VPWR VPWR _4178_/A1 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1437 _3749_/X VGND VGND VPWR VPWR _6728_/D sky130_fd_sc_hd__dlygate4sd3_1
X_5055_ _5085_/B _5118_/A _5055_/C _5055_/D VGND VGND VPWR VPWR _5055_/X sky130_fd_sc_hd__and4bb_1
XFILLER_57_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1448 _6577_/Q VGND VGND VPWR VPWR _4165_/A1 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1459 _6573_/Q VGND VGND VPWR VPWR _4161_/A1 sky130_fd_sc_hd__dlygate4sd3_1
X_4006_ hold169/X hold46/X _4007_/S VGND VGND VPWR VPWR _4006_/X sky130_fd_sc_hd__mux2_1
XFILLER_65_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_290 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5957_ _5979_/A _5977_/A _5981_/B VGND VGND VPWR VPWR _5957_/X sky130_fd_sc_hd__and3_4
XFILLER_71_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4908_ _4703_/A _4676_/B _4886_/Y _4737_/B _4506_/C VGND VGND VPWR VPWR _5016_/B
+ sky130_fd_sc_hd__o221a_1
XFILLER_21_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5888_ _7115_/Q _5612_/A _5612_/B VGND VGND VPWR VPWR _5888_/X sky130_fd_sc_hd__o21a_1
XFILLER_21_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4839_ _4574_/B _4839_/B _4839_/C _4839_/D VGND VGND VPWR VPWR _4839_/X sky130_fd_sc_hd__and4b_1
XFILLER_166_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_181_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_193_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6509_ _7131_/CLK _6509_/D fanout502/X VGND VGND VPWR VPWR _6509_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_134_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_134_498 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold20 hold20/A VGND VGND VPWR VPWR hold20/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_48_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold31 hold31/A VGND VGND VPWR VPWR hold31/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_152_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold42 hold42/A VGND VGND VPWR VPWR hold42/X sky130_fd_sc_hd__buf_6
Xhold53 hold53/A VGND VGND VPWR VPWR hold53/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_130_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold64 hold64/A VGND VGND VPWR VPWR hold64/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_102_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold75 hold75/A VGND VGND VPWR VPWR hold75/X sky130_fd_sc_hd__clkbuf_16
Xhold86 hold86/A VGND VGND VPWR VPWR hold86/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold97 hold97/A VGND VGND VPWR VPWR hold97/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_75_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_6 _5208_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_137_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3170_ _6487_/Q VGND VGND VPWR VPWR _3240_/A sky130_fd_sc_hd__inv_2
XFILLER_66_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6860_ _6988_/CLK _6860_/D fanout518/X VGND VGND VPWR VPWR _6860_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_179_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5811_ _6825_/Q _5927_/A2 _5808_/X _5810_/X VGND VGND VPWR VPWR _5811_/X sky130_fd_sc_hd__a211o_1
XFILLER_50_614 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6791_ _7086_/CLK _6791_/D fanout516/X VGND VGND VPWR VPWR _6791_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_179_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5742_ _6878_/Q _5618_/X _5924_/B2 _6950_/Q VGND VGND VPWR VPWR _5742_/X sky130_fd_sc_hd__a22o_1
X_5673_ _6795_/Q _5926_/B1 _5671_/X _5672_/X VGND VGND VPWR VPWR _5673_/X sky130_fd_sc_hd__a211o_1
XFILLER_148_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4624_ _4617_/B _4634_/A _4390_/A input99/X VGND VGND VPWR VPWR _4778_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_163_527 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold501 _6521_/Q VGND VGND VPWR VPWR hold501/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4555_ _4596_/B _4555_/B VGND VGND VPWR VPWR _4962_/C sky130_fd_sc_hd__nand2_8
Xhold512 _5275_/X VGND VGND VPWR VPWR _6845_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold523 _6861_/Q VGND VGND VPWR VPWR hold523/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold534 _5432_/X VGND VGND VPWR VPWR _6985_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold545 _6801_/Q VGND VGND VPWR VPWR hold545/X sky130_fd_sc_hd__dlygate4sd3_1
X_3506_ _6454_/Q _4002_/A _4190_/A _6603_/Q _3505_/X VGND VGND VPWR VPWR _3518_/A
+ sky130_fd_sc_hd__a221o_1
Xhold556 _4325_/X VGND VGND VPWR VPWR _6718_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_171_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4486_ _4490_/B _4561_/B VGND VGND VPWR VPWR _4489_/B sky130_fd_sc_hd__nor2_2
Xhold567 _6696_/Q VGND VGND VPWR VPWR hold567/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold578 _4028_/X VGND VGND VPWR VPWR _6471_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6225_ _6671_/Q _5951_/X _6285_/A2 _6631_/Q _6224_/X VGND VGND VPWR VPWR _6225_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_89_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_435 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold589 _5200_/X VGND VGND VPWR VPWR _6778_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3437_ hold39/X _3440_/B hold51/X VGND VGND VPWR VPWR _3628_/B sky130_fd_sc_hd__or3b_4
XTAP_850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3368_ _3706_/A _3525_/A VGND VGND VPWR VPWR _5325_/A sky130_fd_sc_hd__nor2_8
X_6156_ _6953_/Q _5978_/X _6282_/B1 _6977_/Q VGND VGND VPWR VPWR _6156_/X sky130_fd_sc_hd__a22o_1
XTAP_861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1201 _6942_/Q VGND VGND VPWR VPWR _5384_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1212 _3976_/X VGND VGND VPWR VPWR _6426_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_112_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1223 _6540_/Q VGND VGND VPWR VPWR _4122_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_97_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5107_ _4988_/A _4588_/B _4594_/X _4721_/B VGND VGND VPWR VPWR _5108_/C sky130_fd_sc_hd__o22a_1
Xhold1234 _4268_/X VGND VGND VPWR VPWR _6670_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3299_ hold74/X _3366_/A VGND VGND VPWR VPWR hold75/A sky130_fd_sc_hd__or2_4
XFILLER_111_192 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6087_ _6918_/Q _5937_/X _5969_/A _6822_/Q _6086_/X VGND VGND VPWR VPWR _6093_/C
+ sky130_fd_sc_hd__a221o_1
Xhold1245 _6814_/Q VGND VGND VPWR VPWR _5240_/A0 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1256 _6353_/X VGND VGND VPWR VPWR _7151_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1267 _6578_/Q VGND VGND VPWR VPWR _4167_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_57_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5038_ _5038_/A _5038_/B _5038_/C VGND VGND VPWR VPWR _5038_/X sky130_fd_sc_hd__and3_1
Xhold1278 _5258_/X VGND VGND VPWR VPWR _6830_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_26_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1289 _6806_/Q VGND VGND VPWR VPWR _5231_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_33 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6989_ _7082_/CLK _6989_/D fanout520/X VGND VGND VPWR VPWR _6989_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_40_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput110 wb_adr_i[1] VGND VGND VPWR VPWR _4679_/A sky130_fd_sc_hd__buf_6
Xinput121 wb_adr_i[2] VGND VGND VPWR VPWR _4596_/B sky130_fd_sc_hd__buf_8
Xinput132 wb_dat_i[0] VGND VGND VPWR VPWR _6324_/B1 sky130_fd_sc_hd__clkbuf_1
XFILLER_76_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput143 wb_dat_i[1] VGND VGND VPWR VPWR _6327_/B1 sky130_fd_sc_hd__clkbuf_1
Xinput154 wb_dat_i[2] VGND VGND VPWR VPWR _6329_/B1 sky130_fd_sc_hd__clkbuf_1
XFILLER_76_555 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput165 wb_sel_i[0] VGND VGND VPWR VPWR _6317_/A2 sky130_fd_sc_hd__clkbuf_1
XFILLER_64_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_279 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_430 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_176_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4340_ _4679_/A _4542_/A _4554_/A _4596_/B VGND VGND VPWR VPWR _4356_/B sky130_fd_sc_hd__o211a_1
X_4271_ hold626/X _4289_/A1 _4272_/S VGND VGND VPWR VPWR _4271_/X sky130_fd_sc_hd__mux2_1
XFILLER_113_435 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3222_ _6919_/Q VGND VGND VPWR VPWR _3222_/Y sky130_fd_sc_hd__inv_2
X_6010_ _6955_/Q _5957_/X _5978_/X _6947_/Q VGND VGND VPWR VPWR _6010_/X sky130_fd_sc_hd__a22o_1
XFILLER_79_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_544 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_352 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6912_ _6945_/CLK _6912_/D fanout506/X VGND VGND VPWR VPWR _6912_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_50_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6843_ _6945_/CLK _6843_/D fanout506/X VGND VGND VPWR VPWR _6843_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_35_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6774_ _7042_/CLK hold70/X fanout523/X VGND VGND VPWR VPWR _7193_/A sky130_fd_sc_hd__dfrtp_1
X_3986_ _3986_/A0 _6354_/A1 _3992_/S VGND VGND VPWR VPWR _3986_/X sky130_fd_sc_hd__mux2_1
XFILLER_50_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5725_ _6869_/Q _5625_/X _5643_/X _6885_/Q VGND VGND VPWR VPWR _5725_/X sky130_fd_sc_hd__a22o_1
XFILLER_148_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_148_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5656_ _6906_/Q _5922_/A2 _5926_/B1 _6794_/Q _5655_/X VGND VGND VPWR VPWR _5656_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_176_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_190_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4607_ _4678_/A _4717_/A VGND VGND VPWR VPWR _4972_/A sky130_fd_sc_hd__or2_4
X_5587_ _7098_/Q _7097_/Q VGND VGND VPWR VPWR _5977_/A sky130_fd_sc_hd__and2b_2
Xhold320 _4234_/X VGND VGND VPWR VPWR _6632_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold331 _6796_/Q VGND VGND VPWR VPWR hold331/X sky130_fd_sc_hd__dlygate4sd3_1
X_4538_ _4575_/A _4629_/B VGND VGND VPWR VPWR _4623_/B sky130_fd_sc_hd__nor2_1
Xhold342 _4294_/X VGND VGND VPWR VPWR _6692_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_144_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold353 _6821_/Q VGND VGND VPWR VPWR hold353/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold364 _4115_/X VGND VGND VPWR VPWR _6534_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_117_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold375 _6836_/Q VGND VGND VPWR VPWR hold375/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_171_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold386 _4242_/X VGND VGND VPWR VPWR _6649_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4469_ _4554_/A _4596_/B _4448_/A VGND VGND VPWR VPWR _4469_/X sky130_fd_sc_hd__or3b_2
Xhold397 _6753_/Q VGND VGND VPWR VPWR hold397/X sky130_fd_sc_hd__dlygate4sd3_1
X_6208_ _6471_/Q _5941_/Y _5980_/Y _6466_/Q _6207_/X VGND VGND VPWR VPWR _6218_/A
+ sky130_fd_sc_hd__a221o_1
X_7188_ _7188_/A VGND VGND VPWR VPWR _7188_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_58_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6139_ _7077_/Q _6289_/A2 _5978_/X _6952_/Q _6138_/X VGND VGND VPWR VPWR _6142_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_133_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1020 _6979_/Q VGND VGND VPWR VPWR _5426_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1031 _5165_/X VGND VGND VPWR VPWR _6752_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_133_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1042 _6931_/Q VGND VGND VPWR VPWR _5372_/A0 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1053 _5398_/X VGND VGND VPWR VPWR _6954_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1064 _6930_/Q VGND VGND VPWR VPWR _5371_/A0 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1075 _6630_/Q VGND VGND VPWR VPWR _4232_/A0 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1086 _5281_/X VGND VGND VPWR VPWR _6850_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_204 _5534_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1097 _6838_/Q VGND VGND VPWR VPWR _5267_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_430 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_215 _3454_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_181_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_174_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_5_csclk clkbuf_3_1_0_csclk/X VGND VGND VPWR VPWR _6698_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_122_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_319 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_544 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3840_ _3856_/S _3845_/S VGND VGND VPWR VPWR _3841_/B sky130_fd_sc_hd__nor2_1
XFILLER_60_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3771_ _6604_/Q _4196_/A _4032_/A _6475_/Q VGND VGND VPWR VPWR _3771_/X sky130_fd_sc_hd__a22o_1
XFILLER_9_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5510_ hold441/X _5519_/A1 _5510_/S VGND VGND VPWR VPWR _5510_/X sky130_fd_sc_hd__mux2_1
XFILLER_9_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6490_ _7058_/CLK _6490_/D fanout524/X VGND VGND VPWR VPWR _7181_/A sky130_fd_sc_hd__dfrtp_1
XFILLER_145_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5441_ _5441_/A0 hold27/X hold35/X VGND VGND VPWR VPWR hold36/A sky130_fd_sc_hd__mux2_1
XFILLER_160_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5372_ _5372_/A0 _5495_/A1 hold42/X VGND VGND VPWR VPWR _5372_/X sky130_fd_sc_hd__mux2_1
X_7111_ _7131_/CLK _7111_/D fanout501/X VGND VGND VPWR VPWR _7111_/Q sky130_fd_sc_hd__dfrtp_1
X_4323_ hold899/X _5189_/A1 _4326_/S VGND VGND VPWR VPWR _4323_/X sky130_fd_sc_hd__mux2_1
XFILLER_141_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_254 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7042_ _7042_/CLK _7042_/D fanout520/X VGND VGND VPWR VPWR _7042_/Q sky130_fd_sc_hd__dfrtp_4
X_4254_ hold571/X _6357_/A1 _4254_/S VGND VGND VPWR VPWR _4254_/X sky130_fd_sc_hd__mux2_1
XFILLER_86_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3205_ _6658_/Q VGND VGND VPWR VPWR _3205_/Y sky130_fd_sc_hd__inv_2
X_4185_ _3625_/X _4185_/A1 _4189_/S VGND VGND VPWR VPWR _6594_/D sky130_fd_sc_hd__mux2_1
XFILLER_28_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_694 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6826_ _6978_/CLK _6826_/D fanout490/X VGND VGND VPWR VPWR _6826_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_51_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_263 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6757_ _6976_/CLK _6757_/D fanout501/X VGND VGND VPWR VPWR _6757_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_149_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3969_ hold140/X hold148/X _6624_/Q VGND VGND VPWR VPWR _3969_/X sky130_fd_sc_hd__mux2_1
XFILLER_10_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5708_ _6812_/Q _5913_/A2 _5922_/A2 _6908_/Q VGND VGND VPWR VPWR _5708_/X sky130_fd_sc_hd__a22o_1
XFILLER_149_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_164_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6688_ _6718_/CLK _6688_/D _6401_/A VGND VGND VPWR VPWR _6688_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_148_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5639_ _5667_/A _5651_/B _5649_/C VGND VGND VPWR VPWR _5639_/X sky130_fd_sc_hd__and3b_4
XFILLER_128_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold150 _3990_/X VGND VGND VPWR VPWR _6439_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold161 _6631_/Q VGND VGND VPWR VPWR hold161/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_132_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold172 _4295_/X VGND VGND VPWR VPWR _6693_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold183 _6981_/Q VGND VGND VPWR VPWR hold183/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold194 _5239_/X VGND VGND VPWR VPWR _6813_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_78_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_169_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_186_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5990_ _6834_/Q _5946_/X _6294_/A2 _7079_/Q _5989_/X VGND VGND VPWR VPWR _6002_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_64_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4941_ _4927_/X _4940_/X _5062_/A VGND VGND VPWR VPWR _4941_/Y sky130_fd_sc_hd__a21boi_1
XFILLER_33_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_178_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4872_ _4721_/B _4671_/B _4630_/B _4678_/A VGND VGND VPWR VPWR _4872_/X sky130_fd_sc_hd__a31o_1
XFILLER_33_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6611_ _6707_/CLK _6611_/D _3940_/B VGND VGND VPWR VPWR _6611_/Q sky130_fd_sc_hd__dfstp_2
X_3823_ _6416_/Q _3826_/A VGND VGND VPWR VPWR _3824_/B sky130_fd_sc_hd__nor2_1
XFILLER_177_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_192_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6542_ _6697_/CLK _6542_/D fanout485/X VGND VGND VPWR VPWR _6542_/Q sky130_fd_sc_hd__dfrtp_2
X_3754_ _3754_/A _3754_/B VGND VGND VPWR VPWR _3754_/X sky130_fd_sc_hd__or2_1
XFILLER_192_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6473_ _6565_/CLK _6473_/D fanout495/X VGND VGND VPWR VPWR _6473_/Q sky130_fd_sc_hd__dfrtp_1
X_3685_ _3749_/A1 _3684_/X _3685_/S VGND VGND VPWR VPWR _3685_/X sky130_fd_sc_hd__mux2_1
XFILLER_146_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5424_ _5424_/A _5511_/B VGND VGND VPWR VPWR _5432_/S sky130_fd_sc_hd__and2_4
XFILLER_161_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_160_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_161_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput200 _3188_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[32] sky130_fd_sc_hd__buf_12
Xoutput211 _3213_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[8] sky130_fd_sc_hd__buf_12
Xoutput222 _3926_/X VGND VGND VPWR VPWR mgmt_gpio_out[1] sky130_fd_sc_hd__buf_12
XFILLER_161_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput233 _7174_/X VGND VGND VPWR VPWR mgmt_gpio_out[2] sky130_fd_sc_hd__buf_12
XFILLER_133_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput244 _7177_/X VGND VGND VPWR VPWR mgmt_gpio_out[5] sky130_fd_sc_hd__buf_12
X_5355_ hold371/X _5532_/A1 _5360_/S VGND VGND VPWR VPWR _5355_/X sky130_fd_sc_hd__mux2_1
Xoutput255 _3944_/Y VGND VGND VPWR VPWR pad_flash_io1_ieb sky130_fd_sc_hd__buf_12
Xoutput266 _6741_/Q VGND VGND VPWR VPWR pll_div[4] sky130_fd_sc_hd__buf_12
Xoutput277 _6433_/Q VGND VGND VPWR VPWR pll_trim[15] sky130_fd_sc_hd__buf_12
X_4306_ hold773/X _6355_/A1 _4308_/S VGND VGND VPWR VPWR _4306_/X sky130_fd_sc_hd__mux2_1
Xoutput288 _6749_/Q VGND VGND VPWR VPWR pll_trim[25] sky130_fd_sc_hd__buf_12
XFILLER_114_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput299 _6753_/Q VGND VGND VPWR VPWR pwr_ctrl_out[2] sky130_fd_sc_hd__buf_12
XFILLER_102_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5286_ hold737/X _5457_/A1 _5288_/S VGND VGND VPWR VPWR _5286_/X sky130_fd_sc_hd__mux2_1
XFILLER_141_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_235 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7025_ _7069_/CLK _7025_/D fanout516/X VGND VGND VPWR VPWR _7025_/Q sky130_fd_sc_hd__dfrtp_2
X_4237_ _4237_/A _6352_/B VGND VGND VPWR VPWR _4242_/S sky130_fd_sc_hd__and2_2
X_4168_ hold961/X _5189_/A1 _4171_/S VGND VGND VPWR VPWR _4168_/X sky130_fd_sc_hd__mux2_1
XFILLER_55_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4099_ _4099_/A0 hold3/X hold8/X VGND VGND VPWR VPWR hold9/A sky130_fd_sc_hd__mux2_1
XFILLER_55_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_252 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6809_ _7070_/CLK _6809_/D fanout507/X VGND VGND VPWR VPWR _6809_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_168_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_600 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_70_csclk clkbuf_3_1_0_csclk/X VGND VGND VPWR VPWR _7063_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_137_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_99 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_152_614 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_155_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_98 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_132_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout460 _4299_/A1 VGND VGND VPWR VPWR _5531_/A1 sky130_fd_sc_hd__buf_4
Xfanout471 hold7/X VGND VGND VPWR VPWR _5511_/B sky130_fd_sc_hd__clkbuf_16
XFILLER_19_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout482 _3263_/Y VGND VGND VPWR VPWR _6396_/B sky130_fd_sc_hd__clkbuf_16
XFILLER_48_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout493 _6401_/A VGND VGND VPWR VPWR _6400_/A sky130_fd_sc_hd__buf_4
XFILLER_120_599 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_631 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_23_csclk _6684_/CLK VGND VGND VPWR VPWR _7079_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_187_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_128_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_174_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_38_csclk clkbuf_3_7_0_csclk/X VGND VGND VPWR VPWR _7060_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_155_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold908 _4207_/X VGND VGND VPWR VPWR _6613_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold919 _6849_/Q VGND VGND VPWR VPWR hold919/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_115_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3470_ _3470_/A _3470_/B _3470_/C _3470_/D VGND VGND VPWR VPWR _3470_/Y sky130_fd_sc_hd__nor4_1
XFILLER_182_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_179 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5140_ _5121_/X _5134_/X _5136_/Y _5102_/X VGND VGND VPWR VPWR _5140_/X sky130_fd_sc_hd__a22o_1
XFILLER_36_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5071_ _5068_/A _5065_/Y _5068_/B _5131_/B _5112_/B VGND VGND VPWR VPWR _5071_/X
+ sky130_fd_sc_hd__o41a_1
X_4022_ hold931/X _6354_/A1 _4025_/S VGND VGND VPWR VPWR _4022_/X sky130_fd_sc_hd__mux2_1
XFILLER_84_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5973_ _5973_/A _5973_/B _5973_/C _5973_/D VGND VGND VPWR VPWR _5973_/Y sky130_fd_sc_hd__nor4_1
XFILLER_64_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4924_ _4985_/A _4924_/B _4935_/B _4921_/Y VGND VGND VPWR VPWR _4924_/X sky130_fd_sc_hd__or4b_1
XFILLER_33_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_178_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4855_ _4965_/A _4962_/C VGND VGND VPWR VPWR _4855_/X sky130_fd_sc_hd__and2_1
XFILLER_138_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3806_ _6946_/Q _5388_/A _5158_/A _6748_/Q VGND VGND VPWR VPWR _3814_/B sky130_fd_sc_hd__a22o_1
X_4786_ _4786_/A VGND VGND VPWR VPWR _4786_/Y sky130_fd_sc_hd__inv_2
XFILLER_193_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6525_ _6527_/CLK _6525_/D fanout524/X VGND VGND VPWR VPWR _6525_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_181_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3737_ _6476_/Q _4032_/A _4291_/A _6691_/Q VGND VGND VPWR VPWR _3737_/X sky130_fd_sc_hd__a22o_1
XFILLER_118_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_655 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6456_ _6696_/CLK _6456_/D fanout495/X VGND VGND VPWR VPWR _6456_/Q sky130_fd_sc_hd__dfrtp_1
X_3668_ _6682_/Q _4279_/A _4291_/A _6692_/Q VGND VGND VPWR VPWR _3668_/X sky130_fd_sc_hd__a22o_1
XFILLER_133_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5407_ _5407_/A0 _5530_/A1 _5414_/S VGND VGND VPWR VPWR _5407_/X sky130_fd_sc_hd__mux2_1
X_6387_ _6400_/A _6399_/B VGND VGND VPWR VPWR _6387_/X sky130_fd_sc_hd__and2_1
XFILLER_133_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3599_ _6745_/Q _5151_/A _3572_/Y input95/X VGND VGND VPWR VPWR _3599_/X sky130_fd_sc_hd__a22o_1
XFILLER_88_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5338_ hold347/X _5515_/A1 _5342_/S VGND VGND VPWR VPWR _5338_/X sky130_fd_sc_hd__mux2_1
XFILLER_142_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_190 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5269_ hold634/X _5545_/A1 _5270_/S VGND VGND VPWR VPWR _5269_/X sky130_fd_sc_hd__mux2_1
XFILLER_102_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7008_ _7069_/CLK _7008_/D fanout516/X VGND VGND VPWR VPWR _7008_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_28_344 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_723 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_140_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_691 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_182_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_341 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4640_ _4692_/C _4640_/B VGND VGND VPWR VPWR _4640_/X sky130_fd_sc_hd__or2_1
XFILLER_187_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4571_ _4692_/A _5022_/B _4568_/X _4570_/X VGND VGND VPWR VPWR _4579_/B sky130_fd_sc_hd__o211a_1
Xmax_cap402 _5645_/X VGND VGND VPWR VPWR _5917_/B1 sky130_fd_sc_hd__buf_12
X_6310_ _3747_/Y _6310_/A1 _6316_/S VGND VGND VPWR VPWR _7134_/D sky130_fd_sc_hd__mux2_1
XFILLER_128_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmax_cap413 _5627_/X VGND VGND VPWR VPWR _5913_/A2 sky130_fd_sc_hd__buf_6
X_3522_ _3523_/A _3560_/B VGND VGND VPWR VPWR _4196_/A sky130_fd_sc_hd__nor2_8
Xhold705 _7005_/Q VGND VGND VPWR VPWR hold705/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_171_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_128_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold716 _5419_/X VGND VGND VPWR VPWR _6973_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold727 _7031_/Q VGND VGND VPWR VPWR hold727/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold738 _5286_/X VGND VGND VPWR VPWR _6855_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6241_ _6687_/Q _5942_/X _5972_/B _6692_/Q _6234_/X VGND VGND VPWR VPWR _6251_/A
+ sky130_fd_sc_hd__a221o_1
Xhold749 _7084_/Q VGND VGND VPWR VPWR hold749/X sky130_fd_sc_hd__dlygate4sd3_1
X_3453_ _7076_/Q _5529_/A _3384_/Y input25/X _3452_/X VGND VGND VPWR VPWR _3454_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_171_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6172_ _6993_/Q _6286_/B1 _5977_/X _6929_/Q _6171_/X VGND VGND VPWR VPWR _6177_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_130_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3384_ _3706_/B _3391_/B VGND VGND VPWR VPWR _3384_/Y sky130_fd_sc_hd__nor2_8
XFILLER_130_127 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5123_ _4721_/B _5026_/A _4788_/A _5122_/X _5106_/A VGND VGND VPWR VPWR _5123_/X
+ sky130_fd_sc_hd__o311a_1
Xhold1405 _6585_/Q VGND VGND VPWR VPWR _4175_/A1 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1416 _6443_/Q VGND VGND VPWR VPWR hold979/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_57_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1427 _7134_/Q VGND VGND VPWR VPWR _6310_/A1 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1438 _6733_/Q VGND VGND VPWR VPWR _3435_/A1 sky130_fd_sc_hd__dlygate4sd3_1
X_5054_ _5081_/B _5054_/B _5054_/C VGND VGND VPWR VPWR _5055_/D sky130_fd_sc_hd__and3_1
Xhold1449 _6638_/Q VGND VGND VPWR VPWR _3872_/B1 sky130_fd_sc_hd__dlygate4sd3_1
X_4005_ hold809/X _6355_/A1 _4007_/S VGND VGND VPWR VPWR _4005_/X sky130_fd_sc_hd__mux2_1
XFILLER_25_303 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_472 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5956_ _5981_/A _5963_/C _5981_/C VGND VGND VPWR VPWR _5956_/X sky130_fd_sc_hd__and3_1
XFILLER_52_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4907_ _4944_/A _4489_/B _4751_/Y _4899_/Y VGND VGND VPWR VPWR _5010_/B sky130_fd_sc_hd__a211o_1
XFILLER_33_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5887_ _6542_/Q _5667_/X _5876_/X _5886_/X _5610_/A VGND VGND VPWR VPWR _5887_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_139_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4838_ _4692_/A _4831_/X _4828_/A VGND VGND VPWR VPWR _4839_/D sky130_fd_sc_hd__a21o_1
XFILLER_193_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4769_ _4943_/A _4515_/B _4720_/C VGND VGND VPWR VPWR _5008_/C sky130_fd_sc_hd__o21ba_1
X_6508_ _7124_/CLK _6508_/D fanout502/X VGND VGND VPWR VPWR _6508_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_193_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6439_ _7034_/CLK _6439_/D fanout488/X VGND VGND VPWR VPWR _6439_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_162_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold10 hold10/A VGND VGND VPWR VPWR hold10/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold21 hold21/A VGND VGND VPWR VPWR hold21/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold32 hold32/A VGND VGND VPWR VPWR hold32/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_76_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold43 hold43/A VGND VGND VPWR VPWR hold43/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold54 hold54/A VGND VGND VPWR VPWR hold54/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_75_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold65 hold65/A VGND VGND VPWR VPWR hold65/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold76 hold76/A VGND VGND VPWR VPWR hold76/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_188_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold87 hold87/A VGND VGND VPWR VPWR hold87/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_28_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold98 hold98/A VGND VGND VPWR VPWR hold98/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_44_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_189_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_667 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_172_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_7 _5208_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_137_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_153_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_112_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5810_ _6905_/Q _5623_/X _5637_/X _6857_/Q _5809_/X VGND VGND VPWR VPWR _5810_/X
+ sky130_fd_sc_hd__a221o_1
X_6790_ _6965_/CLK _6790_/D fanout514/X VGND VGND VPWR VPWR _6790_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_50_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5741_ _6990_/Q _5622_/X _5637_/X _6854_/Q VGND VGND VPWR VPWR _5741_/X sky130_fd_sc_hd__a22o_1
XFILLER_187_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_188_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5672_ _6843_/Q _5632_/X _5639_/X _6803_/Q VGND VGND VPWR VPWR _5672_/X sky130_fd_sc_hd__a22o_1
XFILLER_30_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_175_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_148_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4623_ _4630_/A _4623_/B VGND VGND VPWR VPWR _4784_/A sky130_fd_sc_hd__xnor2_1
XFILLER_163_539 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4554_ _4554_/A _4575_/B VGND VGND VPWR VPWR _4965_/C sky130_fd_sc_hd__or2_4
Xhold502 _4100_/X VGND VGND VPWR VPWR _6521_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold513 _6468_/Q VGND VGND VPWR VPWR hold513/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold524 _5293_/X VGND VGND VPWR VPWR _6861_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3505_ input56/X _5190_/A _5397_/A _6958_/Q VGND VGND VPWR VPWR _3505_/X sky130_fd_sc_hd__a22o_1
Xhold535 _6689_/Q VGND VGND VPWR VPWR hold535/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold546 _5225_/X VGND VGND VPWR VPWR _6801_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_144_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4485_ _4977_/B _4692_/C _4965_/B _4988_/A _4622_/A VGND VGND VPWR VPWR _4648_/C
+ sky130_fd_sc_hd__o32a_1
XFILLER_171_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold557 _6893_/Q VGND VGND VPWR VPWR hold557/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold568 _4299_/X VGND VGND VPWR VPWR _6696_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6224_ _6656_/Q _6288_/A2 _5948_/X _6546_/Q VGND VGND VPWR VPWR _6224_/X sky130_fd_sc_hd__a22o_1
Xhold579 _6664_/Q VGND VGND VPWR VPWR hold579/X sky130_fd_sc_hd__dlygate4sd3_1
X_3436_ _7031_/Q _5478_/A _5235_/A _6815_/Q VGND VGND VPWR VPWR _3436_/X sky130_fd_sc_hd__a22o_1
XFILLER_131_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6155_ _6179_/A1 _5612_/Y _6153_/X _6154_/X VGND VGND VPWR VPWR _7125_/D sky130_fd_sc_hd__o22a_1
XTAP_851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3367_ _3706_/B _3560_/B VGND VGND VPWR VPWR _3984_/A sky130_fd_sc_hd__nor2_8
XTAP_862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1202 _5384_/X VGND VGND VPWR VPWR _6942_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5106_ _5106_/A _5106_/B _5106_/C _5135_/D VGND VGND VPWR VPWR _5106_/Y sky130_fd_sc_hd__nand4_1
XTAP_884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1213 _6742_/Q VGND VGND VPWR VPWR _5152_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_57_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1224 _4122_/X VGND VGND VPWR VPWR _6540_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6086_ _6958_/Q _5957_/X _5978_/X _6950_/Q VGND VGND VPWR VPWR _6086_/X sky130_fd_sc_hd__a22o_1
Xhold1235 _6434_/Q VGND VGND VPWR VPWR _3985_/A0 sky130_fd_sc_hd__dlygate4sd3_1
X_3298_ hold39/X hold50/X VGND VGND VPWR VPWR _3366_/A sky130_fd_sc_hd__nand2_1
Xhold1246 _5240_/X VGND VGND VPWR VPWR _6814_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1257 _6442_/Q VGND VGND VPWR VPWR _3994_/A0 sky130_fd_sc_hd__dlygate4sd3_1
X_5037_ _5037_/A _5090_/A _5037_/C _5037_/D VGND VGND VPWR VPWR _5038_/C sky130_fd_sc_hd__and4_1
Xhold1268 _4167_/X VGND VGND VPWR VPWR _6578_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_73_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1279 _6870_/Q VGND VGND VPWR VPWR _5303_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_604 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6988_ _6988_/CLK _6988_/D fanout518/X VGND VGND VPWR VPWR _6988_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_15_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5939_ _5979_/A _5979_/B _5963_/C VGND VGND VPWR VPWR _5939_/X sky130_fd_sc_hd__and3_4
XFILLER_139_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_683 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_178_182 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_166_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_147_44 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_147_99 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput100 wb_adr_i[10] VGND VGND VPWR VPWR _4336_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_88_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput111 wb_adr_i[20] VGND VGND VPWR VPWR _4544_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_49_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput122 wb_adr_i[30] VGND VGND VPWR VPWR input122/X sky130_fd_sc_hd__clkbuf_1
XFILLER_103_683 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput133 wb_dat_i[10] VGND VGND VPWR VPWR _6330_/B1 sky130_fd_sc_hd__clkbuf_1
XFILLER_48_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput144 wb_dat_i[20] VGND VGND VPWR VPWR _6335_/A2 sky130_fd_sc_hd__clkbuf_1
Xinput155 wb_dat_i[30] VGND VGND VPWR VPWR _6341_/A2 sky130_fd_sc_hd__clkbuf_1
Xinput166 wb_sel_i[1] VGND VGND VPWR VPWR _6348_/B1 sky130_fd_sc_hd__clkbuf_1
XFILLER_76_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_442 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_185_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_145_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_126_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4270_ hold787/X _5505_/A1 _4272_/S VGND VGND VPWR VPWR _4270_/X sky130_fd_sc_hd__mux2_1
XFILLER_113_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_203 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6911_ _6999_/CLK _6911_/D fanout524/X VGND VGND VPWR VPWR _6911_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_63_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6842_ _7041_/CLK _6842_/D fanout520/X VGND VGND VPWR VPWR _6842_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_90_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6773_ _7042_/CLK _6773_/D fanout523/X VGND VGND VPWR VPWR _7192_/A sky130_fd_sc_hd__dfrtp_1
X_3985_ _3985_/A0 _6353_/A1 _3992_/S VGND VGND VPWR VPWR _3985_/X sky130_fd_sc_hd__mux2_1
XFILLER_22_158 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5724_ _6981_/Q _5642_/X _5807_/B1 _6933_/Q _5714_/Y VGND VGND VPWR VPWR _5724_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_31_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5655_ _6866_/Q _5928_/B1 _5627_/X _6810_/Q VGND VGND VPWR VPWR _5655_/X sky130_fd_sc_hd__a22o_1
X_4606_ _4717_/A VGND VGND VPWR VPWR _4606_/Y sky130_fd_sc_hd__inv_2
X_5586_ _7098_/Q _7097_/Q VGND VGND VPWR VPWR _5976_/A sky130_fd_sc_hd__or2_4
XFILLER_191_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold310 _4326_/X VGND VGND VPWR VPWR _6719_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_163_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4537_ _4828_/A _4537_/B VGND VGND VPWR VPWR _4537_/X sky130_fd_sc_hd__and2_1
Xhold321 _6988_/Q VGND VGND VPWR VPWR hold321/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_132_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold332 _5220_/X VGND VGND VPWR VPWR _6796_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold343 _6869_/Q VGND VGND VPWR VPWR hold343/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold354 _5248_/X VGND VGND VPWR VPWR _6821_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold365 _6788_/Q VGND VGND VPWR VPWR hold365/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold376 _5265_/X VGND VGND VPWR VPWR _6836_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4468_ _4640_/B _5022_/B VGND VGND VPWR VPWR _4732_/A sky130_fd_sc_hd__nor2_1
XFILLER_77_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold387 _6529_/Q VGND VGND VPWR VPWR hold387/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold398 _5166_/X VGND VGND VPWR VPWR _6753_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6207_ _6646_/Q _5950_/X _6270_/B1 _6676_/Q _6206_/X VGND VGND VPWR VPWR _6207_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_89_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3419_ _6448_/Q _3993_/A _5397_/A _6960_/Q _3418_/X VGND VGND VPWR VPWR _3419_/X
+ sky130_fd_sc_hd__a221o_2
X_7187_ _7187_/A VGND VGND VPWR VPWR _7187_/X sky130_fd_sc_hd__clkbuf_1
X_4399_ _4429_/B _4399_/B VGND VGND VPWR VPWR _4892_/A sky130_fd_sc_hd__nand2_2
XFILLER_98_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6138_ _6960_/Q _5957_/X _5974_/B _6832_/Q VGND VGND VPWR VPWR _6138_/X sky130_fd_sc_hd__a22o_1
XTAP_681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1010 _6454_/Q VGND VGND VPWR VPWR _4007_/A0 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1021 _5426_/X VGND VGND VPWR VPWR _6979_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_85_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1032 _6743_/Q VGND VGND VPWR VPWR _5153_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_133_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1043 _5372_/X VGND VGND VPWR VPWR _6931_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1054 _6947_/Q VGND VGND VPWR VPWR _5390_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_58_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6069_ _6837_/Q _5946_/X _5962_/X _6893_/Q VGND VGND VPWR VPWR _6069_/X sky130_fd_sc_hd__a22o_1
Xhold1065 _5371_/X VGND VGND VPWR VPWR _6930_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1076 _4232_/X VGND VGND VPWR VPWR _6630_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_73_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1087 _7063_/Q VGND VGND VPWR VPWR _5521_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_205 _5515_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1098 _5267_/X VGND VGND VPWR VPWR _6838_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_216 _5969_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_442 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_166_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_182_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_491 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_189_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3770_ _3952_/A _4112_/B _5253_/A _6826_/Q _3769_/X VGND VGND VPWR VPWR _3777_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_158_631 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_692 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_158_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5440_ hold128/X _5476_/A1 hold35/X VGND VGND VPWR VPWR _5440_/X sky130_fd_sc_hd__mux2_1
XFILLER_66_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5371_ _5371_/A0 _5521_/A1 hold42/X VGND VGND VPWR VPWR _5371_/X sky130_fd_sc_hd__mux2_1
X_7110_ _7131_/CLK _7110_/D fanout499/X VGND VGND VPWR VPWR _7110_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_113_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4322_ _4322_/A0 _5308_/A1 _4326_/S VGND VGND VPWR VPWR _4322_/X sky130_fd_sc_hd__mux2_1
XFILLER_113_211 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7041_ _7041_/CLK _7041_/D fanout520/X VGND VGND VPWR VPWR _7041_/Q sky130_fd_sc_hd__dfrtp_4
X_4253_ hold259/X hold46/X _4254_/S VGND VGND VPWR VPWR _4253_/X sky130_fd_sc_hd__mux2_1
XFILLER_87_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_266 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3204_ _6917_/Q VGND VGND VPWR VPWR _3204_/Y sky130_fd_sc_hd__clkinv_2
X_4184_ _3684_/X _4184_/A1 _4189_/S VGND VGND VPWR VPWR _6593_/D sky130_fd_sc_hd__mux2_1
XFILLER_95_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_3_7_0_wb_clk_i clkbuf_3_7_0_wb_clk_i/A VGND VGND VPWR VPWR _3931_/A1 sky130_fd_sc_hd__clkbuf_8
X_6825_ _7017_/CLK _6825_/D fanout507/X VGND VGND VPWR VPWR _6825_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_23_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_467 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3968_ hold437/X _5534_/A1 _3974_/S VGND VGND VPWR VPWR _3968_/X sky130_fd_sc_hd__mux2_1
X_6756_ _6994_/CLK _6756_/D fanout490/X VGND VGND VPWR VPWR _7173_/A sky130_fd_sc_hd__dfrtp_2
XFILLER_50_275 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5707_ _6844_/Q _5922_/B1 _5705_/X _5706_/X VGND VGND VPWR VPWR _5707_/X sky130_fd_sc_hd__a211o_1
X_6687_ _6689_/CLK _6687_/D fanout510/X VGND VGND VPWR VPWR _6687_/Q sky130_fd_sc_hd__dfstp_1
X_3899_ _4334_/C _4334_/D _3899_/C input116/X VGND VGND VPWR VPWR _3900_/D sky130_fd_sc_hd__or4b_1
XFILLER_164_623 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5638_ _6818_/Q _5636_/X _5918_/B1 _6850_/Q VGND VGND VPWR VPWR _5638_/X sky130_fd_sc_hd__a22o_1
XFILLER_164_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_191_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5569_ _7093_/Q _7092_/Q VGND VGND VPWR VPWR _5645_/B sky130_fd_sc_hd__and2_2
XFILLER_117_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_163_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold140 _7164_/Q VGND VGND VPWR VPWR hold140/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold151 _6747_/Q VGND VGND VPWR VPWR hold151/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold162 _4233_/X VGND VGND VPWR VPWR _6631_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold173 _6782_/Q VGND VGND VPWR VPWR hold173/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold184 _5428_/X VGND VGND VPWR VPWR _6981_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold195 _7017_/Q VGND VGND VPWR VPWR hold195/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_77_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_288 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_684 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_704 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_135_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_92_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4940_ _4991_/A _4940_/B _4940_/C _4940_/D VGND VGND VPWR VPWR _4940_/X sky130_fd_sc_hd__and4b_1
XFILLER_64_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4871_ _4631_/A _4870_/X _4869_/X _4679_/Y _4616_/X VGND VGND VPWR VPWR _4878_/B
+ sky130_fd_sc_hd__o2111a_1
XTAP_2890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_404 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6610_ _6769_/CLK _6610_/D fanout492/X VGND VGND VPWR VPWR _6610_/Q sky130_fd_sc_hd__dfrtp_2
X_3822_ _3867_/A _3825_/B _3824_/A _3165_/A VGND VGND VPWR VPWR _6417_/D sky130_fd_sc_hd__o22a_1
XFILLER_177_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_437 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6541_ _7153_/CLK _6541_/D fanout486/X VGND VGND VPWR VPWR _6541_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_193_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3753_ _6994_/Q _5442_/A _4127_/A _6545_/Q _3752_/X VGND VGND VPWR VPWR _3754_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_192_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6472_ _6683_/CLK _6472_/D fanout509/X VGND VGND VPWR VPWR _6472_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_118_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_146_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3684_ _3684_/A _3684_/B _3684_/C _3683_/Y VGND VGND VPWR VPWR _3684_/X sky130_fd_sc_hd__or4b_4
X_5423_ hold227/X hold27/X _5423_/S VGND VGND VPWR VPWR _5423_/X sky130_fd_sc_hd__mux2_1
XFILLER_133_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput201 _3187_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[33] sky130_fd_sc_hd__buf_12
Xoutput212 _3212_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[9] sky130_fd_sc_hd__buf_12
XFILLER_145_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_173_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput223 _7185_/X VGND VGND VPWR VPWR mgmt_gpio_out[20] sky130_fd_sc_hd__buf_12
Xoutput234 _7195_/X VGND VGND VPWR VPWR mgmt_gpio_out[30] sky130_fd_sc_hd__buf_12
X_5354_ hold980/X _5495_/A1 _5360_/S VGND VGND VPWR VPWR _5354_/X sky130_fd_sc_hd__mux2_1
Xoutput245 _3923_/X VGND VGND VPWR VPWR mgmt_gpio_out[6] sky130_fd_sc_hd__buf_12
Xoutput256 _3944_/A VGND VGND VPWR VPWR pad_flash_io1_oeb sky130_fd_sc_hd__buf_12
Xoutput267 _6735_/Q VGND VGND VPWR VPWR pll_ena sky130_fd_sc_hd__buf_12
X_4305_ hold949/X _6354_/A1 _4308_/S VGND VGND VPWR VPWR _4305_/X sky130_fd_sc_hd__mux2_1
Xoutput278 _6418_/Q VGND VGND VPWR VPWR pll_trim[16] sky130_fd_sc_hd__buf_12
Xoutput289 _6436_/Q VGND VGND VPWR VPWR pll_trim[2] sky130_fd_sc_hd__buf_12
XFILLER_141_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5285_ _5285_/A0 _5465_/A1 _5288_/S VGND VGND VPWR VPWR _5285_/X sky130_fd_sc_hd__mux2_1
XFILLER_114_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7024_ _7060_/CLK _7024_/D fanout521/X VGND VGND VPWR VPWR _7024_/Q sky130_fd_sc_hd__dfrtp_2
X_4236_ hold897/X _4236_/A1 _4236_/S VGND VGND VPWR VPWR _4236_/X sky130_fd_sc_hd__mux2_1
XFILLER_101_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4167_ _4167_/A0 _5308_/A1 _4171_/S VGND VGND VPWR VPWR _4167_/X sky130_fd_sc_hd__mux2_1
X_4098_ _4098_/A0 _6354_/A1 hold8/X VGND VGND VPWR VPWR _4098_/X sky130_fd_sc_hd__mux2_1
XFILLER_82_164 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_4_csclk clkbuf_3_1_0_csclk/X VGND VGND VPWR VPWR _6718_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_169_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_169_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_169_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6808_ _6961_/CLK _6808_/D fanout516/X VGND VGND VPWR VPWR _6808_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_23_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6739_ _7037_/CLK _6739_/D fanout484/X VGND VGND VPWR VPWR _6739_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_137_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_472 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_164_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_155_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_151_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout450 hold45/X VGND VGND VPWR VPWR hold46/A sky130_fd_sc_hd__buf_6
XFILLER_48_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout461 hold90/X VGND VGND VPWR VPWR _4299_/A1 sky130_fd_sc_hd__clkbuf_8
XFILLER_171_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout472 hold7/X VGND VGND VPWR VPWR _5538_/B sky130_fd_sc_hd__buf_4
XFILLER_59_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout483 input99/X VGND VGND VPWR VPWR _4542_/A sky130_fd_sc_hd__buf_8
Xfanout494 fanout496/X VGND VGND VPWR VPWR _6401_/A sky130_fd_sc_hd__buf_6
XFILLER_59_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_754 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_159_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_612 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold909 _6945_/Q VGND VGND VPWR VPWR hold909/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_182_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_183_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_158 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5070_ _5070_/A _5070_/B _5070_/C VGND VGND VPWR VPWR _5131_/B sky130_fd_sc_hd__nand3_1
XFILLER_29_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4021_ _4021_/A0 _6353_/A1 _4025_/S VGND VGND VPWR VPWR _4021_/X sky130_fd_sc_hd__mux2_1
XFILLER_64_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_624 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5972_ _5972_/A _5972_/B _5972_/C _5971_/Y VGND VGND VPWR VPWR _5973_/D sky130_fd_sc_hd__or4b_1
XFILLER_64_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4923_ _4576_/X _4640_/X _4788_/A VGND VGND VPWR VPWR _4929_/B sky130_fd_sc_hd__a21oi_1
XFILLER_178_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4854_ _4854_/A _4854_/B VGND VGND VPWR VPWR _5087_/B sky130_fd_sc_hd__nor2_2
XFILLER_178_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3805_ _7063_/Q _5520_/A _3803_/X _3804_/Y VGND VGND VPWR VPWR _3814_/A sky130_fd_sc_hd__a22o_1
XFILLER_178_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4785_ _4935_/A _4785_/B VGND VGND VPWR VPWR _4786_/A sky130_fd_sc_hd__and2b_1
X_3736_ _3736_/A _3736_/B _3736_/C _3736_/D VGND VGND VPWR VPWR _3746_/C sky130_fd_sc_hd__nor4_1
X_6524_ _6527_/CLK _6524_/D fanout524/X VGND VGND VPWR VPWR _6524_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_109_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6455_ _7038_/CLK _6455_/D fanout490/X VGND VGND VPWR VPWR _6455_/Q sky130_fd_sc_hd__dfrtp_1
X_3667_ _3667_/A _3667_/B _3667_/C wire348/X VGND VGND VPWR VPWR _3684_/B sky130_fd_sc_hd__or4b_1
X_5406_ _5406_/A _5511_/B VGND VGND VPWR VPWR _5414_/S sky130_fd_sc_hd__and2_4
X_6386_ _6400_/A _6401_/B VGND VGND VPWR VPWR _6386_/X sky130_fd_sc_hd__and2_1
X_3598_ _6965_/Q _5406_/A _3384_/Y input23/X _3597_/X VGND VGND VPWR VPWR _3605_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_133_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5337_ _5337_/A0 hold3/X _5342_/S VGND VGND VPWR VPWR hold13/A sky130_fd_sc_hd__mux2_1
XFILLER_102_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_114_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_87_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5268_ hold701/X _5544_/A1 _5270_/S VGND VGND VPWR VPWR _5268_/X sky130_fd_sc_hd__mux2_1
XFILLER_85_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_102_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4219_ hold539/X _6357_/A1 _4219_/S VGND VGND VPWR VPWR _4219_/X sky130_fd_sc_hd__mux2_1
X_7007_ _7029_/CLK _7007_/D fanout522/X VGND VGND VPWR VPWR _7007_/Q sky130_fd_sc_hd__dfrtp_1
X_5199_ _6396_/B hold76/X _5538_/B VGND VGND VPWR VPWR _5207_/S sky130_fd_sc_hd__and3b_4
XFILLER_28_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_141_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_1_1__f__1162_ clkbuf_0__1162_/X VGND VGND VPWR VPWR _6313_/A0 sky130_fd_sc_hd__clkbuf_16
XFILLER_165_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_411 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_147 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_378 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4570_ _4691_/A _4570_/B _4569_/X VGND VGND VPWR VPWR _4570_/X sky130_fd_sc_hd__or3b_1
XFILLER_190_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3521_ _7022_/Q hold18/A _5343_/A _6910_/Q _3520_/X VGND VGND VPWR VPWR _3535_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_155_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmax_cap403 _5643_/X VGND VGND VPWR VPWR _5913_/B1 sky130_fd_sc_hd__buf_12
Xmax_cap414 _5626_/X VGND VGND VPWR VPWR _5924_/B2 sky130_fd_sc_hd__buf_12
Xhold706 _5455_/X VGND VGND VPWR VPWR _7005_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold717 _7023_/Q VGND VGND VPWR VPWR hold717/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold728 _5484_/X VGND VGND VPWR VPWR _7031_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6240_ _6457_/Q _6291_/A2 _6232_/X _6237_/X _6239_/X VGND VGND VPWR VPWR _6252_/B
+ sky130_fd_sc_hd__a2111o_1
XFILLER_6_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3452_ _6967_/Q _5406_/A _5460_/A _7015_/Q VGND VGND VPWR VPWR _3452_/X sky130_fd_sc_hd__a22o_2
Xhold739 _6877_/Q VGND VGND VPWR VPWR hold739/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_170_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6171_ _6809_/Q _5973_/B _5962_/X _6897_/Q VGND VGND VPWR VPWR _6171_/X sky130_fd_sc_hd__a22o_1
XFILLER_131_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3383_ _3503_/A hold82/X VGND VGND VPWR VPWR _5388_/A sky130_fd_sc_hd__nor2_8
XFILLER_124_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5122_ _4640_/B _4588_/B _5026_/B _4581_/A _4523_/A VGND VGND VPWR VPWR _5122_/X
+ sky130_fd_sc_hd__o221a_1
Xhold1406 _6570_/Q VGND VGND VPWR VPWR _4158_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_29_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1417 _3995_/X VGND VGND VPWR VPWR _6443_/D sky130_fd_sc_hd__dlygate4sd3_1
X_5053_ _4501_/B _4965_/C _4967_/X _5052_/X VGND VGND VPWR VPWR _5054_/C sky130_fd_sc_hd__o211a_1
Xhold1428 _7133_/Q VGND VGND VPWR VPWR _6309_/A1 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1439 _3435_/X VGND VGND VPWR VPWR _6733_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_84_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4004_ hold521/X _4299_/A1 _4007_/S VGND VGND VPWR VPWR _4004_/X sky130_fd_sc_hd__mux2_1
XFILLER_38_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_646 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5955_ _5981_/A _5979_/A _5981_/B VGND VGND VPWR VPWR _5955_/X sky130_fd_sc_hd__and3_4
XFILLER_40_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4906_ _4906_/A _5074_/B _4906_/C VGND VGND VPWR VPWR _4914_/A sky130_fd_sc_hd__and3_1
X_5886_ _5886_/A _5886_/B _5886_/C _5885_/Y VGND VGND VPWR VPWR _5886_/X sky130_fd_sc_hd__or4b_1
XFILLER_139_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_166_504 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4837_ _4943_/B _4988_/A _4649_/A _4537_/B VGND VGND VPWR VPWR _4839_/C sky130_fd_sc_hd__a31o_1
XFILLER_193_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_147_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4768_ _4767_/X _4714_/A _4768_/C _5017_/C VGND VGND VPWR VPWR _4770_/B sky130_fd_sc_hd__and4bb_1
X_6507_ _7124_/CLK _6507_/D fanout502/X VGND VGND VPWR VPWR _6507_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_107_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3719_ _3719_/A _5183_/A VGND VGND VPWR VPWR _5158_/A sky130_fd_sc_hd__nor2_2
X_4699_ _4713_/A _5005_/B VGND VGND VPWR VPWR _5017_/B sky130_fd_sc_hd__or2_1
XFILLER_134_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6438_ _7034_/CLK _6438_/D fanout488/X VGND VGND VPWR VPWR _6438_/Q sky130_fd_sc_hd__dfstp_2
X_6369_ _6370_/A _6401_/B VGND VGND VPWR VPWR _6369_/X sky130_fd_sc_hd__and2_1
Xclkbuf_leaf_22_csclk _6684_/CLK VGND VGND VPWR VPWR _7051_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold11 hold11/A VGND VGND VPWR VPWR hold2/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_48_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold22 hold68/X VGND VGND VPWR VPWR hold69/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_29_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold33 hold33/A VGND VGND VPWR VPWR hold33/X sky130_fd_sc_hd__buf_6
Xhold44 hold44/A VGND VGND VPWR VPWR hold44/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_76_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold55 hold55/A VGND VGND VPWR VPWR hold55/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_29_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold66 hold66/A VGND VGND VPWR VPWR hold66/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold77 hold77/A VGND VGND VPWR VPWR hold77/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold88 hold88/A VGND VGND VPWR VPWR hold88/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold99 hold99/A VGND VGND VPWR VPWR hold99/X sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_37_csclk clkbuf_3_7_0_csclk/X VGND VGND VPWR VPWR _7058_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_44_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_679 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_178 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_0_mgmt_gpio_in[4] mgmt_gpio_in[4] VGND VGND VPWR VPWR clkbuf_0_mgmt_gpio_in[4]/X
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_31_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_570 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_8 _5298_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_156 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5740_ _5740_/A _5740_/B VGND VGND VPWR VPWR _5740_/X sky130_fd_sc_hd__or2_1
XFILLER_96_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5671_ _6987_/Q _5622_/X _5920_/A2 _6827_/Q VGND VGND VPWR VPWR _5671_/X sky130_fd_sc_hd__a22o_1
X_4622_ _4622_/A _4965_/A VGND VGND VPWR VPWR _5061_/A sky130_fd_sc_hd__or2_1
XFILLER_135_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4553_ _4746_/A _4575_/B VGND VGND VPWR VPWR _4555_/B sky130_fd_sc_hd__nor2_2
XFILLER_156_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold503 _6433_/Q VGND VGND VPWR VPWR hold503/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold514 _4024_/X VGND VGND VPWR VPWR _6468_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_144_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold525 _6429_/Q VGND VGND VPWR VPWR hold525/X sky130_fd_sc_hd__dlygate4sd3_1
X_3504_ _3523_/A _5183_/B VGND VGND VPWR VPWR _4190_/A sky130_fd_sc_hd__nor2_4
XFILLER_116_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_171_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold536 _4290_/X VGND VGND VPWR VPWR _6689_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4484_ _4622_/A _4988_/A VGND VGND VPWR VPWR _4959_/A sky130_fd_sc_hd__nor2_2
Xhold547 _6713_/Q VGND VGND VPWR VPWR hold547/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_307 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold558 _5329_/X VGND VGND VPWR VPWR _6893_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6223_ _6626_/Q _5973_/A _5957_/X _6706_/Q VGND VGND VPWR VPWR _6223_/X sky130_fd_sc_hd__a22o_1
X_3435_ _3434_/X _3435_/A1 _3749_/S VGND VGND VPWR VPWR _3435_/X sky130_fd_sc_hd__mux2_1
XFILLER_116_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold569 _6965_/Q VGND VGND VPWR VPWR hold569/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_103_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6154_ _6154_/A1 _3878_/Y _5610_/Y VGND VGND VPWR VPWR _6154_/X sky130_fd_sc_hd__o21a_1
XFILLER_131_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3366_ _3366_/A _3440_/B VGND VGND VPWR VPWR _3560_/B sky130_fd_sc_hd__or2_4
XTAP_841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1203 _6710_/Q VGND VGND VPWR VPWR _4316_/A0 sky130_fd_sc_hd__dlygate4sd3_1
X_5105_ _5105_/A _5105_/B _5105_/C VGND VGND VPWR VPWR _5135_/D sky130_fd_sc_hd__and3_1
XTAP_885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1214 _5152_/X VGND VGND VPWR VPWR _6742_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6085_ hold86/A _5955_/X _6294_/B1 _7043_/Q _6084_/X VGND VGND VPWR VPWR _6093_/B
+ sky130_fd_sc_hd__a221o_1
Xhold1225 _6802_/Q VGND VGND VPWR VPWR _5227_/A0 sky130_fd_sc_hd__dlygate4sd3_1
X_3297_ _3503_/A _3719_/A VGND VGND VPWR VPWR _3297_/Y sky130_fd_sc_hd__nor2_2
XTAP_896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1236 _3985_/X VGND VGND VPWR VPWR _6434_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1247 _6418_/Q VGND VGND VPWR VPWR _3960_/A0 sky130_fd_sc_hd__dlygate4sd3_1
X_5036_ _4586_/B _5026_/B _5025_/Y _4513_/A _4585_/X VGND VGND VPWR VPWR _5037_/D
+ sky130_fd_sc_hd__o221a_1
Xhold1258 _3994_/X VGND VGND VPWR VPWR _6442_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1269 _6990_/Q VGND VGND VPWR VPWR _5438_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_432 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6987_ _7082_/CLK hold95/X fanout519/X VGND VGND VPWR VPWR _6987_/Q sky130_fd_sc_hd__dfstp_2
X_5938_ _5979_/A _5978_/B _5963_/C VGND VGND VPWR VPWR _5969_/A sky130_fd_sc_hd__and3_4
XFILLER_15_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_179_695 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5869_ _6621_/Q _5914_/A2 _5633_/X _6667_/Q _5868_/X VGND VGND VPWR VPWR _5872_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_178_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_250 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_193_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_135_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_147_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_651 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput101 wb_adr_i[11] VGND VGND VPWR VPWR _4336_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_103_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput112 wb_adr_i[21] VGND VGND VPWR VPWR _4368_/A sky130_fd_sc_hd__clkbuf_1
Xinput123 wb_adr_i[31] VGND VGND VPWR VPWR input123/X sky130_fd_sc_hd__clkbuf_1
XFILLER_48_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput134 wb_dat_i[11] VGND VGND VPWR VPWR _6332_/B1 sky130_fd_sc_hd__clkbuf_1
Xinput145 wb_dat_i[21] VGND VGND VPWR VPWR _6339_/A2 sky130_fd_sc_hd__clkbuf_1
XFILLER_48_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput156 wb_dat_i[31] VGND VGND VPWR VPWR _6344_/A2 sky130_fd_sc_hd__clkbuf_1
XFILLER_102_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput167 wb_sel_i[2] VGND VGND VPWR VPWR _6318_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_91_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_207 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_646 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_454 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_679 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_240 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_145_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_126_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3220_ _6789_/Q VGND VGND VPWR VPWR _3220_/Y sky130_fd_sc_hd__inv_2
XFILLER_79_351 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_121_492 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6910_ _7043_/CLK _6910_/D _6396_/A VGND VGND VPWR VPWR _6910_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_47_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6841_ _7074_/CLK _6841_/D fanout507/X VGND VGND VPWR VPWR _6841_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_23_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6772_ _7042_/CLK _6772_/D fanout520/X VGND VGND VPWR VPWR _7191_/A sky130_fd_sc_hd__dfrtp_1
X_3984_ _3984_/A _6352_/B VGND VGND VPWR VPWR _3992_/S sky130_fd_sc_hd__and2_2
X_5723_ _6965_/Q _5925_/B1 _5718_/X _5719_/X _5722_/X VGND VGND VPWR VPWR _5723_/X
+ sky130_fd_sc_hd__a2111o_1
X_5654_ _6898_/Q _5918_/A2 _5632_/X _6842_/Q VGND VGND VPWR VPWR _5654_/X sky130_fd_sc_hd__a22o_1
XFILLER_175_142 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4605_ _4609_/B _4617_/A VGND VGND VPWR VPWR _4717_/A sky130_fd_sc_hd__or2_4
XFILLER_191_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5585_ _7098_/Q _7097_/Q VGND VGND VPWR VPWR _5978_/B sky130_fd_sc_hd__nor2_2
XFILLER_163_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold300 _6357_/X VGND VGND VPWR VPWR _7155_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold311 _6844_/Q VGND VGND VPWR VPWR hold311/X sky130_fd_sc_hd__dlygate4sd3_1
X_4536_ _4536_/A VGND VGND VPWR VPWR _4537_/B sky130_fd_sc_hd__clkinv_2
XFILLER_117_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold322 _5436_/X VGND VGND VPWR VPWR _6988_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold333 _7065_/Q VGND VGND VPWR VPWR hold333/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_132_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold344 _5302_/X VGND VGND VPWR VPWR _6869_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_117_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold355 _6908_/Q VGND VGND VPWR VPWR hold355/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold366 _5211_/X VGND VGND VPWR VPWR _6788_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4467_ _4581_/A _4549_/B VGND VGND VPWR VPWR _4774_/A sky130_fd_sc_hd__or2_1
XFILLER_131_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold377 _6996_/Q VGND VGND VPWR VPWR hold377/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_132_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold388 _4109_/X VGND VGND VPWR VPWR _6529_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6206_ _6686_/Q _5942_/X _5979_/X _6451_/Q VGND VGND VPWR VPWR _6206_/X sky130_fd_sc_hd__a22o_1
Xhold399 _6682_/Q VGND VGND VPWR VPWR hold399/X sky130_fd_sc_hd__dlygate4sd3_1
X_3418_ _7016_/Q _5460_/A _5478_/A _7032_/Q VGND VGND VPWR VPWR _3418_/X sky130_fd_sc_hd__a22o_1
X_4398_ _4569_/A _4535_/A VGND VGND VPWR VPWR _4587_/A sky130_fd_sc_hd__nand2_4
X_7186_ _7186_/A VGND VGND VPWR VPWR _7186_/X sky130_fd_sc_hd__clkbuf_1
XTAP_660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1000 _6615_/Q VGND VGND VPWR VPWR _4210_/A0 sky130_fd_sc_hd__dlygate4sd3_1
X_3349_ _3349_/A _3349_/B _3349_/C _3348_/Y VGND VGND VPWR VPWR _3396_/A sky130_fd_sc_hd__or4b_1
XFILLER_98_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6137_ _7069_/Q _6283_/A2 _6290_/B1 _7024_/Q _6136_/X VGND VGND VPWR VPWR _6143_/C
+ sky130_fd_sc_hd__a221o_1
XTAP_671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1011 _4007_/X VGND VGND VPWR VPWR _6454_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1022 _7011_/Q VGND VGND VPWR VPWR _5462_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1033 _5153_/X VGND VGND VPWR VPWR _6743_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1044 _6867_/Q VGND VGND VPWR VPWR _5300_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_73_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6068_ _6068_/A _6068_/B _6068_/C _6067_/Y VGND VGND VPWR VPWR _6068_/X sky130_fd_sc_hd__or4b_1
XFILLER_45_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1055 _5390_/X VGND VGND VPWR VPWR _6947_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_73_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1066 _6834_/Q VGND VGND VPWR VPWR _5263_/A0 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1077 _7006_/Q VGND VGND VPWR VPWR _5456_/A0 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1088 _5521_/X VGND VGND VPWR VPWR _7063_/D sky130_fd_sc_hd__dlygate4sd3_1
X_5019_ _5019_/A _5019_/B VGND VGND VPWR VPWR _5019_/Y sky130_fd_sc_hd__nand2_1
XTAP_2505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1099 _6755_/Q VGND VGND VPWR VPWR _5169_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_206 _5515_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_217 _3952_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_454 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_167_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_127_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_182_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_182_668 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_387 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_571 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_189_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_189_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_172_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_145_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5370_ hold41/X _5511_/B VGND VGND VPWR VPWR hold42/A sky130_fd_sc_hd__and2_4
XFILLER_59_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4321_ _4321_/A _5187_/B VGND VGND VPWR VPWR _4326_/S sky130_fd_sc_hd__and2_2
XFILLER_153_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_113_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_114_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7040_ _7073_/CLK _7040_/D fanout499/X VGND VGND VPWR VPWR _7040_/Q sky130_fd_sc_hd__dfstp_2
X_4252_ hold415/X _5523_/A1 _4254_/S VGND VGND VPWR VPWR _4252_/X sky130_fd_sc_hd__mux2_1
XFILLER_113_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3203_ _6925_/Q VGND VGND VPWR VPWR _3203_/Y sky130_fd_sc_hd__inv_2
XFILLER_113_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4183_ _3747_/Y _4183_/A1 _4189_/S VGND VGND VPWR VPWR _6592_/D sky130_fd_sc_hd__mux2_1
XFILLER_79_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_354 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_527 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6824_ _7050_/CLK _6824_/D fanout515/X VGND VGND VPWR VPWR _6824_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_35_295 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_435 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_479 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6755_ _6769_/CLK _6755_/D _6399_/A VGND VGND VPWR VPWR _6755_/Q sky130_fd_sc_hd__dfrtp_1
X_3967_ hold21/X hold67/X _6624_/Q VGND VGND VPWR VPWR hold68/A sky130_fd_sc_hd__mux2_1
XFILLER_50_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5706_ _6836_/Q _5928_/A2 _5651_/X _6796_/Q VGND VGND VPWR VPWR _5706_/X sky130_fd_sc_hd__a22o_1
XFILLER_149_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6686_ _6686_/CLK _6686_/D fanout492/X VGND VGND VPWR VPWR _6686_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_148_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3898_ _4335_/D _4334_/A _3177_/Y VGND VGND VPWR VPWR _3900_/C sky130_fd_sc_hd__or3b_1
XFILLER_148_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5637_ _5646_/A _5643_/B _5646_/B VGND VGND VPWR VPWR _5637_/X sky130_fd_sc_hd__and3b_4
XFILLER_164_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_148_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_163_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5568_ _6508_/Q _5643_/B VGND VGND VPWR VPWR _5573_/B sky130_fd_sc_hd__nand2_1
XFILLER_2_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold130 _7024_/Q VGND VGND VPWR VPWR hold130/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_2_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold141 hold149/X VGND VGND VPWR VPWR hold141/X sky130_fd_sc_hd__dlygate4sd3_1
X_4519_ _4943_/A _4515_/B _4517_/X _5008_/A _4774_/A VGND VGND VPWR VPWR _4519_/X
+ sky130_fd_sc_hd__o2111a_1
Xhold152 _5157_/X VGND VGND VPWR VPWR _6747_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_105_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5499_ hold157/X hold142/X _5501_/S VGND VGND VPWR VPWR _5499_/X sky130_fd_sc_hd__mux2_1
Xhold163 _6975_/Q VGND VGND VPWR VPWR hold163/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold174 _5204_/X VGND VGND VPWR VPWR _6782_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold185 _6825_/Q VGND VGND VPWR VPWR hold185/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold196 _5468_/X VGND VGND VPWR VPWR _7017_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_120_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7169_ _3939_/A1 _7169_/D _6399_/X VGND VGND VPWR VPWR _7169_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_19_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_343 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_99 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_716 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_127_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_182_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_182_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_210 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4870_ _4965_/A _5005_/A _5021_/B VGND VGND VPWR VPWR _4870_/X sky130_fd_sc_hd__o21a_1
XTAP_2880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3821_ _6416_/Q _3826_/A VGND VGND VPWR VPWR _3824_/A sky130_fd_sc_hd__and2_1
XFILLER_32_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_574 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6540_ _6697_/CLK _6540_/D fanout484/X VGND VGND VPWR VPWR _6540_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_20_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3752_ _6710_/Q _4315_/A _4309_/A _6705_/Q VGND VGND VPWR VPWR _3752_/X sky130_fd_sc_hd__a22o_1
X_6471_ _6696_/CLK _6471_/D fanout495/X VGND VGND VPWR VPWR _6471_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_185_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3683_ _3683_/A _3683_/B _3683_/C _3683_/D VGND VGND VPWR VPWR _3683_/Y sky130_fd_sc_hd__nor4_1
XFILLER_146_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5422_ hold247/X hold114/X _5423_/S VGND VGND VPWR VPWR _5422_/X sky130_fd_sc_hd__mux2_1
XFILLER_145_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput202 _3186_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[34] sky130_fd_sc_hd__buf_12
Xoutput213 _3927_/X VGND VGND VPWR VPWR mgmt_gpio_out[0] sky130_fd_sc_hd__buf_12
XFILLER_133_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput224 _7186_/X VGND VGND VPWR VPWR mgmt_gpio_out[21] sky130_fd_sc_hd__buf_12
X_5353_ _5353_/A0 _5488_/A1 _5360_/S VGND VGND VPWR VPWR _5353_/X sky130_fd_sc_hd__mux2_1
XFILLER_114_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput235 _7196_/X VGND VGND VPWR VPWR mgmt_gpio_out[31] sky130_fd_sc_hd__buf_12
XFILLER_99_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput246 _7178_/X VGND VGND VPWR VPWR mgmt_gpio_out[7] sky130_fd_sc_hd__buf_12
Xoutput257 _6745_/Q VGND VGND VPWR VPWR pll90_sel[0] sky130_fd_sc_hd__buf_12
Xoutput268 _6742_/Q VGND VGND VPWR VPWR pll_sel[0] sky130_fd_sc_hd__buf_12
X_4304_ _4304_/A0 _5488_/A1 _4308_/S VGND VGND VPWR VPWR _4304_/X sky130_fd_sc_hd__mux2_1
Xoutput279 _6419_/Q VGND VGND VPWR VPWR pll_trim[17] sky130_fd_sc_hd__buf_12
XFILLER_114_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5284_ hold763/X _5542_/A1 _5288_/S VGND VGND VPWR VPWR _5284_/X sky130_fd_sc_hd__mux2_1
XFILLER_4_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_298 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7023_ _7031_/CLK _7023_/D fanout522/X VGND VGND VPWR VPWR _7023_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_87_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4235_ hold245/X hold46/X _4236_/S VGND VGND VPWR VPWR _4235_/X sky130_fd_sc_hd__mux2_1
XFILLER_101_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4166_ _4166_/A _5187_/B VGND VGND VPWR VPWR _4171_/S sky130_fd_sc_hd__and2_2
XFILLER_110_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_549 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4097_ _4097_/A0 _5308_/A1 hold8/X VGND VGND VPWR VPWR _4097_/X sky130_fd_sc_hd__mux2_1
XFILLER_82_176 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6807_ _6881_/CLK _6807_/D fanout523/X VGND VGND VPWR VPWR _6807_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_51_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4999_ _5057_/A _4999_/B _4999_/C _4795_/X VGND VGND VPWR VPWR _5000_/A sky130_fd_sc_hd__or4b_1
XFILLER_23_298 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6738_ _7037_/CLK _6738_/D fanout484/X VGND VGND VPWR VPWR _6738_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_11_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_177_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_149_484 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6669_ _6708_/CLK _6669_/D _6401_/A VGND VGND VPWR VPWR _6669_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_109_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_151_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_164_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_132_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout440 _5543_/A1 VGND VGND VPWR VPWR _5465_/A1 sky130_fd_sc_hd__buf_4
XFILLER_59_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout451 _5532_/A1 VGND VGND VPWR VPWR _6355_/A1 sky130_fd_sc_hd__buf_6
Xfanout462 hold94/X VGND VGND VPWR VPWR hold90/A sky130_fd_sc_hd__buf_8
XFILLER_48_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout473 hold6/X VGND VGND VPWR VPWR hold7/A sky130_fd_sc_hd__buf_8
XFILLER_19_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout484 _3940_/B VGND VGND VPWR VPWR fanout484/X sky130_fd_sc_hd__buf_8
Xfanout495 fanout496/X VGND VGND VPWR VPWR fanout495/X sky130_fd_sc_hd__buf_8
XFILLER_171_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_270 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_624 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_182_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_235 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4020_ _4020_/A _6352_/B VGND VGND VPWR VPWR _4025_/S sky130_fd_sc_hd__and2_2
XFILLER_77_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5971_ _5971_/A _5971_/B VGND VGND VPWR VPWR _5971_/Y sky130_fd_sc_hd__nor2_1
XFILLER_65_699 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4922_ _5048_/A _4922_/B VGND VGND VPWR VPWR _5112_/A sky130_fd_sc_hd__nor2_1
XFILLER_45_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4853_ _4942_/C _5087_/A _4852_/Y _4531_/X VGND VGND VPWR VPWR _4853_/X sky130_fd_sc_hd__a31o_1
XFILLER_178_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3804_ _5168_/A _5183_/B VGND VGND VPWR VPWR _3804_/Y sky130_fd_sc_hd__nor2_1
XFILLER_193_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4784_ _4784_/A _4784_/B VGND VGND VPWR VPWR _4785_/B sky130_fd_sc_hd__nor2_1
XFILLER_165_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_opt_2_0_csclk _6684_/CLK VGND VGND VPWR VPWR clkbuf_opt_2_0_csclk/X sky130_fd_sc_hd__clkbuf_16
X_6523_ _6990_/CLK _6523_/D _6396_/A VGND VGND VPWR VPWR _6523_/Q sky130_fd_sc_hd__dfrtp_1
X_3735_ _6600_/Q _4190_/A _4214_/A _6620_/Q _3734_/X VGND VGND VPWR VPWR _3736_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_118_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_146_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_174_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6454_ _6559_/CLK _6454_/D _3264_/A VGND VGND VPWR VPWR _6454_/Q sky130_fd_sc_hd__dfrtp_1
X_3666_ _3666_/A _3666_/B _3666_/C _3666_/D VGND VGND VPWR VPWR _3666_/Y sky130_fd_sc_hd__nor4_1
XFILLER_146_498 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5405_ hold118/X hold27/X _5405_/S VGND VGND VPWR VPWR _5405_/X sky130_fd_sc_hd__mux2_1
X_6385_ _6401_/A _6401_/B VGND VGND VPWR VPWR _6385_/X sky130_fd_sc_hd__and2_1
X_3597_ _6445_/Q _3993_/A _4315_/A _6713_/Q VGND VGND VPWR VPWR _3597_/X sky130_fd_sc_hd__a22o_1
X_5336_ hold947/X _5531_/A1 _5342_/S VGND VGND VPWR VPWR _5336_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_235 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5267_ _5267_/A0 _5543_/A1 _5270_/S VGND VGND VPWR VPWR _5267_/X sky130_fd_sc_hd__mux2_1
X_7006_ _7083_/CLK _7006_/D fanout517/X VGND VGND VPWR VPWR _7006_/Q sky130_fd_sc_hd__dfrtp_1
X_4218_ hold65/X hold46/X _4219_/S VGND VGND VPWR VPWR hold66/A sky130_fd_sc_hd__mux2_1
X_5198_ hold116/X hold27/X _5198_/S VGND VGND VPWR VPWR _5198_/X sky130_fd_sc_hd__mux2_1
XFILLER_55_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4149_ hold249/X hold46/X _4150_/S VGND VGND VPWR VPWR _4149_/X sky130_fd_sc_hd__mux2_1
XFILLER_56_655 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_169_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_149_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_177_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_752 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_192_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_747 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_376 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3520_ _6814_/Q _5235_/A _4208_/A _6618_/Q VGND VGND VPWR VPWR _3520_/X sky130_fd_sc_hd__a22o_1
Xmax_cap404 _5639_/X VGND VGND VPWR VPWR _5926_/A2 sky130_fd_sc_hd__buf_12
XFILLER_6_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmax_cap415 _5625_/X VGND VGND VPWR VPWR _5928_/B1 sky130_fd_sc_hd__buf_12
XFILLER_115_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold707 _6989_/Q VGND VGND VPWR VPWR hold707/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold718 _5475_/X VGND VGND VPWR VPWR _7023_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold729 _6959_/Q VGND VGND VPWR VPWR hold729/X sky130_fd_sc_hd__dlygate4sd3_1
X_3451_ _6439_/Q _3984_/A _5151_/A _6747_/Q _3444_/X VGND VGND VPWR VPWR _3454_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_143_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6170_ _6825_/Q _5969_/A _6290_/A2 _7009_/Q _6169_/X VGND VGND VPWR VPWR _6177_/A
+ sky130_fd_sc_hd__a221o_1
X_3382_ _6937_/Q hold41/A _5307_/A _6881_/Q _3381_/X VGND VGND VPWR VPWR _3395_/B
+ sky130_fd_sc_hd__a221o_1
Xclkbuf_leaf_3_csclk clkbuf_3_1_0_csclk/X VGND VGND VPWR VPWR _6708_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_124_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5121_ _5121_/A _5121_/B _5121_/C VGND VGND VPWR VPWR _5121_/X sky130_fd_sc_hd__and3_1
XFILLER_69_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1407 _7140_/Q VGND VGND VPWR VPWR _6316_/A1 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1418 _6587_/Q VGND VGND VPWR VPWR _4177_/A1 sky130_fd_sc_hd__dlygate4sd3_1
X_5052_ _4719_/B _5043_/X _4972_/X _4868_/A VGND VGND VPWR VPWR _5052_/X sky130_fd_sc_hd__o211a_1
Xhold1429 _6595_/Q VGND VGND VPWR VPWR _4186_/A1 sky130_fd_sc_hd__dlygate4sd3_1
X_4003_ _4003_/A0 _5488_/A1 _4007_/S VGND VGND VPWR VPWR _4003_/X sky130_fd_sc_hd__mux2_1
XFILLER_84_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_154 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_658 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5954_ _5968_/A _5981_/A _5981_/C VGND VGND VPWR VPWR _5972_/B sky130_fd_sc_hd__and3_4
XFILLER_80_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4905_ _4401_/X _4885_/B _5105_/A _4736_/X _5100_/B VGND VGND VPWR VPWR _4906_/C
+ sky130_fd_sc_hd__o2111a_1
X_5885_ _7153_/Q _5614_/X _5630_/X _6707_/Q _5884_/X VGND VGND VPWR VPWR _5885_/Y
+ sky130_fd_sc_hd__a221oi_1
XFILLER_21_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4836_ _4692_/A _4495_/X _5026_/A _4479_/A VGND VGND VPWR VPWR _4836_/X sky130_fd_sc_hd__o22a_1
XFILLER_178_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4767_ _4911_/A _4767_/B VGND VGND VPWR VPWR _4767_/X sky130_fd_sc_hd__or2_1
X_6506_ _7124_/CLK _6506_/D fanout501/X VGND VGND VPWR VPWR _6506_/Q sky130_fd_sc_hd__dfstp_1
X_3718_ _6631_/Q _4231_/A _4261_/A _6666_/Q _3717_/X VGND VGND VPWR VPWR _3726_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_146_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4698_ _4713_/A _4717_/B VGND VGND VPWR VPWR _4714_/A sky130_fd_sc_hd__nor2_1
XFILLER_134_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_161_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6437_ _7034_/CLK _6437_/D fanout488/X VGND VGND VPWR VPWR _6437_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_146_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3649_ _6662_/Q _4255_/A _4267_/A _6672_/Q _3634_/X VGND VGND VPWR VPWR _3667_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_134_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_47 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6368_ _6400_/A _6401_/B VGND VGND VPWR VPWR _6368_/X sky130_fd_sc_hd__and2_1
XFILLER_115_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_88_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5319_ hold335/X _5541_/A1 hold84/A VGND VGND VPWR VPWR _5319_/X sky130_fd_sc_hd__mux2_1
XFILLER_102_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6299_ _6549_/Q _6299_/A2 _5974_/B _6569_/Q VGND VGND VPWR VPWR _6299_/X sky130_fd_sc_hd__a22o_1
Xhold12 hold2/X VGND VGND VPWR VPWR hold12/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_48_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold23 hold23/A VGND VGND VPWR VPWR hold23/X sky130_fd_sc_hd__buf_12
XFILLER_102_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_599 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold34 hold34/A VGND VGND VPWR VPWR hold34/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold45 hold45/A VGND VGND VPWR VPWR hold45/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold56 hold56/A VGND VGND VPWR VPWR hold56/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_29_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold67 hold67/A VGND VGND VPWR VPWR hold67/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_75_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold78 hold78/A VGND VGND VPWR VPWR hold78/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_91_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold89 hold93/X VGND VGND VPWR VPWR hold94/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_90_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_219 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_189_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_207 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_177_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_9 _3339_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_165_582 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_193_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_112_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_168 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5670_ _3182_/Y _5646_/A _5667_/B VGND VGND VPWR VPWR _5670_/Y sky130_fd_sc_hd__a21oi_1
XTAP_1091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_341 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_187_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4621_ _4622_/A _4965_/A VGND VGND VPWR VPWR _4854_/B sky130_fd_sc_hd__nor2_1
XFILLER_30_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4552_ _4622_/A _5043_/B VGND VGND VPWR VPWR _4854_/A sky130_fd_sc_hd__nor2_2
Xhold504 _3983_/X VGND VGND VPWR VPWR _6433_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold515 _6459_/Q VGND VGND VPWR VPWR hold515/X sky130_fd_sc_hd__dlygate4sd3_1
X_3503_ _3503_/A _5183_/B VGND VGND VPWR VPWR _4002_/A sky130_fd_sc_hd__nor2_8
Xhold526 _3979_/X VGND VGND VPWR VPWR _6429_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4483_ _4596_/B _4793_/A VGND VGND VPWR VPWR _4988_/A sky130_fd_sc_hd__nand2_8
XFILLER_116_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold537 _7050_/Q VGND VGND VPWR VPWR hold537/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_171_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold548 _4319_/X VGND VGND VPWR VPWR _6713_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6222_ _6651_/Q _5972_/A _5969_/C _6711_/Q _6221_/X VGND VGND VPWR VPWR _6227_/B
+ sky130_fd_sc_hd__a221o_1
Xhold559 _6681_/Q VGND VGND VPWR VPWR hold559/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_319 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3434_ _6732_/Q _3433_/X _3685_/S VGND VGND VPWR VPWR _3434_/X sky130_fd_sc_hd__mux2_1
XFILLER_143_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6153_ _6792_/Q _6004_/B _6143_/X _6152_/X _5610_/A VGND VGND VPWR VPWR _6153_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_124_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3365_ _6913_/Q _5343_/A _5235_/A _6817_/Q VGND VGND VPWR VPWR _3365_/X sky130_fd_sc_hd__a22o_1
XTAP_842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5104_ _4692_/A _4828_/A _4615_/X _4683_/B _4503_/D VGND VGND VPWR VPWR _5105_/C
+ sky130_fd_sc_hd__o221a_1
XTAP_864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1204 _4316_/X VGND VGND VPWR VPWR _6710_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6084_ _6910_/Q _5972_/A _5974_/B _6830_/Q VGND VGND VPWR VPWR _6084_/X sky130_fd_sc_hd__a22o_1
XTAP_886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1215 _6455_/Q VGND VGND VPWR VPWR _4009_/A0 sky130_fd_sc_hd__dlygate4sd3_1
X_3296_ hold39/X hold74/X hold51/X VGND VGND VPWR VPWR _3719_/A sky130_fd_sc_hd__or3b_4
Xhold1226 _5227_/X VGND VGND VPWR VPWR _6802_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1237 _6655_/Q VGND VGND VPWR VPWR _4250_/A0 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1248 _3960_/X VGND VGND VPWR VPWR _6418_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_57_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5035_ _5121_/A _5089_/B _5035_/C _5087_/D VGND VGND VPWR VPWR _5037_/C sky130_fd_sc_hd__and4_1
Xhold1259 _6660_/Q VGND VGND VPWR VPWR _4256_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_66_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6986_ _7067_/CLK _6986_/D fanout513/X VGND VGND VPWR VPWR _6986_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_81_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5937_ _5978_/B _5981_/B _5981_/C VGND VGND VPWR VPWR _5937_/X sky130_fd_sc_hd__and3_4
XFILLER_179_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5868_ _6647_/Q _5918_/A2 _5645_/X _7036_/Q VGND VGND VPWR VPWR _5868_/X sky130_fd_sc_hd__a22o_1
X_4819_ _4819_/A _5108_/A _4819_/C VGND VGND VPWR VPWR _4820_/B sky130_fd_sc_hd__and3_1
X_5799_ _6792_/Q _5667_/X _5790_/X _5798_/X _5610_/A VGND VGND VPWR VPWR _5799_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_31_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_262 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_490 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput102 wb_adr_i[12] VGND VGND VPWR VPWR _4335_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_76_503 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput113 wb_adr_i[22] VGND VGND VPWR VPWR _3891_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_0_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_163_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput124 wb_adr_i[3] VGND VGND VPWR VPWR _4746_/A sky130_fd_sc_hd__buf_2
XFILLER_193_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput135 wb_dat_i[12] VGND VGND VPWR VPWR _6336_/B1 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput146 wb_dat_i[22] VGND VGND VPWR VPWR _6342_/A2 sky130_fd_sc_hd__clkbuf_1
Xinput157 wb_dat_i[3] VGND VGND VPWR VPWR _6333_/B1 sky130_fd_sc_hd__clkbuf_1
XFILLER_48_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput168 wb_sel_i[3] VGND VGND VPWR VPWR _6320_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_56_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_189_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_110 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_165_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_363 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_83_csclk _6661_/CLK VGND VGND VPWR VPWR _6711_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_94_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6840_ _7050_/CLK _6840_/D fanout515/X VGND VGND VPWR VPWR _6840_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_63_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6771_ _7082_/CLK hold91/X fanout520/X VGND VGND VPWR VPWR _7190_/A sky130_fd_sc_hd__dfrtp_1
X_3983_ hold503/X _5519_/A1 _3983_/S VGND VGND VPWR VPWR _3983_/X sky130_fd_sc_hd__mux2_1
XFILLER_22_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_447 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5722_ _6925_/Q _5633_/X _5720_/X _5721_/X VGND VGND VPWR VPWR _5722_/X sky130_fd_sc_hd__a211o_1
XFILLER_31_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5653_ _6858_/Q _5631_/X _5647_/X _7026_/Q _5652_/X VGND VGND VPWR VPWR _5653_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_176_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_175_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4604_ _4678_/A _4713_/A VGND VGND VPWR VPWR _4973_/A sky130_fd_sc_hd__or2_4
X_5584_ _5609_/B _5964_/A VGND VGND VPWR VPWR _5593_/A sky130_fd_sc_hd__nor2_1
XFILLER_175_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_36_csclk clkbuf_3_7_0_csclk/X VGND VGND VPWR VPWR _6527_/CLK sky130_fd_sc_hd__clkbuf_16
Xhold301 _7062_/Q VGND VGND VPWR VPWR hold301/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4535_ _4535_/A _4944_/B VGND VGND VPWR VPWR _4536_/A sky130_fd_sc_hd__and2_1
Xhold312 _5274_/X VGND VGND VPWR VPWR _6844_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold323 _6860_/Q VGND VGND VPWR VPWR hold323/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold334 _5523_/X VGND VGND VPWR VPWR _7065_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold345 _7068_/Q VGND VGND VPWR VPWR hold345/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_132_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4466_ _4965_/A _5022_/B VGND VGND VPWR VPWR _4525_/A sky130_fd_sc_hd__nor2_1
Xhold356 _5346_/X VGND VGND VPWR VPWR _6908_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold367 _7073_/Q VGND VGND VPWR VPWR hold367/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_117_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold378 _5445_/X VGND VGND VPWR VPWR _6996_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold389 _6438_/Q VGND VGND VPWR VPWR hold389/X sky130_fd_sc_hd__dlygate4sd3_1
X_6205_ _6205_/A1 _6305_/A2 _6203_/X _6204_/X VGND VGND VPWR VPWR _7127_/D sky130_fd_sc_hd__o22a_1
XFILLER_171_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3417_ _5179_/B _3403_/X _3412_/X _3414_/X _3416_/X VGND VGND VPWR VPWR _3433_/C
+ sky130_fd_sc_hd__a2111o_2
X_7185_ _7185_/A VGND VGND VPWR VPWR _7185_/X sky130_fd_sc_hd__clkbuf_1
X_4397_ _4545_/A _4564_/A _4564_/B _4397_/D VGND VGND VPWR VPWR _4535_/A sky130_fd_sc_hd__and4_2
XFILLER_131_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6136_ _7085_/Q _6294_/A2 _5981_/X _6936_/Q VGND VGND VPWR VPWR _6136_/X sky130_fd_sc_hd__a22o_1
XTAP_661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3348_ _3348_/A _3348_/B VGND VGND VPWR VPWR _3348_/Y sky130_fd_sc_hd__nor2_1
XTAP_672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1001 _4210_/X VGND VGND VPWR VPWR _6615_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1012 _6626_/Q VGND VGND VPWR VPWR _4227_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1023 _5462_/X VGND VGND VPWR VPWR _7011_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1034 _6841_/Q VGND VGND VPWR VPWR _5270_/A0 sky130_fd_sc_hd__dlygate4sd3_1
X_6067_ _6067_/A _6067_/B VGND VGND VPWR VPWR _6067_/Y sky130_fd_sc_hd__nor2_1
Xhold1045 _5300_/X VGND VGND VPWR VPWR _6867_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3279_ hold72/X _4882_/B2 _6624_/Q VGND VGND VPWR VPWR hold73/A sky130_fd_sc_hd__mux2_1
Xhold1056 _6818_/Q VGND VGND VPWR VPWR _5245_/A0 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1067 _5263_/X VGND VGND VPWR VPWR _6834_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_45_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5018_ _5018_/A _5135_/C _5018_/C VGND VGND VPWR VPWR _5019_/B sky130_fd_sc_hd__and3_1
XFILLER_73_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_100_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1078 _5456_/X VGND VGND VPWR VPWR _7006_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1089 _6680_/Q VGND VGND VPWR VPWR _4280_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_207 hold8/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_218 _5537_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6969_ _6969_/CLK _6969_/D fanout506/X VGND VGND VPWR VPWR _6969_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_41_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_460 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_346 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_158_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_182_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_530 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_135_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_190_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold890 _5408_/X VGND VGND VPWR VPWR _6963_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_3_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_190_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_190_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_399 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_202 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_173_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_173_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_173_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_145_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_403 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4320_ hold445/X _5534_/A1 _4320_/S VGND VGND VPWR VPWR _4320_/X sky130_fd_sc_hd__mux2_1
XFILLER_126_574 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_736 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4251_ hold563/X _4299_/A1 _4254_/S VGND VGND VPWR VPWR _4251_/X sky130_fd_sc_hd__mux2_1
XFILLER_87_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_141_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_577 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3202_ _6933_/Q VGND VGND VPWR VPWR _3202_/Y sky130_fd_sc_hd__inv_2
XFILLER_141_599 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4182_ _3816_/X _4182_/A1 _4189_/S VGND VGND VPWR VPWR _6591_/D sky130_fd_sc_hd__mux2_1
XFILLER_79_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6823_ _7060_/CLK _6823_/D fanout521/X VGND VGND VPWR VPWR _6823_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_168_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6754_ _7076_/CLK _6754_/D fanout502/X VGND VGND VPWR VPWR _6754_/Q sky130_fd_sc_hd__dfrtp_4
X_3966_ hold541/X _5491_/A1 _3974_/S VGND VGND VPWR VPWR _3966_/X sky130_fd_sc_hd__mux2_1
X_5705_ _6988_/Q _5622_/X _5624_/X _6828_/Q VGND VGND VPWR VPWR _5705_/X sky130_fd_sc_hd__a22o_1
X_6685_ _6708_/CLK _6685_/D fanout492/X VGND VGND VPWR VPWR _6685_/Q sky130_fd_sc_hd__dfrtp_4
X_3897_ _4336_/A _4336_/B _4335_/B _3896_/Y VGND VGND VPWR VPWR _3900_/B sky130_fd_sc_hd__or4b_1
X_5636_ _5646_/A _5643_/B _5648_/C VGND VGND VPWR VPWR _5636_/X sky130_fd_sc_hd__and3b_4
XFILLER_148_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_163_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5567_ _7093_/Q _7092_/Q VGND VGND VPWR VPWR _5643_/B sky130_fd_sc_hd__nor2_4
XFILLER_117_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold120 _6883_/Q VGND VGND VPWR VPWR hold120/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_191_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4518_ _4692_/A _4581_/A VGND VGND VPWR VPWR _5008_/A sky130_fd_sc_hd__or2_1
Xhold131 _5476_/X VGND VGND VPWR VPWR _7024_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold142 hold142/A VGND VGND VPWR VPWR hold142/X sky130_fd_sc_hd__clkbuf_16
Xhold153 _6423_/Q VGND VGND VPWR VPWR hold153/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5498_ _5498_/A0 _5543_/A1 _5501_/S VGND VGND VPWR VPWR _5498_/X sky130_fd_sc_hd__mux2_1
XFILLER_132_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold164 _5421_/X VGND VGND VPWR VPWR _6975_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold175 _7144_/Q VGND VGND VPWR VPWR hold175/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold186 _5252_/X VGND VGND VPWR VPWR _6825_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4449_ _4449_/A _4449_/B _4449_/C VGND VGND VPWR VPWR _4632_/A sky130_fd_sc_hd__and3_1
Xhold197 _6797_/Q VGND VGND VPWR VPWR hold197/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_120_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_36 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7168_ _3939_/A1 _7168_/D _6398_/X VGND VGND VPWR VPWR _7168_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_86_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6119_ _6919_/Q _6288_/A2 _5969_/C _7044_/Q VGND VGND VPWR VPWR _6119_/X sky130_fd_sc_hd__a22o_2
XTAP_480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7099_ _7131_/CLK _7099_/D fanout502/X VGND VGND VPWR VPWR _7099_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_86_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_347 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_712 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_636 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_96_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_491 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_188 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3820_ _6487_/Q _3819_/B _6415_/Q VGND VGND VPWR VPWR _3826_/A sky130_fd_sc_hd__o21a_1
XFILLER_32_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3751_ _6794_/Q _5217_/A _4014_/A _6460_/Q _3750_/X VGND VGND VPWR VPWR _3754_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_185_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6470_ _6696_/CLK _6470_/D fanout495/X VGND VGND VPWR VPWR _6470_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_71_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3682_ _7041_/Q _5493_/A _5478_/A _7028_/Q _3681_/X VGND VGND VPWR VPWR _3683_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_145_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5421_ hold163/X hold142/X _5423_/S VGND VGND VPWR VPWR _5421_/X sky130_fd_sc_hd__mux2_1
XFILLER_146_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_161_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_161_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput203 _3916_/X VGND VGND VPWR VPWR mgmt_gpio_oeb[35] sky130_fd_sc_hd__buf_12
X_5352_ _5352_/A _5529_/B VGND VGND VPWR VPWR _5360_/S sky130_fd_sc_hd__and2_4
Xoutput214 _3920_/X VGND VGND VPWR VPWR mgmt_gpio_out[10] sky130_fd_sc_hd__buf_12
XFILLER_114_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput225 _7187_/X VGND VGND VPWR VPWR mgmt_gpio_out[22] sky130_fd_sc_hd__buf_12
Xoutput236 _3917_/X VGND VGND VPWR VPWR mgmt_gpio_out[32] sky130_fd_sc_hd__buf_12
Xoutput247 _3922_/X VGND VGND VPWR VPWR mgmt_gpio_out[8] sky130_fd_sc_hd__buf_12
XFILLER_99_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4303_ _4303_/A _6352_/B VGND VGND VPWR VPWR _4308_/S sky130_fd_sc_hd__and2_2
Xoutput258 _6746_/Q VGND VGND VPWR VPWR pll90_sel[1] sky130_fd_sc_hd__buf_12
XFILLER_141_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput269 _6743_/Q VGND VGND VPWR VPWR pll_sel[1] sky130_fd_sc_hd__buf_12
X_5283_ _5283_/A0 hold3/X _5288_/S VGND VGND VPWR VPWR _5283_/X sky130_fd_sc_hd__mux2_1
XFILLER_99_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7022_ _7022_/CLK _7022_/D fanout517/X VGND VGND VPWR VPWR _7022_/Q sky130_fd_sc_hd__dfrtp_1
X_4234_ hold319/X _5523_/A1 _4236_/S VGND VGND VPWR VPWR _4234_/X sky130_fd_sc_hd__mux2_1
XFILLER_4_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4165_ _3396_/X _4165_/A1 _4165_/S VGND VGND VPWR VPWR _6577_/D sky130_fd_sc_hd__mux2_1
XFILLER_114_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4096_ _4096_/A _5511_/B VGND VGND VPWR VPWR hold8/A sky130_fd_sc_hd__and2_4
XFILLER_24_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6806_ _6990_/CLK _6806_/D _6396_/A VGND VGND VPWR VPWR _6806_/Q sky130_fd_sc_hd__dfrtp_2
X_4998_ _4988_/A _4495_/X _4806_/X _4997_/X VGND VGND VPWR VPWR _5131_/A sky130_fd_sc_hd__o211ai_1
X_6737_ _7037_/CLK _6737_/D fanout484/X VGND VGND VPWR VPWR _6737_/Q sky130_fd_sc_hd__dfrtp_4
X_3949_ _6643_/Q _3956_/B VGND VGND VPWR VPWR _6637_/D sky130_fd_sc_hd__and2_1
XFILLER_23_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6668_ _6708_/CLK _6668_/D _6401_/A VGND VGND VPWR VPWR _6668_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_149_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5619_ _7095_/Q _7094_/Q VGND VGND VPWR VPWR _5650_/B sky130_fd_sc_hd__and2_2
X_6599_ _6630_/CLK _6599_/D fanout495/X VGND VGND VPWR VPWR _6599_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_192_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_155_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_160_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout430 hold27/X VGND VGND VPWR VPWR _5519_/A1 sky130_fd_sc_hd__buf_6
Xfanout441 _4236_/A1 VGND VGND VPWR VPWR _5543_/A1 sky130_fd_sc_hd__buf_4
Xfanout452 hold3/X VGND VGND VPWR VPWR _5532_/A1 sky130_fd_sc_hd__buf_6
Xfanout463 _5521_/A1 VGND VGND VPWR VPWR _6353_/A1 sky130_fd_sc_hd__buf_6
XFILLER_58_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout485 _3940_/B VGND VGND VPWR VPWR fanout485/X sky130_fd_sc_hd__buf_4
XFILLER_58_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout496 fanout526/X VGND VGND VPWR VPWR fanout496/X sky130_fd_sc_hd__buf_6
XFILLER_73_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_171_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_187_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_129_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_179 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_96_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_347 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5970_ _5940_/B _5979_/B _5981_/C _5948_/X _5962_/X VGND VGND VPWR VPWR _5974_/C
+ sky130_fd_sc_hd__a311o_1
XFILLER_92_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4921_ _4921_/A _5026_/A VGND VGND VPWR VPWR _4921_/Y sky130_fd_sc_hd__nand2_1
XFILLER_33_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_178_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4852_ _4418_/B _4569_/X _4851_/X VGND VGND VPWR VPWR _4852_/Y sky130_fd_sc_hd__a21oi_1
X_3803_ _7159_/Q _6404_/Q _3181_/Y VGND VGND VPWR VPWR _3803_/X sky130_fd_sc_hd__or3b_4
XFILLER_60_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4783_ _4581_/A _4921_/A _5043_/B _4719_/B VGND VGND VPWR VPWR _4818_/A sky130_fd_sc_hd__o22a_1
XFILLER_165_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_159_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6522_ _6990_/CLK _6522_/D _6396_/A VGND VGND VPWR VPWR _6522_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_20_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3734_ _6579_/Q _4166_/A _5187_/A _6769_/Q VGND VGND VPWR VPWR _3734_/X sky130_fd_sc_hd__a22o_1
XFILLER_146_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_158_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6453_ _6632_/CLK _6453_/D _3264_/A VGND VGND VPWR VPWR _6453_/Q sky130_fd_sc_hd__dfrtp_4
X_3665_ _6452_/Q _4002_/A _5487_/A _7036_/Q _3632_/X VGND VGND VPWR VPWR _3666_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_174_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_146_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5404_ hold144/X _5476_/A1 _5405_/S VGND VGND VPWR VPWR _5404_/X sky130_fd_sc_hd__mux2_1
X_6384_ _6401_/A _6401_/B VGND VGND VPWR VPWR _6384_/X sky130_fd_sc_hd__and2_1
X_3596_ _3596_/A _3596_/B _3596_/C _3595_/Y VGND VGND VPWR VPWR _3625_/C sky130_fd_sc_hd__or4b_1
XFILLER_114_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5335_ _5335_/A0 _5530_/A1 _5342_/S VGND VGND VPWR VPWR _5335_/X sky130_fd_sc_hd__mux2_1
XFILLER_88_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5266_ hold761/X _5542_/A1 _5270_/S VGND VGND VPWR VPWR _5266_/X sky130_fd_sc_hd__mux2_1
XFILLER_87_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7005_ _7082_/CLK _7005_/D fanout519/X VGND VGND VPWR VPWR _7005_/Q sky130_fd_sc_hd__dfrtp_4
X_4217_ hold829/X _5505_/A1 _4219_/S VGND VGND VPWR VPWR _4217_/X sky130_fd_sc_hd__mux2_1
X_5197_ hold138/X _5476_/A1 _5198_/S VGND VGND VPWR VPWR _5197_/X sky130_fd_sc_hd__mux2_1
XFILLER_110_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4148_ hold815/X _5505_/A1 _4150_/S VGND VGND VPWR VPWR _4148_/X sky130_fd_sc_hd__mux2_1
XFILLER_56_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_667 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_604 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4079_ _6396_/B hold75/X _4092_/S _4044_/X _5511_/B VGND VGND VPWR VPWR _4095_/S
+ sky130_fd_sc_hd__o221a_4
XFILLER_43_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_165_764 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_192_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_639 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_182_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_388 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_322 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_156_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_156_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_183_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmax_cap405 _5637_/X VGND VGND VPWR VPWR _5918_/B1 sky130_fd_sc_hd__buf_8
XFILLER_128_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmax_cap416 _5624_/X VGND VGND VPWR VPWR _5920_/A2 sky130_fd_sc_hd__buf_8
XFILLER_128_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold708 _5437_/X VGND VGND VPWR VPWR _6989_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold719 _6927_/Q VGND VGND VPWR VPWR hold719/X sky130_fd_sc_hd__dlygate4sd3_1
X_3450_ _6943_/Q _5379_/A _4096_/A _7200_/A _3443_/X VGND VGND VPWR VPWR _3461_/B
+ sky130_fd_sc_hd__a221o_1
X_3381_ _6945_/Q _5379_/A _5262_/A _6841_/Q VGND VGND VPWR VPWR _3381_/X sky130_fd_sc_hd__a22o_1
XFILLER_130_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5120_ _5120_/A _5120_/B VGND VGND VPWR VPWR _5120_/Y sky130_fd_sc_hd__nor2_1
XFILLER_34_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5051_ _4676_/B _4973_/B _5043_/X _4597_/Y _4877_/D VGND VGND VPWR VPWR _5054_/B
+ sky130_fd_sc_hd__o221a_1
Xhold1408 _6593_/Q VGND VGND VPWR VPWR _4184_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_85_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1419 _6584_/Q VGND VGND VPWR VPWR _4174_/A1 sky130_fd_sc_hd__dlygate4sd3_1
X_4002_ _4002_/A _5187_/B VGND VGND VPWR VPWR _4007_/S sky130_fd_sc_hd__and2_4
XFILLER_37_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_291 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5953_ _5959_/A _5953_/B VGND VGND VPWR VPWR _5953_/Y sky130_fd_sc_hd__nor2_8
XFILLER_40_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4904_ _4471_/B _4456_/Y _4748_/A _4703_/A _4903_/X VGND VGND VPWR VPWR _4912_/C
+ sky130_fd_sc_hd__o221a_1
X_5884_ _6580_/Q _5617_/X _5922_/A2 _6652_/Q VGND VGND VPWR VPWR _5884_/X sky130_fd_sc_hd__a22o_2
XFILLER_178_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4835_ _4495_/X _5026_/A _5135_/A VGND VGND VPWR VPWR _5132_/C sky130_fd_sc_hd__o21a_1
XFILLER_138_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_178_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4766_ _5136_/B _4766_/B _4766_/C _4766_/D VGND VGND VPWR VPWR _4770_/A sky130_fd_sc_hd__and4_1
XFILLER_119_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3717_ input12/X _3355_/Y _4014_/A _6461_/Q VGND VGND VPWR VPWR _3717_/X sky130_fd_sc_hd__a22o_1
X_6505_ _6969_/CLK _6505_/D fanout506/X VGND VGND VPWR VPWR _7178_/A sky130_fd_sc_hd__dfrtp_1
XFILLER_181_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_162_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_107_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4697_ _4717_/A _5005_/B VGND VGND VPWR VPWR _4697_/X sky130_fd_sc_hd__or2_1
XFILLER_20_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6436_ _6746_/CLK _6436_/D fanout488/X VGND VGND VPWR VPWR _6436_/Q sky130_fd_sc_hd__dfstp_2
X_3648_ _3648_/A _3648_/B _3648_/C _3647_/Y VGND VGND VPWR VPWR _3684_/A sky130_fd_sc_hd__or4b_1
XFILLER_161_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_162_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_134_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6367_ _6370_/A _6401_/B VGND VGND VPWR VPWR _6367_/X sky130_fd_sc_hd__and2_1
X_3579_ _6861_/Q _5289_/A _3577_/X _3578_/X VGND VGND VPWR VPWR _3579_/X sky130_fd_sc_hd__a211o_1
XFILLER_136_59 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5318_ hold120/X hold90/X hold84/X VGND VGND VPWR VPWR _5318_/X sky130_fd_sc_hd__mux2_1
X_6298_ _6654_/Q _5972_/A _5946_/X _6582_/Q VGND VGND VPWR VPWR _6298_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold13 hold13/A VGND VGND VPWR VPWR hold13/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold24 hold24/A VGND VGND VPWR VPWR hold24/X sky130_fd_sc_hd__dlygate4sd3_1
X_5249_ _5249_/A0 _5465_/A1 _5252_/S VGND VGND VPWR VPWR _5249_/X sky130_fd_sc_hd__mux2_1
XFILLER_29_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold35 hold35/A VGND VGND VPWR VPWR hold35/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_102_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold46 hold46/A VGND VGND VPWR VPWR hold46/X sky130_fd_sc_hd__buf_6
XFILLER_28_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold57 hold57/A VGND VGND VPWR VPWR hold57/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold68 hold68/A VGND VGND VPWR VPWR hold68/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold79 hold79/A VGND VGND VPWR VPWR hold79/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_56_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_456 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_177_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_169_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_177_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_138_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_193_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4620_ _4678_/A _4620_/B VGND VGND VPWR VPWR _4676_/B sky130_fd_sc_hd__or2_4
XFILLER_128_230 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4551_ _4596_/B _4551_/B VGND VGND VPWR VPWR _5043_/B sky130_fd_sc_hd__or2_4
XFILLER_129_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_144_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_190_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3502_ _3502_/A _3502_/B _3502_/C _3502_/D VGND VGND VPWR VPWR _3567_/B sky130_fd_sc_hd__nor4_2
Xhold505 _6559_/Q VGND VGND VPWR VPWR hold505/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold516 _4013_/X VGND VGND VPWR VPWR _6459_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4482_ _4622_/A _4921_/A VGND VGND VPWR VPWR _4915_/A sky130_fd_sc_hd__or2_1
Xhold527 _6515_/Q VGND VGND VPWR VPWR hold527/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold538 _5506_/X VGND VGND VPWR VPWR _7050_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6221_ _6481_/Q _5953_/Y _5955_/X _6716_/Q VGND VGND VPWR VPWR _6221_/X sky130_fd_sc_hd__a22o_1
Xhold549 _6543_/Q VGND VGND VPWR VPWR hold549/X sky130_fd_sc_hd__dlygate4sd3_1
X_3433_ _3433_/A _3433_/B _3433_/C _3432_/Y VGND VGND VPWR VPWR _3433_/X sky130_fd_sc_hd__or4b_4
XFILLER_116_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_171_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6152_ _6152_/A _6152_/B _6152_/C _6004_/B VGND VGND VPWR VPWR _6152_/X sky130_fd_sc_hd__or4b_1
XTAP_821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3364_ _3523_/A _3391_/B VGND VGND VPWR VPWR _5235_/A sky130_fd_sc_hd__nor2_8
XFILLER_106_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5103_ _4721_/B _5005_/B _4734_/X _4906_/A _5018_/A VGND VGND VPWR VPWR _5106_/C
+ sky130_fd_sc_hd__o2111a_1
XTAP_854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_0__1162_ _3567_/Y VGND VGND VPWR VPWR clkbuf_0__1162_/X sky130_fd_sc_hd__clkbuf_16
X_6083_ _7051_/Q _5975_/C _6285_/B1 _7014_/Q _6082_/X VGND VGND VPWR VPWR _6093_/A
+ sky130_fd_sc_hd__a221o_1
XTAP_876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1205 _6465_/Q VGND VGND VPWR VPWR _4021_/A0 sky130_fd_sc_hd__dlygate4sd3_1
X_3295_ hold73/X hold80/X VGND VGND VPWR VPWR hold74/A sky130_fd_sc_hd__or2_1
Xhold1216 _4009_/X VGND VGND VPWR VPWR _6455_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1227 _6962_/Q VGND VGND VPWR VPWR _5407_/A0 sky130_fd_sc_hd__dlygate4sd3_1
X_5034_ _4418_/B _4569_/X _4958_/C _5033_/X VGND VGND VPWR VPWR _5087_/D sky130_fd_sc_hd__a211oi_1
Xhold1238 _4250_/X VGND VGND VPWR VPWR _6655_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_38_431 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1249 _7047_/Q VGND VGND VPWR VPWR _5503_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_38_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6985_ _7074_/CLK _6985_/D fanout505/X VGND VGND VPWR VPWR _6985_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_80_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5936_ _5979_/B _5963_/C _5981_/C VGND VGND VPWR VPWR _5936_/X sky130_fd_sc_hd__and3_4
XFILLER_40_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5867_ _5867_/A1 _6305_/A2 _5865_/X _5866_/X VGND VGND VPWR VPWR _7115_/D sky130_fd_sc_hd__o22a_1
XFILLER_139_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4818_ _4818_/A _4818_/B _4818_/C _4818_/D VGND VGND VPWR VPWR _4819_/C sky130_fd_sc_hd__and4_1
X_5798_ _6808_/Q _5926_/A2 _5794_/X _5795_/X _5797_/X VGND VGND VPWR VPWR _5798_/X
+ sky130_fd_sc_hd__a2111o_4
XFILLER_166_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_193_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_147_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4749_ _4943_/B _4703_/A _4622_/A VGND VGND VPWR VPWR _4883_/C sky130_fd_sc_hd__a21o_1
XFILLER_31_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6419_ _6994_/CLK _6419_/D fanout489/X VGND VGND VPWR VPWR _6419_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_122_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_134_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_13 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_163_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput103 wb_adr_i[13] VGND VGND VPWR VPWR _4335_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_102_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput114 wb_adr_i[23] VGND VGND VPWR VPWR _3891_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_49_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput125 wb_adr_i[4] VGND VGND VPWR VPWR _4614_/A sky130_fd_sc_hd__clkbuf_4
Xinput136 wb_dat_i[13] VGND VGND VPWR VPWR _6338_/B1 sky130_fd_sc_hd__clkbuf_1
Xinput147 wb_dat_i[23] VGND VGND VPWR VPWR _6345_/A2 sky130_fd_sc_hd__clkbuf_1
XFILLER_102_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput158 wb_dat_i[4] VGND VGND VPWR VPWR _6335_/B1 sky130_fd_sc_hd__clkbuf_1
Xinput169 wb_stb_i VGND VGND VPWR VPWR _3894_/D sky130_fd_sc_hd__clkbuf_4
XFILLER_186_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_189_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_2_csclk clkbuf_3_1_0_csclk/X VGND VGND VPWR VPWR _6769_/CLK sky130_fd_sc_hd__clkbuf_16
XPHY_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_185_678 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_184_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_141_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_375 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3982_ hold269/X hold114/X _3983_/S VGND VGND VPWR VPWR _3982_/X sky130_fd_sc_hd__mux2_1
X_6770_ _7082_/CLK _6770_/D fanout520/X VGND VGND VPWR VPWR _7189_/A sky130_fd_sc_hd__dfrtp_1
XFILLER_22_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5721_ _6813_/Q _5913_/A2 _5646_/X _6997_/Q VGND VGND VPWR VPWR _5721_/X sky130_fd_sc_hd__a22o_1
XFILLER_50_459 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_175_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5652_ _6986_/Q _5622_/X _5645_/X _6442_/Q VGND VGND VPWR VPWR _5652_/X sky130_fd_sc_hd__a22o_1
XFILLER_176_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4603_ _4713_/A VGND VGND VPWR VPWR _4603_/Y sky130_fd_sc_hd__inv_2
X_5583_ _7098_/Q _7097_/Q VGND VGND VPWR VPWR _5964_/A sky130_fd_sc_hd__nand2_8
XFILLER_129_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4534_ _4534_/A _4534_/B VGND VGND VPWR VPWR _4534_/X sky130_fd_sc_hd__and2_1
XFILLER_190_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold302 _5519_/X VGND VGND VPWR VPWR _7062_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_144_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold313 _7041_/Q VGND VGND VPWR VPWR hold313/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold324 _5292_/X VGND VGND VPWR VPWR _6860_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_171_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold335 _6884_/Q VGND VGND VPWR VPWR hold335/X sky130_fd_sc_hd__dlygate4sd3_1
X_4465_ _4901_/A _4465_/B VGND VGND VPWR VPWR _5022_/B sky130_fd_sc_hd__or2_4
Xhold346 _5526_/X VGND VGND VPWR VPWR _7068_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold357 _7175_/A VGND VGND VPWR VPWR hold357/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold368 _5532_/X VGND VGND VPWR VPWR _7073_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6204_ _7126_/Q _5612_/A _5612_/B VGND VGND VPWR VPWR _6204_/X sky130_fd_sc_hd__o21a_1
X_3416_ input18/X _3355_/Y _5190_/A input59/X _3415_/X VGND VGND VPWR VPWR _3416_/X
+ sky130_fd_sc_hd__a221o_1
Xhold379 hold379/A VGND VGND VPWR VPWR hold379/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_131_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7184_ _7184_/A VGND VGND VPWR VPWR _7184_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_131_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4396_ _4390_/A _4390_/B _4391_/Y _4395_/X VGND VGND VPWR VPWR _4397_/D sky130_fd_sc_hd__o22a_1
XTAP_640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6135_ _6448_/Q _5601_/Y _5962_/X _6896_/Q _6134_/X VGND VGND VPWR VPWR _6143_/B
+ sky130_fd_sc_hd__a221o_1
X_3347_ _6985_/Q _5424_/A _3343_/Y input51/X _3346_/X VGND VGND VPWR VPWR _3348_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_100_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1002 _6481_/Q VGND VGND VPWR VPWR _4040_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1013 _4227_/X VGND VGND VPWR VPWR _6626_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1024 _6923_/Q VGND VGND VPWR VPWR _5363_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6066_ _7013_/Q _6285_/B1 _6282_/B1 _6973_/Q _6065_/X VGND VGND VPWR VPWR _6067_/B
+ sky130_fd_sc_hd__a221o_1
Xhold1035 _5270_/X VGND VGND VPWR VPWR _6841_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3278_ hold71/X hold78/X _3856_/S VGND VGND VPWR VPWR hold72/A sky130_fd_sc_hd__mux2_1
Xhold1046 _6690_/Q VGND VGND VPWR VPWR _4292_/A0 sky130_fd_sc_hd__dlygate4sd3_1
X_5017_ _5017_/A _5017_/B _5017_/C _5017_/D VGND VGND VPWR VPWR _5018_/C sky130_fd_sc_hd__and4_1
Xhold1057 _5245_/X VGND VGND VPWR VPWR _6818_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_39_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1068 _6750_/Q VGND VGND VPWR VPWR _5162_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_85_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1079 hold1548/X VGND VGND VPWR VPWR _4047_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_208 hold46/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_219 _5533_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6968_ _6969_/CLK _6968_/D fanout506/X VGND VGND VPWR VPWR _6968_/Q sky130_fd_sc_hd__dfrtp_1
X_5919_ _6679_/Q _5649_/X _5919_/B1 _6634_/Q _5918_/X VGND VGND VPWR VPWR _5919_/X
+ sky130_fd_sc_hd__a221o_1
X_6899_ _7056_/CLK _6899_/D fanout504/X VGND VGND VPWR VPWR _6899_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_139_358 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_147_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_542 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_123_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold880 _4120_/X VGND VGND VPWR VPWR _6539_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold891 _7072_/Q VGND VGND VPWR VPWR hold891/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_107_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_172 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_91_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_231 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_189_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_724 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_158_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_100 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_158_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_126_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_415 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_114_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4250_ _4250_/A0 _5308_/A1 _4254_/S VGND VGND VPWR VPWR _4250_/X sky130_fd_sc_hd__mux2_1
XFILLER_113_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3201_ _6941_/Q VGND VGND VPWR VPWR _3201_/Y sky130_fd_sc_hd__inv_2
XFILLER_141_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4181_ _6638_/Q _4181_/B VGND VGND VPWR VPWR _4189_/S sky130_fd_sc_hd__nand2_8
XFILLER_95_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_540 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6822_ _7043_/CLK _6822_/D _6396_/A VGND VGND VPWR VPWR _6822_/Q sky130_fd_sc_hd__dfrtp_2
X_6753_ _7076_/CLK _6753_/D fanout502/X VGND VGND VPWR VPWR _6753_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_50_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3965_ hold44/X hold175/X _6624_/Q VGND VGND VPWR VPWR _3965_/X sky130_fd_sc_hd__mux2_4
X_5704_ _7020_/Q _5929_/B1 _5915_/B1 _6860_/Q VGND VGND VPWR VPWR _5704_/X sky130_fd_sc_hd__a22o_1
XFILLER_188_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6684_ _6684_/CLK _6684_/D fanout510/X VGND VGND VPWR VPWR _6684_/Q sky130_fd_sc_hd__dfrtp_1
X_3896_ _4336_/C _4336_/D _4335_/A VGND VGND VPWR VPWR _3896_/Y sky130_fd_sc_hd__nor3_1
X_5635_ _6922_/Q _5633_/X _5634_/X _6938_/Q VGND VGND VPWR VPWR _5635_/X sky130_fd_sc_hd__a22o_1
XFILLER_12_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5566_ _5566_/A0 _5564_/Y _7092_/Q VGND VGND VPWR VPWR _5566_/X sky130_fd_sc_hd__mux2_1
XFILLER_117_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold110 _5280_/X VGND VGND VPWR VPWR _5288_/S sky130_fd_sc_hd__buf_8
XFILLER_163_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold121 _5318_/X VGND VGND VPWR VPWR _6883_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_117_575 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4517_ _4554_/A _4570_/B _4515_/B _4516_/X VGND VGND VPWR VPWR _4517_/X sky130_fd_sc_hd__o31a_1
Xhold132 _6856_/Q VGND VGND VPWR VPWR hold132/X sky130_fd_sc_hd__dlygate4sd3_1
X_5497_ hold751/X _5542_/A1 _5501_/S VGND VGND VPWR VPWR _5497_/X sky130_fd_sc_hd__mux2_1
Xhold143 _4118_/X VGND VGND VPWR VPWR _6537_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_105_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold154 _3970_/X VGND VGND VPWR VPWR _6423_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold165 _6691_/Q VGND VGND VPWR VPWR hold165/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold176 _3965_/X VGND VGND VPWR VPWR hold45/A sky130_fd_sc_hd__dlygate4sd3_1
X_4448_ _4448_/A _4679_/B VGND VGND VPWR VPWR _4902_/A sky130_fd_sc_hd__nand2_2
XFILLER_171_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold187 _6929_/Q VGND VGND VPWR VPWR hold187/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold198 _5221_/X VGND VGND VPWR VPWR _6797_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_132_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_144_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7167_ _7171_/CLK _7167_/D _6397_/X VGND VGND VPWR VPWR _7167_/Q sky130_fd_sc_hd__dfrtp_1
X_4379_ _4613_/C _4406_/A VGND VGND VPWR VPWR _4569_/A sky130_fd_sc_hd__nor2_2
XTAP_470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6118_ _6118_/A _6118_/B _6118_/C _6117_/Y VGND VGND VPWR VPWR _6118_/X sky130_fd_sc_hd__or4b_1
X_7098_ _7124_/CLK _7098_/D fanout502/X VGND VGND VPWR VPWR _7098_/Q sky130_fd_sc_hd__dfstp_4
XTAP_481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_464 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6049_ _6916_/Q _6288_/A2 _6270_/B1 _6932_/Q VGND VGND VPWR VPWR _6049_/X sky130_fd_sc_hd__a22o_1
XTAP_3027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_592 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_359 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_82_csclk _6661_/CLK VGND VGND VPWR VPWR _6707_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_10_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_155_648 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_185_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_20_csclk clkbuf_3_5_0_csclk/X VGND VGND VPWR VPWR _6559_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_110_239 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_35_csclk clkbuf_3_7_0_csclk/X VGND VGND VPWR VPWR _6887_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_45_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3750_ _7039_/Q _5493_/A _3361_/Y _6442_/Q VGND VGND VPWR VPWR _3750_/X sky130_fd_sc_hd__a22o_1
X_3681_ _7004_/Q _5451_/A _3433_/A _3628_/Y VGND VGND VPWR VPWR _3681_/X sky130_fd_sc_hd__a211o_1
XFILLER_158_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_145_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5420_ _5420_/A0 _5465_/A1 _5423_/S VGND VGND VPWR VPWR _5420_/X sky130_fd_sc_hd__mux2_1
XFILLER_64_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_173_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_145_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5351_ hold855/X _5537_/A1 _5351_/S VGND VGND VPWR VPWR _5351_/X sky130_fd_sc_hd__mux2_1
Xoutput204 _3915_/X VGND VGND VPWR VPWR mgmt_gpio_oeb[36] sky130_fd_sc_hd__buf_12
Xoutput215 _7179_/X VGND VGND VPWR VPWR mgmt_gpio_out[11] sky130_fd_sc_hd__buf_12
XFILLER_126_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput226 _7188_/X VGND VGND VPWR VPWR mgmt_gpio_out[23] sky130_fd_sc_hd__buf_12
Xoutput237 _3918_/X VGND VGND VPWR VPWR mgmt_gpio_out[33] sky130_fd_sc_hd__buf_12
Xoutput248 _3940_/Y VGND VGND VPWR VPWR pad_flash_clk_oeb sky130_fd_sc_hd__buf_12
X_4302_ hold575/X _6357_/A1 _4302_/S VGND VGND VPWR VPWR _4302_/X sky130_fd_sc_hd__mux2_1
Xoutput259 _6747_/Q VGND VGND VPWR VPWR pll90_sel[2] sky130_fd_sc_hd__buf_12
X_5282_ hold939/X _5531_/A1 _5288_/S VGND VGND VPWR VPWR _5282_/X sky130_fd_sc_hd__mux2_1
XFILLER_99_245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7021_ _7029_/CLK _7021_/D fanout525/X VGND VGND VPWR VPWR _7021_/Q sky130_fd_sc_hd__dfrtp_4
X_4233_ hold161/X hold90/X _4236_/S VGND VGND VPWR VPWR _4233_/X sky130_fd_sc_hd__mux2_1
XFILLER_87_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_632 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4164_ _3433_/X _4164_/A1 _4165_/S VGND VGND VPWR VPWR _6576_/D sky130_fd_sc_hd__mux2_1
XFILLER_114_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4095_ hold231/X _4094_/X _4095_/S VGND VGND VPWR VPWR _4095_/X sky130_fd_sc_hd__mux2_1
XFILLER_55_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6805_ _7054_/CLK _6805_/D fanout503/X VGND VGND VPWR VPWR _6805_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_169_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4997_ _4748_/B _4597_/Y _4932_/B VGND VGND VPWR VPWR _4997_/X sky130_fd_sc_hd__o21a_1
XFILLER_23_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6736_ _7037_/CLK _6736_/D fanout484/X VGND VGND VPWR VPWR _6736_/Q sky130_fd_sc_hd__dfstp_2
X_3948_ _3948_/A _3956_/B VGND VGND VPWR VPWR _6638_/D sky130_fd_sc_hd__and2_1
XFILLER_139_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6667_ _6708_/CLK _6667_/D _6401_/A VGND VGND VPWR VPWR _6667_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_164_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3879_ _7088_/Q _7089_/Q _7090_/Q _7091_/Q VGND VGND VPWR VPWR _3880_/B sky130_fd_sc_hd__or4bb_1
XFILLER_176_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5618_ _5646_/A _5645_/B _5646_/B VGND VGND VPWR VPWR _5618_/X sky130_fd_sc_hd__and3b_4
XFILLER_191_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6598_ _7137_/CLK _6598_/D VGND VGND VPWR VPWR _6598_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_124_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5549_ _6509_/Q _6507_/Q _6508_/Q _5612_/A VGND VGND VPWR VPWR _5558_/D sky130_fd_sc_hd__o31a_1
XFILLER_145_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_25 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout431 hold98/X VGND VGND VPWR VPWR hold27/A sky130_fd_sc_hd__buf_8
Xfanout442 _6357_/A1 VGND VGND VPWR VPWR _4236_/A1 sky130_fd_sc_hd__clkbuf_4
Xfanout453 _5523_/A1 VGND VGND VPWR VPWR _5505_/A1 sky130_fd_sc_hd__buf_6
Xfanout464 _5521_/A1 VGND VGND VPWR VPWR _5488_/A1 sky130_fd_sc_hd__buf_6
XFILLER_59_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout475 _3174_/Y VGND VGND VPWR VPWR _5610_/A sky130_fd_sc_hd__buf_12
XFILLER_86_451 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout486 _3940_/B VGND VGND VPWR VPWR fanout486/X sky130_fd_sc_hd__buf_8
XFILLER_171_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout497 fanout499/X VGND VGND VPWR VPWR fanout497/X sky130_fd_sc_hd__buf_8
XFILLER_104_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_478 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_143_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_136_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_3_6_0_wb_clk_i clkbuf_3_7_0_wb_clk_i/A VGND VGND VPWR VPWR _7150_/CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_151_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_684 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_315 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_359 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4920_ _4920_/A _4920_/B VGND VGND VPWR VPWR _4984_/C sky130_fd_sc_hd__nor2_2
X_4851_ _4922_/B _4851_/B _4850_/X VGND VGND VPWR VPWR _4851_/X sky130_fd_sc_hd__or3b_1
XTAP_2690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3802_ _3802_/A _3802_/B _3802_/C _3802_/D VGND VGND VPWR VPWR _3815_/C sky130_fd_sc_hd__nor4_2
XFILLER_159_751 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4782_ _4959_/A _4854_/A VGND VGND VPWR VPWR _5100_/B sky130_fd_sc_hd__nor2_2
X_6521_ _6711_/CLK _6521_/D fanout486/X VGND VGND VPWR VPWR _6521_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_158_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3733_ hold75/X _5183_/A VGND VGND VPWR VPWR _5187_/A sky130_fd_sc_hd__nor2_1
XFILLER_174_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6452_ _7038_/CLK _6452_/D fanout489/X VGND VGND VPWR VPWR _6452_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_174_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3664_ _6964_/Q _5406_/A _5397_/A _6956_/Q _3633_/X VGND VGND VPWR VPWR _3666_/C
+ sky130_fd_sc_hd__a221o_2
XFILLER_106_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5403_ hold729/X _5457_/A1 _5405_/S VGND VGND VPWR VPWR _5403_/X sky130_fd_sc_hd__mux2_1
X_6383_ _6401_/A _6401_/B VGND VGND VPWR VPWR _6383_/X sky130_fd_sc_hd__and2_1
X_3595_ _6909_/Q _5343_/A _4096_/A input64/X _3594_/X VGND VGND VPWR VPWR _3595_/Y
+ sky130_fd_sc_hd__a221oi_4
X_5334_ _5334_/A _5529_/B VGND VGND VPWR VPWR _5342_/S sky130_fd_sc_hd__and2_4
XFILLER_88_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5265_ hold375/X _5523_/A1 _5270_/S VGND VGND VPWR VPWR _5265_/X sky130_fd_sc_hd__mux2_1
X_7004_ _7079_/CLK _7004_/D fanout514/X VGND VGND VPWR VPWR _7004_/Q sky130_fd_sc_hd__dfrtp_1
X_4216_ hold933/X _5189_/A1 _4219_/S VGND VGND VPWR VPWR _4216_/X sky130_fd_sc_hd__mux2_1
X_5196_ hold765/X _5457_/A1 _5198_/S VGND VGND VPWR VPWR _5196_/X sky130_fd_sc_hd__mux2_1
X_4147_ hold925/X _5189_/A1 _4150_/S VGND VGND VPWR VPWR _4147_/X sky130_fd_sc_hd__mux2_1
XFILLER_95_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_679 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4078_ _4078_/A0 _4077_/X _4078_/S VGND VGND VPWR VPWR _4078_/X sky130_fd_sc_hd__mux2_1
XFILLER_55_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6719_ _7155_/CLK _6719_/D _6370_/A VGND VGND VPWR VPWR _6719_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_192_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_180_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_152_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_226 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_570 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_318 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmax_cap406 _5636_/X VGND VGND VPWR VPWR _5927_/A2 sky130_fd_sc_hd__buf_8
XFILLER_7_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmax_cap417 _5623_/X VGND VGND VPWR VPWR _5918_/A2 sky130_fd_sc_hd__buf_12
Xhold709 _6933_/Q VGND VGND VPWR VPWR hold709/X sky130_fd_sc_hd__dlygate4sd3_1
Xmax_cap428 _4223_/B VGND VGND VPWR VPWR _4222_/B sky130_fd_sc_hd__buf_2
XFILLER_109_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_143_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_143_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3380_ _3797_/A _3523_/A VGND VGND VPWR VPWR _5262_/A sky130_fd_sc_hd__nor2_8
XFILLER_124_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5050_ _5050_/A VGND VGND VPWR VPWR _5055_/C sky130_fd_sc_hd__inv_2
XFILLER_27_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1409 _6590_/Q VGND VGND VPWR VPWR _4180_/A1 sky130_fd_sc_hd__dlygate4sd3_1
X_4001_ hold913/X _5537_/A1 _4001_/S VGND VGND VPWR VPWR _4001_/X sky130_fd_sc_hd__mux2_1
XFILLER_111_378 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5952_ _5964_/A _5953_/B VGND VGND VPWR VPWR _5952_/Y sky130_fd_sc_hd__nor2_8
XFILLER_80_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4903_ _4692_/A _4965_/A _4748_/A VGND VGND VPWR VPWR _4903_/X sky130_fd_sc_hd__a21o_1
X_5883_ _6477_/Q _5620_/X _5627_/X _6557_/Q _5882_/X VGND VGND VPWR VPWR _5886_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_61_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4834_ _4513_/A _5026_/A _4515_/X VGND VGND VPWR VPWR _4834_/X sky130_fd_sc_hd__o21a_1
XFILLER_178_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4765_ _4943_/A _4479_/A _4715_/B _4394_/Y VGND VGND VPWR VPWR _4766_/D sky130_fd_sc_hd__o22a_1
XFILLER_193_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_193_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6504_ _6711_/CLK _6504_/D fanout486/X VGND VGND VPWR VPWR _6504_/Q sky130_fd_sc_hd__dfrtp_1
X_3716_ _6615_/Q _4208_/A _3715_/X _3433_/A VGND VGND VPWR VPWR _3716_/X sky130_fd_sc_hd__a211o_1
X_4696_ _4965_/B _4719_/B VGND VGND VPWR VPWR _5008_/B sky130_fd_sc_hd__or2_1
XFILLER_146_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_162_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6435_ _6746_/CLK _6435_/D fanout488/X VGND VGND VPWR VPWR _6435_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_146_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3647_ _7065_/Q _5520_/A _4014_/A _6462_/Q _3646_/X VGND VGND VPWR VPWR _3647_/Y
+ sky130_fd_sc_hd__a221oi_1
XFILLER_162_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6366_ _6400_/A _6401_/B VGND VGND VPWR VPWR _6366_/X sky130_fd_sc_hd__and2_1
X_3578_ _6602_/Q _4190_/A _4202_/A _6612_/Q _3573_/X VGND VGND VPWR VPWR _3578_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_114_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5317_ _5317_/A0 _5521_/A1 hold84/A VGND VGND VPWR VPWR _5317_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_130_632 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6297_ _6719_/Q _5955_/X _5978_/X _6699_/Q _6296_/X VGND VGND VPWR VPWR _6302_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_142_492 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold14 hold14/A VGND VGND VPWR VPWR hold14/X sky130_fd_sc_hd__dlygate4sd3_1
X_5248_ hold353/X _5515_/A1 _5252_/S VGND VGND VPWR VPWR _5248_/X sky130_fd_sc_hd__mux2_1
Xhold25 hold25/A VGND VGND VPWR VPWR hold25/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_75_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold36 hold36/A VGND VGND VPWR VPWR hold36/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_29_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold47 hold47/A VGND VGND VPWR VPWR hold47/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold58 hold58/A VGND VGND VPWR VPWR hold58/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold69 hold69/A VGND VGND VPWR VPWR hold69/X sky130_fd_sc_hd__dlygate4sd3_1
X_5179_ _5179_/A _5179_/B VGND VGND VPWR VPWR _5179_/X sky130_fd_sc_hd__or2_1
XFILLER_56_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_468 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_177_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_152_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_71 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4550_ _4746_/A _4595_/B VGND VGND VPWR VPWR _4551_/B sky130_fd_sc_hd__nand2_1
XFILLER_128_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_128_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3501_ _6878_/Q _5307_/A _4255_/A _6664_/Q _3500_/X VGND VGND VPWR VPWR _3502_/D
+ sky130_fd_sc_hd__a221o_2
Xhold506 _4144_/X VGND VGND VPWR VPWR _6559_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4481_ _4622_/A _4921_/A VGND VGND VPWR VPWR _4481_/Y sky130_fd_sc_hd__nor2_1
Xhold517 _6745_/Q VGND VGND VPWR VPWR hold517/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_143_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold528 _4091_/X VGND VGND VPWR VPWR _6515_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6220_ _6456_/Q _6291_/A2 _5952_/Y _7152_/Q _6219_/X VGND VGND VPWR VPWR _6227_/A
+ sky130_fd_sc_hd__a221o_1
Xhold539 _6623_/Q VGND VGND VPWR VPWR hold539/X sky130_fd_sc_hd__dlygate4sd3_1
X_3432_ _3432_/A _3432_/B _3432_/C _3432_/D VGND VGND VPWR VPWR _3432_/Y sky130_fd_sc_hd__nor4_1
XFILLER_143_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_143_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6151_ _6824_/Q _5969_/A _6148_/X _6150_/X VGND VGND VPWR VPWR _6152_/C sky130_fd_sc_hd__a211o_1
X_3363_ hold75/X _3525_/A VGND VGND VPWR VPWR _5343_/A sky130_fd_sc_hd__nor2_8
XTAP_811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5102_ _5102_/A _5102_/B _5102_/C VGND VGND VPWR VPWR _5102_/X sky130_fd_sc_hd__and3_1
XFILLER_97_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3294_ _3761_/A hold82/X VGND VGND VPWR VPWR _5529_/A sky130_fd_sc_hd__nor2_8
XFILLER_85_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6082_ _7030_/Q _5947_/Y _6290_/B1 _7022_/Q _6081_/X VGND VGND VPWR VPWR _6082_/X
+ sky130_fd_sc_hd__a221o_1
XTAP_866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1206 _4021_/X VGND VGND VPWR VPWR _6465_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1217 _6545_/Q VGND VGND VPWR VPWR _4128_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_85_527 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1228 _5407_/X VGND VGND VPWR VPWR _6962_/D sky130_fd_sc_hd__dlygate4sd3_1
X_5033_ _4569_/A _4573_/A _4946_/C _4930_/C VGND VGND VPWR VPWR _5033_/X sky130_fd_sc_hd__a31o_1
Xhold1239 _6826_/Q VGND VGND VPWR VPWR _5254_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_38_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_443 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_487 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6984_ _6984_/CLK _6984_/D fanout503/X VGND VGND VPWR VPWR _6984_/Q sky130_fd_sc_hd__dfrtp_4
X_5935_ _7100_/Q _7099_/Q VGND VGND VPWR VPWR _5981_/C sky130_fd_sc_hd__nor2_4
X_5866_ _7114_/Q _5612_/A _5612_/B VGND VGND VPWR VPWR _5866_/X sky130_fd_sc_hd__o21a_1
XFILLER_178_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_139_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_354 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4817_ _5065_/A _4817_/B _4817_/C _4817_/D VGND VGND VPWR VPWR _4818_/D sky130_fd_sc_hd__and4_1
X_5797_ _6848_/Q _5922_/B1 _5780_/X _5796_/X VGND VGND VPWR VPWR _5797_/X sky130_fd_sc_hd__a211o_1
XFILLER_178_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_540 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4748_ _4748_/A _4748_/B VGND VGND VPWR VPWR _4748_/X sky130_fd_sc_hd__or2_1
XFILLER_147_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_147_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4679_ _4679_/A _4679_/B VGND VGND VPWR VPWR _4679_/Y sky130_fd_sc_hd__nand2_2
X_6418_ _6994_/CLK _6418_/D fanout489/X VGND VGND VPWR VPWR _6418_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_150_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6349_ _6644_/Q _6320_/A _6348_/X VGND VGND VPWR VPWR _6349_/X sky130_fd_sc_hd__a21o_1
XFILLER_88_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_25 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_759 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput104 wb_adr_i[14] VGND VGND VPWR VPWR _4335_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_88_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput115 wb_adr_i[24] VGND VGND VPWR VPWR _3899_/C sky130_fd_sc_hd__clkbuf_1
Xinput126 wb_adr_i[5] VGND VGND VPWR VPWR _4779_/A sky130_fd_sc_hd__clkbuf_2
Xinput137 wb_dat_i[14] VGND VGND VPWR VPWR _6341_/B1 sky130_fd_sc_hd__clkbuf_1
XFILLER_88_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput148 wb_dat_i[24] VGND VGND VPWR VPWR _6324_/A2 sky130_fd_sc_hd__clkbuf_1
Xinput159 wb_dat_i[5] VGND VGND VPWR VPWR _6339_/B1 sky130_fd_sc_hd__clkbuf_1
XFILLER_102_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_179_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_188_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_370 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_153_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_571 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3981_ hold191/X hold142/X _3983_/S VGND VGND VPWR VPWR _3981_/X sky130_fd_sc_hd__mux2_1
X_5720_ _6909_/Q _5628_/X _5927_/A2 _6821_/Q VGND VGND VPWR VPWR _5720_/X sky130_fd_sc_hd__a22o_1
XFILLER_94_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_176_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5651_ _5646_/A _5651_/B _5651_/C VGND VGND VPWR VPWR _5651_/X sky130_fd_sc_hd__and3b_4
XFILLER_30_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4602_ _4609_/B _4613_/C _4614_/A VGND VGND VPWR VPWR _4713_/A sky130_fd_sc_hd__or3b_4
X_5582_ _7098_/Q _7097_/Q VGND VGND VPWR VPWR _5979_/B sky130_fd_sc_hd__and2_2
XFILLER_175_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_175_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4533_ _4640_/B _4943_/C _4588_/B VGND VGND VPWR VPWR _4534_/B sky130_fd_sc_hd__a21o_1
XFILLER_117_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold303 _6679_/Q VGND VGND VPWR VPWR hold303/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold314 _5496_/X VGND VGND VPWR VPWR _7041_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold325 _6828_/Q VGND VGND VPWR VPWR hold325/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_190_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4464_ _4894_/A _4892_/A VGND VGND VPWR VPWR _4465_/B sky130_fd_sc_hd__or2_1
Xhold336 _5319_/X VGND VGND VPWR VPWR _6884_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold347 _6901_/Q VGND VGND VPWR VPWR hold347/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_171_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold358 _4070_/X VGND VGND VPWR VPWR _6501_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6203_ _6540_/Q _6004_/B _6202_/X _5610_/A VGND VGND VPWR VPWR _6203_/X sky130_fd_sc_hd__o211a_1
XFILLER_116_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold369 _6780_/Q VGND VGND VPWR VPWR hold369/X sky130_fd_sc_hd__dlygate4sd3_1
X_3415_ _7053_/Q _5502_/A _3384_/Y input27/X VGND VGND VPWR VPWR _3415_/X sky130_fd_sc_hd__a22o_1
X_7183_ _7183_/A VGND VGND VPWR VPWR _7183_/X sky130_fd_sc_hd__clkbuf_1
X_4395_ _4409_/B _4707_/C VGND VGND VPWR VPWR _4395_/X sky130_fd_sc_hd__and2_1
XTAP_630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6134_ _6992_/Q _6286_/B1 _6300_/B1 _6880_/Q VGND VGND VPWR VPWR _6134_/X sky130_fd_sc_hd__a22o_1
XTAP_641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3346_ _6993_/Q hold34/A _5415_/A _6977_/Q VGND VGND VPWR VPWR _3346_/X sky130_fd_sc_hd__a22o_1
XTAP_652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1003 _4040_/X VGND VGND VPWR VPWR _6481_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1014 _6749_/Q VGND VGND VPWR VPWR _5160_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_85_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6065_ _6901_/Q _6296_/B1 _5981_/X _6933_/Q VGND VGND VPWR VPWR _6065_/X sky130_fd_sc_hd__a22o_1
Xhold1025 _5363_/X VGND VGND VPWR VPWR _6923_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3277_ _3328_/A hold31/X hold16/X hold58/X VGND VGND VPWR VPWR _3552_/A sky130_fd_sc_hd__or4b_4
Xhold1036 _6541_/Q VGND VGND VPWR VPWR _4123_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_100_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1047 _4292_/X VGND VGND VPWR VPWR _6690_/D sky130_fd_sc_hd__dlygate4sd3_1
X_5016_ _5016_/A _5016_/B _5016_/C VGND VGND VPWR VPWR _5135_/C sky130_fd_sc_hd__and3_1
Xhold1058 _6842_/Q VGND VGND VPWR VPWR _5272_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_38_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1069 _5162_/X VGND VGND VPWR VPWR _6750_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_26_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_209 hold90/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6967_ _7060_/CLK _6967_/D fanout521/X VGND VGND VPWR VPWR _6967_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_41_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5918_ _6649_/Q _5918_/A2 _5918_/B1 _6608_/Q VGND VGND VPWR VPWR _5918_/X sky130_fd_sc_hd__a22o_1
X_6898_ _7056_/CLK _6898_/D fanout504/X VGND VGND VPWR VPWR _6898_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_22_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5849_ _6666_/Q _5633_/X _5634_/X _6686_/Q _5848_/X VGND VGND VPWR VPWR _5850_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_179_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_135_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold870 _4034_/X VGND VGND VPWR VPWR _6476_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold881 _6479_/Q VGND VGND VPWR VPWR hold881/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold892 _5531_/X VGND VGND VPWR VPWR _7072_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_103_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_190_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_189_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_148_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_99_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_99_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_113_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3200_ _6949_/Q VGND VGND VPWR VPWR _3200_/Y sky130_fd_sc_hd__inv_2
X_4180_ _3396_/X _4180_/A1 _4180_/S VGND VGND VPWR VPWR _6590_/D sky130_fd_sc_hd__mux2_1
XFILLER_67_302 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_254 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6821_ _7060_/CLK _6821_/D fanout521/X VGND VGND VPWR VPWR _6821_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_23_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6752_ _7076_/CLK _6752_/D fanout502/X VGND VGND VPWR VPWR _6752_/Q sky130_fd_sc_hd__dfrtp_4
X_3964_ hold817/X _6355_/A1 _3974_/S VGND VGND VPWR VPWR _3964_/X sky130_fd_sc_hd__mux2_1
X_5703_ _6940_/Q _5816_/B1 _5696_/X _5698_/X _5702_/X VGND VGND VPWR VPWR _5703_/X
+ sky130_fd_sc_hd__a2111o_1
XFILLER_176_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6683_ _6683_/CLK _6683_/D fanout509/X VGND VGND VPWR VPWR _6683_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_176_432 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3895_ _3895_/A _3895_/B _3895_/C _3895_/D VGND VGND VPWR VPWR _3901_/C sky130_fd_sc_hd__and4_1
X_5634_ _5646_/A _5645_/B _5651_/B VGND VGND VPWR VPWR _5634_/X sky130_fd_sc_hd__and3_4
XFILLER_136_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5565_ _6506_/Q _6508_/Q VGND VGND VPWR VPWR _5565_/X sky130_fd_sc_hd__or2_1
XFILLER_128_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_163_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold100 _7028_/Q VGND VGND VPWR VPWR hold100/X sky130_fd_sc_hd__dlygate4sd3_1
X_4516_ _4513_/A _4943_/B _4514_/X _4515_/X _4410_/X VGND VGND VPWR VPWR _4516_/X
+ sky130_fd_sc_hd__o2111a_1
Xhold111 _5283_/X VGND VGND VPWR VPWR _6852_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold122 _7019_/Q VGND VGND VPWR VPWR hold122/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_2_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold133 _5287_/X VGND VGND VPWR VPWR _6856_/D sky130_fd_sc_hd__dlygate4sd3_1
X_5496_ hold313/X _5523_/A1 _5501_/S VGND VGND VPWR VPWR _5496_/X sky130_fd_sc_hd__mux2_1
XFILLER_105_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_587 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold144 _6960_/Q VGND VGND VPWR VPWR hold144/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_172_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold155 _6983_/Q VGND VGND VPWR VPWR hold155/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold166 _4293_/X VGND VGND VPWR VPWR _6691_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4447_ _4679_/B VGND VGND VPWR VPWR _4447_/Y sky130_fd_sc_hd__inv_2
Xhold177 _5230_/X VGND VGND VPWR VPWR _6805_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold188 _5369_/X VGND VGND VPWR VPWR _6929_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold199 hold199/A VGND VGND VPWR VPWR hold199/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_144_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7166_ net499_2/A _7166_/D _6396_/X VGND VGND VPWR VPWR hold25/A sky130_fd_sc_hd__dfrtp_1
X_4378_ _4378_/A _4542_/C VGND VGND VPWR VPWR _4406_/A sky130_fd_sc_hd__or2_1
Xclkbuf_leaf_1_csclk clkbuf_3_1_0_csclk/X VGND VGND VPWR VPWR _6686_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6117_ _6117_/A _6117_/B VGND VGND VPWR VPWR _6117_/Y sky130_fd_sc_hd__nor2_1
X_3329_ _3571_/B _5183_/A VGND VGND VPWR VPWR _5208_/A sky130_fd_sc_hd__nor2_8
XTAP_471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7097_ _7124_/CLK _7097_/D fanout501/X VGND VGND VPWR VPWR _7097_/Q sky130_fd_sc_hd__dfstp_4
XTAP_482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6048_ _7004_/Q _6290_/A2 _5962_/X _6892_/Q VGND VGND VPWR VPWR _6048_/X sky130_fd_sc_hd__a22o_1
XTAP_3006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_169_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_460 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_182_446 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_598 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_150_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_699 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_70 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_158_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_471 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3680_ _6828_/Q _5253_/A _4297_/A _6697_/Q _3679_/X VGND VGND VPWR VPWR _3683_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_118_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5350_ hold241/X hold114/X _5351_/S VGND VGND VPWR VPWR _5350_/X sky130_fd_sc_hd__mux2_1
XFILLER_57_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput205 _3914_/X VGND VGND VPWR VPWR mgmt_gpio_oeb[37] sky130_fd_sc_hd__buf_12
Xoutput216 _7180_/X VGND VGND VPWR VPWR mgmt_gpio_out[12] sky130_fd_sc_hd__buf_12
XFILLER_154_671 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput227 _7189_/X VGND VGND VPWR VPWR mgmt_gpio_out[24] sky130_fd_sc_hd__buf_12
X_4301_ hold583/X _5491_/A1 _4302_/S VGND VGND VPWR VPWR _4301_/X sky130_fd_sc_hd__mux2_1
Xoutput238 _7197_/X VGND VGND VPWR VPWR mgmt_gpio_out[34] sky130_fd_sc_hd__buf_12
Xoutput249 _3937_/X VGND VGND VPWR VPWR pad_flash_csb sky130_fd_sc_hd__buf_12
X_5281_ _5281_/A0 _5521_/A1 _5288_/S VGND VGND VPWR VPWR _5281_/X sky130_fd_sc_hd__mux2_1
XFILLER_99_257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7020_ _7022_/CLK hold20/X fanout517/X VGND VGND VPWR VPWR _7020_/Q sky130_fd_sc_hd__dfrtp_2
X_4232_ _4232_/A0 _5521_/A1 _4236_/S VGND VGND VPWR VPWR _4232_/X sky130_fd_sc_hd__mux2_1
XFILLER_101_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_611 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4163_ _3471_/X _4163_/A1 _4165_/S VGND VGND VPWR VPWR _6575_/D sky130_fd_sc_hd__mux2_1
XFILLER_83_603 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4094_ _5207_/A0 hold27/X hold76/X VGND VGND VPWR VPWR _4094_/X sky130_fd_sc_hd__mux2_1
XFILLER_55_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6804_ _6990_/CLK _6804_/D _6396_/A VGND VGND VPWR VPWR _6804_/Q sky130_fd_sc_hd__dfrtp_4
X_4996_ _4587_/A _4547_/X _4939_/C _4995_/X VGND VGND VPWR VPWR _5070_/B sky130_fd_sc_hd__o211a_1
XFILLER_23_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6735_ _7037_/CLK _6735_/D fanout485/X VGND VGND VPWR VPWR _6735_/Q sky130_fd_sc_hd__dfrtp_4
X_3947_ _6403_/Q _3947_/B VGND VGND VPWR VPWR _3947_/X sky130_fd_sc_hd__and2b_4
XFILLER_23_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6666_ _6769_/CLK _6666_/D fanout492/X VGND VGND VPWR VPWR _6666_/Q sky130_fd_sc_hd__dfrtp_1
X_3878_ _6507_/Q _5605_/A VGND VGND VPWR VPWR _3878_/Y sky130_fd_sc_hd__nand2_2
X_5617_ _5646_/A _5649_/C _5648_/C VGND VGND VPWR VPWR _5617_/X sky130_fd_sc_hd__and3b_4
X_6597_ _7137_/CLK _6597_/D VGND VGND VPWR VPWR _6597_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_191_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5548_ _5570_/A _6763_/Q _6509_/Q _3876_/X _5547_/X VGND VGND VPWR VPWR _7087_/D
+ sky130_fd_sc_hd__o311a_1
XFILLER_145_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_37 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5479_ _5479_/A0 _5530_/A1 _5486_/S VGND VGND VPWR VPWR _5479_/X sky130_fd_sc_hd__mux2_1
XFILLER_132_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_408 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout432 _5476_/A1 VGND VGND VPWR VPWR _5545_/A1 sky130_fd_sc_hd__buf_6
Xfanout443 hold23/X VGND VGND VPWR VPWR _6357_/A1 sky130_fd_sc_hd__buf_6
X_7149_ _3931_/A1 _7149_/D _4181_/B VGND VGND VPWR VPWR _7149_/Q sky130_fd_sc_hd__dfrtp_2
Xfanout454 hold3/X VGND VGND VPWR VPWR _5523_/A1 sky130_fd_sc_hd__buf_6
XFILLER_101_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout465 _5521_/A1 VGND VGND VPWR VPWR _5308_/A1 sky130_fd_sc_hd__buf_6
Xfanout476 _5923_/B VGND VGND VPWR VPWR _5667_/A sky130_fd_sc_hd__buf_4
Xfanout487 fanout526/X VGND VGND VPWR VPWR _3940_/B sky130_fd_sc_hd__clkbuf_8
XFILLER_86_463 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_240 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout498 fanout500/X VGND VGND VPWR VPWR fanout498/X sky130_fd_sc_hd__buf_8
XFILLER_58_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_104_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_167_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_155_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_118 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_527 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_161_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4850_ _5088_/B _5081_/B _5089_/A _4850_/D VGND VGND VPWR VPWR _4850_/X sky130_fd_sc_hd__and4_1
XTAP_2680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3801_ _7010_/Q _5460_/A _3984_/A _6434_/Q _3800_/X VGND VGND VPWR VPWR _3802_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_60_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4781_ _4781_/A VGND VGND VPWR VPWR _4988_/B sky130_fd_sc_hd__inv_2
XFILLER_159_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6520_ _7042_/CLK hold9/X fanout519/X VGND VGND VPWR VPWR _7197_/A sky130_fd_sc_hd__dfrtp_1
X_3732_ _6963_/Q _5406_/A _3572_/Y input96/X _3731_/X VGND VGND VPWR VPWR _3736_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_186_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_173_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6451_ _6695_/CLK _6451_/D fanout490/X VGND VGND VPWR VPWR _6451_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_146_435 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3663_ _6916_/Q _5352_/A _4237_/A _6647_/Q _3635_/X VGND VGND VPWR VPWR _3666_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_9_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5402_ _5402_/A0 _5465_/A1 _5405_/S VGND VGND VPWR VPWR _5402_/X sky130_fd_sc_hd__mux2_1
XFILLER_161_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6382_ _6401_/A _6401_/B VGND VGND VPWR VPWR _6382_/X sky130_fd_sc_hd__and2_1
X_3594_ _6563_/Q _4145_/A _4214_/A hold65/A VGND VGND VPWR VPWR _3594_/X sky130_fd_sc_hd__a22o_2
XFILLER_127_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5333_ hold911/X _5537_/A1 _5333_/S VGND VGND VPWR VPWR _5333_/X sky130_fd_sc_hd__mux2_1
XFILLER_161_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5264_ hold873/X _5531_/A1 _5270_/S VGND VGND VPWR VPWR _5264_/X sky130_fd_sc_hd__mux2_1
X_7003_ _7056_/CLK _7003_/D fanout504/X VGND VGND VPWR VPWR _7003_/Q sky130_fd_sc_hd__dfstp_1
X_4215_ _4215_/A0 _5308_/A1 _4219_/S VGND VGND VPWR VPWR _4215_/X sky130_fd_sc_hd__mux2_1
XFILLER_68_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5195_ _5195_/A0 hold23/X _5198_/S VGND VGND VPWR VPWR hold70/A sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_81_csclk _6661_/CLK VGND VGND VPWR VPWR _7037_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_68_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4146_ _4146_/A0 _5308_/A1 _4150_/S VGND VGND VPWR VPWR _4146_/X sky130_fd_sc_hd__mux2_1
XFILLER_18_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_124 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4077_ hold879/X _5537_/A1 _4077_/S VGND VGND VPWR VPWR _4077_/X sky130_fd_sc_hd__mux2_1
XFILLER_71_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_169_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4979_ _4979_/A _4979_/B _4979_/C VGND VGND VPWR VPWR _4979_/X sky130_fd_sc_hd__and3_1
X_6718_ _6718_/CLK _6718_/D fanout496/X VGND VGND VPWR VPWR _6718_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_20_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_137_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_164_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6649_ _7037_/CLK _6649_/D fanout484/X VGND VGND VPWR VPWR _6649_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_166_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_34_csclk clkbuf_3_7_0_csclk/X VGND VGND VPWR VPWR _6881_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_117_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_160_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_49_csclk _7000_/CLK VGND VGND VPWR VPWR _6945_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_47_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_582 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_360 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmax_cap407 _5634_/X VGND VGND VPWR VPWR _5816_/B1 sky130_fd_sc_hd__buf_8
Xmax_cap418 _5620_/X VGND VGND VPWR VPWR _5921_/A2 sky130_fd_sc_hd__buf_12
XFILLER_6_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_143_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_693 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_302 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4000_ hold636/X _5545_/A1 _4001_/S VGND VGND VPWR VPWR _4000_/X sky130_fd_sc_hd__mux2_1
XFILLER_93_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5951_ _5968_/A _5979_/A _5978_/B VGND VGND VPWR VPWR _5951_/X sky130_fd_sc_hd__and3_4
X_4902_ _4902_/A _4902_/B _4902_/C VGND VGND VPWR VPWR _5074_/B sky130_fd_sc_hd__and3_1
XFILLER_52_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5882_ _6606_/Q _5918_/B1 _5648_/X _6717_/Q VGND VGND VPWR VPWR _5882_/X sky130_fd_sc_hd__a22o_1
XFILLER_178_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4833_ _4515_/B _5026_/A _5008_/A VGND VGND VPWR VPWR _4833_/X sky130_fd_sc_hd__o21a_1
XFILLER_178_379 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4764_ _4965_/A _4676_/B _4752_/X _4763_/X _4506_/B VGND VGND VPWR VPWR _4766_/C
+ sky130_fd_sc_hd__o2111a_1
XFILLER_119_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6503_ _7054_/CLK _6503_/D fanout503/X VGND VGND VPWR VPWR _7177_/A sky130_fd_sc_hd__dfrtp_1
X_3715_ _6859_/Q _5289_/A _4127_/A _6546_/Q _3714_/X VGND VGND VPWR VPWR _3715_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_119_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4695_ _4965_/B _4695_/B VGND VGND VPWR VPWR _4723_/B sky130_fd_sc_hd__or2_1
X_6434_ _6746_/CLK _6434_/D fanout488/X VGND VGND VPWR VPWR _6434_/Q sky130_fd_sc_hd__dfstp_2
X_3646_ _6457_/Q _4008_/A _4309_/A _6707_/Q VGND VGND VPWR VPWR _3646_/X sky130_fd_sc_hd__a22o_2
XFILLER_162_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6365_ _6400_/A _6401_/B VGND VGND VPWR VPWR _6365_/X sky130_fd_sc_hd__and2_1
XFILLER_115_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3577_ _6885_/Q hold83/A _5307_/A _6877_/Q _3574_/X VGND VGND VPWR VPWR _3577_/X
+ sky130_fd_sc_hd__a221o_1
X_5316_ hold83/X _5538_/B VGND VGND VPWR VPWR hold84/A sky130_fd_sc_hd__and2_4
XFILLER_115_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6296_ _6629_/Q _6296_/A2 _6296_/B1 _6649_/Q VGND VGND VPWR VPWR _6296_/X sky130_fd_sc_hd__a22o_1
XFILLER_29_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5247_ hold327/X _5541_/A1 _5252_/S VGND VGND VPWR VPWR _5247_/X sky130_fd_sc_hd__mux2_1
XFILLER_88_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold15 hold15/A VGND VGND VPWR VPWR hold15/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold26 hold97/X VGND VGND VPWR VPWR hold98/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold37 hold37/A VGND VGND VPWR VPWR hold37/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_152_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold48 hold48/A VGND VGND VPWR VPWR hold48/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_130_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5178_ _5178_/A0 _5495_/A1 _5178_/S VGND VGND VPWR VPWR _5178_/X sky130_fd_sc_hd__mux2_1
Xhold59 hold59/A VGND VGND VPWR VPWR hold59/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_188_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4129_ _4129_/A0 _6354_/A1 _4132_/S VGND VGND VPWR VPWR _4129_/X sky130_fd_sc_hd__mux2_1
XFILLER_56_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_138_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_177_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_177_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_177_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_490 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_408 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_180_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_124 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_129_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3500_ _3500_/A1 _4077_/S _5511_/A _7059_/Q VGND VGND VPWR VPWR _3500_/X sky130_fd_sc_hd__a22o_2
XFILLER_128_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4480_ _4691_/A _4793_/A VGND VGND VPWR VPWR _4921_/A sky130_fd_sc_hd__nand2_8
Xhold507 _6607_/Q VGND VGND VPWR VPWR hold507/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold518 _5155_/X VGND VGND VPWR VPWR _6745_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold529 _6548_/Q VGND VGND VPWR VPWR hold529/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_183_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3431_ _3431_/A _3431_/B VGND VGND VPWR VPWR _3432_/D sky130_fd_sc_hd__or2_1
XFILLER_143_257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6150_ _6904_/Q _6296_/B1 _6294_/B1 _7045_/Q _6149_/X VGND VGND VPWR VPWR _6150_/X
+ sky130_fd_sc_hd__a221o_1
XTAP_801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3362_ input10/X _3360_/Y _3993_/A _6449_/Q _3359_/X VGND VGND VPWR VPWR _3362_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_112_611 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_97_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5101_ _5101_/A _5101_/B _5101_/C VGND VGND VPWR VPWR _5102_/C sky130_fd_sc_hd__and3_1
XTAP_834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6081_ _7083_/Q _6294_/A2 _5977_/X _6926_/Q VGND VGND VPWR VPWR _6081_/X sky130_fd_sc_hd__a22o_1
XTAP_856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3293_ hold81/X _3354_/A VGND VGND VPWR VPWR hold82/A sky130_fd_sc_hd__or2_4
XTAP_867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1207 _6748_/Q VGND VGND VPWR VPWR _5159_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_85_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5032_ _4403_/A _5021_/X _4950_/X VGND VGND VPWR VPWR _5035_/C sky130_fd_sc_hd__o21ba_1
XTAP_889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1218 _4128_/X VGND VGND VPWR VPWR _6545_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_85_539 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1229 _6619_/Q VGND VGND VPWR VPWR _4215_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_97_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_499 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6983_ _7046_/CLK _6983_/D fanout503/X VGND VGND VPWR VPWR _6983_/Q sky130_fd_sc_hd__dfrtp_4
X_5934_ _7101_/Q _7102_/Q VGND VGND VPWR VPWR _5963_/C sky130_fd_sc_hd__nor2_4
XFILLER_178_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5865_ _6541_/Q _5667_/X _5854_/X _5864_/X _5610_/A VGND VGND VPWR VPWR _5865_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_33_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4816_ _4816_/A _4816_/B _4816_/C _4816_/D VGND VGND VPWR VPWR _4817_/D sky130_fd_sc_hd__and4_1
XFILLER_21_366 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5796_ _6840_/Q _5928_/A2 _5651_/X _6800_/Q VGND VGND VPWR VPWR _5796_/X sky130_fd_sc_hd__a22o_1
XFILLER_193_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_119_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_166_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4747_ _5043_/A _4901_/B _4899_/B VGND VGND VPWR VPWR _5010_/A sky130_fd_sc_hd__a21oi_1
XFILLER_147_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4678_ _4678_/A _4965_/B VGND VGND VPWR VPWR _5005_/B sky130_fd_sc_hd__or2_4
XFILLER_162_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6417_ _7171_/CLK _6417_/D _6373_/X VGND VGND VPWR VPWR _6417_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_107_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3629_ _5183_/A _5183_/B VGND VGND VPWR VPWR _3629_/Y sky130_fd_sc_hd__nor2_2
XFILLER_1_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6348_ _6642_/Q _6318_/B _6348_/B1 _6643_/Q VGND VGND VPWR VPWR _6348_/X sky130_fd_sc_hd__a22o_1
XFILLER_115_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_37 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6279_ _7129_/Q _5612_/A _5612_/B VGND VGND VPWR VPWR _6279_/X sky130_fd_sc_hd__o21a_1
XFILLER_130_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput105 wb_adr_i[15] VGND VGND VPWR VPWR _4335_/C sky130_fd_sc_hd__clkbuf_1
Xinput116 wb_adr_i[25] VGND VGND VPWR VPWR input116/X sky130_fd_sc_hd__clkbuf_1
XFILLER_88_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput127 wb_adr_i[6] VGND VGND VPWR VPWR _4617_/B sky130_fd_sc_hd__buf_4
Xinput138 wb_dat_i[15] VGND VGND VPWR VPWR _6344_/B1 sky130_fd_sc_hd__clkbuf_1
Xinput149 wb_dat_i[25] VGND VGND VPWR VPWR _6327_/A2 sky130_fd_sc_hd__clkbuf_1
XFILLER_56_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_403 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_112_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_683 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_138_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_138_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_574 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_165_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_165_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_352 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_140_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_97_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3980_ hold393/X _5534_/A1 _3983_/S VGND VGND VPWR VPWR _3980_/X sky130_fd_sc_hd__mux2_1
XPHY_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_672 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5650_ _5667_/A _5650_/B _5651_/C VGND VGND VPWR VPWR _5650_/X sky130_fd_sc_hd__and3b_4
XFILLER_30_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_176_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_188_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4601_ _5043_/B _4962_/C VGND VGND VPWR VPWR _4862_/B sky130_fd_sc_hd__and2_1
XFILLER_30_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_175_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5581_ _5565_/X _5609_/B _7097_/Q VGND VGND VPWR VPWR _7097_/D sky130_fd_sc_hd__mux2_1
XFILLER_191_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4532_ _4587_/A _4479_/A _4586_/B _4495_/X _4629_/B VGND VGND VPWR VPWR _4534_/A
+ sky130_fd_sc_hd__a41o_1
XFILLER_191_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold304 _4278_/X VGND VGND VPWR VPWR _6679_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold315 hold315/A VGND VGND VPWR VPWR hold315/X sky130_fd_sc_hd__dlygate4sd3_1
X_4463_ _4885_/A _4456_/Y _4640_/B _4748_/A VGND VGND VPWR VPWR _4463_/X sky130_fd_sc_hd__o22a_1
XFILLER_171_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold326 _5256_/X VGND VGND VPWR VPWR _6828_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold337 _6892_/Q VGND VGND VPWR VPWR hold337/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold348 _5338_/X VGND VGND VPWR VPWR _6901_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6202_ _6202_/A _6202_/B _6202_/C _6004_/B VGND VGND VPWR VPWR _6202_/X sky130_fd_sc_hd__or4b_1
X_3414_ _6928_/Q _5361_/A _3975_/A _6432_/Q _3413_/X VGND VGND VPWR VPWR _3414_/X
+ sky130_fd_sc_hd__a221o_1
Xhold359 _7058_/Q VGND VGND VPWR VPWR hold359/X sky130_fd_sc_hd__dlygate4sd3_1
X_7182_ _7182_/A VGND VGND VPWR VPWR _7182_/X sky130_fd_sc_hd__clkbuf_1
X_4394_ _4888_/A _4592_/A _4617_/B VGND VGND VPWR VPWR _4394_/Y sky130_fd_sc_hd__nand3b_4
XTAP_620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6133_ _6808_/Q _5973_/B _5971_/A _6872_/Q _6132_/X VGND VGND VPWR VPWR _6143_/A
+ sky130_fd_sc_hd__a221o_1
XTAP_631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3345_ _3553_/A hold75/X VGND VGND VPWR VPWR _5415_/A sky130_fd_sc_hd__nor2_8
XTAP_642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1004 _6803_/Q VGND VGND VPWR VPWR _5228_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_100_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6064_ _6941_/Q _5942_/X _5972_/A _6909_/Q _6063_/X VGND VGND VPWR VPWR _6067_/A
+ sky130_fd_sc_hd__a221o_1
XTAP_686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1015 _5160_/X VGND VGND VPWR VPWR _6749_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3276_ hold16/X hold58/X VGND VGND VPWR VPWR _3291_/B sky130_fd_sc_hd__nand2b_1
Xhold1026 _6787_/Q VGND VGND VPWR VPWR _5210_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1037 _4123_/X VGND VGND VPWR VPWR _6541_/D sky130_fd_sc_hd__dlygate4sd3_1
X_5015_ _5073_/B _5074_/C _5015_/C VGND VGND VPWR VPWR _5019_/A sky130_fd_sc_hd__and3_1
XFILLER_100_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1048 _6882_/Q VGND VGND VPWR VPWR _5317_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_85_369 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1059 _5272_/X VGND VGND VPWR VPWR _6842_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_54_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_263 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6966_ _7022_/CLK hold87/X fanout517/X VGND VGND VPWR VPWR hold86/A sky130_fd_sc_hd__dfrtp_2
XFILLER_41_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5917_ _6464_/Q _5642_/X _5917_/B1 _7038_/Q VGND VGND VPWR VPWR _5917_/X sky130_fd_sc_hd__a22o_1
X_6897_ _7032_/CLK _6897_/D fanout506/X VGND VGND VPWR VPWR _6897_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_167_603 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5848_ _7152_/Q _5614_/X _5620_/X _6476_/Q VGND VGND VPWR VPWR _5848_/X sky130_fd_sc_hd__a22o_1
XFILLER_166_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_59 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5779_ _5779_/A1 _6305_/A2 _5777_/X _5778_/X VGND VGND VPWR VPWR _7111_/D sky130_fd_sc_hd__o22a_1
XFILLER_108_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_341 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold860 _5392_/X VGND VGND VPWR VPWR _6949_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_174_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold871 _6603_/Q VGND VGND VPWR VPWR hold871/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold882 _4037_/X VGND VGND VPWR VPWR _6479_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold893 hold893/A VGND VGND VPWR VPWR hold893/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_190_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_157_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_314 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6820_ _7041_/CLK _6820_/D fanout518/X VGND VGND VPWR VPWR _6820_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_35_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6751_ _7076_/CLK _6751_/D fanout502/X VGND VGND VPWR VPWR _6751_/Q sky130_fd_sc_hd__dfrtp_4
X_3963_ hold1/X hold10/X _6624_/Q VGND VGND VPWR VPWR hold11/A sky130_fd_sc_hd__mux2_1
XFILLER_149_603 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_1_1_0_wb_clk_i clkbuf_0_wb_clk_i/X VGND VGND VPWR VPWR clkbuf_1_1_1_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_8
X_5702_ _6820_/Q _5927_/A2 _5699_/X _5701_/X VGND VGND VPWR VPWR _5702_/X sky130_fd_sc_hd__a211o_1
X_6682_ _7038_/CLK _6682_/D fanout490/X VGND VGND VPWR VPWR _6682_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_31_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3894_ input123/X input122/X _3894_/C _3894_/D VGND VGND VPWR VPWR _3895_/D sky130_fd_sc_hd__and4bb_1
XFILLER_148_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5633_ _5646_/A _5651_/B _5651_/C VGND VGND VPWR VPWR _5633_/X sky130_fd_sc_hd__and3_4
XFILLER_12_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5564_ _6506_/Q _6508_/Q VGND VGND VPWR VPWR _5564_/Y sky130_fd_sc_hd__nor2_1
XFILLER_128_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4515_ _4692_/A _4515_/B VGND VGND VPWR VPWR _4515_/X sky130_fd_sc_hd__or2_1
Xhold101 _5481_/X VGND VGND VPWR VPWR _7028_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold112 hold112/A VGND VGND VPWR VPWR hold112/X sky130_fd_sc_hd__dlygate4sd3_1
X_5495_ hold953/X _5495_/A1 _5501_/S VGND VGND VPWR VPWR _5495_/X sky130_fd_sc_hd__mux2_1
Xhold123 _5471_/X VGND VGND VPWR VPWR _7019_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_144_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold134 _6528_/Q VGND VGND VPWR VPWR hold134/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold145 _5404_/X VGND VGND VPWR VPWR _6960_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold156 _5430_/X VGND VGND VPWR VPWR _6983_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4446_ _4575_/A _4789_/B VGND VGND VPWR VPWR _4679_/B sky130_fd_sc_hd__nor2_2
XFILLER_172_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold167 _7066_/Q VGND VGND VPWR VPWR hold167/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold178 _7025_/Q VGND VGND VPWR VPWR hold178/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold189 _7076_/Q VGND VGND VPWR VPWR hold189/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7165_ net499_2/A _7165_/D _6395_/X VGND VGND VPWR VPWR _7165_/Q sky130_fd_sc_hd__dfrtp_1
X_4377_ _4378_/A _4542_/C VGND VGND VPWR VPWR _4419_/B sky130_fd_sc_hd__nor2_1
XFILLER_86_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6116_ _6823_/Q _5969_/A _5975_/C _7052_/Q _6115_/X VGND VGND VPWR VPWR _6117_/B
+ sky130_fd_sc_hd__a221o_1
X_3328_ _3328_/A _3328_/B VGND VGND VPWR VPWR _5183_/A sky130_fd_sc_hd__nand2_8
X_7096_ _7131_/CLK _7096_/D fanout501/X VGND VGND VPWR VPWR _7096_/Q sky130_fd_sc_hd__dfstp_1
XTAP_461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6047_ _7073_/Q _6289_/A2 _6300_/B1 _6876_/Q _6046_/X VGND VGND VPWR VPWR _6052_/B
+ sky130_fd_sc_hd__a221o_1
X_3259_ _6485_/Q _3259_/B VGND VGND VPWR VPWR _3261_/B sky130_fd_sc_hd__nand2_1
XTAP_3007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_203 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6949_ _7083_/CLK _6949_/D fanout517/X VGND VGND VPWR VPWR _6949_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_41_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_179_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_623 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_182_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold690 _5232_/X VGND VGND VPWR VPWR _6807_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_150_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1390 _6805_/Q VGND VGND VPWR VPWR _5230_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_17_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_455 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_146_606 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_499 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput206 _3171_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[3] sky130_fd_sc_hd__buf_12
XFILLER_114_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput217 _3932_/X VGND VGND VPWR VPWR mgmt_gpio_out[13] sky130_fd_sc_hd__buf_12
X_4300_ hold837/X _6355_/A1 _4302_/S VGND VGND VPWR VPWR _4300_/X sky130_fd_sc_hd__mux2_1
XFILLER_99_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_154_683 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput228 _7190_/X VGND VGND VPWR VPWR mgmt_gpio_out[25] sky130_fd_sc_hd__buf_12
Xoutput239 _3919_/X VGND VGND VPWR VPWR mgmt_gpio_out[35] sky130_fd_sc_hd__buf_12
XFILLER_5_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5280_ _5280_/A _5529_/B VGND VGND VPWR VPWR _5280_/X sky130_fd_sc_hd__and2_4
XFILLER_99_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_385 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4231_ _4231_/A hold7/X VGND VGND VPWR VPWR _4236_/S sky130_fd_sc_hd__and2_4
XFILLER_99_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4162_ _6313_/A0 _4162_/A1 _4165_/S VGND VGND VPWR VPWR _6574_/D sky130_fd_sc_hd__mux2_1
XFILLER_67_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4093_ hold285/X _4092_/X _4095_/S VGND VGND VPWR VPWR _4093_/X sky130_fd_sc_hd__mux2_1
XFILLER_67_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_523 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6803_ _6984_/CLK _6803_/D fanout504/X VGND VGND VPWR VPWR _6803_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_23_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4995_ _4594_/X _5005_/A _4687_/B _4615_/B VGND VGND VPWR VPWR _4995_/X sky130_fd_sc_hd__o22a_1
X_6734_ _3939_/A1 _6734_/D _6386_/X VGND VGND VPWR VPWR _6734_/Q sky130_fd_sc_hd__dfrtn_1
X_3946_ _6404_/Q _3946_/B VGND VGND VPWR VPWR _3946_/X sky130_fd_sc_hd__and2b_4
XFILLER_23_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6665_ _6711_/CLK _6665_/D fanout486/X VGND VGND VPWR VPWR _6665_/Q sky130_fd_sc_hd__dfrtp_2
X_3877_ _5570_/A _6763_/Q _3876_/X VGND VGND VPWR VPWR _6506_/D sky130_fd_sc_hd__o21ai_1
XFILLER_139_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_192_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5616_ _7095_/Q _7094_/Q VGND VGND VPWR VPWR _5648_/C sky130_fd_sc_hd__and2b_2
XFILLER_191_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_136_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_192_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6596_ _7137_/CLK _6596_/D VGND VGND VPWR VPWR _6596_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_136_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5547_ _6506_/Q _3876_/A _7087_/Q VGND VGND VPWR VPWR _5547_/X sky130_fd_sc_hd__a21o_1
XFILLER_117_352 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5478_ _5478_/A _5529_/B VGND VGND VPWR VPWR _5486_/S sky130_fd_sc_hd__and2_4
XFILLER_155_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4429_ _4613_/C _4429_/B VGND VGND VPWR VPWR _4430_/C sky130_fd_sc_hd__or2_4
Xfanout422 _5610_/Y VGND VGND VPWR VPWR _5612_/B sky130_fd_sc_hd__buf_6
Xfanout433 hold113/X VGND VGND VPWR VPWR _5476_/A1 sky130_fd_sc_hd__buf_4
X_7148_ _3931_/A1 _7148_/D _4181_/B VGND VGND VPWR VPWR hold96/A sky130_fd_sc_hd__dfrtp_1
Xfanout444 hold69/X VGND VGND VPWR VPWR hold23/A sky130_fd_sc_hd__buf_12
XFILLER_59_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout455 hold3/X VGND VGND VPWR VPWR _5541_/A1 sky130_fd_sc_hd__buf_8
Xfanout466 _5521_/A1 VGND VGND VPWR VPWR _5530_/A1 sky130_fd_sc_hd__buf_6
Xfanout477 _5923_/B VGND VGND VPWR VPWR _5646_/A sky130_fd_sc_hd__buf_4
XFILLER_59_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout488 fanout489/X VGND VGND VPWR VPWR fanout488/X sky130_fd_sc_hd__buf_6
XFILLER_101_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7079_ _7079_/CLK _7079_/D fanout514/X VGND VGND VPWR VPWR _7079_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_46_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout499 fanout500/X VGND VGND VPWR VPWR fanout499/X sky130_fd_sc_hd__buf_4
XFILLER_86_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_154_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_731 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_170_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_355 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_97_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_100 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_420 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3800_ _7026_/Q _5478_/A _3360_/Y input34/X VGND VGND VPWR VPWR _3800_/X sky130_fd_sc_hd__a22o_1
XFILLER_21_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4780_ _4788_/A _4935_/A _4935_/B VGND VGND VPWR VPWR _4781_/A sky130_fd_sc_hd__nor3_1
XFILLER_20_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3731_ _6971_/Q _5415_/A _4321_/A _6716_/Q VGND VGND VPWR VPWR _3731_/X sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_0_csclk _6661_/CLK VGND VGND VPWR VPWR _7153_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_174_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6450_ _7038_/CLK _6450_/D fanout488/X VGND VGND VPWR VPWR _6450_/Q sky130_fd_sc_hd__dfrtp_2
X_3662_ _7073_/Q _5529_/A _4026_/A _6472_/Q _3639_/X VGND VGND VPWR VPWR _3666_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_173_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_146_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_609 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5401_ hold711/X _5542_/A1 _5405_/S VGND VGND VPWR VPWR _5401_/X sky130_fd_sc_hd__mux2_1
X_6381_ _6400_/A _6401_/B VGND VGND VPWR VPWR _6381_/X sky130_fd_sc_hd__and2_1
X_3593_ input55/X _5190_/A _4249_/A _6658_/Q _3575_/X VGND VGND VPWR VPWR _3596_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_173_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5332_ hold233/X hold114/X _5333_/S VGND VGND VPWR VPWR _5332_/X sky130_fd_sc_hd__mux2_1
XFILLER_126_171 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5263_ _5263_/A0 _5521_/A1 _5270_/S VGND VGND VPWR VPWR _5263_/X sky130_fd_sc_hd__mux2_1
XFILLER_87_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7002_ _7055_/CLK _7002_/D fanout504/X VGND VGND VPWR VPWR _7002_/Q sky130_fd_sc_hd__dfstp_1
X_4214_ _4214_/A hold7/X VGND VGND VPWR VPWR _4219_/S sky130_fd_sc_hd__and2_2
X_5194_ hold759/X _5542_/A1 _5198_/S VGND VGND VPWR VPWR _5194_/X sky130_fd_sc_hd__mux2_1
X_4145_ _4145_/A hold7/X VGND VGND VPWR VPWR _4150_/S sky130_fd_sc_hd__and2_2
XFILLER_28_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_434 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4076_ hold373/X _4075_/X _4078_/S VGND VGND VPWR VPWR _4076_/X sky130_fd_sc_hd__mux2_1
XFILLER_55_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_147 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_467 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4978_ _4691_/C _4576_/X _4695_/B _4962_/X VGND VGND VPWR VPWR _4978_/X sky130_fd_sc_hd__o22a_1
X_6717_ _7155_/CLK _6717_/D _6370_/A VGND VGND VPWR VPWR _6717_/Q sky130_fd_sc_hd__dfstp_4
X_3929_ _3220_/Y input2/X input1/X VGND VGND VPWR VPWR _3929_/X sky130_fd_sc_hd__mux2_4
XFILLER_177_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6648_ _7037_/CLK _6648_/D fanout484/X VGND VGND VPWR VPWR _6648_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_137_436 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_192_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6579_ _6708_/CLK _6579_/D fanout492/X VGND VGND VPWR VPWR _6579_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_124_119 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_132_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_174 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_434 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_372 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_331 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_751 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_155_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmax_cap408 _5632_/X VGND VGND VPWR VPWR _5922_/B1 sky130_fd_sc_hd__buf_6
Xmax_cap419 _5618_/X VGND VGND VPWR VPWR _5914_/A2 sky130_fd_sc_hd__buf_8
XFILLER_143_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_206 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_314 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_483 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5950_ _5981_/A _5962_/B _5963_/C VGND VGND VPWR VPWR _5950_/X sky130_fd_sc_hd__and3_4
XFILLER_46_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4901_ _4901_/A _4901_/B _4895_/B VGND VGND VPWR VPWR _4902_/C sky130_fd_sc_hd__or3b_1
XFILLER_80_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5881_ _6611_/Q _5631_/X _5647_/X _6457_/Q _5880_/X VGND VGND VPWR VPWR _5886_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_61_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4832_ _4943_/B _4988_/A VGND VGND VPWR VPWR _4832_/Y sky130_fd_sc_hd__nand2_1
XANTENNA_190 _3950_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4763_ _4763_/A _5007_/B _4763_/C VGND VGND VPWR VPWR _4763_/X sky130_fd_sc_hd__and3_1
XFILLER_159_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6502_ _6969_/CLK _6502_/D fanout506/X VGND VGND VPWR VPWR _7176_/A sky130_fd_sc_hd__dfrtp_1
X_3714_ _6419_/Q _3958_/A _4297_/A _6696_/Q VGND VGND VPWR VPWR _3714_/X sky130_fd_sc_hd__a22o_1
X_4694_ _5043_/A _4703_/B _4630_/B _4715_/B VGND VGND VPWR VPWR _4694_/X sky130_fd_sc_hd__o22a_1
XFILLER_174_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6433_ _6994_/CLK _6433_/D fanout490/X VGND VGND VPWR VPWR _6433_/Q sky130_fd_sc_hd__dfstp_2
X_3645_ input13/X _3355_/Y _5163_/A _6753_/Q _3644_/X VGND VGND VPWR VPWR _3648_/C
+ sky130_fd_sc_hd__a221o_4
XFILLER_20_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6364_ _6400_/A _6401_/B VGND VGND VPWR VPWR _6364_/X sky130_fd_sc_hd__and2_1
X_3576_ _6633_/Q _4231_/A _4208_/A _6617_/Q VGND VGND VPWR VPWR _3576_/X sky130_fd_sc_hd__a22o_1
XFILLER_136_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5315_ _5315_/A0 hold27/X _5315_/S VGND VGND VPWR VPWR hold99/A sky130_fd_sc_hd__mux2_1
X_6295_ _7038_/Q _6295_/A2 wire390/X _6608_/Q _6294_/X VGND VGND VPWR VPWR _6302_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_130_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_142_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5246_ _5246_/A0 _5531_/A1 _5252_/S VGND VGND VPWR VPWR _5246_/X sky130_fd_sc_hd__mux2_1
XFILLER_102_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold16 hold16/A VGND VGND VPWR VPWR hold16/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold27 hold27/A VGND VGND VPWR VPWR hold27/X sky130_fd_sc_hd__buf_8
Xhold38 hold38/A VGND VGND VPWR VPWR hold38/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_29_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5177_ hold251/X hold114/X _5178_/S VGND VGND VPWR VPWR _5177_/X sky130_fd_sc_hd__mux2_1
Xhold49 hold49/A VGND VGND VPWR VPWR hold49/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_84_710 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4128_ _4128_/A0 _6353_/A1 _4132_/S VGND VGND VPWR VPWR _4128_/X sky130_fd_sc_hd__mux2_1
XFILLER_56_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4059_ hold317/X _4058_/X _4061_/S VGND VGND VPWR VPWR _4059_/X sky130_fd_sc_hd__mux2_1
XFILLER_37_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_342 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_138_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_192_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_117_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_153_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_428 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_250 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_61 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_187_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_188_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_172 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_80_csclk _6661_/CLK VGND VGND VPWR VPWR _6746_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_129_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_190_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_171_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_128_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold508 _4200_/X VGND VGND VPWR VPWR _6607_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_128_288 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3430_ _6968_/Q _5406_/A _3360_/Y input9/X _3404_/X VGND VGND VPWR VPWR _3431_/B
+ sky130_fd_sc_hd__a221o_1
Xhold519 _6781_/Q VGND VGND VPWR VPWR hold519/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_143_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3361_ hold75/X _3554_/A VGND VGND VPWR VPWR _3361_/Y sky130_fd_sc_hd__nor2_8
XTAP_802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_623 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5100_ _5100_/A _5100_/B _5100_/C VGND VGND VPWR VPWR _5101_/C sky130_fd_sc_hd__and3_1
XTAP_835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6080_ _6080_/A1 _6305_/A2 _6078_/X _6079_/X VGND VGND VPWR VPWR _7122_/D sky130_fd_sc_hd__o22a_1
XFILLER_97_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3292_ hold39/X hold51/X VGND VGND VPWR VPWR _3354_/A sky130_fd_sc_hd__nand2_1
XFILLER_112_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5031_ _4947_/C _4829_/Y _4951_/X VGND VGND VPWR VPWR _5090_/A sky130_fd_sc_hd__a21oi_2
XTAP_879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1208 _5159_/X VGND VGND VPWR VPWR _6748_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_97_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1219 _6614_/Q VGND VGND VPWR VPWR _4209_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_97_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_111_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6982_ _7067_/CLK _6982_/D fanout513/X VGND VGND VPWR VPWR _6982_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_25_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5933_ _7118_/Q _6305_/A2 _5931_/X _5932_/X VGND VGND VPWR VPWR _7118_/D sky130_fd_sc_hd__o22a_1
Xclkbuf_leaf_33_csclk clkbuf_3_7_0_csclk/X VGND VGND VPWR VPWR _6999_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_33_150 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5864_ _5864_/A _5864_/B _5864_/C _5863_/Y VGND VGND VPWR VPWR _5864_/X sky130_fd_sc_hd__or4b_1
XFILLER_21_312 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4815_ _4394_/Y _4687_/B _4806_/X _5132_/B VGND VGND VPWR VPWR _4816_/D sky130_fd_sc_hd__o211a_1
XFILLER_166_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5795_ _7024_/Q _5929_/B1 _5915_/B1 _6864_/Q VGND VGND VPWR VPWR _5795_/X sky130_fd_sc_hd__a22o_1
XFILLER_21_378 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_159_380 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_48_csclk _7000_/CLK VGND VGND VPWR VPWR _7072_/CLK sky130_fd_sc_hd__clkbuf_16
X_4746_ _4746_/A _4746_/B _4557_/B VGND VGND VPWR VPWR _4746_/X sky130_fd_sc_hd__or3b_1
XFILLER_193_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_174_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_162_512 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4677_ _4707_/B _4677_/B VGND VGND VPWR VPWR _4715_/B sky130_fd_sc_hd__nand2_8
X_6416_ _7171_/CLK _6416_/D _6372_/X VGND VGND VPWR VPWR _6416_/Q sky130_fd_sc_hd__dfrtp_1
X_3628_ _3706_/B _3628_/B VGND VGND VPWR VPWR _3628_/Y sky130_fd_sc_hd__nor2_1
XFILLER_162_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6347_ _6347_/A1 _4221_/X _4222_/X _3903_/A VGND VGND VPWR VPWR _7149_/D sky130_fd_sc_hd__o211a_2
XFILLER_0_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3559_ _7030_/Q _5478_/A _5262_/A _6838_/Q _3558_/X VGND VGND VPWR VPWR _3565_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_142_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6278_ _6543_/Q _6004_/B _6268_/X _6277_/X _5610_/A VGND VGND VPWR VPWR _6278_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_163_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput106 wb_adr_i[16] VGND VGND VPWR VPWR _4334_/B sky130_fd_sc_hd__clkbuf_1
Xinput117 wb_adr_i[26] VGND VGND VPWR VPWR _3895_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_48_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_464 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput128 wb_adr_i[7] VGND VGND VPWR VPWR _4888_/A sky130_fd_sc_hd__buf_4
X_5229_ hold339/X _5523_/A1 _5234_/S VGND VGND VPWR VPWR _5229_/X sky130_fd_sc_hd__mux2_1
Xinput139 wb_dat_i[16] VGND VGND VPWR VPWR _6323_/A2 sky130_fd_sc_hd__clkbuf_1
XFILLER_57_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_183 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_172_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_90 _3943_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_534 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_141_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_180_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_2_3_0_wb_clk_i clkbuf_2_3_0_wb_clk_i/A VGND VGND VPWR VPWR clkbuf_3_7_0_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_97_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_264 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_684 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4600_ _4678_/A _4725_/B VGND VGND VPWR VPWR _4687_/B sky130_fd_sc_hd__or2_2
X_5580_ _5667_/A _5597_/B _5579_/B _5579_/Y VGND VGND VPWR VPWR _7096_/D sky130_fd_sc_hd__o31a_1
XFILLER_30_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4531_ _4435_/Y _4946_/C _6642_/Q VGND VGND VPWR VPWR _4531_/X sky130_fd_sc_hd__a21bo_1
Xhold305 _6829_/Q VGND VGND VPWR VPWR hold305/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold316 _4083_/X VGND VGND VPWR VPWR _6511_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_144_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4462_ _4471_/A _4885_/A VGND VGND VPWR VPWR _4748_/A sky130_fd_sc_hd__or2_2
Xhold327 _6820_/Q VGND VGND VPWR VPWR hold327/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold338 _5328_/X VGND VGND VPWR VPWR _6892_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6201_ _6201_/A _6201_/B _6201_/C _6200_/Y VGND VGND VPWR VPWR _6202_/C sky130_fd_sc_hd__or4b_1
XFILLER_89_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold349 _6885_/Q VGND VGND VPWR VPWR hold349/X sky130_fd_sc_hd__dlygate4sd3_1
X_3413_ _7077_/Q _5529_/A _4077_/S input69/X VGND VGND VPWR VPWR _3413_/X sky130_fd_sc_hd__a22o_2
XFILLER_144_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7181_ _7181_/A VGND VGND VPWR VPWR _7181_/X sky130_fd_sc_hd__clkbuf_1
X_4393_ _4888_/A _4613_/C _4614_/A _4617_/B VGND VGND VPWR VPWR _4707_/C sky130_fd_sc_hd__and4b_4
XTAP_610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3344_ _3719_/A hold33/X VGND VGND VPWR VPWR hold34/A sky130_fd_sc_hd__nor2_8
XFILLER_98_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6132_ _6848_/Q _5939_/X _6290_/A2 _7008_/Q _6131_/X VGND VGND VPWR VPWR _6132_/X
+ sky130_fd_sc_hd__a221o_1
XTAP_621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3275_ _6624_/Q hold15/X VGND VGND VPWR VPWR hold16/A sky130_fd_sc_hd__and2b_1
XFILLER_112_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6063_ _6997_/Q _6282_/A2 _5971_/A _6869_/Q VGND VGND VPWR VPWR _6063_/X sky130_fd_sc_hd__a22o_1
XTAP_676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1005 _5228_/X VGND VGND VPWR VPWR _6803_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1016 _6762_/Q VGND VGND VPWR VPWR _5178_/A0 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1027 _5210_/X VGND VGND VPWR VPWR _6787_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1038 _7152_/Q VGND VGND VPWR VPWR _6354_/A0 sky130_fd_sc_hd__dlygate4sd3_1
X_5014_ _5100_/C _5105_/B _5101_/A _5014_/D VGND VGND VPWR VPWR _5015_/C sky130_fd_sc_hd__and4_1
Xhold1049 _5317_/X VGND VGND VPWR VPWR _6882_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_38_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_562 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_275 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6965_ _6965_/CLK _6965_/D fanout514/X VGND VGND VPWR VPWR _6965_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_81_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5916_ _5916_/A _5916_/B VGND VGND VPWR VPWR _5916_/X sky130_fd_sc_hd__or2_1
XFILLER_22_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6896_ _7032_/CLK _6896_/D fanout506/X VGND VGND VPWR VPWR _6896_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_167_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5847_ _6471_/Q _5622_/X _5631_/X _6610_/Q _5846_/X VGND VGND VPWR VPWR _5850_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_139_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5778_ _5778_/A1 _3878_/Y _5612_/B VGND VGND VPWR VPWR _5778_/X sky130_fd_sc_hd__o21a_1
XFILLER_158_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4729_ _4960_/B _4728_/X _4222_/X _4589_/Y VGND VGND VPWR VPWR _4729_/X sky130_fd_sc_hd__a211o_1
XFILLER_175_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_707 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold850 _4284_/X VGND VGND VPWR VPWR _6684_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_174_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold861 _6462_/Q VGND VGND VPWR VPWR hold861/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold872 _4195_/X VGND VGND VPWR VPWR _6603_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold883 _6618_/Q VGND VGND VPWR VPWR hold883/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold894 _4104_/X VGND VGND VPWR VPWR _6524_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_1_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_190_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_88_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1550 _7180_/A VGND VGND VPWR VPWR hold295/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_57_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_147 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_172_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_141_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6750_ _7010_/CLK _6750_/D fanout498/X VGND VGND VPWR VPWR _6750_/Q sky130_fd_sc_hd__dfstp_2
X_3962_ _3962_/A0 _6354_/A1 _3974_/S VGND VGND VPWR VPWR _3962_/X sky130_fd_sc_hd__mux2_1
X_5701_ _6900_/Q _5623_/X _5637_/X _6852_/Q _5700_/X VGND VGND VPWR VPWR _5701_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_188_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_149_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6681_ _6696_/CLK _6681_/D fanout495/X VGND VGND VPWR VPWR _6681_/Q sky130_fd_sc_hd__dfrtp_1
X_3893_ _3893_/A _3893_/B VGND VGND VPWR VPWR _3895_/C sky130_fd_sc_hd__nor2_1
XFILLER_31_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5632_ _5646_/A _5645_/B _5648_/C VGND VGND VPWR VPWR _5632_/X sky130_fd_sc_hd__and3b_4
XFILLER_136_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_163_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5563_ _5563_/A1 _5559_/A _5562_/Y VGND VGND VPWR VPWR _5563_/X sky130_fd_sc_hd__o21a_1
XFILLER_129_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4514_ _5017_/A _4514_/B _4514_/C _4768_/C VGND VGND VPWR VPWR _4514_/X sky130_fd_sc_hd__and4_1
Xhold102 _6956_/Q VGND VGND VPWR VPWR hold102/X sky130_fd_sc_hd__dlygate4sd3_1
X_5494_ _5494_/A0 _5530_/A1 _5501_/S VGND VGND VPWR VPWR _5494_/X sky130_fd_sc_hd__mux2_1
Xhold113 hold113/A VGND VGND VPWR VPWR hold113/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_117_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold124 _6833_/Q VGND VGND VPWR VPWR hold124/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold135 _4108_/X VGND VGND VPWR VPWR _6528_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_105_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold146 _6757_/Q VGND VGND VPWR VPWR hold146/X sky130_fd_sc_hd__dlygate4sd3_1
X_4445_ _4977_/B _4721_/B VGND VGND VPWR VPWR _4789_/B sky130_fd_sc_hd__or2_4
Xhold157 _7044_/Q VGND VGND VPWR VPWR hold157/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold168 _5524_/X VGND VGND VPWR VPWR _7066_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_171_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold179 _5477_/X VGND VGND VPWR VPWR _7025_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_144_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7164_ net499_2/A _7164_/D _6394_/X VGND VGND VPWR VPWR _7164_/Q sky130_fd_sc_hd__dfrtp_1
X_4376_ _4679_/A _4554_/A _4596_/B _4614_/A VGND VGND VPWR VPWR _4542_/C sky130_fd_sc_hd__and4_2
XTAP_440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6115_ _6887_/Q _6296_/A2 _5955_/X _6967_/Q VGND VGND VPWR VPWR _6115_/X sky130_fd_sc_hd__a22o_1
XTAP_451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3327_ _6849_/Q _5271_/A _5226_/A _6809_/Q VGND VGND VPWR VPWR _3327_/X sky130_fd_sc_hd__a22o_1
XFILLER_100_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7095_ _7131_/CLK _7095_/D fanout501/X VGND VGND VPWR VPWR _7095_/Q sky130_fd_sc_hd__dfrtp_2
XTAP_462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6046_ _6940_/Q _5942_/X _5972_/B _7057_/Q VGND VGND VPWR VPWR _6046_/X sky130_fd_sc_hd__a22o_1
XFILLER_37_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3258_ _3165_/Y _3234_/C _3247_/Y _3257_/X VGND VGND VPWR VPWR _7159_/D sky130_fd_sc_hd__o31ai_1
XTAP_3008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3189_ _6445_/Q VGND VGND VPWR VPWR _3189_/Y sky130_fd_sc_hd__inv_2
XFILLER_94_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_392 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6948_ _6948_/CLK _6948_/D fanout514/X VGND VGND VPWR VPWR _6948_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_169_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6879_ _6881_/CLK _6879_/D fanout524/X VGND VGND VPWR VPWR _6879_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_139_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_167_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_108_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_108_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_162_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_162_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold680 _5537_/X VGND VGND VPWR VPWR _7078_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold691 _6865_/Q VGND VGND VPWR VPWR hold691/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_110_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1380 _6852_/Q VGND VGND VPWR VPWR _5283_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_18_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1391 _7147_/Q VGND VGND VPWR VPWR _3971_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_72_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_351 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_118_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_146_618 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput207 _3217_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[4] sky130_fd_sc_hd__buf_12
XFILLER_160_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput218 _7181_/X VGND VGND VPWR VPWR mgmt_gpio_out[16] sky130_fd_sc_hd__buf_12
Xoutput229 _7191_/X VGND VGND VPWR VPWR mgmt_gpio_out[26] sky130_fd_sc_hd__buf_12
XFILLER_154_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_397 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_194 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4230_ hold865/X _4236_/A1 _4230_/S VGND VGND VPWR VPWR _4230_/X sky130_fd_sc_hd__mux2_1
X_4161_ _3625_/X _4161_/A1 _4165_/S VGND VGND VPWR VPWR _6573_/D sky130_fd_sc_hd__mux2_1
XFILLER_67_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4092_ hold136/X _5476_/A1 _4092_/S VGND VGND VPWR VPWR _4092_/X sky130_fd_sc_hd__mux2_1
XFILLER_82_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6802_ _6978_/CLK _6802_/D fanout490/X VGND VGND VPWR VPWR _6802_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_51_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4994_ _4994_/A _4994_/B VGND VGND VPWR VPWR _5002_/B sky130_fd_sc_hd__or2_1
X_6733_ _3939_/A1 _6733_/D _6385_/X VGND VGND VPWR VPWR _6733_/Q sky130_fd_sc_hd__dfrtn_1
X_3945_ input85/X _3247_/A _6404_/Q VGND VGND VPWR VPWR _3945_/X sky130_fd_sc_hd__mux2_2
XFILLER_149_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_149_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6664_ _6699_/CLK _6664_/D fanout509/X VGND VGND VPWR VPWR _6664_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_31_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3876_ _3876_/A _3876_/B VGND VGND VPWR VPWR _3876_/X sky130_fd_sc_hd__or2_1
XFILLER_177_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5615_ _7092_/Q _7093_/Q VGND VGND VPWR VPWR _5649_/C sky130_fd_sc_hd__and2b_2
X_6595_ _7137_/CLK _6595_/D VGND VGND VPWR VPWR _6595_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_176_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_192_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5546_ hold223/X hold27/X _5546_/S VGND VGND VPWR VPWR _5546_/X sky130_fd_sc_hd__mux2_1
XFILLER_117_364 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_191_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_144_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5477_ hold178/X hold27/X hold19/X VGND VGND VPWR VPWR _5477_/X sky130_fd_sc_hd__mux2_1
XFILLER_144_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_144_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_160_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4428_ _4561_/B _4495_/B VGND VGND VPWR VPWR _4581_/A sky130_fd_sc_hd__or2_4
XFILLER_99_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_2_3__f_mgmt_gpio_in[4] clkbuf_0_mgmt_gpio_in[4]/X VGND VGND VPWR VPWR net499_2/A
+ sky130_fd_sc_hd__clkbuf_16
Xfanout423 _4575_/X VGND VGND VPWR VPWR _4748_/B sky130_fd_sc_hd__buf_6
XFILLER_58_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout434 hold113/X VGND VGND VPWR VPWR hold114/A sky130_fd_sc_hd__clkbuf_16
X_7147_ _3931_/A1 _7147_/D _4181_/B VGND VGND VPWR VPWR _7147_/Q sky130_fd_sc_hd__dfrtp_1
Xfanout445 _5533_/A1 VGND VGND VPWR VPWR _5491_/A1 sky130_fd_sc_hd__buf_8
XFILLER_101_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4359_ _4367_/B _4399_/B VGND VGND VPWR VPWR _4886_/A sky130_fd_sc_hd__nor2_1
XFILLER_86_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout456 hold12/X VGND VGND VPWR VPWR hold3/A sky130_fd_sc_hd__buf_6
Xfanout467 hold588/X VGND VGND VPWR VPWR _5521_/A1 sky130_fd_sc_hd__buf_12
Xfanout478 _7096_/Q VGND VGND VPWR VPWR _5923_/B sky130_fd_sc_hd__buf_12
XFILLER_171_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout489 fanout490/X VGND VGND VPWR VPWR fanout489/X sky130_fd_sc_hd__buf_8
X_7078_ _7078_/CLK _7078_/D fanout507/X VGND VGND VPWR VPWR _7078_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_100_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_318 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6029_ _6029_/A1 _5612_/A _5612_/B VGND VGND VPWR VPWR _6029_/X sky130_fd_sc_hd__o21a_1
XFILLER_58_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_331 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_129_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_367 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_579 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3730_ _7003_/Q _5451_/A _5179_/B _6762_/Q _3729_/X VGND VGND VPWR VPWR _3736_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_13_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_159_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_186_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3661_ _3661_/A _3661_/B _3661_/C _3660_/Y VGND VGND VPWR VPWR _3667_/C sky130_fd_sc_hd__or4b_1
XFILLER_174_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5400_ hold102/X hold3/X _5405_/S VGND VGND VPWR VPWR _5400_/X sky130_fd_sc_hd__mux2_1
XFILLER_62_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6380_ _6400_/A _6401_/B VGND VGND VPWR VPWR _6380_/X sky130_fd_sc_hd__and2_1
XFILLER_173_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3592_ _6853_/Q _3374_/Y _5253_/A _6829_/Q _3591_/X VGND VGND VPWR VPWR _3596_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_127_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5331_ hold699/X _5544_/A1 _5333_/S VGND VGND VPWR VPWR _5331_/X sky130_fd_sc_hd__mux2_1
XFILLER_126_183 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5262_ _5262_/A _5511_/B VGND VGND VPWR VPWR _5270_/S sky130_fd_sc_hd__and2_4
X_7001_ _7050_/CLK _7001_/D fanout515/X VGND VGND VPWR VPWR _7001_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_114_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4213_ hold883/X _4236_/A1 _4213_/S VGND VGND VPWR VPWR _4213_/X sky130_fd_sc_hd__mux2_1
XFILLER_68_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5193_ hold289/X _5541_/A1 _5198_/S VGND VGND VPWR VPWR _5193_/X sky130_fd_sc_hd__mux2_1
XFILLER_96_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4144_ hold505/X _6357_/A1 _4144_/S VGND VGND VPWR VPWR _4144_/X sky130_fd_sc_hd__mux2_1
XFILLER_18_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4075_ hold271/X hold114/X _4112_/B VGND VGND VPWR VPWR _4075_/X sky130_fd_sc_hd__mux2_1
XFILLER_83_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_479 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_3_4_0_csclk clkbuf_3_5_0_csclk/A VGND VGND VPWR VPWR _6684_/CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_24_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4977_ _5022_/A _4977_/B _4947_/B VGND VGND VPWR VPWR _5061_/C sky130_fd_sc_hd__or3b_1
X_6716_ _6769_/CLK _6716_/D _6399_/A VGND VGND VPWR VPWR _6716_/Q sky130_fd_sc_hd__dfrtp_4
X_3928_ _3219_/Y _7157_/Q _6396_/B VGND VGND VPWR VPWR _3928_/X sky130_fd_sc_hd__mux2_2
X_6647_ _7037_/CLK _6647_/D fanout484/X VGND VGND VPWR VPWR _6647_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_50_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3859_ _7158_/Q _3860_/S VGND VGND VPWR VPWR _3859_/Y sky130_fd_sc_hd__nor2_1
XFILLER_166_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6578_ _6686_/CLK _6578_/D fanout492/X VGND VGND VPWR VPWR _6578_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_152_407 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5529_ _5529_/A _5529_/B VGND VGND VPWR VPWR _5537_/S sky130_fd_sc_hd__and2_4
XFILLER_105_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_182_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_132_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_182_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_627 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_343 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_763 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_cap409 _5631_/X VGND VGND VPWR VPWR _5915_/B1 sky130_fd_sc_hd__buf_12
XFILLER_155_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_155_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_143_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_151_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4900_ _5022_/B _4965_/B VGND VGND VPWR VPWR _4912_/B sky130_fd_sc_hd__or2_1
X_5880_ _5667_/B _5879_/X _5644_/X _6452_/Q VGND VGND VPWR VPWR _5880_/X sky130_fd_sc_hd__a2bb2o_1
X_4831_ _4943_/B _4988_/A VGND VGND VPWR VPWR _4831_/X sky130_fd_sc_hd__and2_2
XTAP_2490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_180 _5969_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_191 _3263_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4762_ _4615_/B _4715_/B _4736_/X _4739_/Y _4761_/X VGND VGND VPWR VPWR _4763_/C
+ sky130_fd_sc_hd__o2111a_1
X_6501_ _7033_/CLK _6501_/D fanout503/X VGND VGND VPWR VPWR _7175_/A sky130_fd_sc_hd__dfrtp_1
X_3713_ _3713_/A _3713_/B _3713_/C _3713_/D VGND VGND VPWR VPWR _3747_/A sky130_fd_sc_hd__nor4_2
X_4693_ _4965_/A _4965_/B _4676_/B VGND VGND VPWR VPWR _4706_/A sky130_fd_sc_hd__a21oi_1
XFILLER_146_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6432_ _6994_/CLK _6432_/D fanout489/X VGND VGND VPWR VPWR _6432_/Q sky130_fd_sc_hd__dfstp_2
X_3644_ _7081_/Q _5538_/A _5379_/A _6940_/Q VGND VGND VPWR VPWR _3644_/X sky130_fd_sc_hd__a22o_2
XFILLER_174_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6363_ _6400_/A _6401_/B VGND VGND VPWR VPWR _6363_/X sky130_fd_sc_hd__and2_1
X_3575_ _7058_/Q _5511_/A _4267_/A _6673_/Q VGND VGND VPWR VPWR _3575_/X sky130_fd_sc_hd__a22o_1
X_5314_ hold451/X _5545_/A1 _5315_/S VGND VGND VPWR VPWR _5314_/X sky130_fd_sc_hd__mux2_1
XFILLER_115_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6294_ _6664_/Q _6294_/A2 _6294_/B1 _6714_/Q VGND VGND VPWR VPWR _6294_/X sky130_fd_sc_hd__a22o_1
XFILLER_130_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5245_ _5245_/A0 _5521_/A1 _5252_/S VGND VGND VPWR VPWR _5245_/X sky130_fd_sc_hd__mux2_1
XFILLER_114_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold17 hold32/X VGND VGND VPWR VPWR hold33/A sky130_fd_sc_hd__buf_8
XFILLER_130_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold28 hold28/A VGND VGND VPWR VPWR hold28/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_69_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5176_ hold199/X hold142/X _5178_/S VGND VGND VPWR VPWR _5176_/X sky130_fd_sc_hd__mux2_1
XFILLER_69_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold39 hold39/A VGND VGND VPWR VPWR hold39/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_152_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_571 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_722 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4127_ _4127_/A _6352_/B VGND VGND VPWR VPWR _4132_/S sky130_fd_sc_hd__and2_2
XFILLER_28_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_16 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4058_ hold221/X _5476_/A1 _4103_/B VGND VGND VPWR VPWR _4058_/X sky130_fd_sc_hd__mux2_1
XFILLER_37_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_3_5_0_wb_clk_i clkbuf_3_5_0_wb_clk_i/A VGND VGND VPWR VPWR _7140_/CLK sky130_fd_sc_hd__clkbuf_8
XPHY_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_177_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_177_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_192_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_160_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_262 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_142_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_184 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold509 _6925_/Q VGND VGND VPWR VPWR hold509/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_167_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3360_ hold82/A _5168_/A VGND VGND VPWR VPWR _3360_/Y sky130_fd_sc_hd__nor2_8
XTAP_803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3291_ _3328_/A _3291_/B hold31/X VGND VGND VPWR VPWR _3557_/A sky130_fd_sc_hd__or3b_4
XFILLER_151_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5030_ _5038_/B VGND VGND VPWR VPWR _5124_/A sky130_fd_sc_hd__clkinv_2
XTAP_869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1209 _6705_/Q VGND VGND VPWR VPWR _4310_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_53_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6981_ _6990_/CLK _6981_/D fanout513/X VGND VGND VPWR VPWR _6981_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_19_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5932_ _7117_/Q _5612_/A _5612_/B VGND VGND VPWR VPWR _5932_/X sky130_fd_sc_hd__o21a_1
XFILLER_53_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5863_ _6605_/Q _5918_/B1 _5646_/X _6481_/Q _5862_/X VGND VGND VPWR VPWR _5863_/Y
+ sky130_fd_sc_hd__a221oi_1
XFILLER_80_279 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4814_ _4678_/A _4394_/Y _5043_/B _4495_/X _4921_/A VGND VGND VPWR VPWR _4816_/C
+ sky130_fd_sc_hd__o32a_1
X_5794_ _6936_/Q _5807_/B1 _5791_/X _5793_/X VGND VGND VPWR VPWR _5794_/X sky130_fd_sc_hd__a211o_1
X_4745_ _4901_/B _4745_/B VGND VGND VPWR VPWR _4911_/B sky130_fd_sc_hd__nor2_1
XFILLER_193_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_174_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4676_ _4703_/A _4676_/B VGND VGND VPWR VPWR _4709_/A sky130_fd_sc_hd__nor2_1
XFILLER_174_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6415_ _7171_/CLK _6415_/D _6371_/X VGND VGND VPWR VPWR _6415_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_162_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3627_ _3626_/X _3627_/A1 _3749_/S VGND VGND VPWR VPWR _6730_/D sky130_fd_sc_hd__mux2_1
XFILLER_162_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6346_ _6345_/X _6346_/A1 _6346_/S VGND VGND VPWR VPWR _7148_/D sky130_fd_sc_hd__mux2_1
X_3558_ _7067_/Q _5520_/A _4291_/A _6694_/Q VGND VGND VPWR VPWR _3558_/X sky130_fd_sc_hd__a22o_1
XFILLER_1_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6277_ _6277_/A _6277_/B _6277_/C _5975_/X VGND VGND VPWR VPWR _6277_/X sky130_fd_sc_hd__or4b_2
XFILLER_102_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_130_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3489_ _3489_/A _3489_/B _3489_/C _3489_/D VGND VGND VPWR VPWR _3489_/Y sky130_fd_sc_hd__nor4_1
Xinput107 wb_adr_i[17] VGND VGND VPWR VPWR _4334_/A sky130_fd_sc_hd__clkbuf_1
Xinput118 wb_adr_i[27] VGND VGND VPWR VPWR _3893_/A sky130_fd_sc_hd__clkbuf_1
X_5228_ _5228_/A0 _5531_/A1 _5234_/S VGND VGND VPWR VPWR _5228_/X sky130_fd_sc_hd__mux2_1
Xinput129 wb_adr_i[8] VGND VGND VPWR VPWR _4336_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_69_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5159_ _5159_/A0 _5488_/A1 _5160_/S VGND VGND VPWR VPWR _5159_/X sky130_fd_sc_hd__mux2_1
XFILLER_56_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_2_1_0_csclk clkbuf_2_1_0_csclk/A VGND VGND VPWR VPWR clkbuf_3_3_0_csclk/A
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_72_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_184_148 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_80 user_clock VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_91 _3943_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_153_546 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_180_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_137_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_102_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_416 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_224 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_188_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_318 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_178_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4530_ _4590_/A _4530_/B _4561_/B VGND VGND VPWR VPWR _4946_/C sky130_fd_sc_hd__nor3_2
XFILLER_11_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold306 _5257_/X VGND VGND VPWR VPWR _6829_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4461_ _4542_/A _5025_/A VGND VGND VPWR VPWR _4640_/B sky130_fd_sc_hd__nand2_8
Xhold317 _7187_/A VGND VGND VPWR VPWR hold317/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_144_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_192 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold328 _5247_/X VGND VGND VPWR VPWR _6820_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6200_ _6200_/A _6200_/B VGND VGND VPWR VPWR _6200_/Y sky130_fd_sc_hd__nor2_1
Xhold339 _6804_/Q VGND VGND VPWR VPWR hold339/X sky130_fd_sc_hd__dlygate4sd3_1
X_3412_ _6832_/Q _5253_/A _3409_/X _3411_/X VGND VGND VPWR VPWR _3412_/X sky130_fd_sc_hd__a211o_2
X_7180_ _7180_/A VGND VGND VPWR VPWR _7180_/X sky130_fd_sc_hd__clkbuf_1
X_4392_ _4888_/A _4617_/B VGND VGND VPWR VPWR _4609_/B sky130_fd_sc_hd__nand2b_1
XFILLER_98_611 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6131_ _6944_/Q _5942_/X _6282_/B1 _6976_/Q VGND VGND VPWR VPWR _6131_/X sky130_fd_sc_hd__a22o_1
XTAP_611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3343_ _3571_/A _5183_/B VGND VGND VPWR VPWR _3343_/Y sky130_fd_sc_hd__nor2_4
XFILLER_97_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6062_ _6445_/Q _5601_/Y _6300_/B1 _6877_/Q _6061_/X VGND VGND VPWR VPWR _6068_/C
+ sky130_fd_sc_hd__a221o_1
XTAP_666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3274_ hold14/X _3856_/S _3273_/Y VGND VGND VPWR VPWR hold15/A sky130_fd_sc_hd__a21bo_1
XTAP_677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1006 _6546_/Q VGND VGND VPWR VPWR _4129_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_98_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1017 _5178_/X VGND VGND VPWR VPWR _6762_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5013_ _4692_/A _4965_/A _5022_/B VGND VGND VPWR VPWR _5014_/D sky130_fd_sc_hd__a21o_1
XTAP_699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1028 _6419_/Q VGND VGND VPWR VPWR _3962_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_85_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1039 _6354_/X VGND VGND VPWR VPWR _7152_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_38_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_287 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6964_ _7075_/CLK _6964_/D fanout505/X VGND VGND VPWR VPWR _6964_/Q sky130_fd_sc_hd__dfrtp_4
X_5915_ _6709_/Q _5915_/A2 _5915_/B1 _6613_/Q _5914_/X VGND VGND VPWR VPWR _5916_/B
+ sky130_fd_sc_hd__a221o_1
X_6895_ _6961_/CLK _6895_/D fanout521/X VGND VGND VPWR VPWR _6895_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_179_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5846_ _6696_/Q _5626_/X _5632_/X _6600_/Q VGND VGND VPWR VPWR _5846_/X sky130_fd_sc_hd__a22o_1
XFILLER_166_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5777_ _6791_/Q _5667_/X _5765_/X _5776_/X _3174_/Y VGND VGND VPWR VPWR _5777_/X
+ sky130_fd_sc_hd__o221a_2
XFILLER_166_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4728_ _4959_/C _4854_/A _4728_/C _4942_/B VGND VGND VPWR VPWR _4728_/X sky130_fd_sc_hd__or4b_1
XFILLER_135_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_147_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_108_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4659_ _5043_/B _4962_/C _4678_/A _4721_/B VGND VGND VPWR VPWR _4659_/X sky130_fd_sc_hd__a211o_1
XFILLER_174_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_162_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_600 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold840 _5454_/X VGND VGND VPWR VPWR _7004_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold851 _6866_/Q VGND VGND VPWR VPWR hold851/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_107_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold862 _4017_/X VGND VGND VPWR VPWR _6462_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_190_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold873 _6835_/Q VGND VGND VPWR VPWR hold873/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold884 _4213_/X VGND VGND VPWR VPWR _6618_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6329_ _6642_/Q _6329_/A2 _6329_/B1 _4222_/B VGND VGND VPWR VPWR _6329_/X sky130_fd_sc_hd__a22o_1
XFILLER_115_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold895 _6769_/Q VGND VGND VPWR VPWR hold895/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_76_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_284 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1540 _7176_/A VGND VGND VPWR VPWR hold630/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_29_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1551 _6511_/Q VGND VGND VPWR VPWR hold315/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_29_254 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_141_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_32_csclk clkbuf_3_7_0_csclk/X VGND VGND VPWR VPWR _7031_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_122_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_47_csclk clkbuf_3_6_0_csclk/X VGND VGND VPWR VPWR _7074_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_94_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3961_ hold88/X hold92/X _6624_/Q VGND VGND VPWR VPWR hold93/A sky130_fd_sc_hd__mux2_1
X_5700_ _6868_/Q _5625_/X _5643_/X _6884_/Q VGND VGND VPWR VPWR _5700_/X sky130_fd_sc_hd__a22o_1
XFILLER_31_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6680_ _7038_/CLK _6680_/D fanout490/X VGND VGND VPWR VPWR _6680_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_92_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3892_ _4368_/A _4544_/A VGND VGND VPWR VPWR _4449_/B sky130_fd_sc_hd__nand2_1
X_5631_ _5667_/A _5646_/B _5651_/C VGND VGND VPWR VPWR _5631_/X sky130_fd_sc_hd__and3b_4
XFILLER_148_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_176_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5562_ _7091_/Q _5559_/A _5561_/A VGND VGND VPWR VPWR _5562_/Y sky130_fd_sc_hd__a21boi_1
XFILLER_191_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4513_ _4513_/A _4549_/B VGND VGND VPWR VPWR _4768_/C sky130_fd_sc_hd__or2_1
XFILLER_191_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_144_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5493_ _5493_/A _5529_/B VGND VGND VPWR VPWR _5501_/S sky130_fd_sc_hd__and2_4
Xhold103 _5400_/X VGND VGND VPWR VPWR _6956_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_7_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold114 hold114/A VGND VGND VPWR VPWR hold114/X sky130_fd_sc_hd__clkbuf_16
Xhold125 _5261_/X VGND VGND VPWR VPWR _6833_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_144_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold136 _6784_/Q VGND VGND VPWR VPWR hold136/X sky130_fd_sc_hd__dlygate4sd3_1
X_4444_ _4617_/B _4888_/A _4614_/A _4613_/C VGND VGND VPWR VPWR _4721_/B sky130_fd_sc_hd__or4b_4
Xhold147 _5173_/X VGND VGND VPWR VPWR _6757_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold158 _5499_/X VGND VGND VPWR VPWR _7044_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold169 _6453_/Q VGND VGND VPWR VPWR hold169/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_132_549 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7163_ net499_2/A _7163_/D _6393_/X VGND VGND VPWR VPWR hold21/A sky130_fd_sc_hd__dfrtp_1
XFILLER_113_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4375_ _4614_/A _4409_/B VGND VGND VPWR VPWR _4378_/A sky130_fd_sc_hd__nor2_1
XTAP_430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6114_ _7060_/Q _5972_/B _5962_/X _6895_/Q _6113_/X VGND VGND VPWR VPWR _6117_/A
+ sky130_fd_sc_hd__a221o_1
XTAP_441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3326_ _3531_/A _3487_/A VGND VGND VPWR VPWR _5226_/A sky130_fd_sc_hd__nor2_8
XFILLER_112_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7094_ _7124_/CLK _7094_/D fanout501/X VGND VGND VPWR VPWR _7094_/Q sky130_fd_sc_hd__dfrtp_2
XTAP_452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6045_ _6964_/Q _5955_/X _6294_/B1 _7041_/Q _6044_/X VGND VGND VPWR VPWR _6052_/A
+ sky130_fd_sc_hd__a221o_1
XTAP_496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3257_ _3165_/A _6415_/Q _6485_/Q _3164_/Y VGND VGND VPWR VPWR _3257_/X sky130_fd_sc_hd__a31o_1
XFILLER_86_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3188_ _7042_/Q VGND VGND VPWR VPWR _3188_/Y sky130_fd_sc_hd__inv_2
XTAP_2308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6947_ _7027_/CLK _6947_/D fanout498/X VGND VGND VPWR VPWR _6947_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_169_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_290 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6878_ _7043_/CLK _6878_/D fanout520/X VGND VGND VPWR VPWR _6878_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_179_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5829_ _6578_/Q _5617_/X _5914_/A2 _6619_/Q VGND VGND VPWR VPWR _5829_/X sky130_fd_sc_hd__a22o_1
XFILLER_139_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_163_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold670 _5304_/X VGND VGND VPWR VPWR _6871_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_1_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold681 _6967_/Q VGND VGND VPWR VPWR hold681/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold692 _5297_/X VGND VGND VPWR VPWR _6865_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_134_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1370 hold1545/X VGND VGND VPWR VPWR _5207_/A0 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1381 _7077_/Q VGND VGND VPWR VPWR _5536_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_57_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1392 _6987_/Q VGND VGND VPWR VPWR _5435_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_18_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_185_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput208 _3216_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[5] sky130_fd_sc_hd__buf_12
XFILLER_126_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput219 _7182_/X VGND VGND VPWR VPWR mgmt_gpio_out[17] sky130_fd_sc_hd__buf_12
XFILLER_5_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4160_ _3684_/X _4160_/A1 _4165_/S VGND VGND VPWR VPWR _6572_/D sky130_fd_sc_hd__mux2_1
XFILLER_67_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4091_ hold527/X _4090_/X _4095_/S VGND VGND VPWR VPWR _4091_/X sky130_fd_sc_hd__mux2_1
XFILLER_83_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_488 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6801_ _6928_/CLK _6801_/D fanout501/X VGND VGND VPWR VPWR _6801_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_90_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4993_ _5064_/B _5064_/C VGND VGND VPWR VPWR _4994_/B sky130_fd_sc_hd__nand2_1
X_3944_ _3944_/A VGND VGND VPWR VPWR _3944_/Y sky130_fd_sc_hd__inv_2
X_6732_ _3500_/A1 _6732_/D _6384_/X VGND VGND VPWR VPWR _6732_/Q sky130_fd_sc_hd__dfrtn_1
XFILLER_176_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6663_ _6698_/CLK _6663_/D fanout496/X VGND VGND VPWR VPWR _6663_/Q sky130_fd_sc_hd__dfstp_1
X_3875_ _7088_/Q _7090_/Q _7091_/Q _7089_/Q VGND VGND VPWR VPWR _3876_/B sky130_fd_sc_hd__or4b_1
XFILLER_149_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5614_ _5667_/A _5645_/B _5646_/B VGND VGND VPWR VPWR _5614_/X sky130_fd_sc_hd__and3_4
XFILLER_31_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6594_ _7130_/CLK _6594_/D VGND VGND VPWR VPWR _6594_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_136_107 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5545_ hold644/X _5545_/A1 _5546_/S VGND VGND VPWR VPWR _5545_/X sky130_fd_sc_hd__mux2_1
XFILLER_191_235 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_3_0_0_csclk clkbuf_3_1_0_csclk/A VGND VGND VPWR VPWR _6661_/CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_117_376 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5476_ hold130/X _5476_/A1 hold19/X VGND VGND VPWR VPWR _5476_/X sky130_fd_sc_hd__mux2_1
XFILLER_132_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4427_ _4574_/A _4944_/B VGND VGND VPWR VPWR _4495_/B sky130_fd_sc_hd__nand2_1
XFILLER_120_519 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7146_ _3931_/A1 _7146_/D _4181_/B VGND VGND VPWR VPWR _7146_/Q sky130_fd_sc_hd__dfrtp_1
Xfanout424 _4649_/A VGND VGND VPWR VPWR _5026_/A sky130_fd_sc_hd__buf_8
X_4358_ _4356_/B _4592_/A _4357_/B _4613_/C VGND VGND VPWR VPWR _4399_/B sky130_fd_sc_hd__o2bb2a_1
XFILLER_98_271 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout435 _5526_/A1 VGND VGND VPWR VPWR _5544_/A1 sky130_fd_sc_hd__buf_6
XFILLER_58_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout446 _5533_/A1 VGND VGND VPWR VPWR _4289_/A1 sky130_fd_sc_hd__clkbuf_4
Xfanout457 _4299_/A1 VGND VGND VPWR VPWR _6354_/A1 sky130_fd_sc_hd__buf_6
Xfanout468 _5187_/B VGND VGND VPWR VPWR _6352_/B sky130_fd_sc_hd__buf_6
X_3309_ hold81/X _3366_/A VGND VGND VPWR VPWR _3374_/A sky130_fd_sc_hd__or2_4
X_7077_ _7078_/CLK _7077_/D fanout507/X VGND VGND VPWR VPWR _7077_/Q sky130_fd_sc_hd__dfrtp_1
Xfanout479 hold104/X VGND VGND VPWR VPWR _3856_/S sky130_fd_sc_hd__clkbuf_8
X_4289_ hold598/X _4289_/A1 _4290_/S VGND VGND VPWR VPWR _4289_/X sky130_fd_sc_hd__mux2_1
XFILLER_86_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6028_ _6787_/Q _6004_/B _6027_/X _5610_/A VGND VGND VPWR VPWR _6028_/X sky130_fd_sc_hd__o211a_1
XFILLER_86_499 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_129_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_379 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_104_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_179 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_161_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3660_ _6852_/Q _3374_/Y _5244_/A _6820_/Q _3659_/X VGND VGND VPWR VPWR _3660_/Y
+ sky130_fd_sc_hd__a221oi_1
XFILLER_173_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3591_ _6837_/Q _5262_/A _4166_/A _6581_/Q VGND VGND VPWR VPWR _3591_/X sky130_fd_sc_hd__a22o_1
XFILLER_127_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5330_ hold401/X _5534_/A1 _5333_/S VGND VGND VPWR VPWR _5330_/X sky130_fd_sc_hd__mux2_1
XFILLER_126_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5261_ hold124/X hold27/X _5261_/S VGND VGND VPWR VPWR _5261_/X sky130_fd_sc_hd__mux2_1
XFILLER_142_655 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7000_ _7000_/CLK _7000_/D fanout503/X VGND VGND VPWR VPWR _7000_/Q sky130_fd_sc_hd__dfrtp_1
X_4212_ hold590/X _5491_/A1 _4213_/S VGND VGND VPWR VPWR _4212_/X sky130_fd_sc_hd__mux2_1
XFILLER_87_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_142_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5192_ _5192_/A0 hold90/X _5198_/S VGND VGND VPWR VPWR hold91/A sky130_fd_sc_hd__mux2_1
XFILLER_68_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4143_ hold648/X _4289_/A1 _4144_/S VGND VGND VPWR VPWR _4143_/X sky130_fd_sc_hd__mux2_1
XFILLER_122_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4074_ hold291/X _4073_/X _4078_/S VGND VGND VPWR VPWR _4074_/X sky130_fd_sc_hd__mux2_1
XFILLER_49_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4976_ _5081_/C _4976_/B _4976_/C VGND VGND VPWR VPWR _4979_/C sky130_fd_sc_hd__and3_1
X_6715_ _6769_/CLK _6715_/D _6399_/A VGND VGND VPWR VPWR _6715_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_177_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3927_ _6498_/Q input3/X input1/X VGND VGND VPWR VPWR _3927_/X sky130_fd_sc_hd__mux2_4
XFILLER_137_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6646_ _7037_/CLK _6646_/D fanout484/X VGND VGND VPWR VPWR _6646_/Q sky130_fd_sc_hd__dfrtp_4
X_3858_ _6485_/Q _3858_/B VGND VGND VPWR VPWR _3860_/S sky130_fd_sc_hd__nand2_1
XFILLER_149_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_192_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3789_ _5168_/A _5161_/B VGND VGND VPWR VPWR _3789_/Y sky130_fd_sc_hd__nor2_1
X_6577_ _7140_/CLK _6577_/D VGND VGND VPWR VPWR _6577_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_152_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_600 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5528_ hold656/X _5537_/A1 _5528_/S VGND VGND VPWR VPWR _5528_/X sky130_fd_sc_hd__mux2_1
XFILLER_172_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5459_ hold965/X _5537_/A1 _5459_/S VGND VGND VPWR VPWR _5459_/X sky130_fd_sc_hd__mux2_1
XFILLER_133_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_160_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_422 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7129_ _7130_/CLK _7129_/D fanout488/X VGND VGND VPWR VPWR _7129_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_101_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_639 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_168_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_183_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_176 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_403 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_266 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_439 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_322 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_170 _5406_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4830_ _4959_/A _4959_/C VGND VGND VPWR VPWR _5087_/A sky130_fd_sc_hd__nor2_1
XFILLER_60_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_181 _5973_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_192 _7200_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4761_ _4748_/A _4901_/B _4501_/X _4760_/X VGND VGND VPWR VPWR _4761_/X sky130_fd_sc_hd__o211a_1
XTAP_1790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3712_ _3712_/A _3712_/B _3712_/C _3711_/Y VGND VGND VPWR VPWR _3713_/D sky130_fd_sc_hd__or4b_1
X_6500_ _7054_/CLK _6500_/D fanout503/X VGND VGND VPWR VPWR _7174_/A sky130_fd_sc_hd__dfrtp_1
XFILLER_119_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_174_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4692_ _4692_/A _4977_/B _4692_/C VGND VGND VPWR VPWR _4930_/C sky130_fd_sc_hd__nor3_2
XFILLER_174_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6431_ _6994_/CLK _6431_/D fanout489/X VGND VGND VPWR VPWR _6431_/Q sky130_fd_sc_hd__dfstp_1
X_3643_ _6652_/Q hold62/A _4208_/A _6616_/Q _3642_/X VGND VGND VPWR VPWR _3648_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_134_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6362_ _6400_/A _6399_/B VGND VGND VPWR VPWR _6362_/X sky130_fd_sc_hd__and2_1
X_3574_ _6845_/Q _5271_/A _5334_/A _6901_/Q VGND VGND VPWR VPWR _3574_/X sky130_fd_sc_hd__a22o_1
XFILLER_127_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5313_ hold757/X _5457_/A1 _5315_/S VGND VGND VPWR VPWR _5313_/X sky130_fd_sc_hd__mux2_1
XFILLER_154_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6293_ _6293_/A _6293_/B _6293_/C _6292_/Y VGND VGND VPWR VPWR _6293_/X sky130_fd_sc_hd__or4b_1
XFILLER_88_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5244_ _5244_/A _5511_/B VGND VGND VPWR VPWR _5252_/S sky130_fd_sc_hd__and2_4
XFILLER_114_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold18 hold18/A VGND VGND VPWR VPWR hold18/X sky130_fd_sc_hd__dlygate4sd3_1
X_5175_ hold383/X _5532_/A1 _5178_/S VGND VGND VPWR VPWR _5175_/X sky130_fd_sc_hd__mux2_1
Xhold29 hold29/A VGND VGND VPWR VPWR hold29/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_130_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_263 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4126_ hold471/X _5534_/A1 _4126_/S VGND VGND VPWR VPWR _4126_/X sky130_fd_sc_hd__mux2_1
XFILLER_96_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_734 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4057_ hold638/X _4056_/X _4061_/S VGND VGND VPWR VPWR _4057_/X sky130_fd_sc_hd__mux2_1
XFILLER_45_28 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_34 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4959_ _4959_/A _4959_/B _4959_/C _5087_/B VGND VGND VPWR VPWR _4959_/X sky130_fd_sc_hd__or4b_1
XFILLER_177_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6629_ _6632_/CLK _6629_/D _3264_/A VGND VGND VPWR VPWR _6629_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_137_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_192_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_193_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_655 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_142_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3290_ _3503_/A _3797_/A VGND VGND VPWR VPWR _5406_/A sky130_fd_sc_hd__nor2_8
XFILLER_111_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6980_ _7079_/CLK _6980_/D fanout514/X VGND VGND VPWR VPWR _6980_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_53_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_93_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5931_ _6544_/Q _5667_/X _5920_/X _5930_/X _5610_/A VGND VGND VPWR VPWR _5931_/X
+ sky130_fd_sc_hd__o221a_2
XFILLER_80_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5862_ _6646_/Q _5918_/A2 _5922_/A2 _6651_/Q VGND VGND VPWR VPWR _5862_/X sky130_fd_sc_hd__a22o_1
XFILLER_61_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4813_ _4933_/B _4813_/B _4813_/C _4813_/D VGND VGND VPWR VPWR _4816_/B sky130_fd_sc_hd__and4_1
XFILLER_33_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5793_ _6904_/Q _5623_/X _5637_/X _6856_/Q _5792_/X VGND VGND VPWR VPWR _5793_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_166_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4744_ _4717_/A _4715_/B _4410_/X VGND VGND VPWR VPWR _4772_/B sky130_fd_sc_hd__o21a_1
XFILLER_159_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4675_ _4678_/A _4901_/B VGND VGND VPWR VPWR _4717_/B sky130_fd_sc_hd__or2_4
XFILLER_135_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3626_ _3686_/A1 _3625_/X _3685_/S VGND VGND VPWR VPWR _3626_/X sky130_fd_sc_hd__mux2_1
X_6414_ _3500_/A1 _6414_/D _6370_/X VGND VGND VPWR VPWR _6414_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_162_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3557_ _3557_/A _3628_/B VGND VGND VPWR VPWR _4291_/A sky130_fd_sc_hd__nor2_8
XFILLER_115_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6345_ _6642_/Q _6345_/A2 _6345_/B1 _4222_/B _6344_/X VGND VGND VPWR VPWR _6345_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_103_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6276_ _6607_/Q wire390/X _6273_/X _6275_/X VGND VGND VPWR VPWR _6277_/C sky130_fd_sc_hd__a211o_1
X_3488_ input48/X _4103_/B _5145_/A _6741_/Q _3486_/X VGND VGND VPWR VPWR _3489_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_130_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5227_ _5227_/A0 _5488_/A1 _5234_/S VGND VGND VPWR VPWR _5227_/X sky130_fd_sc_hd__mux2_1
Xinput108 wb_adr_i[18] VGND VGND VPWR VPWR _4334_/D sky130_fd_sc_hd__clkbuf_1
Xinput119 wb_adr_i[28] VGND VGND VPWR VPWR _3893_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_69_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_583 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5158_ _5158_/A _6352_/B VGND VGND VPWR VPWR _5160_/S sky130_fd_sc_hd__and2_1
XFILLER_29_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4109_ hold387/X _5526_/A1 _4111_/S VGND VGND VPWR VPWR _4109_/X sky130_fd_sc_hd__mux2_1
XFILLER_29_469 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5089_ _5089_/A _5089_/B _5089_/C VGND VGND VPWR VPWR _5090_/B sky130_fd_sc_hd__and3_1
XFILLER_56_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_112_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_169_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_169_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_169_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_184_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_177_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_70 _6690_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_122_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_81 user_clock VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_126_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_92 _3943_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_153_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_192_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_141_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_133_260 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_236 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_175_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_188_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_129_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4460_ _4679_/A _4542_/A VGND VGND VPWR VPWR _4629_/B sky130_fd_sc_hd__nand2_4
Xhold307 _6654_/Q VGND VGND VPWR VPWR hold307/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_7_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold318 _4059_/X VGND VGND VPWR VPWR _6496_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3411_ _6792_/Q _5208_/A _3343_/Y input50/X _3410_/X VGND VGND VPWR VPWR _3411_/X
+ sky130_fd_sc_hd__a221o_1
Xhold329 _6868_/Q VGND VGND VPWR VPWR hold329/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_144_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4391_ _4542_/C _4383_/C _4888_/A VGND VGND VPWR VPWR _4391_/Y sky130_fd_sc_hd__a21boi_1
X_6130_ _6154_/A1 _5612_/Y _6128_/X _6129_/X VGND VGND VPWR VPWR _7124_/D sky130_fd_sc_hd__o22a_1
X_3342_ _3440_/A _3401_/B VGND VGND VPWR VPWR _5183_/B sky130_fd_sc_hd__or2_4
XFILLER_98_623 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6061_ _6989_/Q _6286_/B1 _6284_/B1 _6861_/Q VGND VGND VPWR VPWR _6061_/X sky130_fd_sc_hd__a22o_1
X_3273_ _3856_/S _6414_/Q VGND VGND VPWR VPWR _3273_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_39_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1007 _4129_/X VGND VGND VPWR VPWR _6546_/D sky130_fd_sc_hd__dlygate4sd3_1
X_5012_ _5043_/A _4470_/A _5061_/A _4746_/X _4912_/B VGND VGND VPWR VPWR _5101_/A
+ sky130_fd_sc_hd__o2111a_1
Xhold1018 _6519_/Q VGND VGND VPWR VPWR _4098_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1029 _3962_/X VGND VGND VPWR VPWR _6419_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_66_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6963_ _7072_/CLK _6963_/D fanout504/X VGND VGND VPWR VPWR _6963_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_53_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5914_ _6623_/Q _5914_/A2 _5634_/X _6689_/Q VGND VGND VPWR VPWR _5914_/X sky130_fd_sc_hd__a22o_1
XFILLER_22_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6894_ _7039_/CLK _6894_/D fanout498/X VGND VGND VPWR VPWR _6894_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_179_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5845_ _5845_/A1 _6305_/A2 _5843_/X _5844_/X VGND VGND VPWR VPWR _7114_/D sky130_fd_sc_hd__o22a_1
XFILLER_22_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5776_ _6975_/Q _5644_/X _5766_/X _5770_/X _5775_/X VGND VGND VPWR VPWR _5776_/X
+ sky130_fd_sc_hd__a2111o_1
XFILLER_158_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4727_ _4691_/A _4595_/B _4439_/Y _4930_/C _4726_/X VGND VGND VPWR VPWR _4728_/C
+ sky130_fd_sc_hd__a311o_1
XFILLER_147_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4658_ _4701_/A _4861_/B _4616_/X _4657_/X VGND VGND VPWR VPWR _4658_/X sky130_fd_sc_hd__o211a_1
XFILLER_190_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput90 spimemio_flash_io2_oeb VGND VGND VPWR VPWR input90/X sky130_fd_sc_hd__dlymetal6s2s_1
X_3609_ _7021_/Q hold18/A _4121_/A _6543_/Q _3608_/X VGND VGND VPWR VPWR _3614_/B
+ sky130_fd_sc_hd__a221o_1
Xhold830 _4217_/X VGND VGND VPWR VPWR _6621_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold841 _6873_/Q VGND VGND VPWR VPWR hold841/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_1_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold852 _5299_/X VGND VGND VPWR VPWR _6866_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_162_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4589_ _4534_/X _4580_/X _4531_/X VGND VGND VPWR VPWR _4589_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_89_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold863 _7153_/Q VGND VGND VPWR VPWR hold863/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold874 _5264_/X VGND VGND VPWR VPWR _6835_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_103_411 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6328_ _6327_/X _6328_/A1 _6346_/S VGND VGND VPWR VPWR _7142_/D sky130_fd_sc_hd__mux2_1
Xhold885 _6569_/Q VGND VGND VPWR VPWR hold885/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold896 _5189_/X VGND VGND VPWR VPWR _6769_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_131_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6259_ _6558_/Q _6259_/A2 _5973_/B _6553_/Q VGND VGND VPWR VPWR _6259_/X sky130_fd_sc_hd__a22o_1
XFILLER_131_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_296 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1530 _6527_/Q VGND VGND VPWR VPWR hold769/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1541 _6498_/Q VGND VGND VPWR VPWR hold1541/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1552 _6533_/Q VGND VGND VPWR VPWR hold984/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_123_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3960_ _3960_/A0 _5488_/A1 _3974_/S VGND VGND VPWR VPWR _3960_/X sky130_fd_sc_hd__mux2_1
XFILLER_51_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_189_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3891_ _3891_/A _3891_/B VGND VGND VPWR VPWR _4499_/B sky130_fd_sc_hd__or2_2
XFILLER_149_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5630_ _5667_/A _5648_/C _5651_/C VGND VGND VPWR VPWR _5630_/X sky130_fd_sc_hd__and3_4
XFILLER_85_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5561_ _5561_/A _5561_/B _5561_/C VGND VGND VPWR VPWR _7090_/D sky130_fd_sc_hd__and3_1
XFILLER_191_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4512_ _4943_/B _4586_/B _4510_/X _4511_/X VGND VGND VPWR VPWR _4514_/C sky130_fd_sc_hd__o211a_1
XFILLER_129_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5492_ hold423/X _5534_/A1 _5492_/S VGND VGND VPWR VPWR _5492_/X sky130_fd_sc_hd__mux2_1
XFILLER_156_171 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold104 _6488_/Q VGND VGND VPWR VPWR hold104/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_144_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold115 _5536_/X VGND VGND VPWR VPWR _7077_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_105_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold126 hold126/A VGND VGND VPWR VPWR hold126/X sky130_fd_sc_hd__dlygate4sd3_1
X_4443_ _4542_/A _5048_/A VGND VGND VPWR VPWR _4656_/A sky130_fd_sc_hd__nand2_1
Xhold137 _5206_/X VGND VGND VPWR VPWR _6784_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_144_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold148 _7146_/Q VGND VGND VPWR VPWR hold148/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold159 _6919_/Q VGND VGND VPWR VPWR hold159/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_113_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7162_ net499_2/A _7162_/D _6392_/X VGND VGND VPWR VPWR hold44/A sky130_fd_sc_hd__dfrtp_1
X_4374_ _4679_/A _4554_/A _4596_/B VGND VGND VPWR VPWR _4409_/B sky130_fd_sc_hd__and3_2
XFILLER_113_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3325_ hold81/A hold39/X hold51/A VGND VGND VPWR VPWR hold40/A sky130_fd_sc_hd__or3b_4
X_6113_ _6839_/Q _5946_/X _5971_/A _6871_/Q VGND VGND VPWR VPWR _6113_/X sky130_fd_sc_hd__a22o_1
X_7093_ _7124_/CLK _7093_/D fanout501/X VGND VGND VPWR VPWR _7093_/Q sky130_fd_sc_hd__dfstp_1
XTAP_431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6044_ _6980_/Q _6176_/A2 _5974_/B _6828_/Q VGND VGND VPWR VPWR _6044_/X sky130_fd_sc_hd__a22o_1
X_3256_ _3247_/A _3256_/A1 _3256_/S VGND VGND VPWR VPWR _7160_/D sky130_fd_sc_hd__mux2_1
XTAP_486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3187_ _7050_/Q VGND VGND VPWR VPWR _3187_/Y sky130_fd_sc_hd__inv_2
XFILLER_27_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_512 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6946_ _6978_/CLK _6946_/D fanout500/X VGND VGND VPWR VPWR _6946_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_54_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_9 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6877_ _7029_/CLK _6877_/D fanout517/X VGND VGND VPWR VPWR _6877_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_169_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5828_ _5828_/A _5828_/B VGND VGND VPWR VPWR _5828_/X sky130_fd_sc_hd__or2_1
XFILLER_139_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5759_ _6991_/Q _5622_/X _5624_/X _6831_/Q VGND VGND VPWR VPWR _5759_/X sky130_fd_sc_hd__a22o_1
XFILLER_108_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_135_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_163_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_162_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_190_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold660 _6857_/Q VGND VGND VPWR VPWR hold660/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold671 _6999_/Q VGND VGND VPWR VPWR hold671/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold682 _5412_/X VGND VGND VPWR VPWR _6967_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold693 _7060_/Q VGND VGND VPWR VPWR hold693/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_77_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1360 hold1360/A VGND VGND VPWR VPWR wb_dat_o[30] sky130_fd_sc_hd__buf_12
XFILLER_18_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1371 _7193_/A VGND VGND VPWR VPWR _5195_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_27_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1382 _6612_/Q VGND VGND VPWR VPWR _4206_/A0 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1393 _6575_/Q VGND VGND VPWR VPWR hold1393/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_159_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_283 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_126_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_160 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput209 _3215_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[6] sky130_fd_sc_hd__buf_12
XFILLER_126_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4090_ hold395/X _5526_/A1 hold76/X VGND VGND VPWR VPWR _4090_/X sky130_fd_sc_hd__mux2_1
XFILLER_191_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_556 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6800_ _7086_/CLK _6800_/D fanout515/X VGND VGND VPWR VPWR _6800_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_91_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4992_ _4513_/A _4988_/A _4748_/B _4973_/A _4817_/B VGND VGND VPWR VPWR _5064_/C
+ sky130_fd_sc_hd__o221a_1
XFILLER_51_548 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6731_ _3500_/A1 _6731_/D _6383_/X VGND VGND VPWR VPWR _6731_/Q sky130_fd_sc_hd__dfrtn_1
X_3943_ _6403_/Q _3943_/B VGND VGND VPWR VPWR _3944_/A sky130_fd_sc_hd__or2_2
XFILLER_189_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6662_ _6689_/CLK _6662_/D fanout509/X VGND VGND VPWR VPWR _6662_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_31_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3874_ _7090_/Q _7091_/Q VGND VGND VPWR VPWR _5607_/C sky130_fd_sc_hd__nor2_1
X_5613_ _7094_/Q _7095_/Q VGND VGND VPWR VPWR _5646_/B sky130_fd_sc_hd__and2b_2
X_6593_ _7130_/CLK _6593_/D VGND VGND VPWR VPWR _6593_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_191_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_191_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5544_ hold749/X _5544_/A1 _5546_/S VGND VGND VPWR VPWR _5544_/X sky130_fd_sc_hd__mux2_1
XFILLER_145_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5475_ hold717/X _5544_/A1 hold19/X VGND VGND VPWR VPWR _5475_/X sky130_fd_sc_hd__mux2_1
XFILLER_160_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_160_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4426_ _4409_/B _4707_/C _4391_/Y _4402_/B VGND VGND VPWR VPWR _4561_/B sky130_fd_sc_hd__a211o_2
XFILLER_99_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_160_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7145_ _3931_/A1 _7145_/D _6308_/B VGND VGND VPWR VPWR hold67/A sky130_fd_sc_hd__dfrtp_1
XFILLER_113_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout425 _4469_/X VGND VGND VPWR VPWR _4901_/B sky130_fd_sc_hd__buf_6
X_4357_ _4357_/A _4357_/B VGND VGND VPWR VPWR _4429_/B sky130_fd_sc_hd__or2_1
XFILLER_98_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout436 _5526_/A1 VGND VGND VPWR VPWR _5457_/A1 sky130_fd_sc_hd__buf_2
Xfanout447 hold45/X VGND VGND VPWR VPWR _5533_/A1 sky130_fd_sc_hd__buf_6
Xfanout458 _4299_/A1 VGND VGND VPWR VPWR _5189_/A1 sky130_fd_sc_hd__buf_6
X_3308_ _6969_/Q _5406_/A _5529_/A _7078_/Q _3307_/X VGND VGND VPWR VPWR _3349_/A
+ sky130_fd_sc_hd__a221o_1
X_7076_ _7076_/CLK _7076_/D fanout502/X VGND VGND VPWR VPWR _7076_/Q sky130_fd_sc_hd__dfrtp_4
Xfanout469 hold6/X VGND VGND VPWR VPWR _5187_/B sky130_fd_sc_hd__clkbuf_8
XFILLER_100_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4288_ hold805/X _5505_/A1 _4290_/S VGND VGND VPWR VPWR _4288_/X sky130_fd_sc_hd__mux2_1
XFILLER_74_607 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6027_ _6027_/A _6027_/B _6027_/C _6004_/B VGND VGND VPWR VPWR _6027_/X sky130_fd_sc_hd__or4b_1
X_3239_ _3856_/S _6485_/Q VGND VGND VPWR VPWR _3819_/B sky130_fd_sc_hd__or2_1
XFILLER_27_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6929_ _7017_/CLK _6929_/D fanout515/X VGND VGND VPWR VPWR _6929_/Q sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_31_csclk clkbuf_3_7_0_csclk/X VGND VGND VPWR VPWR _7029_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_168_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_167_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_46_csclk clkbuf_opt_3_0_csclk/X VGND VGND VPWR VPWR _7075_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_89_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_135_185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold490 _5376_/X VGND VGND VPWR VPWR _6935_/D sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_1_0_0_wb_clk_i clkbuf_0_wb_clk_i/X VGND VGND VPWR VPWR clkbuf_1_0_1_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_77_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_380 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_640 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1190 _4140_/X VGND VGND VPWR VPWR _6555_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_161_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_173_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3590_ _6628_/Q _4225_/A _4237_/A _6648_/Q _3589_/X VGND VGND VPWR VPWR _3596_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_127_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_612 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5260_ hold483/X _5545_/A1 _5261_/S VGND VGND VPWR VPWR _5260_/X sky130_fd_sc_hd__mux2_1
XFILLER_48_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_667 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4211_ hold825/X _5505_/A1 _4213_/S VGND VGND VPWR VPWR _4211_/X sky130_fd_sc_hd__mux2_1
XFILLER_141_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5191_ hold793/X _5521_/A1 _5198_/S VGND VGND VPWR VPWR _5191_/X sky130_fd_sc_hd__mux2_1
X_4142_ hold783/X _5505_/A1 _4144_/S VGND VGND VPWR VPWR _4142_/X sky130_fd_sc_hd__mux2_1
XFILLER_68_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4073_ _4118_/A0 hold142/X _4077_/S VGND VGND VPWR VPWR _4073_/X sky130_fd_sc_hd__mux2_1
XFILLER_110_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_183 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4975_ _4631_/X _4973_/B _4972_/X _4973_/X _4974_/X VGND VGND VPWR VPWR _4976_/C
+ sky130_fd_sc_hd__o2111a_1
X_6714_ _6718_/CLK _6714_/D fanout496/X VGND VGND VPWR VPWR _6714_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_149_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3926_ _3925_/X _3947_/B _6403_/Q VGND VGND VPWR VPWR _3926_/X sky130_fd_sc_hd__mux2_4
XFILLER_177_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6645_ _7037_/CLK _6645_/D fanout485/X VGND VGND VPWR VPWR _6645_/Q sky130_fd_sc_hd__dfrtp_2
X_3857_ _3856_/X _3857_/A1 _3857_/S VGND VGND VPWR VPWR _6407_/D sky130_fd_sc_hd__mux2_1
XFILLER_20_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6576_ _7140_/CLK _6576_/D VGND VGND VPWR VPWR _6576_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_166_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3788_ _6914_/Q _5352_/A _5325_/A _6890_/Q _3787_/X VGND VGND VPWR VPWR _3792_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_118_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_118_664 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5527_ hold608/X _5545_/A1 _5528_/S VGND VGND VPWR VPWR _5527_/X sky130_fd_sc_hd__mux2_1
XFILLER_192_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5458_ hold594/X _5545_/A1 _5459_/S VGND VGND VPWR VPWR _5458_/X sky130_fd_sc_hd__mux2_1
XFILLER_132_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4409_ _4542_/A _4409_/B VGND VGND VPWR VPWR _4943_/A sky130_fd_sc_hd__nand2b_4
XFILLER_160_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5389_ _5389_/A0 _5488_/A1 _5396_/S VGND VGND VPWR VPWR _5389_/X sky130_fd_sc_hd__mux2_1
XFILLER_87_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7128_ _7130_/CLK _7128_/D fanout488/X VGND VGND VPWR VPWR _7128_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_59_434 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7059_ _7059_/CLK _7059_/D fanout517/X VGND VGND VPWR VPWR _7059_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_55_651 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_155_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_171_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_183_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_710 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_278 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_375 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_643 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_160 hold23/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_171 _5511_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_182 _5950_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_193 input46/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_175 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4760_ _4640_/B _4748_/A _4748_/X _4503_/D VGND VGND VPWR VPWR _4760_/X sky130_fd_sc_hd__o211a_1
XTAP_1791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3711_ _3711_/A _3711_/B _3711_/C _3711_/D VGND VGND VPWR VPWR _3711_/Y sky130_fd_sc_hd__nor4_1
XFILLER_186_350 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4691_ _4691_/A _4692_/C _4691_/C _4555_/B VGND VGND VPWR VPWR _4723_/C sky130_fd_sc_hd__or4b_1
X_6430_ _7034_/CLK _6430_/D fanout489/X VGND VGND VPWR VPWR _6430_/Q sky130_fd_sc_hd__dfrtp_4
X_3642_ _6601_/Q _4190_/A _4145_/A _6562_/Q VGND VGND VPWR VPWR _3642_/X sky130_fd_sc_hd__a22o_1
XFILLER_146_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6361_ _6399_/A _6401_/B VGND VGND VPWR VPWR _6361_/X sky130_fd_sc_hd__and2_1
XFILLER_162_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3573_ input38/X hold76/A _4291_/A _6693_/Q VGND VGND VPWR VPWR _3573_/X sky130_fd_sc_hd__a22o_1
XFILLER_127_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5312_ _5312_/A0 _5465_/A1 _5315_/S VGND VGND VPWR VPWR _5312_/X sky130_fd_sc_hd__mux2_1
XFILLER_114_122 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6292_ _6292_/A _6292_/B VGND VGND VPWR VPWR _6292_/Y sky130_fd_sc_hd__nor2_1
X_5243_ hold853/X _5537_/A1 _5243_/S VGND VGND VPWR VPWR _5243_/X sky130_fd_sc_hd__mux2_1
XFILLER_88_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_114_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold19 hold19/A VGND VGND VPWR VPWR hold19/X sky130_fd_sc_hd__dlygate4sd3_1
X_5174_ hold217/X _5533_/A1 _5178_/S VGND VGND VPWR VPWR _5174_/X sky130_fd_sc_hd__mux2_1
XFILLER_68_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4125_ hold549/X _5491_/A1 _4126_/S VGND VGND VPWR VPWR _4125_/X sky130_fd_sc_hd__mux2_1
XFILLER_56_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_275 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4056_ hold387/X _5526_/A1 _4103_/B VGND VGND VPWR VPWR _4056_/X sky130_fd_sc_hd__mux2_1
XFILLER_37_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_632 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4958_ _4958_/A _4958_/B _4958_/C _5121_/A VGND VGND VPWR VPWR _4959_/B sky130_fd_sc_hd__or4b_1
XFILLER_184_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3909_ _3948_/A _3869_/X _3908_/B _6635_/Q VGND VGND VPWR VPWR _6640_/D sky130_fd_sc_hd__a22o_1
X_4889_ _4894_/B _4892_/B VGND VGND VPWR VPWR _4889_/X sky130_fd_sc_hd__or2_1
XFILLER_137_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6628_ _6718_/CLK _6628_/D _6401_/A VGND VGND VPWR VPWR _6628_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_20_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_192_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6559_ _6559_/CLK _6559_/D fanout509/X VGND VGND VPWR VPWR _6559_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_146_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_192_397 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_667 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_129_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5930_ _5930_/A _5930_/B _5930_/C _5929_/Y VGND VGND VPWR VPWR _5930_/X sky130_fd_sc_hd__or4b_1
XFILLER_19_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_172 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_179_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5861_ _6626_/Q _5913_/B1 _5926_/B1 _6546_/Q _5860_/X VGND VGND VPWR VPWR _5864_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_92_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4812_ _4812_/A _4812_/B _4812_/C _4812_/D VGND VGND VPWR VPWR _4813_/D sky130_fd_sc_hd__and4_1
XFILLER_34_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5792_ _6872_/Q _5625_/X _5643_/X _6888_/Q VGND VGND VPWR VPWR _5792_/X sky130_fd_sc_hd__a22o_1
XFILLER_21_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4743_ _4407_/X _4573_/A _4714_/C VGND VGND VPWR VPWR _4743_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_187_692 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_186_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4674_ _5043_/A _4615_/X _4631_/X _4901_/B VGND VGND VPWR VPWR _5116_/A sky130_fd_sc_hd__o22a_1
X_6413_ _3500_/A1 _6413_/D _6369_/X VGND VGND VPWR VPWR hold14/A sky130_fd_sc_hd__dfrtp_1
X_3625_ _3625_/A _3625_/B _3625_/C _3624_/X VGND VGND VPWR VPWR _3625_/X sky130_fd_sc_hd__or4b_4
XFILLER_135_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6344_ _6644_/Q _6344_/A2 _6344_/B1 _6643_/Q VGND VGND VPWR VPWR _6344_/X sky130_fd_sc_hd__a22o_1
X_3556_ _6790_/Q _5208_/A _4285_/A _6689_/Q _3555_/X VGND VGND VPWR VPWR _3565_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_142_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_143_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6275_ _6703_/Q _5975_/C _5980_/Y _6468_/Q _6274_/X VGND VGND VPWR VPWR _6275_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_170_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3487_ _3487_/A _5183_/A VGND VGND VPWR VPWR _5145_/A sky130_fd_sc_hd__nor2_8
X_5226_ _5226_/A _5511_/B VGND VGND VPWR VPWR _5234_/S sky130_fd_sc_hd__and2_4
Xinput109 wb_adr_i[19] VGND VGND VPWR VPWR _4334_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_102_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5157_ hold151/X hold142/X _5157_/S VGND VGND VPWR VPWR _5157_/X sky130_fd_sc_hd__mux2_1
XFILLER_69_595 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4108_ hold134/X hold23/X _4111_/S VGND VGND VPWR VPWR _4108_/X sky130_fd_sc_hd__mux2_1
XFILLER_56_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5088_ _4958_/A _5088_/B _5088_/C VGND VGND VPWR VPWR _5089_/C sky130_fd_sc_hd__and3b_1
XFILLER_44_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4039_ _4039_/A0 _5308_/A1 _4043_/S VGND VGND VPWR VPWR _4039_/X sky130_fd_sc_hd__mux2_1
XFILLER_56_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_169_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_60 _5948_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_71 _6405_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_392 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_82 user_clock VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_193_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_93 _3943_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_126_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_137_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_106_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_464 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_153_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_148_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_707 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_183_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold308 _4248_/X VGND VGND VPWR VPWR _6654_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold319 _6632_/Q VGND VGND VPWR VPWR hold319/X sky130_fd_sc_hd__dlygate4sd3_1
X_3410_ _7008_/Q _5451_/A _3374_/Y _6856_/Q VGND VGND VPWR VPWR _3410_/X sky130_fd_sc_hd__a22o_1
X_4390_ _4390_/A _4390_/B VGND VGND VPWR VPWR _4402_/B sky130_fd_sc_hd__nor2_1
XFILLER_124_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3341_ _3503_/A _3374_/A VGND VGND VPWR VPWR _5424_/A sky130_fd_sc_hd__nor2_8
XTAP_602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_140_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6060_ _6917_/Q _5937_/X _6296_/A2 _6885_/Q _6059_/X VGND VGND VPWR VPWR _6068_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_140_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3272_ hold57/X _6726_/Q _6624_/Q VGND VGND VPWR VPWR hold58/A sky130_fd_sc_hd__mux2_1
XTAP_657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1008 _6461_/Q VGND VGND VPWR VPWR _4016_/A0 sky130_fd_sc_hd__dlygate4sd3_1
X_5011_ _4672_/B _5005_/B _4748_/X _4912_/C _4463_/X VGND VGND VPWR VPWR _5105_/B
+ sky130_fd_sc_hd__o2111a_1
XTAP_679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1019 _4098_/X VGND VGND VPWR VPWR _6519_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_38_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6962_ _7055_/CLK _6962_/D fanout504/X VGND VGND VPWR VPWR _6962_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_53_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5913_ _6559_/Q _5913_/A2 _5913_/B1 _6629_/Q _5912_/X VGND VGND VPWR VPWR _5916_/A
+ sky130_fd_sc_hd__a221o_1
X_6893_ _7080_/CLK _6893_/D fanout514/X VGND VGND VPWR VPWR _6893_/Q sky130_fd_sc_hd__dfrtp_4
X_5844_ _7113_/Q _5612_/A _5612_/B VGND VGND VPWR VPWR _5844_/X sky130_fd_sc_hd__o21a_1
XFILLER_61_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5775_ _6447_/Q _5917_/B1 _5771_/X _5772_/X _5774_/X VGND VGND VPWR VPWR _5775_/X
+ sky130_fd_sc_hd__a2111o_1
XFILLER_166_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_159_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4726_ _5068_/A _4851_/B _4726_/C _4725_/X VGND VGND VPWR VPWR _4726_/X sky130_fd_sc_hd__or4b_1
XFILLER_175_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_175_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_175_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_175_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4657_ _4328_/Y _4575_/B _4703_/B _4676_/B _4962_/C VGND VGND VPWR VPWR _4657_/X
+ sky130_fd_sc_hd__o32a_1
XFILLER_174_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput80 spi_sck VGND VGND VPWR VPWR input80/X sky130_fd_sc_hd__dlymetal6s2s_1
X_3608_ _6997_/Q _5442_/A _4020_/A _6468_/Q VGND VGND VPWR VPWR _3608_/X sky130_fd_sc_hd__a22o_1
Xhold820 _4228_/X VGND VGND VPWR VPWR _6627_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_174_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput91 spimemio_flash_io3_do VGND VGND VPWR VPWR input91/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold831 _6542_/Q VGND VGND VPWR VPWR hold831/X sky130_fd_sc_hd__dlygate4sd3_1
X_4588_ _4921_/A _4588_/B VGND VGND VPWR VPWR _4920_/A sky130_fd_sc_hd__nor2_1
Xhold842 _5306_/X VGND VGND VPWR VPWR _6873_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold853 _6817_/Q VGND VGND VPWR VPWR hold853/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold864 _6355_/X VGND VGND VPWR VPWR _7153_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_162_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6327_ _6644_/Q _6327_/A2 _6327_/B1 _4222_/B _6326_/X VGND VGND VPWR VPWR _6327_/X
+ sky130_fd_sc_hd__a221o_1
Xhold875 _6666_/Q VGND VGND VPWR VPWR hold875/X sky130_fd_sc_hd__dlygate4sd3_1
X_3539_ _6474_/Q _4026_/A _4267_/A _6674_/Q VGND VGND VPWR VPWR _3539_/X sky130_fd_sc_hd__a22o_1
Xmgmt_gpio_15_buff_inst _3930_/X VGND VGND VPWR VPWR mgmt_gpio_out[15] sky130_fd_sc_hd__clkbuf_8
XFILLER_131_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold886 _4156_/X VGND VGND VPWR VPWR _6569_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_130_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold897 _6634_/Q VGND VGND VPWR VPWR hold897/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_107_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6258_ _6713_/Q _6294_/B1 _5976_/Y _6478_/Q _6257_/X VGND VGND VPWR VPWR _6268_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_76_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_467 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_264 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5209_ _5209_/A0 _5530_/A1 _5216_/S VGND VGND VPWR VPWR _5209_/X sky130_fd_sc_hd__mux2_1
X_6189_ _6680_/Q _5949_/X _5980_/Y _6465_/Q VGND VGND VPWR VPWR _6189_/X sky130_fd_sc_hd__a22o_1
Xhold1520 _7115_/Q VGND VGND VPWR VPWR _5867_/A1 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1531 _7117_/Q VGND VGND VPWR VPWR _5911_/A1 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1542 _7183_/A VGND VGND VPWR VPWR hold493/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1553 _7182_/A VGND VGND VPWR VPWR hold275/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_123_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_165_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_148_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_264 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_543 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_189_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_188_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_188_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3890_ _3891_/A _3891_/B VGND VGND VPWR VPWR _4449_/A sky130_fd_sc_hd__nor2_1
XFILLER_43_292 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_149_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5560_ _7088_/Q _7089_/Q _5558_/D _7090_/Q VGND VGND VPWR VPWR _5561_/C sky130_fd_sc_hd__a31o_1
XFILLER_78_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4511_ _4549_/B _4586_/B _4495_/X _4943_/A _5135_/A VGND VGND VPWR VPWR _4511_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_191_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5491_ hold479/X _5491_/A1 _5492_/S VGND VGND VPWR VPWR _5491_/X sky130_fd_sc_hd__mux2_1
XFILLER_156_183 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold105 _3856_/S VGND VGND VPWR VPWR hold105/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_117_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4442_ _4789_/A _4862_/A VGND VGND VPWR VPWR _5100_/A sky130_fd_sc_hd__or2_1
Xhold116 _7196_/A VGND VGND VPWR VPWR hold116/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold127 _4105_/X VGND VGND VPWR VPWR _6525_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold138 _7195_/A VGND VGND VPWR VPWR hold138/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold149 _3969_/X VGND VGND VPWR VPWR hold149/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_144_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7161_ net499_2/A _7161_/D _6391_/X VGND VGND VPWR VPWR hold1/A sky130_fd_sc_hd__dfrtp_1
X_4373_ _4345_/C _4888_/B _4373_/C VGND VGND VPWR VPWR _4737_/B sky130_fd_sc_hd__nand3b_4
XFILLER_98_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_171_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6112_ _6847_/Q _5939_/X _6283_/A2 _7068_/Q _6111_/X VGND VGND VPWR VPWR _6118_/C
+ sky130_fd_sc_hd__a221o_1
XTAP_421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3324_ hold75/X _3531_/A VGND VGND VPWR VPWR _5271_/A sky130_fd_sc_hd__nor2_8
XTAP_432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7092_ _7131_/CLK _7092_/D fanout501/X VGND VGND VPWR VPWR _7092_/Q sky130_fd_sc_hd__dfrtp_2
XTAP_443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6043_ _6043_/A _6043_/B _6043_/C _6042_/Y VGND VGND VPWR VPWR _6043_/X sky130_fd_sc_hd__or4b_1
XTAP_476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3255_ _3256_/A1 _3255_/A1 _3256_/S VGND VGND VPWR VPWR _7161_/D sky130_fd_sc_hd__mux2_1
XTAP_487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3186_ _7058_/Q VGND VGND VPWR VPWR _3186_/Y sky130_fd_sc_hd__inv_2
XFILLER_27_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6945_ _6945_/CLK _6945_/D fanout506/X VGND VGND VPWR VPWR _6945_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_35_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_2_2_0_wb_clk_i clkbuf_2_3_0_wb_clk_i/A VGND VGND VPWR VPWR clkbuf_3_5_0_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_22_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6876_ _7082_/CLK hold4/X fanout520/X VGND VGND VPWR VPWR _6876_/Q sky130_fd_sc_hd__dfrtp_4
X_5827_ _6665_/Q _5633_/X _5918_/B1 _6604_/Q _5826_/X VGND VGND VPWR VPWR _5828_/B
+ sky130_fd_sc_hd__a221o_1
X_5758_ _3222_/Y _5646_/A _5667_/B VGND VGND VPWR VPWR _5758_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_154_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4709_ _4709_/A _4709_/B _4709_/C _4708_/X VGND VGND VPWR VPWR _4711_/B sky130_fd_sc_hd__or4b_1
XFILLER_147_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_163_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5689_ _6787_/Q _5667_/X _5678_/X _5688_/X _5610_/A VGND VGND VPWR VPWR _5689_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_135_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_162_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_190_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold650 _6767_/Q VGND VGND VPWR VPWR hold650/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold661 _5288_/X VGND VGND VPWR VPWR _6857_/D sky130_fd_sc_hd__dlygate4sd3_1
Xmax_cap380 _5952_/Y VGND VGND VPWR VPWR _6290_/A2 sky130_fd_sc_hd__buf_12
XFILLER_162_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold672 _5448_/X VGND VGND VPWR VPWR _6999_/D sky130_fd_sc_hd__dlygate4sd3_1
Xmax_cap391 _5959_/Y VGND VGND VPWR VPWR _5971_/A sky130_fd_sc_hd__buf_12
Xhold683 _6823_/Q VGND VGND VPWR VPWR hold683/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold694 _5517_/X VGND VGND VPWR VPWR _7060_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_1_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_131_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1350 hold1350/A VGND VGND VPWR VPWR wb_dat_o[0] sky130_fd_sc_hd__buf_12
Xhold1361 _6312_/A1 VGND VGND VPWR VPWR hold1361/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_17_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1372 hold1482/X VGND VGND VPWR VPWR _5200_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1383 _6653_/Q VGND VGND VPWR VPWR _4247_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1394 _6577_/Q VGND VGND VPWR VPWR hold1394/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_84_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_404 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_186_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_295 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_173_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_1_0__f__1162_ clkbuf_0__1162_/X VGND VGND VPWR VPWR _4186_/A0 sky130_fd_sc_hd__clkbuf_16
XFILLER_114_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_175_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_191_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4991_ _4991_/A _4991_/B VGND VGND VPWR VPWR _4994_/A sky130_fd_sc_hd__or2_1
XFILLER_91_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6730_ _3939_/A1 _6730_/D _6382_/X VGND VGND VPWR VPWR _6730_/Q sky130_fd_sc_hd__dfrtn_1
X_3942_ _3942_/A VGND VGND VPWR VPWR _3942_/Y sky130_fd_sc_hd__inv_2
XFILLER_189_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6661_ _6661_/CLK _6661_/D fanout490/X VGND VGND VPWR VPWR _6661_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_176_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3873_ _6644_/Q _3869_/X _3873_/B1 VGND VGND VPWR VPWR _6644_/D sky130_fd_sc_hd__a21o_1
XFILLER_31_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5612_ _5612_/A _5612_/B VGND VGND VPWR VPWR _5612_/Y sky130_fd_sc_hd__nand2_2
X_6592_ _7130_/CLK _6592_/D VGND VGND VPWR VPWR _6592_/Q sky130_fd_sc_hd__dfxtp_1
X_5543_ _5543_/A0 _5543_/A1 _5546_/S VGND VGND VPWR VPWR _5543_/X sky130_fd_sc_hd__mux2_1
XFILLER_117_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5474_ _5474_/A0 _5543_/A1 hold19/X VGND VGND VPWR VPWR _5474_/X sky130_fd_sc_hd__mux2_1
XFILLER_105_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_144_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4425_ _4535_/A _4946_/A _4947_/A VGND VGND VPWR VPWR _4425_/X sky130_fd_sc_hd__and3_1
XFILLER_144_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_99_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7144_ _3931_/A1 _7144_/D _6308_/B VGND VGND VPWR VPWR _7144_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_98_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_160_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4356_ _4630_/A _4356_/B VGND VGND VPWR VPWR _4367_/B sky130_fd_sc_hd__xnor2_1
Xfanout426 _4469_/X VGND VGND VPWR VPWR _4703_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_48_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout437 hold142/X VGND VGND VPWR VPWR _5526_/A1 sky130_fd_sc_hd__clkbuf_8
X_3307_ _6929_/Q _3297_/Y _4092_/S input42/X _3306_/X VGND VGND VPWR VPWR _3307_/X
+ sky130_fd_sc_hd__a221o_1
Xfanout448 _5515_/A1 VGND VGND VPWR VPWR _5542_/A1 sky130_fd_sc_hd__buf_6
X_7075_ _7075_/CLK _7075_/D fanout505/X VGND VGND VPWR VPWR _7075_/Q sky130_fd_sc_hd__dfrtp_2
Xfanout459 _4299_/A1 VGND VGND VPWR VPWR _5495_/A1 sky130_fd_sc_hd__buf_6
X_4287_ hold998/X _5189_/A1 _4290_/S VGND VGND VPWR VPWR _4287_/X sky130_fd_sc_hd__mux2_1
X_6026_ _6026_/A _6026_/B _6026_/C _6025_/Y VGND VGND VPWR VPWR _6027_/C sky130_fd_sc_hd__or4b_1
X_3238_ _7169_/Q _7168_/Q VGND VGND VPWR VPWR _3828_/B sky130_fd_sc_hd__nor2_1
XFILLER_74_619 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3169_ _6635_/Q VGND VGND VPWR VPWR _6306_/B sky130_fd_sc_hd__inv_2
XTAP_2118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6928_ _6928_/CLK _6928_/D fanout501/X VGND VGND VPWR VPWR _6928_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_23_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6859_ _7056_/CLK _6859_/D fanout504/X VGND VGND VPWR VPWR _6859_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_13_10 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_183_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_129_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_135_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_112 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold480 _5491_/X VGND VGND VPWR VPWR _7037_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_2_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold491 _6441_/Q VGND VGND VPWR VPWR hold491/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_145_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_295 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1180 _5479_/X VGND VGND VPWR VPWR _7026_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1191 _6946_/Q VGND VGND VPWR VPWR _5389_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_73_652 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_173_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_186_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_624 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_181_292 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4210_ _4210_/A0 _5189_/A1 _4213_/S VGND VGND VPWR VPWR _4210_/X sky130_fd_sc_hd__mux2_1
XFILLER_142_679 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5190_ _5190_/A _5538_/B VGND VGND VPWR VPWR _5198_/S sky130_fd_sc_hd__and2_2
XFILLER_141_178 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4141_ hold935/X _5189_/A1 _4144_/S VGND VGND VPWR VPWR _4141_/X sky130_fd_sc_hd__mux2_1
XFILLER_95_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_110_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4072_ hold630/X _4071_/X _4078_/S VGND VGND VPWR VPWR _4072_/X sky130_fd_sc_hd__mux2_1
XFILLER_83_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_660 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4974_ _4965_/A _4965_/B _4965_/C _4597_/Y VGND VGND VPWR VPWR _4974_/X sky130_fd_sc_hd__a31o_1
X_3925_ _3924_/X input38/X _6405_/Q VGND VGND VPWR VPWR _3925_/X sky130_fd_sc_hd__mux2_1
X_6713_ _6718_/CLK _6713_/D fanout496/X VGND VGND VPWR VPWR _6713_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_149_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6644_ _3931_/A1 _6644_/D _6308_/B VGND VGND VPWR VPWR _6644_/Q sky130_fd_sc_hd__dfrtp_4
X_3856_ _3166_/Y _3247_/A _3856_/S VGND VGND VPWR VPWR _3856_/X sky130_fd_sc_hd__mux2_1
XFILLER_50_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6575_ _7140_/CLK _6575_/D VGND VGND VPWR VPWR _6575_/Q sky130_fd_sc_hd__dfxtp_1
X_3787_ input93/X _3300_/Y _3317_/Y _5511_/A _7055_/Q VGND VGND VPWR VPWR _3787_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_118_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5526_ hold345/X _5526_/A1 _5528_/S VGND VGND VPWR VPWR _5526_/X sky130_fd_sc_hd__mux2_1
XFILLER_117_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_118_687 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5457_ hold721/X _5457_/A1 _5459_/S VGND VGND VPWR VPWR _5457_/X sky130_fd_sc_hd__mux2_1
XFILLER_105_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4408_ _4542_/A _4409_/B VGND VGND VPWR VPWR _4573_/A sky130_fd_sc_hd__and2b_2
XFILLER_182_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5388_ _5388_/A _5529_/B VGND VGND VPWR VPWR _5396_/S sky130_fd_sc_hd__and2_4
XFILLER_87_700 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_571 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7127_ _7130_/CLK _7127_/D fanout488/X VGND VGND VPWR VPWR _7127_/Q sky130_fd_sc_hd__dfrtp_1
X_4339_ _4679_/A _4542_/A VGND VGND VPWR VPWR _4575_/B sky130_fd_sc_hd__or2_2
XFILLER_115_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7058_ _7058_/CLK _7058_/D fanout522/X VGND VGND VPWR VPWR _7058_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_86_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6009_ _6819_/Q _5969_/A _5951_/X _7072_/Q _6008_/X VGND VGND VPWR VPWR _6009_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_55_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_171_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_156_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_156_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_124_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_722 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_370 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_387 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_150 _5532_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_655 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_161 hold23/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_172 _4261_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_183 _5972_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_194 input45/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3710_ input35/X _3360_/Y _4196_/A _6605_/Q _3709_/X VGND VGND VPWR VPWR _3711_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_147_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4690_ _5043_/A _4719_/B VGND VGND VPWR VPWR _4718_/A sky130_fd_sc_hd__nor2_1
XFILLER_159_576 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3641_ _6611_/Q _4202_/A _4261_/A _6667_/Q _3640_/X VGND VGND VPWR VPWR _3648_/A
+ sky130_fd_sc_hd__a221o_1
X_6360_ _6399_/A _6399_/B VGND VGND VPWR VPWR _6360_/X sky130_fd_sc_hd__and2_1
XFILLER_60_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3572_ _3797_/A _5183_/A VGND VGND VPWR VPWR _3572_/Y sky130_fd_sc_hd__nor2_2
X_5311_ hold739/X _5542_/A1 _5315_/S VGND VGND VPWR VPWR _5311_/X sky130_fd_sc_hd__mux2_1
X_6291_ _6459_/Q _6291_/A2 _5975_/C _6704_/Q _6290_/X VGND VGND VPWR VPWR _6292_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_142_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_170_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5242_ hold209/X hold114/X _5243_/S VGND VGND VPWR VPWR _5242_/X sky130_fd_sc_hd__mux2_1
XFILLER_114_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_102_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_30_csclk clkbuf_3_7_0_csclk/X VGND VGND VPWR VPWR _7042_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_69_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5173_ hold146/X hold23/X _5178_/S VGND VGND VPWR VPWR _5173_/X sky130_fd_sc_hd__mux2_1
XFILLER_69_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4124_ hold831/X _6355_/A1 _4126_/S VGND VGND VPWR VPWR _4124_/X sky130_fd_sc_hd__mux2_1
XFILLER_68_287 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput1 debug_mode VGND VGND VPWR VPWR input1/X sky130_fd_sc_hd__clkbuf_2
X_4055_ hold287/X _4054_/X _4061_/S VGND VGND VPWR VPWR _4055_/X sky130_fd_sc_hd__mux2_1
XFILLER_37_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_45_csclk clkbuf_3_6_0_csclk/X VGND VGND VPWR VPWR _6948_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_37_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_460 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4957_ _4489_/B _4832_/Y _4947_/X _4956_/Y _4920_/A VGND VGND VPWR VPWR _4958_/B
+ sky130_fd_sc_hd__a2111o_1
XFILLER_52_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3908_ _6635_/Q _3908_/B VGND VGND VPWR VPWR _3908_/Y sky130_fd_sc_hd__nand2_1
XFILLER_165_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4888_ _4888_/A _4888_/B _4895_/A VGND VGND VPWR VPWR _4892_/B sky130_fd_sc_hd__or3b_4
XFILLER_20_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3839_ _3838_/X _3839_/A1 _3857_/S VGND VGND VPWR VPWR _6413_/D sky130_fd_sc_hd__mux2_1
X_6627_ _6633_/CLK _6627_/D _6370_/A VGND VGND VPWR VPWR _6627_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_137_248 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_343 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6558_ _6698_/CLK _6558_/D fanout495/X VGND VGND VPWR VPWR _6558_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_192_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5509_ hold203/X hold114/X _5510_/S VGND VGND VPWR VPWR _5509_/X sky130_fd_sc_hd__mux2_1
XFILLER_145_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6489_ _7171_/CLK _6489_/D _6378_/X VGND VGND VPWR VPWR _6489_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_106_679 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_168_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_183_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_183_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_109_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_136_270 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_238 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5860_ _6551_/Q _5639_/X _5647_/X _6456_/Q VGND VGND VPWR VPWR _5860_/X sky130_fd_sc_hd__a22o_1
XFILLER_179_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4811_ _4921_/A _4988_/B _4795_/X _4810_/X _5110_/A VGND VGND VPWR VPWR _4812_/D
+ sky130_fd_sc_hd__o2111a_1
XTAP_2290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5791_ _6984_/Q _5642_/X _5644_/X _6976_/Q _5782_/Y VGND VGND VPWR VPWR _5791_/X
+ sky130_fd_sc_hd__a221o_2
XFILLER_61_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4742_ _4549_/B _4515_/B _4972_/A _4703_/A VGND VGND VPWR VPWR _4742_/X sky130_fd_sc_hd__o22a_1
XFILLER_147_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_187_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4673_ _5043_/A _4678_/A VGND VGND VPWR VPWR _4673_/Y sky130_fd_sc_hd__nor2_1
XFILLER_174_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6412_ _3500_/A1 _6412_/D _6368_/X VGND VGND VPWR VPWR hold56/A sky130_fd_sc_hd__dfrtp_1
X_3624_ _3624_/A _3624_/B _3624_/C VGND VGND VPWR VPWR _3624_/X sky130_fd_sc_hd__and3_1
XFILLER_174_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_174_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6343_ _6342_/X _6343_/A1 _6346_/S VGND VGND VPWR VPWR _7147_/D sky130_fd_sc_hd__mux2_1
X_3555_ _6709_/Q _4309_/A _4020_/A _6469_/Q VGND VGND VPWR VPWR _3555_/X sky130_fd_sc_hd__a22o_1
XFILLER_127_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6274_ _6548_/Q _5948_/X _5971_/B _6612_/Q VGND VGND VPWR VPWR _6274_/X sky130_fd_sc_hd__a22o_1
XFILLER_88_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3486_ _7043_/Q _5493_/A _4321_/A _6719_/Q VGND VGND VPWR VPWR _3486_/X sky130_fd_sc_hd__a22o_1
XFILLER_142_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5225_ hold545/X _5519_/A1 _5225_/S VGND VGND VPWR VPWR _5225_/X sky130_fd_sc_hd__mux2_1
X_5156_ hold469/X _5534_/A1 _5157_/S VGND VGND VPWR VPWR _5156_/X sky130_fd_sc_hd__mux2_1
XFILLER_96_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4107_ hold769/X _5542_/A1 _4111_/S VGND VGND VPWR VPWR _4107_/X sky130_fd_sc_hd__mux2_1
XFILLER_29_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5087_ _5087_/A _5087_/B _5087_/C _5087_/D VGND VGND VPWR VPWR _5121_/B sky130_fd_sc_hd__and4_1
X_4038_ _4038_/A hold7/X VGND VGND VPWR VPWR _4043_/S sky130_fd_sc_hd__and2_4
XFILLER_25_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5989_ _6898_/Q _5950_/X _5972_/B _7055_/Q VGND VGND VPWR VPWR _5989_/X sky130_fd_sc_hd__a22o_1
XPHY_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_50 _5369_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_61 _5975_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_72 _6406_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_193_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_21 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_83 user_clock VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_94 _3943_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_153_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_180_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput190 _3197_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[23] sky130_fd_sc_hd__buf_12
XFILLER_153_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_178_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_129_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_156_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_674 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold309 _6719_/Q VGND VGND VPWR VPWR hold309/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_109_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3340_ _6425_/Q _3958_/A _3339_/Y input33/X _3334_/X VGND VGND VPWR VPWR _3348_/A
+ sky130_fd_sc_hd__a221o_2
Xclkbuf_3_4_0_wb_clk_i clkbuf_3_5_0_wb_clk_i/A VGND VGND VPWR VPWR _7137_/CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_125_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_152_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3271_ hold56/X _3856_/S hold14/X VGND VGND VPWR VPWR hold57/A sky130_fd_sc_hd__a21o_1
XFILLER_98_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5010_ _5010_/A _5010_/B VGND VGND VPWR VPWR _5074_/C sky130_fd_sc_hd__nor2_1
XTAP_669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1009 _4016_/X VGND VGND VPWR VPWR _6461_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_23_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_319 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6961_ _6961_/CLK _6961_/D fanout521/X VGND VGND VPWR VPWR _6961_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_81_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5912_ _7155_/Q _5912_/A2 _5912_/B1 _6459_/Q VGND VGND VPWR VPWR _5912_/X sky130_fd_sc_hd__a22o_1
XFILLER_34_430 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6892_ _7083_/CLK _6892_/D fanout517/X VGND VGND VPWR VPWR _6892_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_34_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5843_ _6540_/Q _5667_/X _5832_/X _5842_/X _5610_/A VGND VGND VPWR VPWR _5843_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_21_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5774_ _6839_/Q _5928_/A2 _5926_/A2 _6807_/Q _5773_/X VGND VGND VPWR VPWR _5774_/X
+ sky130_fd_sc_hd__a221o_1
X_4725_ _4789_/B _4725_/B VGND VGND VPWR VPWR _4725_/X sky130_fd_sc_hd__or2_1
XFILLER_135_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4656_ _4656_/A _4902_/A _4656_/C _4656_/D VGND VGND VPWR VPWR _4664_/C sky130_fd_sc_hd__and4_1
XFILLER_174_151 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput70 mgmt_gpio_in[7] VGND VGND VPWR VPWR _3953_/B sky130_fd_sc_hd__clkbuf_4
X_3607_ _6429_/Q _3975_/A _4297_/A _6698_/Q _3606_/X VGND VGND VPWR VPWR _3614_/A
+ sky130_fd_sc_hd__a221o_1
Xinput81 spi_sdo VGND VGND VPWR VPWR input81/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold810 _4005_/X VGND VGND VPWR VPWR _6452_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold821 _6552_/Q VGND VGND VPWR VPWR hold821/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4587_ _4587_/A _5026_/A VGND VGND VPWR VPWR _4933_/A sky130_fd_sc_hd__or2_1
XFILLER_190_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold832 _4124_/X VGND VGND VPWR VPWR _6542_/D sky130_fd_sc_hd__dlygate4sd3_1
Xinput92 spimemio_flash_io3_oeb VGND VGND VPWR VPWR input92/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold843 _6477_/Q VGND VGND VPWR VPWR hold843/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_190_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold854 _5243_/X VGND VGND VPWR VPWR _6817_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3538_ _3761_/A _3538_/B VGND VGND VPWR VPWR _4267_/A sky130_fd_sc_hd__nor2_4
X_6326_ _6642_/Q _6326_/A2 _6326_/B1 _6643_/Q VGND VGND VPWR VPWR _6326_/X sky130_fd_sc_hd__a22o_1
Xhold865 _6629_/Q VGND VGND VPWR VPWR hold865/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold876 _4263_/X VGND VGND VPWR VPWR _6666_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold887 _6706_/Q VGND VGND VPWR VPWR hold887/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_131_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold898 _4236_/X VGND VGND VPWR VPWR _6634_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6257_ _6658_/Q _6288_/A2 _5952_/Y _7154_/Q _6256_/X VGND VGND VPWR VPWR _6257_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_67_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3469_ _7023_/Q hold18/A _5190_/A input57/X _3468_/X VGND VGND VPWR VPWR _3470_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_131_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5208_ _5208_/A _5529_/B VGND VGND VPWR VPWR _5216_/S sky130_fd_sc_hd__and2_4
XFILLER_103_479 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_190_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6188_ _6475_/Q _5976_/Y _5979_/X _6450_/Q _6185_/X VGND VGND VPWR VPWR _6202_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_130_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1510 _6641_/Q VGND VGND VPWR VPWR _3168_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1521 _6721_/Q VGND VGND VPWR VPWR _4882_/B2 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_69_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1532 _7126_/Q VGND VGND VPWR VPWR _6180_/A1 sky130_fd_sc_hd__dlygate4sd3_1
X_5139_ _5120_/B _5138_/X _6726_/Q _4222_/X VGND VGND VPWR VPWR _5139_/X sky130_fd_sc_hd__a2bb2o_1
Xhold1543 _7100_/Q VGND VGND VPWR VPWR _5595_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_96_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1554 _7185_/A VGND VGND VPWR VPWR hold287/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_45_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_514 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_357 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_240 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_180_176 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_555 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_322 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4510_ _4510_/A _4510_/B _4510_/C VGND VGND VPWR VPWR _4510_/X sky130_fd_sc_hd__and3_1
XFILLER_117_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5490_ hold779/X _6355_/A1 _5492_/S VGND VGND VPWR VPWR _5490_/X sky130_fd_sc_hd__mux2_1
Xhold106 _3267_/X VGND VGND VPWR VPWR hold106/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_156_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4441_ _4789_/A _4862_/A VGND VGND VPWR VPWR _5048_/A sky130_fd_sc_hd__nor2_1
Xhold117 _5198_/X VGND VGND VPWR VPWR _6777_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_144_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold128 _6992_/Q VGND VGND VPWR VPWR hold128/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold139 _5197_/X VGND VGND VPWR VPWR _6776_/D sky130_fd_sc_hd__dlygate4sd3_1
X_7160_ net499_2/A _7160_/D _6390_/X VGND VGND VPWR VPWR hold88/A sky130_fd_sc_hd__dfrtp_1
X_4372_ _4346_/A _4346_/B _4545_/A VGND VGND VPWR VPWR _4885_/A sky130_fd_sc_hd__o21ai_4
XFILLER_98_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_171_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6111_ _6799_/Q _6299_/A2 _5974_/B _6831_/Q VGND VGND VPWR VPWR _6111_/X sky130_fd_sc_hd__a22o_1
X_3323_ _6921_/Q _5352_/A _3975_/A _6433_/Q _3322_/X VGND VGND VPWR VPWR _3349_/B
+ sky130_fd_sc_hd__a221o_1
XTAP_411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7091_ _7124_/CLK _7091_/D fanout502/X VGND VGND VPWR VPWR _7091_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_112_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6042_ _6042_/A _6042_/B VGND VGND VPWR VPWR _6042_/Y sky130_fd_sc_hd__nor2_1
XFILLER_98_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3254_ _3255_/A1 _3254_/A1 _3256_/S VGND VGND VPWR VPWR _7162_/D sky130_fd_sc_hd__mux2_1
XTAP_466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3185_ _7066_/Q VGND VGND VPWR VPWR _3185_/Y sky130_fd_sc_hd__inv_2
XFILLER_26_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6944_ _7072_/CLK _6944_/D fanout506/X VGND VGND VPWR VPWR _6944_/Q sky130_fd_sc_hd__dfrtp_1
X_6875_ _7011_/CLK _6875_/D fanout500/X VGND VGND VPWR VPWR _6875_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_167_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5826_ _6625_/Q _5913_/B1 _5649_/X _6675_/Q VGND VGND VPWR VPWR _5826_/X sky130_fd_sc_hd__a22o_1
XFILLER_22_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_499 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5757_ _5757_/A1 _6305_/A2 _5755_/X _5756_/X VGND VGND VPWR VPWR _7110_/D sky130_fd_sc_hd__o22a_1
X_4708_ _4717_/B _4715_/B _5005_/B _4394_/Y VGND VGND VPWR VPWR _4708_/X sky130_fd_sc_hd__a31o_1
X_5688_ _6835_/Q _5617_/X _5683_/X _5687_/X VGND VGND VPWR VPWR _5688_/X sky130_fd_sc_hd__a211o_1
XFILLER_147_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4639_ _4962_/C _4630_/B _4456_/Y VGND VGND VPWR VPWR _4639_/X sky130_fd_sc_hd__o21a_1
XFILLER_190_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold640 _6473_/Q VGND VGND VPWR VPWR hold640/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_78_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold651 _5186_/X VGND VGND VPWR VPWR _6767_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold662 _6763_/Q VGND VGND VPWR VPWR _5179_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_1_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmax_cap370 _3374_/A VGND VGND VPWR VPWR _3571_/B sky130_fd_sc_hd__buf_12
Xmax_cap381 _5951_/X VGND VGND VPWR VPWR _6289_/A2 sky130_fd_sc_hd__buf_12
Xhold673 _6847_/Q VGND VGND VPWR VPWR hold673/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_1_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6309_ _3816_/X _6309_/A1 _6316_/S VGND VGND VPWR VPWR _7133_/D sky130_fd_sc_hd__mux2_1
Xhold684 _5250_/X VGND VGND VPWR VPWR _6823_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold695 _6447_/Q VGND VGND VPWR VPWR hold695/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_77_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_55 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1340 hold1340/A VGND VGND VPWR VPWR wb_dat_o[12] sky130_fd_sc_hd__buf_12
XFILLER_45_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1351 _4184_/A1 VGND VGND VPWR VPWR hold1351/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_91_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1362 hold1362/A VGND VGND VPWR VPWR wb_dat_o[27] sky130_fd_sc_hd__buf_12
XFILLER_84_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1373 _7190_/A VGND VGND VPWR VPWR _5192_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_150_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_175_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1384 _6876_/Q VGND VGND VPWR VPWR _5310_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_84_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1395 _6572_/Q VGND VGND VPWR VPWR hold1395/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_186_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_159_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_622 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_474 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xnet499_2 net499_2/A VGND VGND VPWR VPWR _3935_/B sky130_fd_sc_hd__inv_2
X_4990_ _4581_/A _4547_/X _4989_/X VGND VGND VPWR VPWR _4991_/B sky130_fd_sc_hd__o21ai_1
XFILLER_91_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3941_ _6404_/Q _3941_/B VGND VGND VPWR VPWR _3942_/A sky130_fd_sc_hd__nand2b_1
XFILLER_51_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_189_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_149_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6660_ _6695_/CLK _6660_/D fanout490/X VGND VGND VPWR VPWR _6660_/Q sky130_fd_sc_hd__dfrtp_1
X_3872_ _6643_/Q _3869_/X _3872_/B1 VGND VGND VPWR VPWR _6643_/D sky130_fd_sc_hd__a21o_1
XFILLER_32_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_189_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5611_ _5612_/A _5612_/B VGND VGND VPWR VPWR _5611_/X sky130_fd_sc_hd__and2_2
XFILLER_149_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_176_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6591_ _7130_/CLK _6591_/D VGND VGND VPWR VPWR _6591_/Q sky130_fd_sc_hd__dfxtp_1
X_5542_ hold713/X _5542_/A1 _5546_/S VGND VGND VPWR VPWR _5542_/X sky130_fd_sc_hd__mux2_1
XFILLER_192_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_129_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5473_ hold733/X _5542_/A1 hold19/X VGND VGND VPWR VPWR _5473_/X sky130_fd_sc_hd__mux2_1
XFILLER_144_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4424_ _4535_/A _4946_/A VGND VGND VPWR VPWR _4828_/A sky130_fd_sc_hd__nand2_4
X_7143_ _7150_/CLK _7143_/D _6308_/B VGND VGND VPWR VPWR hold10/A sky130_fd_sc_hd__dfrtp_1
X_4355_ _4679_/A _4542_/A _4554_/A _4596_/B _4614_/A VGND VGND VPWR VPWR _4357_/B
+ sky130_fd_sc_hd__o2111a_1
XFILLER_113_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout427 _4631_/A VGND VGND VPWR VPWR _4678_/A sky130_fd_sc_hd__buf_6
XFILLER_86_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3306_ _7017_/Q _5460_/A hold18/A _7025_/Q VGND VGND VPWR VPWR _3306_/X sky130_fd_sc_hd__a22o_1
X_7074_ _7074_/CLK _7074_/D fanout505/X VGND VGND VPWR VPWR _7074_/Q sky130_fd_sc_hd__dfrtp_4
Xfanout438 hold141/X VGND VGND VPWR VPWR hold142/A sky130_fd_sc_hd__buf_8
X_4286_ _4286_/A0 _5308_/A1 _4290_/S VGND VGND VPWR VPWR _4286_/X sky130_fd_sc_hd__mux2_1
Xfanout449 hold46/X VGND VGND VPWR VPWR _5515_/A1 sky130_fd_sc_hd__buf_8
XFILLER_113_596 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_382 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6025_ _6025_/A _6025_/B VGND VGND VPWR VPWR _6025_/Y sky130_fd_sc_hd__nor2_1
X_3237_ _6415_/Q _3259_/B VGND VGND VPWR VPWR _3867_/A sky130_fd_sc_hd__nand2_2
XFILLER_39_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_374 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3168_ _3168_/A VGND VGND VPWR VPWR _3903_/A sky130_fd_sc_hd__inv_2
XTAP_2108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6927_ _7031_/CLK _6927_/D fanout522/X VGND VGND VPWR VPWR _6927_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_23_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6858_ _7055_/CLK _6858_/D fanout504/X VGND VGND VPWR VPWR _6858_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_13_22 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5809_ _6873_/Q _5625_/X _5643_/X _6889_/Q VGND VGND VPWR VPWR _5809_/X sky130_fd_sc_hd__a22o_1
X_6789_ _6789_/CLK _6789_/D fanout497/X VGND VGND VPWR VPWR _6789_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_167_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_163_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_135_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_136_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_647 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold470 _5156_/X VGND VGND VPWR VPWR _6746_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold481 _6512_/Q VGND VGND VPWR VPWR hold481/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold492 _3992_/X VGND VGND VPWR VPWR _6441_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_2_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_131_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1170 _4274_/X VGND VGND VPWR VPWR _6675_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_85_491 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1181 _6994_/Q VGND VGND VPWR VPWR _5443_/A0 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1192 _5389_/X VGND VGND VPWR VPWR _6946_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_146_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_186_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_141_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4140_ _4140_/A0 _5308_/A1 _4144_/S VGND VGND VPWR VPWR _4140_/X sky130_fd_sc_hd__mux2_1
XFILLER_110_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4071_ hold379/X _5534_/A1 _4077_/S VGND VGND VPWR VPWR _4071_/X sky130_fd_sc_hd__mux2_1
XFILLER_49_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_491 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4973_ _4973_/A _4973_/B VGND VGND VPWR VPWR _4973_/X sky130_fd_sc_hd__or2_1
X_6712_ _6718_/CLK _6712_/D _6401_/A VGND VGND VPWR VPWR _6712_/Q sky130_fd_sc_hd__dfstp_1
X_3924_ _6499_/Q _6734_/Q _6399_/B VGND VGND VPWR VPWR _3924_/X sky130_fd_sc_hd__mux2_1
XFILLER_189_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_189_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6643_ _7150_/CLK _6643_/D _6308_/B VGND VGND VPWR VPWR _6643_/Q sky130_fd_sc_hd__dfrtp_4
X_3855_ _3857_/A1 _3854_/Y _3853_/X VGND VGND VPWR VPWR _6408_/D sky130_fd_sc_hd__a21o_1
XFILLER_164_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3786_ _7047_/Q _5502_/A _3572_/Y input98/X _3785_/X VGND VGND VPWR VPWR _3792_/B
+ sky130_fd_sc_hd__a221o_1
X_6574_ _7137_/CLK _6574_/D VGND VGND VPWR VPWR _6574_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_117_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5525_ _5525_/A0 _5543_/A1 _5528_/S VGND VGND VPWR VPWR _5525_/X sky130_fd_sc_hd__mux2_1
XFILLER_118_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5456_ _5456_/A0 _5543_/A1 _5459_/S VGND VGND VPWR VPWR _5456_/X sky130_fd_sc_hd__mux2_1
XFILLER_132_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4407_ _4472_/A _4946_/A VGND VGND VPWR VPWR _4407_/X sky130_fd_sc_hd__and2b_1
X_5387_ hold909/X _5537_/A1 _5387_/S VGND VGND VPWR VPWR _5387_/X sky130_fd_sc_hd__mux2_1
XFILLER_99_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_160_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7126_ _7131_/CLK _7126_/D fanout501/X VGND VGND VPWR VPWR _7126_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_99_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_113_371 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4338_ _4679_/A _4542_/A VGND VGND VPWR VPWR _4595_/B sky130_fd_sc_hd__nor2_1
XFILLER_113_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4269_ hold959/X _5189_/A1 _4272_/S VGND VGND VPWR VPWR _4269_/X sky130_fd_sc_hd__mux2_1
X_7057_ _7079_/CLK _7057_/D fanout514/X VGND VGND VPWR VPWR _7057_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_46_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6008_ _7080_/Q _6294_/A2 _6294_/B1 _7040_/Q VGND VGND VPWR VPWR _6008_/X sky130_fd_sc_hd__a22o_1
XFILLER_54_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_78 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_183_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_734 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_172_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_93_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_140 _5918_/B1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_151 _5505_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_162 hold23/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_173 _5142_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_184 _5972_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_195 input43/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_159_588 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3640_ _6836_/Q _5262_/A _4166_/A _6580_/Q VGND VGND VPWR VPWR _3640_/X sky130_fd_sc_hd__a22o_1
X_3571_ _3571_/A _3571_/B VGND VGND VPWR VPWR _5163_/A sky130_fd_sc_hd__nor2_8
XFILLER_115_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_400 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5310_ _5310_/A0 hold3/X _5315_/S VGND VGND VPWR VPWR hold4/A sky130_fd_sc_hd__mux2_1
XFILLER_53_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6290_ _7155_/Q _6290_/A2 _6290_/B1 _6469_/Q VGND VGND VPWR VPWR _6290_/X sky130_fd_sc_hd__a22o_1
XFILLER_5_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5241_ hold685/X _5544_/A1 _5243_/S VGND VGND VPWR VPWR _5241_/X sky130_fd_sc_hd__mux2_1
XFILLER_142_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5172_ _5179_/B _5529_/B VGND VGND VPWR VPWR _5178_/S sky130_fd_sc_hd__and2_2
X_4123_ _4123_/A0 _6354_/A1 _4126_/S VGND VGND VPWR VPWR _4123_/X sky130_fd_sc_hd__mux2_1
XFILLER_29_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput2 debug_oeb VGND VGND VPWR VPWR input2/X sky130_fd_sc_hd__clkbuf_1
X_4054_ hold134/X hold23/X _4103_/B VGND VGND VPWR VPWR _4054_/X sky130_fd_sc_hd__mux2_1
XFILLER_68_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_opt_1_0_csclk _7000_/CLK VGND VGND VPWR VPWR clkbuf_opt_1_0_csclk/X sky130_fd_sc_hd__clkbuf_16
XFILLER_71_409 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4956_ _4581_/A _5026_/B _4955_/X VGND VGND VPWR VPWR _4956_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_189_190 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_199 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3907_ _3240_/A _3867_/Y _3858_/B _3856_/S VGND VGND VPWR VPWR _6487_/D sky130_fd_sc_hd__a2bb2o_1
XFILLER_177_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4887_ _4888_/A _4888_/B _4886_/Y _4742_/X VGND VGND VPWR VPWR _5008_/D sky130_fd_sc_hd__o31a_1
XFILLER_192_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6626_ _6686_/CLK _6626_/D fanout492/X VGND VGND VPWR VPWR _6626_/Q sky130_fd_sc_hd__dfrtp_2
X_3838_ hold56/A _3856_/S _3837_/X VGND VGND VPWR VPWR _3838_/X sky130_fd_sc_hd__a21o_1
XFILLER_192_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6557_ _6689_/CLK _6557_/D fanout509/X VGND VGND VPWR VPWR _6557_/Q sky130_fd_sc_hd__dfrtp_4
X_3769_ input43/X _3343_/Y _4267_/A _6670_/Q VGND VGND VPWR VPWR _3769_/X sky130_fd_sc_hd__a22o_1
XFILLER_4_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5508_ hold439/X _5526_/A1 _5510_/S VGND VGND VPWR VPWR _5508_/X sky130_fd_sc_hd__mux2_1
XFILLER_193_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6488_ _7171_/CLK _6488_/D _6377_/X VGND VGND VPWR VPWR _6488_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_105_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5439_ hold723/X _5457_/A1 hold35/X VGND VGND VPWR VPWR _5439_/X sky130_fd_sc_hd__mux2_1
XFILLER_105_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7109_ _7123_/CLK _7109_/D fanout497/X VGND VGND VPWR VPWR _7109_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_47_428 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_472 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_136_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_183_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_183_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_707 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_179_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4810_ _4678_/A _4725_/B _4615_/B _4587_/A _4640_/B VGND VGND VPWR VPWR _4810_/X
+ sky130_fd_sc_hd__o32a_1
XTAP_2291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5790_ _6944_/Q _5816_/B1 _5784_/X _5789_/X VGND VGND VPWR VPWR _5790_/X sky130_fd_sc_hd__a211o_1
XFILLER_33_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_159_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4741_ _4901_/B _4973_/A _4768_/C VGND VGND VPWR VPWR _4741_/X sky130_fd_sc_hd__o21a_1
XFILLER_193_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4672_ _4703_/A _4672_/B VGND VGND VPWR VPWR _4672_/X sky130_fd_sc_hd__or2_1
X_6411_ _3500_/A1 _6411_/D _6367_/X VGND VGND VPWR VPWR hold29/A sky130_fd_sc_hd__dfrtp_1
XFILLER_135_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3623_ _3623_/A _3623_/B _3623_/C _3623_/D VGND VGND VPWR VPWR _3624_/C sky130_fd_sc_hd__nor4_1
XFILLER_174_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6342_ _6642_/Q _6342_/A2 _6342_/B1 _4222_/B _6341_/X VGND VGND VPWR VPWR _6342_/X
+ sky130_fd_sc_hd__a221o_1
X_3554_ _3554_/A _3554_/B VGND VGND VPWR VPWR _4020_/A sky130_fd_sc_hd__nor2_8
XFILLER_155_591 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6273_ _6563_/Q _5969_/A _5957_/X _6708_/Q VGND VGND VPWR VPWR _6273_/X sky130_fd_sc_hd__a22o_1
X_3485_ _3503_/A _5161_/B VGND VGND VPWR VPWR _4321_/A sky130_fd_sc_hd__nor2_8
XFILLER_103_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_639 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5224_ hold642/X _5545_/A1 _5225_/S VGND VGND VPWR VPWR _5224_/X sky130_fd_sc_hd__mux2_1
XFILLER_102_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5155_ hold517/X _5491_/A1 _5157_/S VGND VGND VPWR VPWR _5155_/X sky130_fd_sc_hd__mux2_1
XFILLER_29_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4106_ hold293/X _5541_/A1 _4111_/S VGND VGND VPWR VPWR _4106_/X sky130_fd_sc_hd__mux2_1
X_5086_ _5118_/B _5118_/C _5085_/X _5119_/A VGND VGND VPWR VPWR _5086_/X sky130_fd_sc_hd__o31a_1
XFILLER_84_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4037_ hold881/X _4236_/A1 _4037_/S VGND VGND VPWR VPWR _4037_/X sky130_fd_sc_hd__mux2_1
XFILLER_37_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5988_ _6842_/Q _5939_/X _5955_/X _6962_/Q _5987_/X VGND VGND VPWR VPWR _6002_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_12_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_486 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4939_ _5064_/A _4939_/B _4939_/C VGND VGND VPWR VPWR _4940_/D sky130_fd_sc_hd__and3_1
XFILLER_178_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_40 _4285_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_51 _5369_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_177_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_193_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_62 _6103_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_73 _6406_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6609_ _6769_/CLK _6609_/D fanout492/X VGND VGND VPWR VPWR _6609_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_126_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_84 user_clock VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_192_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_33 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_95 _3943_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_153_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_192_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_33 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_161_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput180 _3207_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[14] sky130_fd_sc_hd__buf_12
XFILLER_121_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_21 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput191 _3196_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[24] sky130_fd_sc_hd__buf_12
XFILLER_0_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_203 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_686 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_388 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_44_csclk clkbuf_3_6_0_csclk/X VGND VGND VPWR VPWR _7080_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_109_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_140_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3270_ hold30/X _3270_/A1 _6624_/Q VGND VGND VPWR VPWR hold31/A sky130_fd_sc_hd__mux2_2
XTAP_626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_59_csclk clkbuf_3_2_0_csclk/X VGND VGND VPWR VPWR _7046_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_97_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6960_ _6961_/CLK _6960_/D fanout521/X VGND VGND VPWR VPWR _6960_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_81_515 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5911_ _5911_/A1 _6305_/A2 _5909_/X _5910_/X VGND VGND VPWR VPWR _7117_/D sky130_fd_sc_hd__o22a_1
X_6891_ _6976_/CLK _6891_/D fanout497/X VGND VGND VPWR VPWR _6891_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_34_442 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5842_ _5842_/A _5842_/B _5842_/C _5841_/Y VGND VGND VPWR VPWR _5842_/X sky130_fd_sc_hd__or4b_1
XFILLER_61_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5773_ _7023_/Q _5929_/B1 _5915_/B1 _6863_/Q VGND VGND VPWR VPWR _5773_/X sky130_fd_sc_hd__a22o_1
XFILLER_21_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4724_ _4732_/B _4724_/B _4724_/C _4723_/X VGND VGND VPWR VPWR _4726_/C sky130_fd_sc_hd__or4b_1
XFILLER_187_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4655_ _4862_/A _4649_/A _4962_/C _4972_/A VGND VGND VPWR VPWR _4656_/D sky130_fd_sc_hd__o22a_1
XFILLER_135_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_190_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold800 _4276_/X VGND VGND VPWR VPWR _6677_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3606_ _6981_/Q _5424_/A _4014_/A _6463_/Q VGND VGND VPWR VPWR _3606_/X sky130_fd_sc_hd__a22o_1
Xinput60 mgmt_gpio_in[31] VGND VGND VPWR VPWR input60/X sky130_fd_sc_hd__clkbuf_2
Xhold811 _6457_/Q VGND VGND VPWR VPWR hold811/X sky130_fd_sc_hd__dlygate4sd3_1
Xinput71 mgmt_gpio_in[8] VGND VGND VPWR VPWR input71/X sky130_fd_sc_hd__clkbuf_2
XFILLER_190_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput82 spi_sdoenb VGND VGND VPWR VPWR input82/X sky130_fd_sc_hd__dlymetal6s2s_1
X_4586_ _4640_/B _4586_/B VGND VGND VPWR VPWR _5132_/B sky130_fd_sc_hd__or2_1
Xinput93 trap VGND VGND VPWR VPWR input93/X sky130_fd_sc_hd__buf_4
Xhold822 _4136_/X VGND VGND VPWR VPWR _6552_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold833 _6606_/Q VGND VGND VPWR VPWR hold833/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold844 _4035_/X VGND VGND VPWR VPWR _6477_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6325_ _6324_/X _6325_/A1 _6346_/S VGND VGND VPWR VPWR _7141_/D sky130_fd_sc_hd__mux2_1
Xhold855 _6913_/Q VGND VGND VPWR VPWR hold855/X sky130_fd_sc_hd__dlygate4sd3_1
X_3537_ _3552_/A _3761_/B VGND VGND VPWR VPWR _4026_/A sky130_fd_sc_hd__nor2_4
XFILLER_116_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_143_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold866 _4230_/X VGND VGND VPWR VPWR _6629_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold877 _6676_/Q VGND VGND VPWR VPWR hold877/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_88_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold888 _4311_/X VGND VGND VPWR VPWR _6706_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold899 _6716_/Q VGND VGND VPWR VPWR hold899/X sky130_fd_sc_hd__dlygate4sd3_1
X_6256_ _6718_/Q _5955_/X _5977_/X _6668_/Q VGND VGND VPWR VPWR _6256_/X sky130_fd_sc_hd__a22o_1
XFILLER_115_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3468_ _7084_/Q _5538_/A _5397_/A _6959_/Q VGND VGND VPWR VPWR _3468_/X sky130_fd_sc_hd__a22o_1
XFILLER_130_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5207_ _5207_/A0 hold27/X _5207_/S VGND VGND VPWR VPWR hold77/A sky130_fd_sc_hd__mux2_1
X_6187_ _6604_/Q wire390/X _6270_/B1 _6675_/Q _6186_/X VGND VGND VPWR VPWR _6187_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_69_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1500 _7107_/Q VGND VGND VPWR VPWR _5691_/A1 sky130_fd_sc_hd__dlygate4sd3_1
X_3399_ _3398_/X _3399_/A1 _3749_/S VGND VGND VPWR VPWR _6734_/D sky130_fd_sc_hd__mux2_1
Xhold1511 _4224_/X VGND VGND VPWR VPWR _6624_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1522 _6720_/Q VGND VGND VPWR VPWR _4730_/B2 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_29_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1533 _6509_/Q VGND VGND VPWR VPWR _3889_/B2 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_57_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5138_ _5084_/X _5138_/B _5138_/C VGND VGND VPWR VPWR _5138_/X sky130_fd_sc_hd__and3b_1
Xhold1544 _7095_/Q VGND VGND VPWR VPWR _5578_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_84_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1555 _6760_/Q VGND VGND VPWR VPWR hold199/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_123_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5069_ _4479_/A _4988_/A _4748_/B _4676_/B _4813_/C VGND VGND VPWR VPWR _5070_/C
+ sky130_fd_sc_hd__o221a_1
XFILLER_72_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_420 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_122 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_369 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_285 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_567 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_180_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_180_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_592 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_129_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_156_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4440_ _4977_/B _4680_/A VGND VGND VPWR VPWR _4862_/A sky130_fd_sc_hd__or2_4
Xhold107 _3268_/X VGND VGND VPWR VPWR _3328_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_171_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_172_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold118 _6961_/Q VGND VGND VPWR VPWR hold118/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_172_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold129 _5440_/X VGND VGND VPWR VPWR _6992_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_171_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4371_ _4368_/A _4544_/A _3891_/A _3891_/B _4707_/B VGND VGND VPWR VPWR _4545_/A
+ sky130_fd_sc_hd__a41o_4
XFILLER_171_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6110_ _6815_/Q _5936_/X _6289_/A2 _7076_/Q _6109_/X VGND VGND VPWR VPWR _6118_/B
+ sky130_fd_sc_hd__a221o_1
X_3322_ _6801_/Q _5217_/A _5493_/A _7046_/Q VGND VGND VPWR VPWR _3322_/X sky130_fd_sc_hd__a22o_1
XTAP_401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7090_ _7131_/CLK _7090_/D fanout502/X VGND VGND VPWR VPWR _7090_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_98_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6041_ _6868_/Q _5971_/A _6285_/B1 _7012_/Q _6040_/X VGND VGND VPWR VPWR _6042_/B
+ sky130_fd_sc_hd__a221o_1
XTAP_456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_575 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3253_ _3254_/A1 hold21/A _3256_/S VGND VGND VPWR VPWR _3253_/X sky130_fd_sc_hd__mux2_1
XFILLER_39_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_112_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3184_ _7074_/Q VGND VGND VPWR VPWR _3184_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_27_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_228 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6943_ _7029_/CLK _6943_/D fanout522/X VGND VGND VPWR VPWR _6943_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_19_291 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_179_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6874_ _7063_/CLK _6874_/D fanout504/X VGND VGND VPWR VPWR _6874_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_179_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_179_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5825_ _6609_/Q _5631_/X _5634_/X _6685_/Q _5824_/X VGND VGND VPWR VPWR _5828_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_50_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5756_ _5756_/A1 _5612_/A _5612_/B VGND VGND VPWR VPWR _5756_/X sky130_fd_sc_hd__o21a_1
X_4707_ _4884_/A _4707_/B _4707_/C VGND VGND VPWR VPWR _4709_/C sky130_fd_sc_hd__and3_1
X_5687_ _6939_/Q _5634_/X _5684_/X _5686_/X VGND VGND VPWR VPWR _5687_/X sky130_fd_sc_hd__a211o_1
XFILLER_135_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_162_100 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4638_ _4799_/B _4638_/B VGND VGND VPWR VPWR _4984_/A sky130_fd_sc_hd__or2_1
XFILLER_190_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold630 hold630/A VGND VGND VPWR VPWR hold630/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold641 _4030_/X VGND VGND VPWR VPWR _6473_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4569_ _4569_/A _4946_/C VGND VGND VPWR VPWR _4569_/X sky130_fd_sc_hd__and2_1
Xmax_cap360 _3361_/Y VGND VGND VPWR VPWR _3993_/A sky130_fd_sc_hd__buf_8
Xhold652 _7079_/Q VGND VGND VPWR VPWR hold652/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold663 _5179_/X VGND VGND VPWR VPWR hold663/X sky130_fd_sc_hd__dlygate4sd3_1
Xmax_cap371 hold33/X VGND VGND VPWR VPWR _3563_/A sky130_fd_sc_hd__buf_12
Xmax_cap382 _5949_/X VGND VGND VPWR VPWR _6283_/A2 sky130_fd_sc_hd__buf_12
X_6308_ _6636_/Q _6308_/B VGND VGND VPWR VPWR _6316_/S sky130_fd_sc_hd__nand2_8
Xhold674 _5277_/X VGND VGND VPWR VPWR _6847_/D sky130_fd_sc_hd__dlygate4sd3_1
Xmax_cap393 _5950_/X VGND VGND VPWR VPWR _6296_/B1 sky130_fd_sc_hd__buf_12
Xhold685 _6815_/Q VGND VGND VPWR VPWR hold685/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_131_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_143_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold696 _3999_/X VGND VGND VPWR VPWR _6447_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_467 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_255 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6239_ _6682_/Q _5949_/X _5980_/Y _6467_/Q VGND VGND VPWR VPWR _6239_/X sky130_fd_sc_hd__a22o_1
XFILLER_76_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_67 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_640 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1330 hold1330/A VGND VGND VPWR VPWR wb_dat_o[14] sky130_fd_sc_hd__buf_12
Xhold1341 _4185_/A1 VGND VGND VPWR VPWR hold1341/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1352 hold1352/A VGND VGND VPWR VPWR wb_dat_o[2] sky130_fd_sc_hd__buf_12
XFILLER_85_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1363 _6309_/A1 VGND VGND VPWR VPWR hold1363/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_18_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_526 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1374 _6531_/Q VGND VGND VPWR VPWR _4111_/A0 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1385 _6993_/Q VGND VGND VPWR VPWR _5441_/A0 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1396 _6439_/Q VGND VGND VPWR VPWR _3990_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_185_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_154_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_154_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_122 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_643 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3940_ _6403_/Q _3940_/B VGND VGND VPWR VPWR _3940_/Y sky130_fd_sc_hd__nor2_1
XFILLER_16_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_149_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3871_ _6642_/Q _3869_/X _3871_/B1 VGND VGND VPWR VPWR _6642_/D sky130_fd_sc_hd__a21o_1
XFILLER_177_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5610_ _5610_/A _6508_/Q VGND VGND VPWR VPWR _5610_/Y sky130_fd_sc_hd__nand2_1
XFILLER_177_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6590_ _7137_/CLK _6590_/D VGND VGND VPWR VPWR _6590_/Q sky130_fd_sc_hd__dfxtp_1
X_5541_ hold277/X _5541_/A1 _5546_/S VGND VGND VPWR VPWR _5541_/X sky130_fd_sc_hd__mux2_1
XFILLER_145_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5472_ _5472_/A0 hold3/X hold19/X VGND VGND VPWR VPWR hold20/A sky130_fd_sc_hd__mux2_1
XFILLER_184_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4423_ _4574_/A _4946_/A VGND VGND VPWR VPWR _4490_/B sky130_fd_sc_hd__nand2_1
XFILLER_132_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_160_615 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7142_ _3931_/A1 _7142_/D _6308_/B VGND VGND VPWR VPWR hold92/A sky130_fd_sc_hd__dfrtp_1
XFILLER_125_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4354_ _4614_/A _4356_/B VGND VGND VPWR VPWR _4357_/A sky130_fd_sc_hd__nor2_1
XFILLER_98_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_113_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3305_ hold33/A _3706_/A VGND VGND VPWR VPWR hold18/A sky130_fd_sc_hd__nor2_8
X_7073_ _7073_/CLK _7073_/D fanout498/X VGND VGND VPWR VPWR _7073_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_59_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout439 hold23/X VGND VGND VPWR VPWR _5534_/A1 sky130_fd_sc_hd__buf_12
X_4285_ _4285_/A hold7/X VGND VGND VPWR VPWR _4290_/S sky130_fd_sc_hd__and2_2
X_6024_ _6843_/Q _5939_/X _5953_/Y _6995_/Q _6023_/X VGND VGND VPWR VPWR _6025_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_140_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3236_ _6417_/Q _6416_/Q _6415_/Q VGND VGND VPWR VPWR _3858_/B sky130_fd_sc_hd__and3_2
XFILLER_67_651 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3167_ _6638_/Q VGND VGND VPWR VPWR _3167_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_39_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6926_ _7059_/CLK _6926_/D fanout517/X VGND VGND VPWR VPWR _6926_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_54_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6857_ _7070_/CLK _6857_/D fanout507/X VGND VGND VPWR VPWR _6857_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_23_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5808_ _6929_/Q _5633_/X _5646_/X _7001_/Q VGND VGND VPWR VPWR _5808_/X sky130_fd_sc_hd__a22o_1
XFILLER_167_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6788_ _7073_/CLK _6788_/D fanout497/X VGND VGND VPWR VPWR _6788_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_13_34 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_707 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5739_ _6814_/Q _5913_/A2 _5816_/B1 _6942_/Q _5738_/X VGND VGND VPWR VPWR _5740_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_129_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_145_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold460 _4314_/X VGND VGND VPWR VPWR _6709_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_151_659 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold471 _6544_/Q VGND VGND VPWR VPWR hold471/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_145_44 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold482 _4085_/X VGND VGND VPWR VPWR _6512_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_150_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold493 hold493/A VGND VGND VPWR VPWR hold493/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_38_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1160 _5366_/X VGND VGND VPWR VPWR _6926_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1171 _6645_/Q VGND VGND VPWR VPWR _4238_/A0 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1182 _5443_/X VGND VGND VPWR VPWR _6994_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1193 _6604_/Q VGND VGND VPWR VPWR _4197_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_2_2__f_mgmt_gpio_in[4] clkbuf_0_mgmt_gpio_in[4]/X VGND VGND VPWR VPWR _3500_/A1
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_141_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_150_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4070_ hold357/X _4069_/X _4078_/S VGND VGND VPWR VPWR _4070_/X sky130_fd_sc_hd__mux2_1
XFILLER_96_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4972_ _4972_/A _4973_/B VGND VGND VPWR VPWR _4972_/X sky130_fd_sc_hd__or2_1
XFILLER_51_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6711_ _6711_/CLK _6711_/D _3940_/B VGND VGND VPWR VPWR _6711_/Q sky130_fd_sc_hd__dfrtp_1
X_3923_ _6504_/Q input77/X _3950_/B VGND VGND VPWR VPWR _3923_/X sky130_fd_sc_hd__mux2_4
XFILLER_149_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_149_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6642_ _7150_/CLK _6642_/D _6308_/B VGND VGND VPWR VPWR _6642_/Q sky130_fd_sc_hd__dfrtp_4
X_3854_ hold71/A _3842_/B _3857_/S VGND VGND VPWR VPWR _3854_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_20_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_165_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6573_ _7140_/CLK _6573_/D VGND VGND VPWR VPWR _6573_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_118_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3785_ _7002_/Q _5451_/A _4321_/A _6715_/Q VGND VGND VPWR VPWR _3785_/X sky130_fd_sc_hd__a22o_1
XFILLER_164_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5524_ hold167/X hold46/X _5528_/S VGND VGND VPWR VPWR _5524_/X sky130_fd_sc_hd__mux2_1
XFILLER_118_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_145_431 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_155 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5455_ hold705/X _5542_/A1 _5459_/S VGND VGND VPWR VPWR _5455_/X sky130_fd_sc_hd__mux2_1
XFILLER_145_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_160_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4406_ _4406_/A _4416_/B VGND VGND VPWR VPWR _4946_/A sky130_fd_sc_hd__and2_2
XFILLER_160_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5386_ hold213/X hold114/X _5387_/S VGND VGND VPWR VPWR _5386_/X sky130_fd_sc_hd__mux2_1
XFILLER_99_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7125_ _7131_/CLK _7125_/D fanout501/X VGND VGND VPWR VPWR _7125_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_101_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4337_ _4337_/A _4337_/B _4337_/C VGND VGND VPWR VPWR _4541_/B sky130_fd_sc_hd__and3_1
XFILLER_113_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7056_ _7056_/CLK _7056_/D fanout504/X VGND VGND VPWR VPWR _7056_/Q sky130_fd_sc_hd__dfstp_1
X_4268_ _4268_/A0 _5308_/A1 _4272_/S VGND VGND VPWR VPWR _4268_/X sky130_fd_sc_hd__mux2_1
X_6007_ _6899_/Q _5950_/X _5952_/Y _7003_/Q _6006_/X VGND VGND VPWR VPWR _6007_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_74_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3219_ _6797_/Q VGND VGND VPWR VPWR _3219_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_86_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4199_ hold833/X _6355_/A1 _4201_/S VGND VGND VPWR VPWR _4199_/X sky130_fd_sc_hd__mux2_1
XFILLER_54_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6909_ _7060_/CLK _6909_/D fanout521/X VGND VGND VPWR VPWR _6909_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_23_584 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_168_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_124_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold290 _5193_/X VGND VGND VPWR VPWR _6772_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_2_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_172_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_26 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_130 _3917_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_141 _5915_/B1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_152 _5530_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_163 hold23/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_174 _3959_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_185 _5969_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_196 _3952_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_147_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_174_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3570_ _6548_/Q _4127_/A _4303_/A _6703_/Q VGND VGND VPWR VPWR _3570_/X sky130_fd_sc_hd__a22o_1
XFILLER_155_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_142_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_114_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5240_ _5240_/A0 _5465_/A1 _5243_/S VGND VGND VPWR VPWR _5240_/X sky130_fd_sc_hd__mux2_1
XFILLER_46_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5171_ _3797_/A _5168_/A _5488_/A1 _5171_/B1 _6352_/B VGND VGND VPWR VPWR _5171_/X
+ sky130_fd_sc_hd__o311a_1
XFILLER_96_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4122_ _4122_/A0 _6353_/A1 _4126_/S VGND VGND VPWR VPWR _4122_/X sky130_fd_sc_hd__mux2_1
XFILLER_110_331 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_598 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4053_ hold604/X _4052_/X _4061_/S VGND VGND VPWR VPWR _4053_/X sky130_fd_sc_hd__mux2_1
Xinput3 debug_out VGND VGND VPWR VPWR input3/X sky130_fd_sc_hd__clkbuf_1
XFILLER_83_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4955_ _4950_/X _4955_/B _4955_/C _4955_/D VGND VGND VPWR VPWR _4955_/X sky130_fd_sc_hd__and4b_1
X_3906_ _3856_/S _3867_/A _3859_/Y _3164_/Y VGND VGND VPWR VPWR _6488_/D sky130_fd_sc_hd__a22o_1
X_4886_ _4886_/A _4895_/A VGND VGND VPWR VPWR _4886_/Y sky130_fd_sc_hd__nand2_1
X_6625_ _7153_/CLK _6625_/D fanout486/X VGND VGND VPWR VPWR _6625_/Q sky130_fd_sc_hd__dfrtp_1
X_3837_ _3856_/S _3837_/B _3837_/C VGND VGND VPWR VPWR _3837_/X sky130_fd_sc_hd__and3b_1
XFILLER_165_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6556_ _6630_/CLK _6556_/D fanout495/X VGND VGND VPWR VPWR _6556_/Q sky130_fd_sc_hd__dfrtp_4
X_3768_ _3768_/A _3768_/B VGND VGND VPWR VPWR _3778_/C sky130_fd_sc_hd__or2_1
XFILLER_180_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5507_ hold585/X _6357_/A1 _5510_/S VGND VGND VPWR VPWR _5507_/X sky130_fd_sc_hd__mux2_1
XFILLER_118_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6487_ _3939_/A1 _6487_/D _6376_/X VGND VGND VPWR VPWR _6487_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_118_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3699_ _7056_/Q _5511_/A _4202_/A _6610_/Q _3698_/X VGND VGND VPWR VPWR _3712_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_105_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_160_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_161_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5438_ _5438_/A0 _5465_/A1 hold35/X VGND VGND VPWR VPWR _5438_/X sky130_fd_sc_hd__mux2_1
Xoutput340 hold1365/X VGND VGND VPWR VPWR hold1366/A sky130_fd_sc_hd__buf_12
XFILLER_105_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_160_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5369_ hold187/X hold27/X _5369_/S VGND VGND VPWR VPWR _5369_/X sky130_fd_sc_hd__mux2_1
XFILLER_114_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7108_ _7123_/CLK _7108_/D fanout497/X VGND VGND VPWR VPWR _7108_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_113_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7039_ _7039_/CLK _7039_/D fanout498/X VGND VGND VPWR VPWR _7039_/Q sky130_fd_sc_hd__dfstp_1
XTAP_1002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_329 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_129_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_167_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_183_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_152_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_128 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4740_ _4587_/A _4549_/B _4684_/Y VGND VGND VPWR VPWR _4740_/X sky130_fd_sc_hd__o21ba_1
XTAP_1591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4671_ _4977_/B _4671_/B _4725_/B VGND VGND VPWR VPWR _4724_/C sky130_fd_sc_hd__nor3_1
XFILLER_186_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6410_ _3500_/A1 _6410_/D _6366_/X VGND VGND VPWR VPWR hold48/A sky130_fd_sc_hd__dfrtp_1
X_3622_ _7029_/Q _5478_/A _4321_/A _6718_/Q _3621_/X VGND VGND VPWR VPWR _3623_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_134_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6341_ _6644_/Q _6341_/A2 _6341_/B1 _6643_/Q VGND VGND VPWR VPWR _6341_/X sky130_fd_sc_hd__a22o_1
X_3553_ _3553_/A _3554_/B VGND VGND VPWR VPWR _4309_/A sky130_fd_sc_hd__nor2_8
XFILLER_155_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6272_ _6483_/Q _5953_/Y _5973_/C hold65/A _6271_/X VGND VGND VPWR VPWR _6277_/B
+ sky130_fd_sc_hd__a221o_1
X_3484_ _6918_/Q _5352_/A hold83/A _6886_/Q _3483_/X VGND VGND VPWR VPWR _3489_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_142_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5223_ hold675/X _5544_/A1 _5225_/S VGND VGND VPWR VPWR _5223_/X sky130_fd_sc_hd__mux2_1
X_5154_ hold803/X _6355_/A1 _5157_/S VGND VGND VPWR VPWR _5154_/X sky130_fd_sc_hd__mux2_1
XFILLER_57_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4105_ hold126/X hold90/X _4111_/S VGND VGND VPWR VPWR _4105_/X sky130_fd_sc_hd__mux2_1
XFILLER_110_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5085_ _5085_/A _5085_/B _5082_/X _5083_/X VGND VGND VPWR VPWR _5085_/X sky130_fd_sc_hd__or4bb_1
XFILLER_84_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4036_ hold602/X _4289_/A1 _4037_/S VGND VGND VPWR VPWR _4036_/X sky130_fd_sc_hd__mux2_1
XFILLER_37_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5987_ _6802_/Q _5973_/B _5959_/Y _6866_/Q VGND VGND VPWR VPWR _5987_/X sky130_fd_sc_hd__a22o_1
XFILLER_24_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_498 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4938_ _4962_/C _4615_/X _4812_/B _4828_/X VGND VGND VPWR VPWR _4939_/C sky130_fd_sc_hd__o211a_1
XANTENNA_30 _3461_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_178_684 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_41 _4020_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4869_ _4692_/C _4861_/B _4686_/X VGND VGND VPWR VPWR _4869_/X sky130_fd_sc_hd__o21a_1
XFILLER_20_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_52 _5459_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_63 _6789_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6608_ _6707_/CLK _6608_/D fanout486/X VGND VGND VPWR VPWR _6608_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA_74 _7157_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_85 user_clock VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_96 _3943_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_193_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6539_ _6969_/CLK _6539_/D fanout506/X VGND VGND VPWR VPWR _6539_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_4_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_192_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_134_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_161_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_307 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput181 _3206_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[15] sky130_fd_sc_hd__buf_12
Xoutput192 _3195_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[25] sky130_fd_sc_hd__buf_12
XFILLER_153_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_153_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_169_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_169_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_178_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_183 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_116_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_184_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_171_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_140_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5910_ _7116_/Q _5612_/A _5612_/B VGND VGND VPWR VPWR _5910_/X sky130_fd_sc_hd__o21a_1
XFILLER_19_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6890_ _7039_/CLK _6890_/D fanout498/X VGND VGND VPWR VPWR _6890_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_34_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_179_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5841_ _6565_/Q _5920_/A2 _5646_/X _6480_/Q _5840_/X VGND VGND VPWR VPWR _5841_/Y
+ sky130_fd_sc_hd__a221oi_1
XFILLER_34_454 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5772_ _6815_/Q _5913_/A2 _5927_/A2 _6823_/Q VGND VGND VPWR VPWR _5772_/X sky130_fd_sc_hd__a22o_1
XFILLER_21_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4723_ _4722_/X _4723_/B _4723_/C _5081_/A VGND VGND VPWR VPWR _4723_/X sky130_fd_sc_hd__and4b_1
XFILLER_30_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4654_ _4594_/X _4861_/B _4671_/B VGND VGND VPWR VPWR _4656_/C sky130_fd_sc_hd__a21o_1
X_3605_ _3605_/A _3605_/B _3605_/C _3605_/D VGND VGND VPWR VPWR _3624_/A sky130_fd_sc_hd__nor4_1
Xinput50 mgmt_gpio_in[22] VGND VGND VPWR VPWR input50/X sky130_fd_sc_hd__clkbuf_2
XFILLER_190_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput61 mgmt_gpio_in[32] VGND VGND VPWR VPWR input61/X sky130_fd_sc_hd__clkbuf_4
Xhold801 _6707_/Q VGND VGND VPWR VPWR hold801/X sky130_fd_sc_hd__dlygate4sd3_1
Xinput72 mgmt_gpio_in[9] VGND VGND VPWR VPWR input72/X sky130_fd_sc_hd__dlymetal6s2s_1
X_4585_ _4586_/B _5026_/A VGND VGND VPWR VPWR _4585_/X sky130_fd_sc_hd__or2_1
XFILLER_128_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold812 _4011_/X VGND VGND VPWR VPWR _6457_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_174_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold823 _6547_/Q VGND VGND VPWR VPWR hold823/X sky130_fd_sc_hd__dlygate4sd3_1
Xinput83 spimemio_flash_clk VGND VGND VPWR VPWR input83/X sky130_fd_sc_hd__buf_2
Xinput94 uart_enabled VGND VGND VPWR VPWR _3950_/B sky130_fd_sc_hd__clkbuf_1
Xhold834 _4199_/X VGND VGND VPWR VPWR _6606_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6324_ _6644_/Q _6324_/A2 _6324_/B1 _4222_/B _6323_/X VGND VGND VPWR VPWR _6324_/X
+ sky130_fd_sc_hd__a221o_1
X_3536_ hold33/X _5183_/B VGND VGND VPWR VPWR _5487_/A sky130_fd_sc_hd__nor2_4
Xhold845 _6472_/Q VGND VGND VPWR VPWR hold845/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold856 _5351_/X VGND VGND VPWR VPWR _6913_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold867 _6551_/Q VGND VGND VPWR VPWR hold867/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold878 _4275_/X VGND VGND VPWR VPWR _6676_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_88_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6255_ _6255_/A1 _6305_/A2 _6253_/X _6254_/X VGND VGND VPWR VPWR _7129_/D sky130_fd_sc_hd__o22a_1
Xhold889 _6963_/Q VGND VGND VPWR VPWR hold889/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_88_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3467_ _6871_/Q _5298_/A _5511_/A _7060_/Q _3466_/X VGND VGND VPWR VPWR _3470_/C
+ sky130_fd_sc_hd__a221o_1
X_5206_ hold136/X _5476_/A1 _5207_/S VGND VGND VPWR VPWR _5206_/X sky130_fd_sc_hd__mux2_1
X_6186_ _6715_/Q _5955_/X _5975_/C _6700_/Q VGND VGND VPWR VPWR _6186_/X sky130_fd_sc_hd__a22o_1
X_3398_ _3435_/A1 _3396_/X _3685_/S VGND VGND VPWR VPWR _3398_/X sky130_fd_sc_hd__mux2_1
Xhold1501 _7114_/Q VGND VGND VPWR VPWR _5845_/A1 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1512 _7128_/Q VGND VGND VPWR VPWR _6230_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_69_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5137_ _4745_/B _5043_/X _5054_/B _4868_/D _4974_/X VGND VGND VPWR VPWR _5138_/C
+ sky130_fd_sc_hd__o2111a_1
Xhold1523 _7091_/Q VGND VGND VPWR VPWR _5563_/A1 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1534 _6783_/Q VGND VGND VPWR VPWR hold395/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_57_546 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1545 _6785_/Q VGND VGND VPWR VPWR hold1545/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1556 _6523_/Q VGND VGND VPWR VPWR hold407/A sky130_fd_sc_hd__dlygate4sd3_1
X_5068_ _5068_/A _5068_/B VGND VGND VPWR VPWR _5112_/C sky130_fd_sc_hd__nor2_1
XFILLER_84_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_376 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4019_ hold994/X _4236_/A1 _4019_/S VGND VGND VPWR VPWR _4019_/X sky130_fd_sc_hd__mux2_1
XFILLER_37_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_432 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_334 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_507 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_304 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_193_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_180_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_402 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_171_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold108 _3533_/A VGND VGND VPWR VPWR _3390_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_156_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold119 _5405_/X VGND VGND VPWR VPWR _6961_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_172_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4370_ _4499_/B _4449_/C VGND VGND VPWR VPWR _4631_/A sky130_fd_sc_hd__or2_2
XFILLER_125_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3321_ _3563_/A _3571_/B VGND VGND VPWR VPWR _5493_/A sky130_fd_sc_hd__nor2_8
XFILLER_125_584 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6040_ _6796_/Q _6299_/A2 _5977_/X _6924_/Q VGND VGND VPWR VPWR _6040_/X sky130_fd_sc_hd__a22o_1
XTAP_446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3252_ _3252_/A0 _3252_/A1 _3256_/S VGND VGND VPWR VPWR _7164_/D sky130_fd_sc_hd__mux2_1
XTAP_457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3183_ _7082_/Q VGND VGND VPWR VPWR _3183_/Y sky130_fd_sc_hd__inv_2
XFILLER_27_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6942_ _6988_/CLK _6942_/D fanout513/X VGND VGND VPWR VPWR _6942_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_19_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6873_ _7072_/CLK _6873_/D fanout505/X VGND VGND VPWR VPWR _6873_/Q sky130_fd_sc_hd__dfrtp_1
X_5824_ _6555_/Q _5627_/X _5926_/B1 _6545_/Q VGND VGND VPWR VPWR _5824_/X sky130_fd_sc_hd__a22o_1
X_5755_ _6790_/Q _5667_/X _5744_/X _5754_/X _5610_/A VGND VGND VPWR VPWR _5755_/X
+ sky130_fd_sc_hd__o221a_4
X_4706_ _4706_/A _4706_/B _4706_/C _4705_/X VGND VGND VPWR VPWR _4709_/B sky130_fd_sc_hd__or4b_1
X_5686_ _7011_/Q _5620_/X _5630_/X _6955_/Q _5685_/X VGND VGND VPWR VPWR _5686_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_148_676 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_148_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4637_ _4637_/A VGND VGND VPWR VPWR _4638_/B sky130_fd_sc_hd__inv_2
XFILLER_162_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_190_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold620 _7016_/Q VGND VGND VPWR VPWR hold620/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold631 _4072_/X VGND VGND VPWR VPWR _6502_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4568_ _4542_/A _4575_/A _4862_/A _5088_/B _4566_/Y VGND VGND VPWR VPWR _4568_/X
+ sky130_fd_sc_hd__o311a_1
XFILLER_190_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmax_cap350 hold61/X VGND VGND VPWR VPWR _3525_/A sky130_fd_sc_hd__buf_12
Xhold642 _6800_/Q VGND VGND VPWR VPWR hold642/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_150_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmax_cap361 _3297_/Y VGND VGND VPWR VPWR _5361_/A sky130_fd_sc_hd__buf_8
XFILLER_104_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold653 _5539_/X VGND VGND VPWR VPWR _7079_/D sky130_fd_sc_hd__dlygate4sd3_1
Xmax_cap372 hold33/X VGND VGND VPWR VPWR _3554_/A sky130_fd_sc_hd__buf_12
XFILLER_162_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold664 hold664/A VGND VGND VPWR VPWR _6763_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3519_ _3525_/A _3628_/B VGND VGND VPWR VPWR _4208_/A sky130_fd_sc_hd__nor2_8
X_6307_ _6307_/A1 _3908_/Y _6306_/Y _3903_/B _6636_/Q VGND VGND VPWR VPWR _7132_/D
+ sky130_fd_sc_hd__a32o_1
Xmax_cap383 _5943_/Y VGND VGND VPWR VPWR _6176_/A2 sky130_fd_sc_hd__buf_6
Xhold675 _6799_/Q VGND VGND VPWR VPWR hold675/X sky130_fd_sc_hd__dlygate4sd3_1
Xmax_cap394 _5948_/X VGND VGND VPWR VPWR _6299_/A2 sky130_fd_sc_hd__buf_12
XFILLER_89_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold686 _5241_/X VGND VGND VPWR VPWR _6815_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4499_ _4544_/A _4499_/B _4368_/A VGND VGND VPWR VPWR _4691_/C sky130_fd_sc_hd__or3b_4
XFILLER_104_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold697 _7179_/A VGND VGND VPWR VPWR hold697/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_131_543 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6238_ _6477_/Q _5976_/Y _5979_/X _6452_/Q _6235_/X VGND VGND VPWR VPWR _6252_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_89_479 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_103_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6169_ _6961_/Q _5957_/X _5974_/B _6833_/Q VGND VGND VPWR VPWR _6169_/X sky130_fd_sc_hd__a22o_1
XTAP_991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1320 hold1320/A VGND VGND VPWR VPWR wb_dat_o[7] sky130_fd_sc_hd__buf_12
XFILLER_134_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1331 _4173_/A1 VGND VGND VPWR VPWR hold1331/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_85_652 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1342 hold1342/A VGND VGND VPWR VPWR wb_dat_o[3] sky130_fd_sc_hd__buf_12
XFILLER_45_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1353 _4180_/A1 VGND VGND VPWR VPWR hold1353/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1364 hold1364/A VGND VGND VPWR VPWR wb_dat_o[24] sky130_fd_sc_hd__buf_12
XFILLER_85_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1375 _7197_/A VGND VGND VPWR VPWR _4099_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1386 _6881_/Q VGND VGND VPWR VPWR _5315_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_45_538 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1397 _6576_/Q VGND VGND VPWR VPWR hold1397/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_43_csclk clkbuf_3_6_0_csclk/X VGND VGND VPWR VPWR _7086_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_2836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_159_21 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_58_csclk clkbuf_3_2_0_csclk/X VGND VGND VPWR VPWR _6928_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_43_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_126_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_175_31 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_181_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_318 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_565 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_727 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_191_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_655 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3870_ hold5/A _6402_/Q _6396_/B VGND VGND VPWR VPWR _3956_/B sky130_fd_sc_hd__o21ai_1
XFILLER_177_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5540_ hold255/X hold90/X _5546_/S VGND VGND VPWR VPWR _5540_/X sky130_fd_sc_hd__mux2_1
XFILLER_192_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_145_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5471_ hold122/X hold90/X hold19/X VGND VGND VPWR VPWR _5471_/X sky130_fd_sc_hd__mux2_1
XFILLER_172_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4422_ _4894_/B _4885_/A _4737_/B _4573_/A VGND VGND VPWR VPWR _4503_/D sky130_fd_sc_hd__or4b_2
XFILLER_160_627 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7141_ _3931_/A1 _7141_/D _6308_/B VGND VGND VPWR VPWR _7141_/Q sky130_fd_sc_hd__dfrtp_1
X_4353_ _4345_/C _4351_/Y _4888_/B VGND VGND VPWR VPWR _4894_/A sky130_fd_sc_hd__o21ai_4
X_3304_ _3440_/A hold74/X VGND VGND VPWR VPWR _3706_/A sky130_fd_sc_hd__or2_4
X_7072_ _7072_/CLK _7072_/D fanout505/X VGND VGND VPWR VPWR _7072_/Q sky130_fd_sc_hd__dfstp_1
Xfanout429 _5519_/A1 VGND VGND VPWR VPWR _5537_/A1 sky130_fd_sc_hd__buf_6
X_4284_ hold849/X _6357_/A1 _4284_/S VGND VGND VPWR VPWR _4284_/X sky130_fd_sc_hd__mux2_1
XFILLER_101_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6023_ _6811_/Q _6259_/A2 _5972_/A _6907_/Q VGND VGND VPWR VPWR _6023_/X sky130_fd_sc_hd__a22o_1
X_3235_ _3245_/B VGND VGND VPWR VPWR _3235_/Y sky130_fd_sc_hd__inv_2
XFILLER_67_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3166_ hold78/A VGND VGND VPWR VPWR _3166_/Y sky130_fd_sc_hd__inv_2
XFILLER_67_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_611 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6925_ _7069_/CLK _6925_/D fanout516/X VGND VGND VPWR VPWR _6925_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_82_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6856_ _7058_/CLK _6856_/D fanout521/X VGND VGND VPWR VPWR _6856_/Q sky130_fd_sc_hd__dfrtp_4
X_5807_ _6985_/Q _5642_/X _5807_/B1 _6937_/Q _5802_/Y VGND VGND VPWR VPWR _5807_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_50_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6787_ _7011_/CLK _6787_/D fanout500/X VGND VGND VPWR VPWR _6787_/Q sky130_fd_sc_hd__dfstp_1
X_3999_ hold695/X _5544_/A1 _4001_/S VGND VGND VPWR VPWR _3999_/X sky130_fd_sc_hd__mux2_1
XFILLER_13_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_183_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5738_ _6982_/Q _5642_/X _5807_/B1 _6934_/Q VGND VGND VPWR VPWR _5738_/X sky130_fd_sc_hd__a22o_1
XFILLER_136_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_175_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5669_ _5690_/A1 _5611_/X _5668_/X VGND VGND VPWR VPWR _7106_/D sky130_fd_sc_hd__a21o_1
XFILLER_136_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold450 _4025_/X VGND VGND VPWR VPWR _6469_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold461 _6848_/Q VGND VGND VPWR VPWR hold461/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold472 _4126_/X VGND VGND VPWR VPWR _6544_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold483 _6832_/Q VGND VGND VPWR VPWR hold483/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_145_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold494 _4051_/X VGND VGND VPWR VPWR _6492_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_1_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_161_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1150 _5294_/X VGND VGND VPWR VPWR _6862_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1161 _6998_/Q VGND VGND VPWR VPWR _5447_/A0 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1172 _4238_/X VGND VGND VPWR VPWR _6645_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_45_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1183 _6890_/Q VGND VGND VPWR VPWR _5326_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1194 _4197_/X VGND VGND VPWR VPWR _6604_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_154_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_186_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_186_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_318 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_2_1_0_wb_clk_i clkbuf_2_1_0_wb_clk_i/A VGND VGND VPWR VPWR clkbuf_3_3_0_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_96_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_630 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_568 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_611 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4971_ _5048_/A _5068_/A _4971_/C VGND VGND VPWR VPWR _4976_/B sky130_fd_sc_hd__nor3_1
XFILLER_51_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6710_ _6711_/CLK _6710_/D _3940_/B VGND VGND VPWR VPWR _6710_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_32_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3922_ _6510_/Q _3263_/C _6406_/Q VGND VGND VPWR VPWR _3922_/X sky130_fd_sc_hd__mux2_1
X_3853_ _3166_/Y _3857_/S _3842_/B hold71/A VGND VGND VPWR VPWR _3853_/X sky130_fd_sc_hd__o211a_1
X_6641_ _7150_/CLK _6641_/D _6308_/B VGND VGND VPWR VPWR _6641_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_165_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3784_ _6986_/Q hold34/A _4202_/A _6609_/Q _3783_/X VGND VGND VPWR VPWR _3792_/A
+ sky130_fd_sc_hd__a221o_1
X_6572_ _7140_/CLK _6572_/D VGND VGND VPWR VPWR _6572_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_192_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5523_ hold333/X _5523_/A1 _5528_/S VGND VGND VPWR VPWR _5523_/X sky130_fd_sc_hd__mux2_1
XFILLER_157_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_173_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_145_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5454_ hold839/X _5505_/A1 _5459_/S VGND VGND VPWR VPWR _5454_/X sky130_fd_sc_hd__mux2_1
XFILLER_117_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4405_ _4613_/C _4542_/C _4435_/B VGND VGND VPWR VPWR _4416_/B sky130_fd_sc_hd__o21a_1
XFILLER_132_126 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5385_ hold665/X _5544_/A1 _5387_/S VGND VGND VPWR VPWR _5385_/X sky130_fd_sc_hd__mux2_1
XFILLER_160_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7124_ _7124_/CLK _7124_/D fanout502/X VGND VGND VPWR VPWR _7124_/Q sky130_fd_sc_hd__dfrtp_1
X_4336_ _4336_/A _4336_/B _4336_/C _4336_/D VGND VGND VPWR VPWR _4337_/C sky130_fd_sc_hd__and4_1
XFILLER_141_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7055_ _7055_/CLK _7055_/D fanout504/X VGND VGND VPWR VPWR _7055_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_86_224 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4267_ _4267_/A hold7/X VGND VGND VPWR VPWR _4272_/S sky130_fd_sc_hd__and2_2
X_6006_ _6915_/Q _6288_/A2 _5977_/X _6923_/Q VGND VGND VPWR VPWR _6006_/X sky130_fd_sc_hd__a22o_1
X_3218_ _6805_/Q VGND VGND VPWR VPWR _3218_/Y sky130_fd_sc_hd__inv_2
XFILLER_27_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4198_ hold986/X _6354_/A1 _4201_/S VGND VGND VPWR VPWR _4198_/X sky130_fd_sc_hd__mux2_1
XFILLER_54_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6908_ _7043_/CLK _6908_/D fanout520/X VGND VGND VPWR VPWR _6908_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_70_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6839_ _6961_/CLK _6839_/D fanout522/X VGND VGND VPWR VPWR _6839_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_23_596 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_183_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_136_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold280 _3996_/X VGND VGND VPWR VPWR _6444_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold291 _7177_/A VGND VGND VPWR VPWR hold291/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_120 input21/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_131 _6741_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_142 _5921_/A2 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_153 _5521_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_164 hold23/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_175 _4120_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_186 _5977_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_197 _6441_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_174_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5170_ _5170_/A _5170_/B VGND VGND VPWR VPWR _5170_/X sky130_fd_sc_hd__or2_1
XFILLER_96_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4121_ _4121_/A _6352_/B VGND VGND VPWR VPWR _4126_/S sky130_fd_sc_hd__and2_2
XFILLER_96_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4052_ hold769/X _5515_/A1 _4103_/B VGND VGND VPWR VPWR _4052_/X sky130_fd_sc_hd__mux2_1
XFILLER_49_471 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput4 mask_rev_in[0] VGND VGND VPWR VPWR input4/X sky130_fd_sc_hd__clkbuf_1
XFILLER_83_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_176 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4954_ _4513_/A _4515_/B _5026_/B VGND VGND VPWR VPWR _4955_/D sky130_fd_sc_hd__a21o_1
XFILLER_177_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_179 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3905_ _7159_/Q _6485_/Q _3858_/B _3905_/B1 VGND VGND VPWR VPWR _6489_/D sky130_fd_sc_hd__a31o_1
X_4885_ _4885_/A _4885_/B VGND VGND VPWR VPWR _4895_/A sky130_fd_sc_hd__nor2_2
XFILLER_20_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_165_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6624_ _7150_/CLK _6624_/D _6308_/B VGND VGND VPWR VPWR _6624_/Q sky130_fd_sc_hd__dfrtp_4
X_3836_ hold56/A hold29/A _3845_/S hold14/A VGND VGND VPWR VPWR _3837_/C sky130_fd_sc_hd__a31o_1
XFILLER_137_207 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3767_ _6685_/Q _4285_/A _3629_/Y _6767_/Q _3766_/X VGND VGND VPWR VPWR _3768_/B
+ sky130_fd_sc_hd__a221o_1
X_6555_ _6630_/CLK _6555_/D fanout495/X VGND VGND VPWR VPWR _6555_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_118_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_443 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5506_ hold537/X _5515_/A1 _5510_/S VGND VGND VPWR VPWR _5506_/X sky130_fd_sc_hd__mux2_1
X_6486_ _7171_/CLK _6486_/D _6375_/X VGND VGND VPWR VPWR _6486_/Q sky130_fd_sc_hd__dfrtp_1
X_3698_ _7080_/Q _5538_/A _5502_/A _7048_/Q VGND VGND VPWR VPWR _3698_/X sky130_fd_sc_hd__a22o_1
Xoutput330 hold1363/X VGND VGND VPWR VPWR hold1364/A sky130_fd_sc_hd__buf_12
X_5437_ hold707/X _5542_/A1 hold35/X VGND VGND VPWR VPWR _5437_/X sky130_fd_sc_hd__mux2_1
Xoutput341 hold1333/X VGND VGND VPWR VPWR hold1334/A sky130_fd_sc_hd__buf_12
XFILLER_161_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5368_ hold273/X hold114/X _5369_/S VGND VGND VPWR VPWR _5368_/X sky130_fd_sc_hd__mux2_1
XFILLER_99_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7107_ _7131_/CLK _7107_/D fanout497/X VGND VGND VPWR VPWR _7107_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_99_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4319_ hold547/X _5491_/A1 _4320_/S VGND VGND VPWR VPWR _4319_/X sky130_fd_sc_hd__mux2_1
X_5299_ hold851/X _5521_/A1 _5306_/S VGND VGND VPWR VPWR _5299_/X sky130_fd_sc_hd__mux2_1
XFILLER_101_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7038_ _7038_/CLK _7038_/D fanout489/X VGND VGND VPWR VPWR _7038_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_75_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_295 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4670_ _4977_/B _4692_/C _4725_/B _4223_/B VGND VGND VPWR VPWR _4960_/B sky130_fd_sc_hd__o31a_1
XFILLER_187_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3621_ _7074_/Q _5529_/A _4196_/A _6607_/Q _3620_/X VGND VGND VPWR VPWR _3621_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_128_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_186_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3552_ _3552_/A hold53/A VGND VGND VPWR VPWR _4285_/A sky130_fd_sc_hd__nor2_8
X_6340_ _6339_/X _6340_/A1 _6346_/S VGND VGND VPWR VPWR _7146_/D sky130_fd_sc_hd__mux2_1
XFILLER_143_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6271_ _6653_/Q _5972_/A _6285_/A2 _6633_/Q VGND VGND VPWR VPWR _6271_/X sky130_fd_sc_hd__a22o_1
XFILLER_170_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3483_ hold86/A _5406_/A hold76/A _3954_/B VGND VGND VPWR VPWR _3483_/X sky130_fd_sc_hd__a22o_1
XFILLER_142_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_143_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5222_ _5222_/A0 _5465_/A1 _5225_/S VGND VGND VPWR VPWR _5222_/X sky130_fd_sc_hd__mux2_1
X_5153_ _5153_/A0 _6354_/A1 _5157_/S VGND VGND VPWR VPWR _5153_/X sky130_fd_sc_hd__mux2_1
XFILLER_84_503 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4104_ hold893/X _5521_/A1 _4111_/S VGND VGND VPWR VPWR _4104_/X sky130_fd_sc_hd__mux2_1
XFILLER_29_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5084_ _5085_/A _5085_/B _5083_/X VGND VGND VPWR VPWR _5084_/X sky130_fd_sc_hd__or3b_1
X_4035_ hold843/X _6355_/A1 _4037_/S VGND VGND VPWR VPWR _4035_/X sky130_fd_sc_hd__mux2_1
XFILLER_84_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_444 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5986_ _6954_/Q _5957_/X _5971_/B _6858_/Q _5985_/X VGND VGND VPWR VPWR _6002_/A
+ sky130_fd_sc_hd__a221o_1
XPHY_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_169_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_178_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4937_ _4988_/A _4791_/B _5070_/A _4934_/X _4936_/X VGND VGND VPWR VPWR _4939_/B
+ sky130_fd_sc_hd__o2111a_1
XFILLER_33_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_20 _5388_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_31 _3461_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4868_ _4868_/A _4960_/C _4868_/C _4868_/D VGND VGND VPWR VPWR _4878_/A sky130_fd_sc_hd__and4_1
XFILLER_178_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_42 _3648_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_53 _5528_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6607_ _6707_/CLK _6607_/D fanout485/X VGND VGND VPWR VPWR _6607_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA_64 _6789_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_75 _7126_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3819_ _6487_/Q _3819_/B VGND VGND VPWR VPWR _3825_/B sky130_fd_sc_hd__nor2_2
XFILLER_165_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_86 input93/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4799_ _4799_/A _4799_/B VGND VGND VPWR VPWR _4984_/B sky130_fd_sc_hd__or2_1
XANTENNA_97 _3943_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6538_ _6711_/CLK _6538_/D fanout486/X VGND VGND VPWR VPWR _6538_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_21_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6469_ _6697_/CLK _6469_/D fanout489/X VGND VGND VPWR VPWR _6469_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_79_319 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput171 _3952_/X VGND VGND VPWR VPWR debug_in sky130_fd_sc_hd__buf_12
Xoutput182 _3204_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[16] sky130_fd_sc_hd__buf_12
XFILLER_121_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput193 _3194_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[26] sky130_fd_sc_hd__buf_12
XFILLER_0_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_238 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_591 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_188_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_178_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_138 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_396 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_463 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5840_ _6560_/Q _5636_/X _5642_/X _6460_/Q VGND VGND VPWR VPWR _5840_/X sky130_fd_sc_hd__a22o_1
XFILLER_34_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5771_ _6967_/Q _5925_/B1 _5650_/X _6895_/Q VGND VGND VPWR VPWR _5771_/X sky130_fd_sc_hd__a22o_1
X_4722_ _4707_/B _4721_/Y _4720_/X _4689_/Y VGND VGND VPWR VPWR _4722_/X sky130_fd_sc_hd__a211o_1
XFILLER_147_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4653_ _5043_/B _4575_/X _4676_/B VGND VGND VPWR VPWR _4664_/B sky130_fd_sc_hd__a21o_1
Xinput40 mgmt_gpio_in[13] VGND VGND VPWR VPWR input40/X sky130_fd_sc_hd__clkbuf_1
X_3604_ _6740_/Q _5145_/A _4008_/A _6458_/Q _3603_/X VGND VGND VPWR VPWR _3605_/D
+ sky130_fd_sc_hd__a221o_1
Xinput51 mgmt_gpio_in[23] VGND VGND VPWR VPWR input51/X sky130_fd_sc_hd__buf_2
Xhold802 _4312_/X VGND VGND VPWR VPWR _6707_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4584_ _4943_/A _4789_/B VGND VGND VPWR VPWR _4724_/B sky130_fd_sc_hd__nor2_1
Xinput62 mgmt_gpio_in[33] VGND VGND VPWR VPWR input62/X sky130_fd_sc_hd__buf_2
Xinput73 pad_flash_io0_di VGND VGND VPWR VPWR _3946_/B sky130_fd_sc_hd__clkbuf_1
Xhold813 _6567_/Q VGND VGND VPWR VPWR hold813/X sky130_fd_sc_hd__dlygate4sd3_1
Xinput84 spimemio_flash_csb VGND VGND VPWR VPWR input84/X sky130_fd_sc_hd__buf_2
Xhold824 _4130_/X VGND VGND VPWR VPWR _6547_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6323_ _6642_/Q _6323_/A2 _6323_/B1 _6643_/Q VGND VGND VPWR VPWR _6323_/X sky130_fd_sc_hd__a22o_1
Xinput95 usr1_vcc_pwrgood VGND VGND VPWR VPWR input95/X sky130_fd_sc_hd__buf_2
Xhold835 _6580_/Q VGND VGND VPWR VPWR hold835/X sky130_fd_sc_hd__dlygate4sd3_1
X_3535_ _3535_/A _3535_/B _3535_/C _3535_/D VGND VGND VPWR VPWR _3566_/B sky130_fd_sc_hd__nor4_1
Xhold846 _4029_/X VGND VGND VPWR VPWR _6472_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold857 _6997_/Q VGND VGND VPWR VPWR hold857/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold868 _4135_/X VGND VGND VPWR VPWR _6551_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6254_ _7128_/Q _5612_/A _5612_/B VGND VGND VPWR VPWR _6254_/X sky130_fd_sc_hd__o21a_1
Xhold879 _6539_/Q VGND VGND VPWR VPWR hold879/X sky130_fd_sc_hd__dlygate4sd3_1
X_3466_ _6807_/Q _5226_/A _5262_/A _6839_/Q VGND VGND VPWR VPWR _3466_/X sky130_fd_sc_hd__a22o_1
XFILLER_115_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5205_ hold395/X _5526_/A1 _5207_/S VGND VGND VPWR VPWR _5205_/X sky130_fd_sc_hd__mux2_1
X_6185_ _6705_/Q _5957_/X _5978_/X _6695_/Q VGND VGND VPWR VPWR _6185_/X sky130_fd_sc_hd__a22o_1
X_3397_ _7170_/Q _6487_/Q VGND VGND VPWR VPWR _3749_/S sky130_fd_sc_hd__nand2_4
Xhold1502 hold48/A VGND VGND VPWR VPWR _3849_/A1 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1513 _7129_/Q VGND VGND VPWR VPWR _6255_/A1 sky130_fd_sc_hd__dlygate4sd3_1
X_5136_ _4711_/A _5136_/B _5136_/C _5136_/D VGND VGND VPWR VPWR _5136_/Y sky130_fd_sc_hd__nand4b_1
Xhold1524 _5563_/X VGND VGND VPWR VPWR _7091_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_69_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1535 _6524_/Q VGND VGND VPWR VPWR hold893/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1546 _6508_/Q VGND VGND VPWR VPWR _5566_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_57_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1557 _7110_/Q VGND VGND VPWR VPWR _5778_/A1 sky130_fd_sc_hd__dlygate4sd3_1
X_5067_ _5067_/A _5067_/B _5067_/C _4821_/C VGND VGND VPWR VPWR _5068_/B sky130_fd_sc_hd__or4b_2
XFILLER_84_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_219 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4018_ hold265/X hold46/X _4019_/S VGND VGND VPWR VPWR _4018_/X sky130_fd_sc_hd__mux2_1
XFILLER_53_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_764 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5969_ _5969_/A _5969_/B _5969_/C VGND VGND VPWR VPWR _5969_/Y sky130_fd_sc_hd__nor3_1
XFILLER_12_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_519 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_316 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_106_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_371 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_164_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_180_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_180_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_528 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_414 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_169_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_313 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_110 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_171_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold109 _3374_/Y VGND VGND VPWR VPWR _5280_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_171_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3320_ _3719_/A _3531_/A VGND VGND VPWR VPWR _5217_/A sky130_fd_sc_hd__nor2_8
XFILLER_152_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_680 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_125_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3251_ _3252_/A1 hold112/A _3256_/S VGND VGND VPWR VPWR _7165_/D sky130_fd_sc_hd__mux2_1
XTAP_436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3182_ _6915_/Q VGND VGND VPWR VPWR _3182_/Y sky130_fd_sc_hd__inv_2
XFILLER_66_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6941_ _7029_/CLK _6941_/D fanout519/X VGND VGND VPWR VPWR _6941_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_47_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6872_ _6999_/CLK _6872_/D fanout524/X VGND VGND VPWR VPWR _6872_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_50_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_263 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5823_ _5823_/A1 _6305_/A2 _5821_/X _5822_/X VGND VGND VPWR VPWR _5823_/X sky130_fd_sc_hd__o22a_1
XFILLER_50_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_179_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5754_ _5754_/A _5754_/B _5754_/C _5753_/Y VGND VGND VPWR VPWR _5754_/X sky130_fd_sc_hd__or4b_2
X_4705_ _4615_/B _4717_/B _4694_/X _5116_/A VGND VGND VPWR VPWR _4705_/X sky130_fd_sc_hd__o211a_1
X_5685_ _7003_/Q _5614_/X _5914_/A2 _6875_/Q VGND VGND VPWR VPWR _5685_/X sky130_fd_sc_hd__a22o_1
XFILLER_30_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4636_ _4921_/A _4636_/B VGND VGND VPWR VPWR _4637_/A sky130_fd_sc_hd__nor2_1
XFILLER_135_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold610 _6920_/Q VGND VGND VPWR VPWR hold610/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold621 _5467_/X VGND VGND VPWR VPWR _7016_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4567_ _4943_/A _4862_/A VGND VGND VPWR VPWR _5068_/A sky130_fd_sc_hd__nor2_4
Xhold632 _6824_/Q VGND VGND VPWR VPWR hold632/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_563 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold643 _5224_/X VGND VGND VPWR VPWR _6800_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_190_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold654 _6663_/Q VGND VGND VPWR VPWR hold654/X sky130_fd_sc_hd__dlygate4sd3_1
Xmax_cap362 _3761_/A VGND VGND VPWR VPWR _3571_/A sky130_fd_sc_hd__buf_12
X_6306_ _6641_/Q _6306_/B VGND VGND VPWR VPWR _6306_/Y sky130_fd_sc_hd__nand2_1
Xmax_cap373 _3553_/A VGND VGND VPWR VPWR _3503_/A sky130_fd_sc_hd__buf_12
X_3518_ _3518_/A _3518_/B _3518_/C _3518_/D VGND VGND VPWR VPWR _3566_/A sky130_fd_sc_hd__nor4_1
Xhold665 _6943_/Q VGND VGND VPWR VPWR hold665/X sky130_fd_sc_hd__dlygate4sd3_1
Xmax_cap384 _5941_/Y VGND VGND VPWR VPWR _6286_/B1 sky130_fd_sc_hd__buf_8
XFILLER_89_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold676 _5223_/X VGND VGND VPWR VPWR _6799_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_103_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4498_ _4894_/B _4892_/A _4885_/A _4417_/B _4737_/B VGND VGND VPWR VPWR _4503_/C
+ sky130_fd_sc_hd__a2111o_1
Xmax_cap395 _5973_/A VGND VGND VPWR VPWR _6296_/A2 sky130_fd_sc_hd__buf_8
XFILLER_143_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold687 _7015_/Q VGND VGND VPWR VPWR hold687/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold698 _4087_/X VGND VGND VPWR VPWR _6513_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6237_ _6606_/Q wire390/X _6270_/B1 _6677_/Q _6236_/X VGND VGND VPWR VPWR _6237_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_77_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_131_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3449_ input31/X _3339_/Y _5520_/A _7068_/Q _3448_/X VGND VGND VPWR VPWR _3461_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_131_577 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6168_ _6168_/A _6168_/B _6168_/C _6167_/Y VGND VGND VPWR VPWR _6168_/X sky130_fd_sc_hd__or4b_1
XTAP_981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_491 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1310 hold1310/A VGND VGND VPWR VPWR wb_dat_o[23] sky130_fd_sc_hd__buf_12
XTAP_992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1321 _4178_/A1 VGND VGND VPWR VPWR hold1321/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1332 hold1332/A VGND VGND VPWR VPWR wb_dat_o[8] sky130_fd_sc_hd__buf_12
Xhold1343 _4183_/A1 VGND VGND VPWR VPWR hold1343/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_111_290 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5119_ _5119_/A _5119_/B VGND VGND VPWR VPWR _5120_/B sky130_fd_sc_hd__nand2_1
XFILLER_84_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1354 hold1354/A VGND VGND VPWR VPWR wb_dat_o[15] sky130_fd_sc_hd__buf_12
X_6099_ _6846_/Q _5939_/X _6300_/B1 _6878_/Q VGND VGND VPWR VPWR _6099_/X sky130_fd_sc_hd__a22o_1
XFILLER_45_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1365 _4186_/A1 VGND VGND VPWR VPWR hold1365/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_84_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1376 _6537_/Q VGND VGND VPWR VPWR _4118_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_85_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1387 _6937_/Q VGND VGND VPWR VPWR _5378_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1398 _6573_/Q VGND VGND VPWR VPWR hold1398/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_3_3_0_wb_clk_i clkbuf_3_3_0_wb_clk_i/A VGND VGND VPWR VPWR _7131_/CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_53_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_159_33 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_166_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_43 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_191_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_712 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5470_ _5470_/A0 _5521_/A1 hold19/X VGND VGND VPWR VPWR _5470_/X sky130_fd_sc_hd__mux2_1
XFILLER_157_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_144_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4421_ _4587_/A _4692_/A VGND VGND VPWR VPWR _5007_/A sky130_fd_sc_hd__or2_1
XFILLER_172_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7140_ _7140_/CLK _7140_/D VGND VGND VPWR VPWR _7140_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_160_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4352_ _4888_/A _4352_/B VGND VGND VPWR VPWR _4373_/C sky130_fd_sc_hd__or2_1
XFILLER_125_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3303_ hold82/A _3554_/A VGND VGND VPWR VPWR _5460_/A sky130_fd_sc_hd__nor2_8
XFILLER_99_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7071_ _7071_/CLK _7071_/D fanout505/X VGND VGND VPWR VPWR _7071_/Q sky130_fd_sc_hd__dfstp_1
X_4283_ hold263/X hold46/X _4284_/S VGND VGND VPWR VPWR _4283_/X sky130_fd_sc_hd__mux2_1
X_6022_ _6443_/Q _6295_/A2 _5973_/C _6875_/Q _6021_/X VGND VGND VPWR VPWR _6025_/A
+ sky130_fd_sc_hd__a221o_1
X_3234_ _3817_/C _3259_/B _3234_/C _6485_/Q VGND VGND VPWR VPWR _3245_/B sky130_fd_sc_hd__and4bb_1
XFILLER_86_439 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_322 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3165_ _3165_/A VGND VGND VPWR VPWR _3165_/Y sky130_fd_sc_hd__inv_2
XFILLER_66_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_623 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6924_ _7073_/CLK _6924_/D fanout498/X VGND VGND VPWR VPWR _6924_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_81_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6855_ _6999_/CLK _6855_/D fanout523/X VGND VGND VPWR VPWR _6855_/Q sky130_fd_sc_hd__dfrtp_2
X_5806_ _6841_/Q _5928_/A2 _5804_/X _5805_/X VGND VGND VPWR VPWR _5806_/X sky130_fd_sc_hd__a211o_1
X_6786_ _7039_/CLK _6786_/D fanout497/X VGND VGND VPWR VPWR _6786_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_50_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3998_ _3998_/A0 _5465_/A1 _4001_/S VGND VGND VPWR VPWR _3998_/X sky130_fd_sc_hd__mux2_1
X_5737_ _6886_/Q _5643_/X _5912_/B1 _7030_/Q _5736_/X VGND VGND VPWR VPWR _5740_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_182_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5668_ _5661_/X _5666_/X _5667_/X _6786_/Q _5609_/Y VGND VGND VPWR VPWR _5668_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_135_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4619_ _4678_/A _4620_/B VGND VGND VPWR VPWR _4619_/Y sky130_fd_sc_hd__nor2_1
XFILLER_190_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5599_ _5940_/B _7102_/Q VGND VGND VPWR VPWR _5981_/B sky130_fd_sc_hd__nor2_4
XFILLER_123_308 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_500 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold440 _5508_/X VGND VGND VPWR VPWR _7052_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_2_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold451 _6880_/Q VGND VGND VPWR VPWR hold451/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_150_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold462 _5278_/X VGND VGND VPWR VPWR _6848_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold473 _6808_/Q VGND VGND VPWR VPWR hold473/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_145_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold484 _5260_/X VGND VGND VPWR VPWR _6832_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold495 _6703_/Q VGND VGND VPWR VPWR hold495/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_143_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_145_79 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_631 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1140 _5290_/X VGND VGND VPWR VPWR _6858_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_85_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_303 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1151 _6810_/Q VGND VGND VPWR VPWR _5236_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_58_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1162 _5447_/X VGND VGND VPWR VPWR _6998_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1173 _6460_/Q VGND VGND VPWR VPWR _4015_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1184 _5326_/X VGND VGND VPWR VPWR _6890_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_173_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1195 _6922_/Q VGND VGND VPWR VPWR _5362_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_8 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_623 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_431 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4970_ _4678_/A _5021_/A _4869_/X VGND VGND VPWR VPWR _4971_/C sky130_fd_sc_hd__o21ai_1
XFILLER_17_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3921_ _6511_/Q _3939_/A1 _6405_/Q VGND VGND VPWR VPWR _3921_/X sky130_fd_sc_hd__mux2_1
X_6640_ _7150_/CLK _6640_/D _6308_/B VGND VGND VPWR VPWR _6640_/Q sky130_fd_sc_hd__dfrtp_1
X_3852_ _3851_/X _3852_/A1 _3857_/S VGND VGND VPWR VPWR _6409_/D sky130_fd_sc_hd__mux2_1
XFILLER_20_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6571_ _7137_/CLK _6571_/D VGND VGND VPWR VPWR _6571_/Q sky130_fd_sc_hd__dfxtp_1
X_3783_ _6578_/Q _4166_/A _4121_/A _6540_/Q VGND VGND VPWR VPWR _3783_/X sky130_fd_sc_hd__a22o_1
X_5522_ hold969/X _5531_/A1 _5528_/S VGND VGND VPWR VPWR _5522_/X sky130_fd_sc_hd__mux2_1
XFILLER_118_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5453_ hold927/X _5531_/A1 _5459_/S VGND VGND VPWR VPWR _5453_/X sky130_fd_sc_hd__mux2_1
XFILLER_133_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_42_csclk clkbuf_3_6_0_csclk/X VGND VGND VPWR VPWR _7050_/CLK sky130_fd_sc_hd__clkbuf_16
X_4404_ _4472_/A _4613_/C _4419_/B VGND VGND VPWR VPWR _4513_/A sky130_fd_sc_hd__or3b_4
XFILLER_160_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5384_ _5384_/A0 _5465_/A1 _5387_/S VGND VGND VPWR VPWR _5384_/X sky130_fd_sc_hd__mux2_1
XFILLER_172_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7123_ _7123_/CLK _7123_/D fanout499/X VGND VGND VPWR VPWR _7123_/Q sky130_fd_sc_hd__dfrtp_1
X_4335_ _4335_/A _4335_/B _4335_/C _4335_/D VGND VGND VPWR VPWR _4337_/B sky130_fd_sc_hd__and4_1
X_7054_ _7054_/CLK _7054_/D fanout503/X VGND VGND VPWR VPWR _7054_/Q sky130_fd_sc_hd__dfrtp_1
X_4266_ hold475/X _5534_/A1 _4266_/S VGND VGND VPWR VPWR _4266_/X sky130_fd_sc_hd__mux2_1
XFILLER_86_236 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6005_ _5609_/Y _6003_/X _6004_/X _5611_/X _6029_/A1 VGND VGND VPWR VPWR _7119_/D
+ sky130_fd_sc_hd__a32o_1
Xclkbuf_leaf_57_csclk clkbuf_3_2_0_csclk/X VGND VGND VPWR VPWR _7076_/CLK sky130_fd_sc_hd__clkbuf_16
X_3217_ _6821_/Q VGND VGND VPWR VPWR _3217_/Y sky130_fd_sc_hd__clkinv_2
X_4197_ _4197_/A0 _6353_/A1 _4201_/S VGND VGND VPWR VPWR _4197_/X sky130_fd_sc_hd__mux2_1
XFILLER_94_280 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6907_ _7046_/CLK _6907_/D fanout500/X VGND VGND VPWR VPWR _6907_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_168_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6838_ _7022_/CLK _6838_/D fanout517/X VGND VGND VPWR VPWR _6838_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_156_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6769_ _6769_/CLK _6769_/D fanout492/X VGND VGND VPWR VPWR _6769_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_7_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_183_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_108_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_163_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold270 _3982_/X VGND VGND VPWR VPWR _6432_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_151_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold281 _6964_/Q VGND VGND VPWR VPWR hold281/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold292 _4074_/X VGND VGND VPWR VPWR _6503_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_77_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_110 _3950_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_121 _3894_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_132 _6744_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_143 _5914_/A2 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_154 _5923_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_165 hold90/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_176 _5234_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_187 _6252_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_198 _6270_/B1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_186_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_436 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_683 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4120_ hold879/X _5537_/A1 _4120_/S VGND VGND VPWR VPWR _4120_/X sky130_fd_sc_hd__mux2_1
XFILLER_96_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4051_ hold493/X _4050_/X _4061_/S VGND VGND VPWR VPWR _4051_/X sky130_fd_sc_hd__mux2_1
XFILLER_96_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput5 mask_rev_in[10] VGND VGND VPWR VPWR input5/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_49_483 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_155 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4953_ _4479_/A _4586_/B _4495_/X _5026_/B VGND VGND VPWR VPWR _4955_/C sky130_fd_sc_hd__a31o_1
XFILLER_177_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3904_ _3164_/Y _3904_/A2 _6485_/Q _3858_/B _3904_/B1 VGND VGND VPWR VPWR _6486_/D
+ sky130_fd_sc_hd__a41o_1
X_4884_ _4884_/A _4944_/A VGND VGND VPWR VPWR _4885_/B sky130_fd_sc_hd__nor2_2
XFILLER_177_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6623_ _6633_/CLK _6623_/D _6370_/A VGND VGND VPWR VPWR _6623_/Q sky130_fd_sc_hd__dfrtp_2
X_3835_ _3834_/X _3835_/A1 _3857_/S VGND VGND VPWR VPWR _6414_/D sky130_fd_sc_hd__mux2_1
XFILLER_20_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_137_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6554_ _6632_/CLK _6554_/D fanout509/X VGND VGND VPWR VPWR _6554_/Q sky130_fd_sc_hd__dfrtp_1
X_3766_ _6470_/Q _4026_/A _4303_/A _6700_/Q VGND VGND VPWR VPWR _3766_/X sky130_fd_sc_hd__a22o_1
XFILLER_20_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5505_ hold628/X _5505_/A1 _5510_/S VGND VGND VPWR VPWR _5505_/X sky130_fd_sc_hd__mux2_1
XFILLER_192_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_455 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6485_ _3939_/A1 _6485_/D _6374_/X VGND VGND VPWR VPWR _6485_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_145_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3697_ _3697_/A _3697_/B VGND VGND VPWR VPWR _3712_/A sky130_fd_sc_hd__or2_1
XFILLER_118_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5436_ hold321/X _5523_/A1 hold35/X VGND VGND VPWR VPWR _5436_/X sky130_fd_sc_hd__mux2_1
Xoutput320 hold1353/X VGND VGND VPWR VPWR hold1354/A sky130_fd_sc_hd__buf_12
Xoutput331 hold1355/X VGND VGND VPWR VPWR hold1356/A sky130_fd_sc_hd__buf_12
Xoutput342 hold1327/X VGND VGND VPWR VPWR hold1328/A sky130_fd_sc_hd__buf_12
XFILLER_160_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5367_ hold719/X _5544_/A1 _5369_/S VGND VGND VPWR VPWR _5367_/X sky130_fd_sc_hd__mux2_1
XFILLER_87_512 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7106_ _7123_/CLK _7106_/D fanout497/X VGND VGND VPWR VPWR _7106_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_59_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4318_ hold403/X _5532_/A1 _4320_/S VGND VGND VPWR VPWR _4318_/X sky130_fd_sc_hd__mux2_1
X_5298_ _5298_/A _5511_/B VGND VGND VPWR VPWR _5306_/S sky130_fd_sc_hd__and2_4
X_7037_ _7037_/CLK _7037_/D fanout485/X VGND VGND VPWR VPWR _7037_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_101_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_14 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4249_ _4249_/A hold7/X VGND VGND VPWR VPWR _4254_/S sky130_fd_sc_hd__and2_2
XFILLER_19_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_659 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_11 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_180 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_11 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_151_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_183_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_650 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_132_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_191 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3620_ _3263_/C _4112_/B _4255_/A _6663_/Q VGND VGND VPWR VPWR _3620_/X sky130_fd_sc_hd__a22o_1
XFILLER_127_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_128_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3551_ _6894_/Q _5325_/A _5442_/A _6998_/Q _3550_/X VGND VGND VPWR VPWR _3565_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_155_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6270_ _6458_/Q _6291_/A2 _6270_/B1 _6678_/Q _6269_/X VGND VGND VPWR VPWR _6277_/A
+ sky130_fd_sc_hd__a221o_1
X_3482_ _6806_/Q _5226_/A _4231_/A _6634_/Q _3480_/X VGND VGND VPWR VPWR _3489_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_115_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5221_ hold197/X _5533_/A1 _5225_/S VGND VGND VPWR VPWR _5221_/X sky130_fd_sc_hd__mux2_1
XFILLER_88_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_288 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5152_ _5152_/A0 _6353_/A1 _5157_/S VGND VGND VPWR VPWR _5152_/X sky130_fd_sc_hd__mux2_1
X_4103_ _6396_/B _4103_/B _5538_/B VGND VGND VPWR VPWR _4111_/S sky130_fd_sc_hd__and3b_4
XFILLER_110_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_515 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_375 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5083_ _4551_/B _4676_/B _4668_/X VGND VGND VPWR VPWR _5083_/X sky130_fd_sc_hd__o21a_1
XFILLER_111_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4034_ hold869/X _5189_/A1 _4037_/S VGND VGND VPWR VPWR _4034_/X sky130_fd_sc_hd__mux2_1
XFILLER_110_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5985_ _6882_/Q _5973_/A _5952_/Y _7002_/Q VGND VGND VPWR VPWR _5985_/X sky130_fd_sc_hd__a22o_1
XFILLER_169_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_456 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4936_ _4862_/B _4631_/X _4935_/X _4788_/A VGND VGND VPWR VPWR _4936_/X sky130_fd_sc_hd__o22a_1
XFILLER_33_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_177_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_10 _3339_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_21 _3384_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4867_ _4901_/B _4597_/Y _4745_/B _4748_/B VGND VGND VPWR VPWR _4868_/D sky130_fd_sc_hd__o22a_1
XANTENNA_32 _3461_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_43 _3648_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_54 _5617_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6606_ _6697_/CLK _6606_/D fanout485/X VGND VGND VPWR VPWR _6606_/Q sky130_fd_sc_hd__dfstp_2
X_3818_ _3818_/A1 _3749_/S _3816_/X _3817_/X VGND VGND VPWR VPWR _6727_/D sky130_fd_sc_hd__a22o_1
XFILLER_193_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_65 _6925_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_177_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_76 user_clock VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4798_ _4788_/A _4638_/B _4665_/C VGND VGND VPWR VPWR _4929_/A sky130_fd_sc_hd__o21ai_1
XANTENNA_87 _3943_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_165_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_98 _3943_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6537_ _7054_/CLK _6537_/D fanout503/X VGND VGND VPWR VPWR _6537_/Q sky130_fd_sc_hd__dfrtp_1
X_3749_ _3748_/X _3749_/A1 _3749_/S VGND VGND VPWR VPWR _3749_/X sky130_fd_sc_hd__mux2_1
XFILLER_119_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_180_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_192_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_146_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6468_ _6707_/CLK _6468_/D fanout484/X VGND VGND VPWR VPWR _6468_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_133_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5419_ hold715/X _5542_/A1 _5423_/S VGND VGND VPWR VPWR _5419_/X sky130_fd_sc_hd__mux2_1
XFILLER_161_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6399_ _6399_/A _6399_/B VGND VGND VPWR VPWR _6399_/X sky130_fd_sc_hd__and2_1
XFILLER_121_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput172 _7173_/X VGND VGND VPWR VPWR irq[0] sky130_fd_sc_hd__buf_12
Xoutput183 _3203_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[17] sky130_fd_sc_hd__buf_12
Xoutput194 _3193_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[27] sky130_fd_sc_hd__buf_12
XFILLER_153_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_178_98 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_171_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_171_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_294 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5770_ _6911_/Q _5628_/X _5767_/X _5769_/X VGND VGND VPWR VPWR _5770_/X sky130_fd_sc_hd__a211o_1
XFILLER_15_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4721_ _4965_/A _4721_/B VGND VGND VPWR VPWR _4721_/Y sky130_fd_sc_hd__nor2_1
X_4652_ _4639_/X _4641_/X _4985_/B _4788_/A VGND VGND VPWR VPWR _4664_/A sky130_fd_sc_hd__a31o_1
XFILLER_174_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput30 mask_rev_in[4] VGND VGND VPWR VPWR input30/X sky130_fd_sc_hd__clkbuf_2
X_3603_ _7013_/Q _5460_/A hold34/A _6989_/Q VGND VGND VPWR VPWR _3603_/X sky130_fd_sc_hd__a22o_2
Xinput41 mgmt_gpio_in[14] VGND VGND VPWR VPWR input41/X sky130_fd_sc_hd__clkbuf_1
XFILLER_162_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4583_ _4789_/B _4748_/B VGND VGND VPWR VPWR _4732_/B sky130_fd_sc_hd__nor2_1
Xinput52 mgmt_gpio_in[24] VGND VGND VPWR VPWR input52/X sky130_fd_sc_hd__buf_2
Xinput63 mgmt_gpio_in[34] VGND VGND VPWR VPWR _3951_/A sky130_fd_sc_hd__clkbuf_8
Xhold803 _6744_/Q VGND VGND VPWR VPWR hold803/X sky130_fd_sc_hd__dlygate4sd3_1
Xinput74 pad_flash_io1_di VGND VGND VPWR VPWR _3947_/B sky130_fd_sc_hd__dlymetal6s2s_1
Xhold814 _4154_/X VGND VGND VPWR VPWR _6567_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6322_ _6322_/A _6322_/B _6317_/X VGND VGND VPWR VPWR _6346_/S sky130_fd_sc_hd__or3b_4
Xhold825 _6616_/Q VGND VGND VPWR VPWR hold825/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3534_ _6846_/Q _5271_/A _4202_/A _6613_/Q _3532_/X VGND VGND VPWR VPWR _3535_/D
+ sky130_fd_sc_hd__a221o_1
Xinput85 spimemio_flash_io0_do VGND VGND VPWR VPWR input85/X sky130_fd_sc_hd__buf_2
XFILLER_155_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput96 usr1_vdd_pwrgood VGND VGND VPWR VPWR input96/X sky130_fd_sc_hd__buf_2
Xhold836 _4169_/X VGND VGND VPWR VPWR _6580_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold847 _6969_/Q VGND VGND VPWR VPWR hold847/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold858 _5446_/X VGND VGND VPWR VPWR _6997_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6253_ _6542_/Q _6004_/B _6252_/X _5610_/A VGND VGND VPWR VPWR _6253_/X sky130_fd_sc_hd__o211a_1
Xhold869 _6476_/Q VGND VGND VPWR VPWR hold869/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_170_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3465_ _6423_/Q _3958_/A _4112_/B _3950_/A _3464_/X VGND VGND VPWR VPWR _3470_/B
+ sky130_fd_sc_hd__a221o_2
XFILLER_89_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5204_ hold173/X hold23/X _5207_/S VGND VGND VPWR VPWR _5204_/X sky130_fd_sc_hd__mux2_1
X_6184_ _6560_/Q _5969_/A _5951_/X _6670_/Q _6183_/X VGND VGND VPWR VPWR _6184_/X
+ sky130_fd_sc_hd__a221o_1
X_3396_ _3396_/A _3396_/B _3395_/Y VGND VGND VPWR VPWR _3396_/X sky130_fd_sc_hd__or3b_4
Xhold1503 _7110_/Q VGND VGND VPWR VPWR _5757_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_97_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5135_ _5135_/A _5135_/B _5135_/C _5135_/D VGND VGND VPWR VPWR _5136_/D sky130_fd_sc_hd__and4_1
XFILLER_111_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1514 _6538_/Q VGND VGND VPWR VPWR hold271/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1525 hold78/A VGND VGND VPWR VPWR _3857_/A1 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1536 _6526_/Q VGND VGND VPWR VPWR hold293/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1547 _5566_/X VGND VGND VPWR VPWR _7092_/D sky130_fd_sc_hd__dlygate4sd3_1
X_5066_ _4862_/A _5026_/A _4902_/B _4934_/X VGND VGND VPWR VPWR _5067_/C sky130_fd_sc_hd__o211ai_1
Xhold1558 _7132_/Q VGND VGND VPWR VPWR _6307_/A1 sky130_fd_sc_hd__dlygate4sd3_1
X_4017_ hold861/X _5505_/A1 _4019_/S VGND VGND VPWR VPWR _4017_/X sky130_fd_sc_hd__mux2_1
XFILLER_25_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5968_ _5968_/A _5978_/B _5981_/C VGND VGND VPWR VPWR _5969_/C sky130_fd_sc_hd__and3_4
X_4919_ _4799_/B _4640_/X _4659_/X VGND VGND VPWR VPWR _4920_/B sky130_fd_sc_hd__o21ai_1
X_5899_ _6653_/Q _5922_/A2 _5636_/X _6563_/Q VGND VGND VPWR VPWR _5899_/X sky130_fd_sc_hd__a22o_1
XFILLER_166_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_148_13 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_46 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_68 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_165_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_12 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_161_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_180_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_189_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_156_122 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_464 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_172_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_140_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3250_ hold112/A _3250_/A1 _3256_/S VGND VGND VPWR VPWR _7166_/D sky130_fd_sc_hd__mux2_1
XTAP_437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3181_ _6755_/Q VGND VGND VPWR VPWR _3181_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_14_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6940_ _6965_/CLK _6940_/D fanout514/X VGND VGND VPWR VPWR _6940_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_94_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_592 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_348 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6871_ _6999_/CLK _6871_/D fanout523/X VGND VGND VPWR VPWR _6871_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_179_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5822_ _7112_/Q _3878_/Y _5612_/B VGND VGND VPWR VPWR _5822_/X sky130_fd_sc_hd__o21a_1
XFILLER_179_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5753_ _6830_/Q _5624_/X _5926_/A2 _6806_/Q _5752_/X VGND VGND VPWR VPWR _5753_/Y
+ sky130_fd_sc_hd__a221oi_1
X_4704_ _4884_/A _4619_/Y _4683_/Y _4703_/Y VGND VGND VPWR VPWR _4706_/C sky130_fd_sc_hd__a211o_1
XFILLER_147_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5684_ _6947_/Q _5626_/X _5647_/X _7027_/Q VGND VGND VPWR VPWR _5684_/X sky130_fd_sc_hd__a22o_1
XFILLER_30_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_175_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4635_ _4784_/A _4924_/B _4784_/B VGND VGND VPWR VPWR _4636_/B sky130_fd_sc_hd__or3b_1
XFILLER_190_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_147_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_190_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_175_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold600 _6483_/Q VGND VGND VPWR VPWR hold600/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold611 _5359_/X VGND VGND VPWR VPWR _6920_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4566_ _4947_/C _4566_/B VGND VGND VPWR VPWR _4566_/Y sky130_fd_sc_hd__nand2_1
Xhold622 _6553_/Q VGND VGND VPWR VPWR hold622/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold633 _5251_/X VGND VGND VPWR VPWR _6824_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6305_ _6305_/A1 _6305_/A2 _6303_/X _6304_/X VGND VGND VPWR VPWR _7131_/D sky130_fd_sc_hd__o22a_1
Xmax_cap352 _4077_/S VGND VGND VPWR VPWR _4112_/B sky130_fd_sc_hd__buf_12
Xhold644 _7085_/Q VGND VGND VPWR VPWR hold644/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_150_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmax_cap363 _3557_/A VGND VGND VPWR VPWR _3761_/A sky130_fd_sc_hd__buf_12
X_3517_ _6684_/Q _4279_/A _4139_/A _6559_/Q _3514_/X VGND VGND VPWR VPWR _3518_/D
+ sky130_fd_sc_hd__a221o_1
Xhold655 _4259_/X VGND VGND VPWR VPWR _6663_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_575 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xmax_cap374 _3552_/A VGND VGND VPWR VPWR _3553_/A sky130_fd_sc_hd__buf_12
XFILLER_103_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold666 _5385_/X VGND VGND VPWR VPWR _6943_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4497_ _5043_/A _4862_/A VGND VGND VPWR VPWR _4526_/C sky130_fd_sc_hd__nor2_1
Xmax_cap385 _5937_/X VGND VGND VPWR VPWR _6288_/A2 sky130_fd_sc_hd__buf_12
Xhold677 _6953_/Q VGND VGND VPWR VPWR hold677/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_131_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmax_cap396 _5936_/X VGND VGND VPWR VPWR _6259_/A2 sky130_fd_sc_hd__buf_12
XFILLER_103_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold688 _5466_/X VGND VGND VPWR VPWR _7015_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6236_ _6717_/Q _5955_/X _5975_/C _6702_/Q VGND VGND VPWR VPWR _6236_/X sky130_fd_sc_hd__a22o_1
Xhold699 _6895_/Q VGND VGND VPWR VPWR hold699/X sky130_fd_sc_hd__dlygate4sd3_1
X_3448_ input49/X _4103_/B hold34/A _6991_/Q VGND VGND VPWR VPWR _3448_/X sky130_fd_sc_hd__a22o_1
XFILLER_131_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6167_ _6167_/A _6167_/B VGND VGND VPWR VPWR _6167_/Y sky130_fd_sc_hd__nor2_1
XFILLER_134_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3379_ _3552_/A _3391_/B VGND VGND VPWR VPWR _5379_/A sky130_fd_sc_hd__nor2_8
Xhold1300 _4101_/X VGND VGND VPWR VPWR _6522_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1311 hold1397/X VGND VGND VPWR VPWR hold1311/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1322 hold1322/A VGND VGND VPWR VPWR wb_dat_o[13] sky130_fd_sc_hd__buf_12
XTAP_993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5118_ _5118_/A _5118_/B _5118_/C VGND VGND VPWR VPWR _5119_/B sky130_fd_sc_hd__nor3_1
Xhold1333 _4187_/A1 VGND VGND VPWR VPWR hold1333/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1344 hold1344/A VGND VGND VPWR VPWR wb_dat_o[1] sky130_fd_sc_hd__buf_12
X_6098_ _6446_/Q _5601_/Y _6296_/A2 _6886_/Q VGND VGND VPWR VPWR _6098_/X sky130_fd_sc_hd__a22o_1
Xhold1355 _6310_/A1 VGND VGND VPWR VPWR hold1355/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1366 hold1366/A VGND VGND VPWR VPWR wb_dat_o[4] sky130_fd_sc_hd__buf_12
Xhold1377 _7154_/Q VGND VGND VPWR VPWR _6356_/A0 sky130_fd_sc_hd__dlygate4sd3_1
X_5049_ _4745_/B _4973_/B _5043_/X _4973_/A _4877_/B VGND VGND VPWR VPWR _5050_/A
+ sky130_fd_sc_hd__o221ai_1
XTAP_2805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1388 _6889_/Q VGND VGND VPWR VPWR _5324_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1399 _7138_/Q VGND VGND VPWR VPWR _6314_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_84_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_58 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_147 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_191_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_191_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_140_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_707 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_177_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4420_ _4513_/A _4692_/A VGND VGND VPWR VPWR _5017_/A sky130_fd_sc_hd__or2_1
XFILLER_129_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4351_ _4888_/A _4352_/B VGND VGND VPWR VPWR _4351_/Y sky130_fd_sc_hd__nor2_2
XFILLER_125_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3302_ hold31/X hold16/X hold58/A _3268_/X VGND VGND VPWR VPWR hold32/A sky130_fd_sc_hd__or4bb_4
X_7070_ _7070_/CLK _7070_/D fanout507/X VGND VGND VPWR VPWR _7070_/Q sky130_fd_sc_hd__dfrtp_1
X_4282_ hold399/X _5532_/A1 _4284_/S VGND VGND VPWR VPWR _4282_/X sky130_fd_sc_hd__mux2_1
X_6021_ _6979_/Q _5943_/Y _6299_/A2 _6795_/Q VGND VGND VPWR VPWR _6021_/X sky130_fd_sc_hd__a22o_1
X_3233_ _6416_/Q _6415_/Q VGND VGND VPWR VPWR _3234_/C sky130_fd_sc_hd__nand2b_1
XFILLER_101_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_1_1_1_csclk clkbuf_1_1_1_csclk/A VGND VGND VPWR VPWR clkbuf_2_3_0_csclk/A
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_39_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3164_ _7159_/Q VGND VGND VPWR VPWR _3164_/Y sky130_fd_sc_hd__inv_2
XFILLER_104_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6923_ _7011_/CLK _6923_/D fanout500/X VGND VGND VPWR VPWR _6923_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_35_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_510 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6854_ _6990_/CLK _6854_/D _6396_/A VGND VGND VPWR VPWR _6854_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_22_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5805_ _6849_/Q _5922_/B1 _5651_/X _6801_/Q _5803_/X VGND VGND VPWR VPWR _5805_/X
+ sky130_fd_sc_hd__a221o_1
X_6785_ _7022_/CLK hold77/X fanout517/X VGND VGND VPWR VPWR _6785_/Q sky130_fd_sc_hd__dfrtp_1
X_3997_ hold703/X _5542_/A1 _4001_/S VGND VGND VPWR VPWR _3997_/X sky130_fd_sc_hd__mux2_1
X_5736_ _7006_/Q _5912_/A2 _5922_/A2 _6910_/Q VGND VGND VPWR VPWR _5736_/X sky130_fd_sc_hd__a22o_1
X_5667_ _5667_/A _5667_/B VGND VGND VPWR VPWR _5667_/X sky130_fd_sc_hd__or2_4
XFILLER_136_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_135_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4618_ _4678_/A _4721_/B VGND VGND VPWR VPWR _4695_/B sky130_fd_sc_hd__or2_4
X_5598_ _5598_/A _5598_/B VGND VGND VPWR VPWR _7101_/D sky130_fd_sc_hd__and2_1
XFILLER_190_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold430 _5184_/X VGND VGND VPWR VPWR _6765_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_151_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_163_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold441 _7054_/Q VGND VGND VPWR VPWR hold441/X sky130_fd_sc_hd__dlygate4sd3_1
X_4549_ _4622_/A _4549_/B VGND VGND VPWR VPWR _4959_/C sky130_fd_sc_hd__nor2_2
XFILLER_104_512 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold452 _5314_/X VGND VGND VPWR VPWR _6880_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_2_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold463 _6484_/Q VGND VGND VPWR VPWR hold463/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold474 _5233_/X VGND VGND VPWR VPWR _6808_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold485 _6648_/Q VGND VGND VPWR VPWR hold485/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold496 _4307_/X VGND VGND VPWR VPWR _6703_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6219_ _6579_/Q _5946_/X _5959_/Y _6615_/Q VGND VGND VPWR VPWR _6219_/X sky130_fd_sc_hd__a22o_1
XFILLER_104_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7199_ _7199_/A VGND VGND VPWR VPWR _7199_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_58_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1130 _5429_/X VGND VGND VPWR VPWR _6982_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1141 _7043_/Q VGND VGND VPWR VPWR _5498_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_73_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1152 _5236_/X VGND VGND VPWR VPWR _6810_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_73_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_161_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_315 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1163 _6560_/Q VGND VGND VPWR VPWR _4146_/A0 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1174 _4015_/X VGND VGND VPWR VPWR _6460_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1185 _6737_/Q VGND VGND VPWR VPWR _5146_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1196 _5362_/X VGND VGND VPWR VPWR _6922_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_543 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_407 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_91_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3920_ _6512_/Q _3247_/A _6406_/Q VGND VGND VPWR VPWR _3920_/X sky130_fd_sc_hd__mux2_1
XFILLER_32_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3851_ hold71/A _6488_/Q _3844_/Y _3850_/X VGND VGND VPWR VPWR _3851_/X sky130_fd_sc_hd__a22o_1
XFILLER_149_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_576 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6570_ _7137_/CLK _6570_/D VGND VGND VPWR VPWR _6570_/Q sky130_fd_sc_hd__dfxtp_1
X_3782_ input61/X _4096_/A _3493_/Y _3780_/X _3781_/X VGND VGND VPWR VPWR _3782_/X
+ sky130_fd_sc_hd__a2111o_1
X_5521_ _5521_/A0 _5521_/A1 _5528_/S VGND VGND VPWR VPWR _5521_/X sky130_fd_sc_hd__mux2_1
XFILLER_173_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5452_ _5452_/A0 _5530_/A1 _5459_/S VGND VGND VPWR VPWR _5452_/X sky130_fd_sc_hd__mux2_1
XFILLER_172_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_117_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4403_ _4403_/A _4495_/A VGND VGND VPWR VPWR _4472_/A sky130_fd_sc_hd__or2_1
XFILLER_133_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5383_ hold741/X _5542_/A1 _5387_/S VGND VGND VPWR VPWR _5383_/X sky130_fd_sc_hd__mux2_1
X_7122_ _7123_/CLK _7122_/D fanout499/X VGND VGND VPWR VPWR _7122_/Q sky130_fd_sc_hd__dfrtp_1
X_4334_ _4334_/A _4334_/B _4334_/C _4334_/D VGND VGND VPWR VPWR _4337_/A sky130_fd_sc_hd__and4_1
XFILLER_125_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7053_ _7054_/CLK _7053_/D fanout503/X VGND VGND VPWR VPWR _7053_/Q sky130_fd_sc_hd__dfrtp_2
X_4265_ hold624/X _4289_/A1 _4266_/S VGND VGND VPWR VPWR _4265_/X sky130_fd_sc_hd__mux2_1
XFILLER_99_598 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6004_ _6786_/Q _6004_/B VGND VGND VPWR VPWR _6004_/X sky130_fd_sc_hd__or2_1
XFILLER_86_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3216_ _6829_/Q VGND VGND VPWR VPWR _3216_/Y sky130_fd_sc_hd__inv_2
XFILLER_101_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4196_ _4196_/A _6352_/B VGND VGND VPWR VPWR _4201_/S sky130_fd_sc_hd__and2_2
XFILLER_27_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_292 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6906_ _7011_/CLK _6906_/D fanout500/X VGND VGND VPWR VPWR _6906_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_54_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_690 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6837_ _7058_/CLK _6837_/D fanout521/X VGND VGND VPWR VPWR _6837_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_50_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6768_ _6769_/CLK _6768_/D fanout492/X VGND VGND VPWR VPWR _6768_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_149_751 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5719_ _6445_/Q _5917_/B1 _5650_/X _6893_/Q VGND VGND VPWR VPWR _5719_/X sky130_fd_sc_hd__a22o_1
X_6699_ _6699_/CLK _6699_/D fanout510/X VGND VGND VPWR VPWR _6699_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_108_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_163_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold260 _4253_/X VGND VGND VPWR VPWR _6658_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold271 hold271/A VGND VGND VPWR VPWR hold271/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold282 _5409_/X VGND VGND VPWR VPWR _6964_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold293 hold293/A VGND VGND VPWR VPWR hold293/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_49_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_105_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_100_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_100 _3943_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_111 _7199_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_122 _3894_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_133 _6440_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_144 _5519_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_155 _5923_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_166 _5288_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_177 _5528_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_188 _6805_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_199 _6294_/A2 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_146_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_186_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_155_710 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_423 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_448 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_110_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_695 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4050_ hold293/X _5541_/A1 _4103_/B VGND VGND VPWR VPWR _4050_/X sky130_fd_sc_hd__mux2_1
XFILLER_110_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput6 mask_rev_in[11] VGND VGND VPWR VPWR input6/X sky130_fd_sc_hd__clkbuf_1
XFILLER_76_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_318 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4952_ _4587_/A _4828_/A _4537_/B _5026_/B VGND VGND VPWR VPWR _4955_/B sky130_fd_sc_hd__a31o_1
XFILLER_17_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3903_ _3903_/A _3903_/B VGND VGND VPWR VPWR _6635_/D sky130_fd_sc_hd__nand2_1
X_4883_ _4883_/A _4915_/A _4883_/C VGND VGND VPWR VPWR _5020_/B sky130_fd_sc_hd__and3_1
XFILLER_177_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3834_ _3273_/Y hold15/A _3837_/B VGND VGND VPWR VPWR _3834_/X sky130_fd_sc_hd__mux2_1
X_6622_ _7155_/CLK hold66/X _6370_/A VGND VGND VPWR VPWR hold65/A sky130_fd_sc_hd__dfrtp_1
XFILLER_20_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_165_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6553_ _6708_/CLK _6553_/D _6400_/A VGND VGND VPWR VPWR _6553_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_192_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3765_ _6930_/Q hold41/A _4231_/A _6630_/Q _3764_/X VGND VGND VPWR VPWR _3768_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_158_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5504_ hold971/X _5531_/A1 _5510_/S VGND VGND VPWR VPWR _5504_/X sky130_fd_sc_hd__mux2_1
XFILLER_173_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6484_ _6632_/CLK _6484_/D fanout509/X VGND VGND VPWR VPWR _6484_/Q sky130_fd_sc_hd__dfrtp_1
X_3696_ _6891_/Q _5325_/A _4303_/A _6701_/Q _3695_/X VGND VGND VPWR VPWR _3697_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_118_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_146_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xpad_flashh_clk_buff_inst _3939_/X VGND VGND VPWR VPWR pad_flash_clk sky130_fd_sc_hd__clkbuf_8
X_5435_ _5435_/A0 hold90/X hold35/X VGND VGND VPWR VPWR hold95/A sky130_fd_sc_hd__mux2_1
XFILLER_10_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput310 _3947_/X VGND VGND VPWR VPWR spimemio_flash_io1_di sky130_fd_sc_hd__buf_12
Xoutput321 hold1335/X VGND VGND VPWR VPWR hold1336/A sky130_fd_sc_hd__buf_12
XFILLER_133_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput332 hold1345/X VGND VGND VPWR VPWR hold1346/A sky130_fd_sc_hd__buf_12
XFILLER_126_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput343 hold1319/X VGND VGND VPWR VPWR hold1320/A sky130_fd_sc_hd__buf_12
X_5366_ _5366_/A0 _5543_/A1 _5369_/S VGND VGND VPWR VPWR _5366_/X sky130_fd_sc_hd__mux2_1
XFILLER_87_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4317_ hold977/X _6354_/A1 _4320_/S VGND VGND VPWR VPWR _4317_/X sky130_fd_sc_hd__mux2_1
X_7105_ _7131_/CLK _7105_/D fanout501/X VGND VGND VPWR VPWR _7105_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_87_524 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5297_ hold691/X _5537_/A1 _5297_/S VGND VGND VPWR VPWR _5297_/X sky130_fd_sc_hd__mux2_1
XFILLER_101_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7036_ _7037_/CLK _7036_/D fanout485/X VGND VGND VPWR VPWR _7036_/Q sky130_fd_sc_hd__dfstp_2
X_4248_ hold307/X _6357_/A1 hold63/X VGND VGND VPWR VPWR _4248_/X sky130_fd_sc_hd__mux2_1
XFILLER_142_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_410 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4179_ _3433_/X _4179_/A1 _4180_/S VGND VGND VPWR VPWR _6589_/D sky130_fd_sc_hd__mux2_1
XFILLER_67_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_34 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_156_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_167_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_528 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_149_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_183_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_183_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_183_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_41_csclk clkbuf_3_6_0_csclk/X VGND VGND VPWR VPWR _7017_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_2273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_186_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_119_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_56_csclk _7000_/CLK VGND VGND VPWR VPWR _7054_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_186_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3550_ input30/X _3339_/Y _4008_/A _6459_/Q VGND VGND VPWR VPWR _3550_/X sky130_fd_sc_hd__a22o_1
XFILLER_155_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3481_ hold61/X _3554_/B VGND VGND VPWR VPWR _4231_/A sky130_fd_sc_hd__nor2_8
XFILLER_115_459 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5220_ hold331/X _5523_/A1 _5225_/S VGND VGND VPWR VPWR _5220_/X sky130_fd_sc_hd__mux2_1
XFILLER_44_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5151_ _5151_/A _6352_/B VGND VGND VPWR VPWR _5157_/S sky130_fd_sc_hd__and2_2
XFILLER_170_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4102_ hold407/X _5526_/A1 hold8/X VGND VGND VPWR VPWR _4102_/X sky130_fd_sc_hd__mux2_1
XFILLER_96_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5082_ _4972_/A _5043_/X _5055_/C _4877_/C _4973_/X VGND VGND VPWR VPWR _5082_/X
+ sky130_fd_sc_hd__o2111a_1
XFILLER_96_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4033_ _4033_/A0 _6353_/A1 _4037_/S VGND VGND VPWR VPWR _4033_/X sky130_fd_sc_hd__mux2_1
XFILLER_49_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5984_ _7010_/Q _5976_/Y _5979_/X _6970_/Q VGND VGND VPWR VPWR _5984_/X sky130_fd_sc_hd__a22o_1
XFILLER_24_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4935_ _4935_/A _4935_/B _4921_/Y VGND VGND VPWR VPWR _4935_/X sky130_fd_sc_hd__or3b_1
Xclkbuf_3_7_0_csclk clkbuf_3_7_0_csclk/A VGND VGND VPWR VPWR clkbuf_3_7_0_csclk/X
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA_11 _5424_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_22 _5520_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4866_ _4901_/B _4719_/B _4695_/B _4748_/B VGND VGND VPWR VPWR _4868_/C sky130_fd_sc_hd__o22a_1
XFILLER_20_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_33 _3461_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6605_ _6707_/CLK _6605_/D fanout485/X VGND VGND VPWR VPWR _6605_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_20_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_44 _3648_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_177_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3817_ _7170_/Q _6487_/Q _3817_/C VGND VGND VPWR VPWR _3817_/X sky130_fd_sc_hd__and3_1
XANTENNA_55 _5622_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4797_ _4479_/A _4640_/B _4725_/B _4703_/B VGND VGND VPWR VPWR _4813_/C sky130_fd_sc_hd__o22a_1
XANTENNA_66 _6933_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_165_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_77 user_clock VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_88 _3943_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6536_ _6969_/CLK _6536_/D fanout506/X VGND VGND VPWR VPWR _6536_/Q sky130_fd_sc_hd__dfrtp_1
X_3748_ _6727_/Q _3747_/Y _3817_/C VGND VGND VPWR VPWR _3748_/X sky130_fd_sc_hd__mux2_1
XANTENNA_99 _3943_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_118_264 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_192_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6467_ _7037_/CLK _6467_/D fanout484/X VGND VGND VPWR VPWR _6467_/Q sky130_fd_sc_hd__dfstp_4
X_3679_ _7020_/Q hold18/A hold41/A _6932_/Q VGND VGND VPWR VPWR _3679_/X sky130_fd_sc_hd__a22o_1
XFILLER_134_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5418_ hold283/X _5541_/A1 _5423_/S VGND VGND VPWR VPWR _5418_/X sky130_fd_sc_hd__mux2_1
X_6398_ _6399_/A _6399_/B VGND VGND VPWR VPWR _6398_/X sky130_fd_sc_hd__and2_1
XFILLER_161_587 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput173 _3953_/X VGND VGND VPWR VPWR irq[1] sky130_fd_sc_hd__buf_12
XFILLER_0_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5349_ hold667/X _5544_/A1 _5351_/S VGND VGND VPWR VPWR _5349_/X sky130_fd_sc_hd__mux2_1
Xoutput184 _3202_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[18] sky130_fd_sc_hd__buf_12
Xoutput195 _3192_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[28] sky130_fd_sc_hd__buf_12
XFILLER_99_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7019_ _7022_/CLK _7019_/D fanout525/X VGND VGND VPWR VPWR _7019_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_28_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_262 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_168_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_169_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_440 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4720_ _4720_/A _4720_/B _4720_/C _5008_/B VGND VGND VPWR VPWR _4720_/X sky130_fd_sc_hd__or4b_2
XTAP_1391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4651_ _4788_/A _4985_/B VGND VGND VPWR VPWR _5057_/A sky130_fd_sc_hd__nor2_1
XFILLER_187_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput20 mask_rev_in[24] VGND VGND VPWR VPWR input20/X sky130_fd_sc_hd__clkbuf_2
X_3602_ _6949_/Q _5388_/A _4273_/A _6678_/Q _3601_/X VGND VGND VPWR VPWR _3605_/C
+ sky130_fd_sc_hd__a221o_1
Xinput31 mask_rev_in[5] VGND VGND VPWR VPWR input31/X sky130_fd_sc_hd__clkbuf_4
XFILLER_174_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4582_ _4862_/A _4748_/B VGND VGND VPWR VPWR _4851_/B sky130_fd_sc_hd__nor2_1
Xinput42 mgmt_gpio_in[15] VGND VGND VPWR VPWR input42/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_116_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput53 mgmt_gpio_in[25] VGND VGND VPWR VPWR input53/X sky130_fd_sc_hd__buf_2
Xinput64 mgmt_gpio_in[35] VGND VGND VPWR VPWR input64/X sky130_fd_sc_hd__buf_2
Xinput75 porb VGND VGND VPWR VPWR input75/X sky130_fd_sc_hd__clkbuf_1
Xhold804 _5154_/X VGND VGND VPWR VPWR _6744_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3533_ _3533_/A _3761_/B VGND VGND VPWR VPWR _4202_/A sky130_fd_sc_hd__nor2_4
X_6321_ _6642_/Q _6318_/Y _6320_/Y _6644_/Q _4222_/X VGND VGND VPWR VPWR _6322_/A
+ sky130_fd_sc_hd__a221o_1
Xhold815 _6562_/Q VGND VGND VPWR VPWR hold815/X sky130_fd_sc_hd__dlygate4sd3_1
Xinput86 spimemio_flash_io0_oeb VGND VGND VPWR VPWR _3941_/B sky130_fd_sc_hd__clkbuf_4
Xhold826 _4211_/X VGND VGND VPWR VPWR _6616_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold837 _6697_/Q VGND VGND VPWR VPWR hold837/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput97 usr2_vcc_pwrgood VGND VGND VPWR VPWR input97/X sky130_fd_sc_hd__buf_2
Xhold848 _5414_/X VGND VGND VPWR VPWR _6969_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6252_ _6252_/A _6252_/B _6252_/C _6004_/B VGND VGND VPWR VPWR _6252_/X sky130_fd_sc_hd__or4b_1
XFILLER_115_245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3464_ _6983_/Q _5424_/A _3360_/Y input8/X VGND VGND VPWR VPWR _3464_/X sky130_fd_sc_hd__a22o_1
Xhold859 _6949_/Q VGND VGND VPWR VPWR hold859/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_115_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_587 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5203_ hold519/X _5515_/A1 _5207_/S VGND VGND VPWR VPWR _5203_/X sky130_fd_sc_hd__mux2_1
X_6183_ _6660_/Q _6294_/A2 _5969_/C _6710_/Q VGND VGND VPWR VPWR _6183_/X sky130_fd_sc_hd__a22o_1
X_3395_ _3395_/A _3395_/B _3395_/C _3395_/D VGND VGND VPWR VPWR _3395_/Y sky130_fd_sc_hd__nor4_1
XFILLER_97_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5134_ _5134_/A _5134_/B _5133_/X VGND VGND VPWR VPWR _5134_/X sky130_fd_sc_hd__or3b_1
XFILLER_57_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1504 _6417_/Q VGND VGND VPWR VPWR _3165_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1515 _6403_/Q VGND VGND VPWR VPWR _3863_/B1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_97_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1526 _6525_/Q VGND VGND VPWR VPWR hold126/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1537 _7093_/Q VGND VGND VPWR VPWR _5572_/B1 sky130_fd_sc_hd__dlygate4sd3_1
X_5065_ _5065_/A _5065_/B _5065_/C VGND VGND VPWR VPWR _5065_/Y sky130_fd_sc_hd__nand3_1
Xhold1548 _7181_/A VGND VGND VPWR VPWR hold1548/X sky130_fd_sc_hd__dlygate4sd3_1
X_4016_ _4016_/A0 _6354_/A1 _4019_/S VGND VGND VPWR VPWR _4016_/X sky130_fd_sc_hd__mux2_1
XFILLER_37_251 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5967_ _7099_/Q _5981_/A _5963_/C _5939_/X _5951_/X VGND VGND VPWR VPWR _5969_/B
+ sky130_fd_sc_hd__a311o_1
XFILLER_40_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4918_ _4513_/A _5026_/A _4713_/A _4861_/B _4817_/C VGND VGND VPWR VPWR _5064_/A
+ sky130_fd_sc_hd__o221a_1
X_5898_ _6718_/Q _5648_/X _5919_/B1 _6633_/Q VGND VGND VPWR VPWR _5898_/X sky130_fd_sc_hd__a22o_1
XFILLER_193_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_193_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4849_ _4588_/B _4831_/X _4847_/X _4848_/Y VGND VGND VPWR VPWR _4850_/D sky130_fd_sc_hd__o211a_1
XFILLER_148_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_166_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6519_ _6711_/CLK _6519_/D fanout486/X VGND VGND VPWR VPWR _6519_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_107_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_543 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_164_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_313 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_240 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_189_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_189_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_189_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_630 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3180_ _6914_/Q VGND VGND VPWR VPWR _3180_/Y sky130_fd_sc_hd__inv_2
XFILLER_93_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6870_ _6988_/CLK _6870_/D _6396_/A VGND VGND VPWR VPWR _6870_/Q sky130_fd_sc_hd__dfrtp_1
X_5821_ _6793_/Q _5667_/X _5812_/X _5820_/X _3174_/Y VGND VGND VPWR VPWR _5821_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_22_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5752_ _6446_/Q _5917_/B1 _5925_/B1 hold86/A VGND VGND VPWR VPWR _5752_/X sky130_fd_sc_hd__a22o_1
X_4703_ _4703_/A _4703_/B VGND VGND VPWR VPWR _4703_/Y sky130_fd_sc_hd__nor2_1
XFILLER_187_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5683_ _6907_/Q _5922_/A2 _5679_/X _5682_/X VGND VGND VPWR VPWR _5683_/X sky130_fd_sc_hd__a211o_1
XFILLER_148_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4634_ _4634_/A _4634_/B VGND VGND VPWR VPWR _4784_/B sky130_fd_sc_hd__or2_1
XFILLER_147_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold601 _4042_/X VGND VGND VPWR VPWR _6483_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4565_ _4943_/B _4565_/B VGND VGND VPWR VPWR _4566_/B sky130_fd_sc_hd__nor2_1
Xhold612 _6952_/Q VGND VGND VPWR VPWR hold612/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold623 _4137_/X VGND VGND VPWR VPWR _6553_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6304_ _6507_/Q _7130_/Q _5611_/X VGND VGND VPWR VPWR _6304_/X sky130_fd_sc_hd__a21o_1
Xhold634 _6840_/Q VGND VGND VPWR VPWR hold634/X sky130_fd_sc_hd__dlygate4sd3_1
Xmax_cap353 _3343_/Y VGND VGND VPWR VPWR _4103_/B sky130_fd_sc_hd__buf_8
X_3516_ _3531_/A hold53/A VGND VGND VPWR VPWR _4139_/A sky130_fd_sc_hd__nor2_4
Xhold645 _5545_/X VGND VGND VPWR VPWR _7085_/D sky130_fd_sc_hd__dlygate4sd3_1
Xmax_cap364 _5980_/Y VGND VGND VPWR VPWR _6290_/B1 sky130_fd_sc_hd__buf_12
Xhold656 _7070_/Q VGND VGND VPWR VPWR hold656/X sky130_fd_sc_hd__dlygate4sd3_1
X_4496_ _4692_/A _4586_/B VGND VGND VPWR VPWR _5135_/A sky130_fd_sc_hd__or2_1
XFILLER_131_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmax_cap375 _5981_/X VGND VGND VPWR VPWR _6270_/B1 sky130_fd_sc_hd__buf_12
XFILLER_116_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold667 _6911_/Q VGND VGND VPWR VPWR hold667/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_143_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xmax_cap386 _5971_/B VGND VGND VPWR VPWR _6284_/B1 sky130_fd_sc_hd__buf_8
Xhold678 _5396_/X VGND VGND VPWR VPWR _6953_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_cap397 _5651_/X VGND VGND VPWR VPWR _5926_/B1 sky130_fd_sc_hd__buf_12
X_6235_ _6707_/Q _5957_/X _5978_/X _6697_/Q VGND VGND VPWR VPWR _6235_/X sky130_fd_sc_hd__a22o_1
XFILLER_89_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3447_ _6447_/Q _3993_/A _5307_/A _6879_/Q _3446_/X VGND VGND VPWR VPWR _3471_/B
+ sky130_fd_sc_hd__a221o_1
Xhold689 _6807_/Q VGND VGND VPWR VPWR hold689/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_134_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6166_ _6921_/Q _5937_/X _5975_/C _7054_/Q _6165_/X VGND VGND VPWR VPWR _6167_/B
+ sky130_fd_sc_hd__a221o_1
X_3378_ hold61/X _3391_/B VGND VGND VPWR VPWR _5307_/A sky130_fd_sc_hd__nor2_8
XTAP_961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1301 _6822_/Q VGND VGND VPWR VPWR _5249_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1312 hold1312/A VGND VGND VPWR VPWR wb_dat_o[22] sky130_fd_sc_hd__buf_12
XTAP_994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1323 _4174_/A1 VGND VGND VPWR VPWR hold1323/X sky130_fd_sc_hd__dlygate4sd3_1
X_5117_ _4719_/B _4973_/B _5114_/X _5138_/B _4868_/C VGND VGND VPWR VPWR _5120_/A
+ sky130_fd_sc_hd__o2111a_1
Xhold1334 hold1334/A VGND VGND VPWR VPWR wb_dat_o[5] sky130_fd_sc_hd__buf_12
XFILLER_111_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6097_ _6798_/Q _6299_/A2 _6282_/B1 _6974_/Q _6096_/X VGND VGND VPWR VPWR _6102_/B
+ sky130_fd_sc_hd__a221o_1
Xhold1345 _6311_/A1 VGND VGND VPWR VPWR hold1345/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1356 hold1356/A VGND VGND VPWR VPWR wb_dat_o[25] sky130_fd_sc_hd__buf_12
Xhold1367 _6313_/A1 VGND VGND VPWR VPWR hold1367/X sky130_fd_sc_hd__dlygate4sd3_1
X_5048_ _5048_/A _5068_/A _5047_/X VGND VGND VPWR VPWR _5118_/A sky130_fd_sc_hd__or3b_1
XFILLER_72_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1378 _6900_/Q VGND VGND VPWR VPWR _5337_/A0 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1389 _6902_/Q VGND VGND VPWR VPWR _5339_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6999_ _6999_/CLK _6999_/D fanout523/X VGND VGND VPWR VPWR _6999_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_13_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_179_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_159_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_335 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_177_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4350_ _4352_/B _4350_/B VGND VGND VPWR VPWR _4888_/B sky130_fd_sc_hd__or2_4
XFILLER_153_660 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3301_ _3571_/A hold75/X VGND VGND VPWR VPWR hold76/A sky130_fd_sc_hd__nor2_8
X_4281_ hold559/X _4299_/A1 _4284_/S VGND VGND VPWR VPWR _4281_/X sky130_fd_sc_hd__mux2_1
XFILLER_99_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6020_ _6987_/Q _5941_/Y _5962_/X _6891_/Q _6019_/X VGND VGND VPWR VPWR _6026_/C
+ sky130_fd_sc_hd__a221o_1
X_3232_ _6417_/Q _6416_/Q VGND VGND VPWR VPWR _3259_/B sky130_fd_sc_hd__and2_1
XFILLER_67_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_302 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6922_ _7010_/CLK _6922_/D fanout498/X VGND VGND VPWR VPWR _6922_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_82_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6853_ _7058_/CLK _6853_/D fanout521/X VGND VGND VPWR VPWR _6853_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_50_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5804_ _6993_/Q _5622_/X _5624_/X _6833_/Q VGND VGND VPWR VPWR _5804_/X sky130_fd_sc_hd__a22o_1
X_6784_ _7058_/CLK _6784_/D fanout521/X VGND VGND VPWR VPWR _6784_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_22_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3996_ hold279/X _5541_/A1 _4001_/S VGND VGND VPWR VPWR _3996_/X sky130_fd_sc_hd__mux2_1
XFILLER_10_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5735_ _5756_/A1 _6305_/A2 _5733_/X _5734_/X VGND VGND VPWR VPWR _5735_/X sky130_fd_sc_hd__o22a_1
XFILLER_148_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5666_ _6994_/Q _5646_/X _5662_/X _5665_/X _5638_/X VGND VGND VPWR VPWR _5666_/X
+ sky130_fd_sc_hd__a2111o_1
XFILLER_108_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4617_ _4617_/A _4617_/B _4888_/A VGND VGND VPWR VPWR _4620_/B sky130_fd_sc_hd__or3b_4
XFILLER_190_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5597_ _7101_/Q _5597_/B _5596_/B VGND VGND VPWR VPWR _5598_/B sky130_fd_sc_hd__or3b_1
XFILLER_116_340 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold420 _5377_/X VGND VGND VPWR VPWR _6936_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold431 _6549_/Q VGND VGND VPWR VPWR hold431/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_190_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4548_ _4622_/A _4943_/B _4581_/A _4547_/X _4546_/X VGND VGND VPWR VPWR _4548_/X
+ sky130_fd_sc_hd__o221a_1
Xhold442 _5510_/X VGND VGND VPWR VPWR _7054_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold453 _6980_/Q VGND VGND VPWR VPWR hold453/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold464 _4043_/X VGND VGND VPWR VPWR _6484_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold475 _6669_/Q VGND VGND VPWR VPWR hold475/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_1_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold486 _4241_/X VGND VGND VPWR VPWR _6648_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4479_ _4479_/A _4549_/B VGND VGND VPWR VPWR _4506_/C sky130_fd_sc_hd__or2_1
Xhold497 _6740_/Q VGND VGND VPWR VPWR hold497/X sky130_fd_sc_hd__dlygate4sd3_1
X_6218_ _6218_/A _6218_/B _6218_/C _6217_/Y VGND VGND VPWR VPWR _6218_/X sky130_fd_sc_hd__or4b_1
X_7198_ _7198_/A VGND VGND VPWR VPWR _7198_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_161_14 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6149_ _6912_/Q _5972_/A _5977_/X _6928_/Q VGND VGND VPWR VPWR _6149_/X sky130_fd_sc_hd__a22o_1
XFILLER_85_430 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1120 _5483_/X VGND VGND VPWR VPWR _7030_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1131 _6934_/Q VGND VGND VPWR VPWR _5375_/A0 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1142 _5498_/X VGND VGND VPWR VPWR _7043_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1153 _6938_/Q VGND VGND VPWR VPWR _5380_/A0 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1164 _4146_/X VGND VGND VPWR VPWR _6560_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_161_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1175 _6700_/Q VGND VGND VPWR VPWR _4304_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1186 _5146_/X VGND VGND VPWR VPWR _6737_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1197 hold1549/X VGND VGND VPWR VPWR _4113_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_72_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_371 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_135_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_141_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_91_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_177_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3850_ hold71/A hold78/A hold37/A VGND VGND VPWR VPWR _3850_/X sky130_fd_sc_hd__a21o_1
XFILLER_32_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3781_ _7071_/Q _5529_/A _5538_/A _7079_/Q VGND VGND VPWR VPWR _3781_/X sky130_fd_sc_hd__a22o_1
X_5520_ _5520_/A _5538_/B VGND VGND VPWR VPWR _5528_/S sky130_fd_sc_hd__and2_4
XFILLER_74_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_185_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5451_ _5451_/A hold6/X VGND VGND VPWR VPWR _5459_/S sky130_fd_sc_hd__and2_4
XFILLER_160_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4402_ _4888_/A _4402_/B VGND VGND VPWR VPWR _4495_/A sky130_fd_sc_hd__nand2b_1
XFILLER_172_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5382_ hold425/X _5541_/A1 _5387_/S VGND VGND VPWR VPWR _5382_/X sky130_fd_sc_hd__mux2_1
X_7121_ _7123_/CLK _7121_/D fanout499/X VGND VGND VPWR VPWR _7121_/Q sky130_fd_sc_hd__dfrtp_1
X_4333_ _4575_/A _4746_/B VGND VGND VPWR VPWR _5043_/A sky130_fd_sc_hd__or2_4
XFILLER_141_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4264_ hold409/X _5532_/A1 _4266_/S VGND VGND VPWR VPWR _4264_/X sky130_fd_sc_hd__mux2_1
XFILLER_101_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7052_ _7069_/CLK _7052_/D fanout516/X VGND VGND VPWR VPWR _7052_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_87_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6003_ _6003_/A _6003_/B _6003_/C _6004_/B VGND VGND VPWR VPWR _6003_/X sky130_fd_sc_hd__or4b_1
X_3215_ _6837_/Q VGND VGND VPWR VPWR _3215_/Y sky130_fd_sc_hd__inv_2
XFILLER_140_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4195_ hold871/X _4236_/A1 _4195_/S VGND VGND VPWR VPWR _4195_/X sky130_fd_sc_hd__mux2_1
XFILLER_39_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6905_ _7032_/CLK _6905_/D fanout506/X VGND VGND VPWR VPWR _6905_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_24_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6836_ _7059_/CLK _6836_/D fanout517/X VGND VGND VPWR VPWR _6836_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_10_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6767_ _7079_/CLK _6767_/D fanout514/X VGND VGND VPWR VPWR _6767_/Q sky130_fd_sc_hd__dfrtp_4
X_3979_ hold525/X _5491_/A1 _3983_/S VGND VGND VPWR VPWR _3979_/X sky130_fd_sc_hd__mux2_1
XFILLER_149_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5718_ _7021_/Q _5929_/B1 _5915_/B1 _6861_/Q _5717_/X VGND VGND VPWR VPWR _5718_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_164_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6698_ _6698_/CLK _6698_/D _6401_/A VGND VGND VPWR VPWR _6698_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_108_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_163_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5649_ _5667_/A _5651_/B _5649_/C VGND VGND VPWR VPWR _5649_/X sky130_fd_sc_hd__and3_4
XFILLER_151_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold250 _4149_/X VGND VGND VPWR VPWR _6563_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold261 _6602_/Q VGND VGND VPWR VPWR hold261/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_151_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold272 _4119_/X VGND VGND VPWR VPWR _6538_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold283 _6972_/Q VGND VGND VPWR VPWR hold283/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold294 _4106_/X VGND VGND VPWR VPWR _6526_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_151 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_100_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_124 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_101 _3943_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_112 _3951_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_123 _3894_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_134 _6294_/B1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_145 _5526_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_156 _5923_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_167 hold142/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_178 _5629_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_544 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_189 _6821_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_1_0_csclk clkbuf_0_csclk/X VGND VGND VPWR VPWR clkbuf_1_1_1_csclk/A sky130_fd_sc_hd__clkbuf_8
XFILLER_155_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_435 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_630 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_490 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput7 mask_rev_in[12] VGND VGND VPWR VPWR input7/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_64_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4951_ _4489_/B _4832_/Y _4947_/X _4920_/A VGND VGND VPWR VPWR _4951_/X sky130_fd_sc_hd__a211o_1
XFILLER_17_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3902_ _6306_/B _3908_/B VGND VGND VPWR VPWR _3903_/B sky130_fd_sc_hd__or2_1
XFILLER_32_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4882_ _4881_/X _4853_/X _5040_/B _4882_/B2 VGND VGND VPWR VPWR _6721_/D sky130_fd_sc_hd__o2bb2a_1
XFILLER_32_352 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6621_ _6633_/CLK _6621_/D _6370_/A VGND VGND VPWR VPWR _6621_/Q sky130_fd_sc_hd__dfstp_1
X_3833_ hold14/A hold56/A hold29/A _3845_/S VGND VGND VPWR VPWR _3837_/B sky130_fd_sc_hd__nand4_1
X_6552_ _6633_/CLK _6552_/D _6370_/A VGND VGND VPWR VPWR _6552_/Q sky130_fd_sc_hd__dfstp_1
X_3764_ _6842_/Q _5271_/A _5262_/A _6834_/Q VGND VGND VPWR VPWR _3764_/X sky130_fd_sc_hd__a22o_1
X_5503_ _5503_/A0 _5530_/A1 _5510_/S VGND VGND VPWR VPWR _5503_/X sky130_fd_sc_hd__mux2_1
X_6483_ _6718_/CLK _6483_/D _6401_/A VGND VGND VPWR VPWR _6483_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_146_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3695_ _6743_/Q _5151_/A _5487_/A _7035_/Q VGND VGND VPWR VPWR _3695_/X sky130_fd_sc_hd__a22o_1
XFILLER_133_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput300 _6754_/Q VGND VGND VPWR VPWR pwr_ctrl_out[3] sky130_fd_sc_hd__buf_12
X_5434_ _5434_/A0 _5521_/A1 hold35/X VGND VGND VPWR VPWR _5434_/X sky130_fd_sc_hd__mux2_1
Xoutput311 _7199_/X VGND VGND VPWR VPWR spimemio_flash_io2_di sky130_fd_sc_hd__buf_12
XFILLER_105_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput322 hold1337/X VGND VGND VPWR VPWR hold1338/A sky130_fd_sc_hd__buf_12
XFILLER_133_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput333 hold1361/X VGND VGND VPWR VPWR hold1362/A sky130_fd_sc_hd__buf_12
Xoutput344 hold1331/X VGND VGND VPWR VPWR hold1332/A sky130_fd_sc_hd__buf_12
XFILLER_126_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5365_ hold509/X _5515_/A1 _5369_/S VGND VGND VPWR VPWR _5365_/X sky130_fd_sc_hd__mux2_1
XFILLER_160_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7104_ _7124_/CLK _7104_/D fanout501/X VGND VGND VPWR VPWR _7104_/Q sky130_fd_sc_hd__dfrtp_1
Xclkbuf_3_3_0_csclk clkbuf_3_3_0_csclk/A VGND VGND VPWR VPWR _7000_/CLK sky130_fd_sc_hd__clkbuf_8
X_4316_ _4316_/A0 _6353_/A1 _4320_/S VGND VGND VPWR VPWR _4316_/X sky130_fd_sc_hd__mux2_1
XFILLER_99_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5296_ hold447/X _5545_/A1 _5297_/S VGND VGND VPWR VPWR _5296_/X sky130_fd_sc_hd__mux2_1
XFILLER_87_536 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7035_ _7037_/CLK _7035_/D fanout485/X VGND VGND VPWR VPWR _7035_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_75_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4247_ _4247_/A0 hold46/X hold63/X VGND VGND VPWR VPWR hold64/A sky130_fd_sc_hd__mux2_1
XFILLER_101_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4178_ _3471_/X _4178_/A1 _4180_/S VGND VGND VPWR VPWR _6588_/D sky130_fd_sc_hd__mux2_1
XFILLER_27_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_422 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_2_0_0_wb_clk_i clkbuf_2_1_0_wb_clk_i/A VGND VGND VPWR VPWR clkbuf_3_1_0_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_11_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6819_ _7074_/CLK _6819_/D fanout504/X VGND VGND VPWR VPWR _6819_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_23_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_167_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_183_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_435 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_137_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_611 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_455 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_159_368 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_530 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3480_ _6654_/Q hold62/A _4297_/A _6699_/Q VGND VGND VPWR VPWR _3480_/X sky130_fd_sc_hd__a22o_1
XFILLER_143_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5150_ hold413/X _5534_/A1 _5150_/S VGND VGND VPWR VPWR _5150_/X sky130_fd_sc_hd__mux2_1
XFILLER_37_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_644 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4101_ _4101_/A0 _5465_/A1 hold8/X VGND VGND VPWR VPWR _4101_/X sky130_fd_sc_hd__mux2_1
XFILLER_69_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5081_ _5081_/A _5081_/B _5081_/C _5081_/D VGND VGND VPWR VPWR _5118_/C sky130_fd_sc_hd__nand4_1
XFILLER_57_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4032_ _4032_/A hold7/X VGND VGND VPWR VPWR _4037_/S sky130_fd_sc_hd__and2_4
XFILLER_49_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5983_ _6810_/Q _6259_/A2 _6285_/A2 _6890_/Q VGND VGND VPWR VPWR _5983_/X sky130_fd_sc_hd__a22o_1
X_4934_ input99/X _4679_/Y _4924_/X _4902_/A VGND VGND VPWR VPWR _4934_/X sky130_fd_sc_hd__o211a_1
XFILLER_177_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4865_ _4965_/B _4962_/C _4556_/A VGND VGND VPWR VPWR _4960_/C sky130_fd_sc_hd__a21o_1
XANTENNA_12 _5415_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_23 _3396_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6604_ _6707_/CLK _6604_/D fanout485/X VGND VGND VPWR VPWR _6604_/Q sky130_fd_sc_hd__dfrtp_2
XANTENNA_34 _3471_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_193_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3816_ _3816_/A _3816_/B _3815_/X VGND VGND VPWR VPWR _3816_/X sky130_fd_sc_hd__or3b_4
XANTENNA_45 _3648_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_56 _5667_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4796_ _4515_/B _4921_/A _5043_/B _4972_/A VGND VGND VPWR VPWR _4818_/B sky130_fd_sc_hd__o22a_1
XANTENNA_67 _6797_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_192_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_78 user_clock VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6535_ _7054_/CLK _6535_/D fanout503/X VGND VGND VPWR VPWR _6535_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA_89 _3943_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3747_ _3747_/A _3747_/B VGND VGND VPWR VPWR _3747_/Y sky130_fd_sc_hd__nand2_4
XFILLER_146_552 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_319 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6466_ _7037_/CLK _6466_/D fanout484/X VGND VGND VPWR VPWR _6466_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_118_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_173_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3678_ _6868_/Q _5298_/A _5307_/A _6876_/Q _3677_/X VGND VGND VPWR VPWR _3683_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_173_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5417_ hold955/X _5495_/A1 _5423_/S VGND VGND VPWR VPWR _5417_/X sky130_fd_sc_hd__mux2_1
X_6397_ _6399_/A _6399_/B VGND VGND VPWR VPWR _6397_/X sky130_fd_sc_hd__and2_1
Xoutput174 _3954_/X VGND VGND VPWR VPWR irq[2] sky130_fd_sc_hd__buf_12
XFILLER_114_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5348_ _5348_/A0 _5465_/A1 _5351_/S VGND VGND VPWR VPWR _5348_/X sky130_fd_sc_hd__mux2_1
Xoutput185 _3201_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[19] sky130_fd_sc_hd__buf_12
Xoutput196 _3191_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[29] sky130_fd_sc_hd__buf_12
XFILLER_99_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5279_ hold919/X _5537_/A1 _5279_/S VGND VGND VPWR VPWR _5279_/X sky130_fd_sc_hd__mux2_1
XFILLER_102_666 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7018_ _7079_/CLK _7018_/D fanout514/X VGND VGND VPWR VPWR _7018_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_28_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_188_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_141_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_178_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_137_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_152_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_555 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_452 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_400 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_179_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_650 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_132 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_154 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_187_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4650_ _4799_/B _4985_/B VGND VGND VPWR VPWR _4665_/C sky130_fd_sc_hd__or2_1
Xinput10 mask_rev_in[15] VGND VGND VPWR VPWR input10/X sky130_fd_sc_hd__dlymetal6s2s_1
X_3601_ _6478_/Q _4032_/A _6352_/A _7154_/Q VGND VGND VPWR VPWR _3601_/X sky130_fd_sc_hd__a22o_1
XFILLER_147_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput21 mask_rev_in[25] VGND VGND VPWR VPWR input21/X sky130_fd_sc_hd__clkbuf_2
Xinput32 mask_rev_in[6] VGND VGND VPWR VPWR input32/X sky130_fd_sc_hd__dlymetal6s2s_1
X_4581_ _4581_/A _4640_/B VGND VGND VPWR VPWR _4581_/X sky130_fd_sc_hd__or2_1
Xinput43 mgmt_gpio_in[16] VGND VGND VPWR VPWR input43/X sky130_fd_sc_hd__clkbuf_4
XFILLER_174_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput54 mgmt_gpio_in[26] VGND VGND VPWR VPWR input54/X sky130_fd_sc_hd__clkbuf_2
X_6320_ _6320_/A _6320_/B VGND VGND VPWR VPWR _6320_/Y sky130_fd_sc_hd__nand2_1
Xhold805 _6687_/Q VGND VGND VPWR VPWR hold805/X sky130_fd_sc_hd__dlygate4sd3_1
X_3532_ _6822_/Q _5244_/A _4133_/A _6554_/Q VGND VGND VPWR VPWR _3532_/X sky130_fd_sc_hd__a22o_1
Xinput65 mgmt_gpio_in[36] VGND VGND VPWR VPWR _7199_/A sky130_fd_sc_hd__buf_4
Xinput76 qspi_enabled VGND VGND VPWR VPWR _3915_/S sky130_fd_sc_hd__clkbuf_8
Xhold816 _4148_/X VGND VGND VPWR VPWR _6562_/D sky130_fd_sc_hd__dlygate4sd3_1
Xinput87 spimemio_flash_io1_do VGND VGND VPWR VPWR _7198_/A sky130_fd_sc_hd__clkbuf_4
Xhold827 _6601_/Q VGND VGND VPWR VPWR hold827/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_155_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput98 usr2_vdd_pwrgood VGND VGND VPWR VPWR input98/X sky130_fd_sc_hd__buf_2
Xhold838 _4300_/X VGND VGND VPWR VPWR _6697_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6251_ _6251_/A _6251_/B _6251_/C _6250_/Y VGND VGND VPWR VPWR _6252_/C sky130_fd_sc_hd__or4b_4
Xhold849 _6684_/Q VGND VGND VPWR VPWR hold849/X sky130_fd_sc_hd__dlygate4sd3_1
X_3463_ _6927_/Q _5361_/A _5451_/A _7007_/Q _3462_/X VGND VGND VPWR VPWR _3470_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_115_257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5202_ hold369/X _5541_/A1 _5207_/S VGND VGND VPWR VPWR _5202_/X sky130_fd_sc_hd__mux2_1
XFILLER_143_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6182_ _6645_/Q _5950_/X _5952_/Y _7151_/Q _6181_/X VGND VGND VPWR VPWR _6182_/X
+ sky130_fd_sc_hd__a221o_1
X_3394_ _6961_/Q _5397_/A _5253_/A _6833_/Q _3393_/X VGND VGND VPWR VPWR _3395_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_97_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5133_ _4495_/X _5026_/B _5038_/A _5132_/X VGND VGND VPWR VPWR _5133_/X sky130_fd_sc_hd__o211a_1
XFILLER_97_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1505 _7167_/Q VGND VGND VPWR VPWR _3242_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1516 _7127_/Q VGND VGND VPWR VPWR _6205_/A1 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1527 _7116_/Q VGND VGND VPWR VPWR _5889_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_97_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1538 _6536_/Q VGND VGND VPWR VPWR hold379/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_111_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5064_ _5064_/A _5064_/B _5064_/C VGND VGND VPWR VPWR _5065_/C sky130_fd_sc_hd__and3_1
Xhold1549 _6532_/Q VGND VGND VPWR VPWR hold1549/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_38_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4015_ _4015_/A0 _5488_/A1 _4019_/S VGND VGND VPWR VPWR _4015_/X sky130_fd_sc_hd__mux2_1
XFILLER_38_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_263 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5966_ _5968_/A _5977_/A _5981_/C VGND VGND VPWR VPWR _5975_/C sky130_fd_sc_hd__and3_4
XFILLER_80_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4917_ _4495_/X _5026_/A _4861_/B _4394_/Y _4805_/X VGND VGND VPWR VPWR _4940_/B
+ sky130_fd_sc_hd__o221a_1
X_5897_ _6478_/Q _5620_/X _5892_/X _5895_/X _5896_/X VGND VGND VPWR VPWR _5897_/X
+ sky130_fd_sc_hd__a2111o_1
XFILLER_32_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4848_ _4563_/B _4566_/B _4947_/C VGND VGND VPWR VPWR _4848_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_165_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_165_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4779_ _4779_/A _4784_/A VGND VGND VPWR VPWR _4935_/B sky130_fd_sc_hd__nand2_1
XFILLER_181_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6518_ _6769_/CLK _6518_/D _6399_/A VGND VGND VPWR VPWR _6518_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_146_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_596 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6449_ _7032_/CLK _6449_/D fanout506/X VGND VGND VPWR VPWR _6449_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_134_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_40_csclk clkbuf_3_6_0_csclk/X VGND VGND VPWR VPWR _7069_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_164_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_2_0_0_csclk clkbuf_2_1_0_csclk/A VGND VGND VPWR VPWR clkbuf_3_1_0_csclk/A
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_130_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_506 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_189_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_263 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_211 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_169_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_172_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_174 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_678 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5820_ _6449_/Q _5917_/B1 _5817_/X _5818_/X _5819_/X VGND VGND VPWR VPWR _5820_/X
+ sky130_fd_sc_hd__a2111o_1
XFILLER_50_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5751_ _7014_/Q _5921_/A2 _5927_/A2 _6822_/Q _5750_/X VGND VGND VPWR VPWR _5754_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_15_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_148_614 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4702_ _4686_/B _4681_/X _4686_/X _4631_/A VGND VGND VPWR VPWR _4706_/B sky130_fd_sc_hd__a22oi_1
X_5682_ _6443_/Q _5645_/X _5680_/X _5681_/X VGND VGND VPWR VPWR _5682_/X sky130_fd_sc_hd__a211o_1
XFILLER_147_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_187_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4633_ input99/X _4542_/C _4779_/A VGND VGND VPWR VPWR _4634_/B sky130_fd_sc_hd__a21oi_1
XFILLER_175_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4564_ _4564_/A _4564_/B _4632_/A VGND VGND VPWR VPWR _4947_/C sky130_fd_sc_hd__and3_1
Xhold602 _6478_/Q VGND VGND VPWR VPWR hold602/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_118_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold613 _5395_/X VGND VGND VPWR VPWR _6952_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_162_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold624 _6668_/Q VGND VGND VPWR VPWR hold624/X sky130_fd_sc_hd__dlygate4sd3_1
X_6303_ _6544_/Q _6004_/B _6293_/X _6302_/X _5610_/A VGND VGND VPWR VPWR _6303_/X
+ sky130_fd_sc_hd__o221a_4
X_3515_ _3557_/A hold52/X VGND VGND VPWR VPWR _4279_/A sky130_fd_sc_hd__nor2_8
Xhold635 _5269_/X VGND VGND VPWR VPWR _6840_/D sky130_fd_sc_hd__dlygate4sd3_1
Xmax_cap354 _3533_/A VGND VGND VPWR VPWR _3523_/A sky130_fd_sc_hd__buf_12
Xhold646 _6568_/Q VGND VGND VPWR VPWR hold646/X sky130_fd_sc_hd__dlygate4sd3_1
X_4495_ _4495_/A _4495_/B VGND VGND VPWR VPWR _4495_/X sky130_fd_sc_hd__or2_4
Xmax_cap365 _5976_/Y VGND VGND VPWR VPWR _6285_/B1 sky130_fd_sc_hd__buf_8
Xhold657 _5528_/X VGND VGND VPWR VPWR _7070_/D sky130_fd_sc_hd__dlygate4sd3_1
Xmax_cap376 _5979_/X VGND VGND VPWR VPWR _6282_/B1 sky130_fd_sc_hd__buf_12
XFILLER_104_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_171_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold668 _5349_/X VGND VGND VPWR VPWR _6911_/D sky130_fd_sc_hd__dlygate4sd3_1
Xmax_cap387 _5973_/C VGND VGND VPWR VPWR _6300_/B1 sky130_fd_sc_hd__buf_8
Xhold679 _7078_/Q VGND VGND VPWR VPWR hold679/X sky130_fd_sc_hd__dlygate4sd3_1
X_6234_ _6562_/Q _5969_/A _6289_/A2 _6672_/Q _6233_/X VGND VGND VPWR VPWR _6234_/X
+ sky130_fd_sc_hd__a221o_1
Xmax_cap398 _5650_/X VGND VGND VPWR VPWR _5919_/B1 sky130_fd_sc_hd__buf_8
X_3446_ _6855_/Q _3374_/Y _5253_/A _6831_/Q VGND VGND VPWR VPWR _3446_/X sky130_fd_sc_hd__a22o_1
XFILLER_143_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6165_ _6841_/Q _5946_/X _5971_/A _6873_/Q VGND VGND VPWR VPWR _6165_/X sky130_fd_sc_hd__a22o_1
XTAP_951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3377_ _3553_/A hold40/X VGND VGND VPWR VPWR hold41/A sky130_fd_sc_hd__nor2_8
XFILLER_134_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1302 _5249_/X VGND VGND VPWR VPWR _6822_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1313 hold1398/X VGND VGND VPWR VPWR hold1313/X sky130_fd_sc_hd__dlygate4sd3_1
X_5116_ _5116_/A _5116_/B _5116_/C VGND VGND VPWR VPWR _5138_/B sky130_fd_sc_hd__and3_1
XTAP_984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1324 hold1324/A VGND VGND VPWR VPWR wb_dat_o[9] sky130_fd_sc_hd__buf_12
X_6096_ _6814_/Q _5936_/X _5942_/X _6942_/Q VGND VGND VPWR VPWR _6096_/X sky130_fd_sc_hd__a22o_1
Xhold1335 _4158_/A1 VGND VGND VPWR VPWR hold1335/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_57_347 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1346 hold1346/A VGND VGND VPWR VPWR wb_dat_o[26] sky130_fd_sc_hd__buf_12
XFILLER_27_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1357 _4162_/A1 VGND VGND VPWR VPWR hold1357/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1368 hold1368/A VGND VGND VPWR VPWR wb_dat_o[28] sky130_fd_sc_hd__buf_12
X_5047_ _4789_/B _5043_/B _4862_/X _5046_/X VGND VGND VPWR VPWR _5047_/X sky130_fd_sc_hd__o211a_1
XFILLER_26_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1379 _7020_/Q VGND VGND VPWR VPWR _5472_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_572 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6998_ _6998_/CLK _6998_/D fanout513/X VGND VGND VPWR VPWR _6998_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_41_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5949_ _5968_/A _5979_/B _5981_/C VGND VGND VPWR VPWR _5949_/X sky130_fd_sc_hd__and3_4
XFILLER_43_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_159_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_178_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_104_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_347 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_734 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_185_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_172_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_160_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_715 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3300_ hold75/A VGND VGND VPWR VPWR _3300_/Y sky130_fd_sc_hd__inv_2
XFILLER_98_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4280_ _4280_/A0 _5488_/A1 _4284_/S VGND VGND VPWR VPWR _4280_/X sky130_fd_sc_hd__mux2_1
XFILLER_140_322 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3231_ _3247_/A _7170_/Q _3231_/S VGND VGND VPWR VPWR _7170_/D sky130_fd_sc_hd__mux2_1
XFILLER_101_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_580 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6921_ _7054_/CLK _6921_/D fanout503/X VGND VGND VPWR VPWR _6921_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_47_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6852_ _7041_/CLK _6852_/D fanout520/X VGND VGND VPWR VPWR _6852_/Q sky130_fd_sc_hd__dfrtp_2
X_5803_ _7025_/Q _5929_/B1 _5915_/B1 _6865_/Q VGND VGND VPWR VPWR _5803_/X sky130_fd_sc_hd__a22o_1
XFILLER_22_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6783_ _7083_/CLK _6783_/D fanout517/X VGND VGND VPWR VPWR _6783_/Q sky130_fd_sc_hd__dfrtp_1
X_3995_ hold979/X _5495_/A1 _4001_/S VGND VGND VPWR VPWR _3995_/X sky130_fd_sc_hd__mux2_1
X_5734_ _7108_/Q _5612_/A _5612_/B VGND VGND VPWR VPWR _5734_/X sky130_fd_sc_hd__o21a_1
XFILLER_50_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_176_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5665_ _6882_/Q _5913_/B1 _5663_/X _5664_/X VGND VGND VPWR VPWR _5665_/X sky130_fd_sc_hd__a211o_1
XFILLER_176_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_148_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_148_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4616_ _5005_/A _4615_/B _4594_/X VGND VGND VPWR VPWR _4616_/X sky130_fd_sc_hd__a21o_1
X_5596_ _5940_/B _5596_/B VGND VGND VPWR VPWR _5598_/A sky130_fd_sc_hd__or2_1
XFILLER_163_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold410 _4264_/X VGND VGND VPWR VPWR _6667_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_135_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_191_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4547_ _4640_/B _4988_/A VGND VGND VPWR VPWR _4547_/X sky130_fd_sc_hd__and2_2
Xhold421 _6904_/Q VGND VGND VPWR VPWR hold421/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold432 _4132_/X VGND VGND VPWR VPWR _6549_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_352 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold443 _6921_/Q VGND VGND VPWR VPWR hold443/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold454 _5427_/X VGND VGND VPWR VPWR _6980_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_1_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold465 _7000_/Q VGND VGND VPWR VPWR hold465/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_145_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold476 _4266_/X VGND VGND VPWR VPWR _6669_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4478_ _4587_/A _4943_/A VGND VGND VPWR VPWR _4506_/B sky130_fd_sc_hd__or2_1
Xhold487 _6791_/Q VGND VGND VPWR VPWR hold487/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold498 _5149_/X VGND VGND VPWR VPWR _6740_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6217_ _6217_/A _6217_/B VGND VGND VPWR VPWR _6217_/Y sky130_fd_sc_hd__nor2_1
XFILLER_104_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3429_ _6888_/Q hold83/A _5298_/A _6872_/Q _3428_/X VGND VGND VPWR VPWR _3431_/A
+ sky130_fd_sc_hd__a221o_1
X_7197_ _7197_/A VGND VGND VPWR VPWR _7197_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_57_100 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6148_ _7000_/Q _6282_/A2 _5955_/X _6968_/Q VGND VGND VPWR VPWR _6148_/X sky130_fd_sc_hd__a22o_1
XTAP_781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1110 _4191_/X VGND VGND VPWR VPWR _6599_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1121 _6665_/Q VGND VGND VPWR VPWR _4262_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1132 _5375_/X VGND VGND VPWR VPWR _6934_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1143 _6715_/Q VGND VGND VPWR VPWR _4322_/A0 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1154 _5380_/X VGND VGND VPWR VPWR _6938_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6079_ _6507_/Q _6079_/A2 _5611_/X VGND VGND VPWR VPWR _6079_/X sky130_fd_sc_hd__a21o_1
XFILLER_57_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1165 _7071_/Q VGND VGND VPWR VPWR _5530_/A0 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1176 _4304_/X VGND VGND VPWR VPWR _6700_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_72_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1187 _6854_/Q VGND VGND VPWR VPWR _5285_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_57_199 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1198 _4113_/X VGND VGND VPWR VPWR _6532_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_26_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_158_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_182_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_186_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_467 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3780_ _6818_/Q _5244_/A _4145_/A _6560_/Q _3779_/X VGND VGND VPWR VPWR _3780_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_158_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_185_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5450_ hold219/X hold27/X _5450_/S VGND VGND VPWR VPWR _5450_/X sky130_fd_sc_hd__mux2_1
XFILLER_67_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_145_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4401_ _4885_/A _4401_/B VGND VGND VPWR VPWR _4401_/X sky130_fd_sc_hd__or2_1
X_5381_ hold988/X _5495_/A1 _5387_/S VGND VGND VPWR VPWR _5381_/X sky130_fd_sc_hd__mux2_1
XFILLER_160_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_3_2_0_wb_clk_i clkbuf_3_3_0_wb_clk_i/A VGND VGND VPWR VPWR _7124_/CLK sky130_fd_sc_hd__clkbuf_8
X_7120_ _7123_/CLK _7120_/D fanout499/X VGND VGND VPWR VPWR _7120_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_5_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4332_ _4575_/A _4746_/B VGND VGND VPWR VPWR _4884_/A sky130_fd_sc_hd__nor2_2
XFILLER_141_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7051_ _7051_/CLK _7051_/D fanout514/X VGND VGND VPWR VPWR _7051_/Q sky130_fd_sc_hd__dfrtp_1
X_4263_ hold875/X _5189_/A1 _4266_/S VGND VGND VPWR VPWR _4263_/X sky130_fd_sc_hd__mux2_1
XFILLER_87_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6002_ _6002_/A _6002_/B _6002_/C _6001_/Y VGND VGND VPWR VPWR _6003_/C sky130_fd_sc_hd__or4b_1
XFILLER_141_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3214_ _6845_/Q VGND VGND VPWR VPWR _3214_/Y sky130_fd_sc_hd__inv_2
X_4194_ hold261/X hold46/X _4195_/S VGND VGND VPWR VPWR _4194_/X sky130_fd_sc_hd__mux2_1
XFILLER_67_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_131_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6904_ _6999_/CLK _6904_/D fanout523/X VGND VGND VPWR VPWR _6904_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_82_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6835_ _7072_/CLK _6835_/D fanout504/X VGND VGND VPWR VPWR _6835_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_11_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6766_ _6948_/CLK _6766_/D fanout514/X VGND VGND VPWR VPWR _6766_/Q sky130_fd_sc_hd__dfrtp_2
X_3978_ hold807/X _6355_/A1 _3983_/S VGND VGND VPWR VPWR _3978_/X sky130_fd_sc_hd__mux2_1
X_5717_ _6797_/Q _5651_/X _5715_/X _5716_/X VGND VGND VPWR VPWR _5717_/X sky130_fd_sc_hd__a211o_1
XFILLER_149_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6697_ _6697_/CLK _6697_/D fanout486/X VGND VGND VPWR VPWR _6697_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_109_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_2_1__f_mgmt_gpio_in[4] clkbuf_0_mgmt_gpio_in[4]/X VGND VGND VPWR VPWR _3939_/A1
+ sky130_fd_sc_hd__clkbuf_16
X_5648_ _5667_/A _5649_/C _5648_/C VGND VGND VPWR VPWR _5648_/X sky130_fd_sc_hd__and3_4
XFILLER_136_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_296 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_447 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5579_ _5667_/A _5579_/B VGND VGND VPWR VPWR _5579_/Y sky130_fd_sc_hd__nand2_1
XFILLER_117_683 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold240 _5212_/X VGND VGND VPWR VPWR _6789_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold251 _6761_/Q VGND VGND VPWR VPWR hold251/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold262 _4194_/X VGND VGND VPWR VPWR _6602_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold273 _6928_/Q VGND VGND VPWR VPWR hold273/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold284 _5418_/X VGND VGND VPWR VPWR _6972_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold295 hold295/A VGND VGND VPWR VPWR hold295/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_49_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_626 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_102 _3943_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_113 _3951_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_124 _3894_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_135 _6294_/B1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_146 _5534_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_121_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_157 _6396_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_168 hold142/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_179 _5632_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_127_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_170_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_642 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput8 mask_rev_in[13] VGND VGND VPWR VPWR input8/X sky130_fd_sc_hd__clkbuf_1
XFILLER_64_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4950_ _4574_/A _4949_/X _4574_/B VGND VGND VPWR VPWR _4950_/X sky130_fd_sc_hd__a21o_1
X_3901_ _4449_/A _4449_/B _3901_/C _3901_/D VGND VGND VPWR VPWR _3908_/B sky130_fd_sc_hd__and4_1
X_4881_ _5040_/B _4881_/B _4881_/C _4881_/D VGND VGND VPWR VPWR _4881_/X sky130_fd_sc_hd__and4_1
XFILLER_189_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6620_ _6630_/CLK _6620_/D fanout495/X VGND VGND VPWR VPWR _6620_/Q sky130_fd_sc_hd__dfrtp_1
X_3832_ hold48/A _3847_/B VGND VGND VPWR VPWR _3845_/S sky130_fd_sc_hd__and2_1
X_6551_ _6769_/CLK _6551_/D fanout492/X VGND VGND VPWR VPWR _6551_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_158_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3763_ _6866_/Q _5298_/A _5190_/A input52/X _3762_/X VGND VGND VPWR VPWR _3778_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_146_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5502_ _5502_/A _5538_/B VGND VGND VPWR VPWR _5510_/S sky130_fd_sc_hd__and2_4
XFILLER_146_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_192_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6482_ _6632_/CLK _6482_/D fanout509/X VGND VGND VPWR VPWR _6482_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_145_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3694_ _6443_/Q _3361_/Y _4249_/A _6656_/Q _3693_/X VGND VGND VPWR VPWR _3697_/A
+ sky130_fd_sc_hd__a221o_1
X_5433_ hold34/X _5538_/B VGND VGND VPWR VPWR hold35/A sky130_fd_sc_hd__and2_4
Xoutput301 _3803_/X VGND VGND VPWR VPWR reset sky130_fd_sc_hd__buf_12
XFILLER_133_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput312 _7200_/X VGND VGND VPWR VPWR spimemio_flash_io3_di sky130_fd_sc_hd__buf_12
Xoutput323 hold1305/X VGND VGND VPWR VPWR hold1306/A sky130_fd_sc_hd__buf_12
X_5364_ hold361/X _5532_/A1 _5369_/S VGND VGND VPWR VPWR _5364_/X sky130_fd_sc_hd__mux2_1
Xoutput334 hold1367/X VGND VGND VPWR VPWR hold1368/A sky130_fd_sc_hd__buf_12
Xoutput345 hold1323/X VGND VGND VPWR VPWR hold1324/A sky130_fd_sc_hd__buf_12
XFILLER_126_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7103_ _7131_/CLK _7103_/D fanout501/X VGND VGND VPWR VPWR _7103_/Q sky130_fd_sc_hd__dfrtp_1
X_4315_ _4315_/A _6352_/B VGND VGND VPWR VPWR _4320_/S sky130_fd_sc_hd__and2_2
XFILLER_141_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5295_ hold747/X _5457_/A1 _5297_/S VGND VGND VPWR VPWR _5295_/X sky130_fd_sc_hd__mux2_1
XFILLER_59_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7034_ _7034_/CLK _7034_/D fanout488/X VGND VGND VPWR VPWR _7034_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_87_548 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4246_ hold618/X _5505_/A1 hold63/X VGND VGND VPWR VPWR _4246_/X sky130_fd_sc_hd__mux2_1
XFILLER_19_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4177_ _4186_/A0 _4177_/A1 _4180_/S VGND VGND VPWR VPWR _6587_/D sky130_fd_sc_hd__mux2_1
XFILLER_83_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_434 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6818_ _7041_/CLK _6818_/D fanout518/X VGND VGND VPWR VPWR _6818_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_149_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6749_ _7010_/CLK _6749_/D fanout498/X VGND VGND VPWR VPWR _6749_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_149_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_191_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_504 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_623 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_92_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_415 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_187_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_174_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_380 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_542 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_115_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4100_ hold501/X _5491_/A1 hold8/X VGND VGND VPWR VPWR _4100_/X sky130_fd_sc_hd__mux2_1
XFILLER_110_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5080_ _4862_/A _5026_/A _4965_/C _4789_/B VGND VGND VPWR VPWR _5081_/D sky130_fd_sc_hd__o22a_1
XFILLER_111_656 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4031_ hold573/X _6357_/A1 _4031_/S VGND VGND VPWR VPWR _4031_/X sky130_fd_sc_hd__mux2_1
XFILLER_2_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5982_ _6946_/Q _5978_/X _6270_/B1 _6930_/Q VGND VGND VPWR VPWR _5982_/X sky130_fd_sc_hd__a22o_1
XFILLER_18_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4933_ _4933_/A _4933_/B _4933_/C VGND VGND VPWR VPWR _5070_/A sky130_fd_sc_hd__and3_1
XFILLER_33_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4864_ _4748_/B _4719_/B _4972_/A _4901_/B VGND VGND VPWR VPWR _4868_/A sky130_fd_sc_hd__o22a_1
XFILLER_178_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_13 _5451_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_509 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3815_ _3782_/X _3815_/B _3815_/C _3815_/D VGND VGND VPWR VPWR _3815_/X sky130_fd_sc_hd__and4b_1
XANTENNA_24 _3433_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6603_ _6632_/CLK _6603_/D _3264_/A VGND VGND VPWR VPWR _6603_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_177_155 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_35 hold62/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_165_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_46 _3755_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4795_ _4456_/Y _5021_/B _4788_/A VGND VGND VPWR VPWR _4795_/X sky130_fd_sc_hd__a21o_1
XANTENNA_57 _5844_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6534_ _7054_/CLK _6534_/D fanout503/X VGND VGND VPWR VPWR _6534_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA_68 _6482_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_146_520 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3746_ _3716_/X _3746_/B _3746_/C _3746_/D VGND VGND VPWR VPWR _3747_/B sky130_fd_sc_hd__and4b_1
XFILLER_118_222 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_79 user_clock VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_146_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_180_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6465_ _6707_/CLK _6465_/D fanout484/X VGND VGND VPWR VPWR _6465_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_134_715 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3677_ _6444_/Q _3993_/A _4020_/A _6467_/Q VGND VGND VPWR VPWR _3677_/X sky130_fd_sc_hd__a22o_1
XFILLER_146_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5416_ _5416_/A0 _5488_/A1 _5423_/S VGND VGND VPWR VPWR _5416_/X sky130_fd_sc_hd__mux2_1
XFILLER_133_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6396_ _6396_/A _6396_/B VGND VGND VPWR VPWR _6396_/X sky130_fd_sc_hd__and2_1
XFILLER_114_450 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5347_ hold351/X _5515_/A1 _5351_/S VGND VGND VPWR VPWR _5347_/X sky130_fd_sc_hd__mux2_1
Xoutput175 _3929_/X VGND VGND VPWR VPWR mgmt_gpio_oeb[0] sky130_fd_sc_hd__buf_12
Xoutput186 _3928_/X VGND VGND VPWR VPWR mgmt_gpio_oeb[1] sky130_fd_sc_hd__buf_12
Xoutput197 _3218_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[2] sky130_fd_sc_hd__buf_12
XFILLER_87_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5278_ hold461/X _5545_/A1 _5279_/S VGND VGND VPWR VPWR _5278_/X sky130_fd_sc_hd__mux2_1
XFILLER_75_518 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7017_ _7017_/CLK _7017_/D fanout515/X VGND VGND VPWR VPWR _7017_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_102_678 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4229_ hold553/X _5491_/A1 _4230_/S VGND VGND VPWR VPWR _4229_/X sky130_fd_sc_hd__mux2_1
XFILLER_56_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_111 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_183_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_149_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_152_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_152_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_464 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_412 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_231 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_275 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_147_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_159_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3600_ _7042_/Q _5493_/A _5179_/B _6758_/Q _3599_/X VGND VGND VPWR VPWR _3605_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_159_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput11 mask_rev_in[16] VGND VGND VPWR VPWR input11/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_30_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput22 mask_rev_in[26] VGND VGND VPWR VPWR input22/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_128_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4580_ _4537_/X _4540_/Y _4548_/X _4559_/X _4579_/X VGND VGND VPWR VPWR _4580_/X
+ sky130_fd_sc_hd__o2111a_1
Xinput33 mask_rev_in[7] VGND VGND VPWR VPWR input33/X sky130_fd_sc_hd__clkbuf_1
XFILLER_162_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput44 mgmt_gpio_in[17] VGND VGND VPWR VPWR input44/X sky130_fd_sc_hd__clkbuf_4
X_3531_ _3531_/A _3628_/B VGND VGND VPWR VPWR _4133_/A sky130_fd_sc_hd__nor2_4
Xinput55 mgmt_gpio_in[27] VGND VGND VPWR VPWR input55/X sky130_fd_sc_hd__buf_2
XFILLER_155_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput66 mgmt_gpio_in[37] VGND VGND VPWR VPWR _7200_/A sky130_fd_sc_hd__buf_4
Xinput77 ser_tx VGND VGND VPWR VPWR input77/X sky130_fd_sc_hd__clkbuf_1
Xhold806 _4288_/X VGND VGND VPWR VPWR _6687_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold817 _6420_/Q VGND VGND VPWR VPWR hold817/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold828 _4193_/X VGND VGND VPWR VPWR _6601_/D sky130_fd_sc_hd__dlygate4sd3_1
Xinput88 spimemio_flash_io1_oeb VGND VGND VPWR VPWR _3943_/B sky130_fd_sc_hd__clkbuf_4
X_6250_ _6250_/A _6250_/B VGND VGND VPWR VPWR _6250_/Y sky130_fd_sc_hd__nor2_1
XFILLER_115_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold839 _7004_/Q VGND VGND VPWR VPWR hold839/X sky130_fd_sc_hd__dlygate4sd3_1
Xinput99 wb_adr_i[0] VGND VGND VPWR VPWR input99/X sky130_fd_sc_hd__clkbuf_4
X_3462_ _6919_/Q _5352_/A _5179_/B _3439_/X VGND VGND VPWR VPWR _3462_/X sky130_fd_sc_hd__a22o_2
X_5201_ hold207/X hold90/X _5207_/S VGND VGND VPWR VPWR _5201_/X sky130_fd_sc_hd__mux2_1
XFILLER_115_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6181_ _6655_/Q _6288_/A2 _5977_/X _6665_/Q VGND VGND VPWR VPWR _6181_/X sky130_fd_sc_hd__a22o_1
X_3393_ _7070_/Q _5520_/A _5511_/A _7062_/Q VGND VGND VPWR VPWR _3393_/X sky130_fd_sc_hd__a22o_1
XFILLER_130_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5132_ _4911_/A _5132_/B _5132_/C VGND VGND VPWR VPWR _5132_/X sky130_fd_sc_hd__and3b_1
Xhold1506 _7132_/Q VGND VGND VPWR VPWR hold1506/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_29_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1517 _6506_/Q VGND VGND VPWR VPWR _3172_/A sky130_fd_sc_hd__dlygate4sd3_1
X_5063_ _4515_/B _4988_/A _4748_/B _4972_/A VGND VGND VPWR VPWR _5065_/B sky130_fd_sc_hd__o22a_1
Xhold1528 _7094_/Q VGND VGND VPWR VPWR _5575_/A1 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1539 _7089_/Q VGND VGND VPWR VPWR _5557_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_96_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4014_ _4014_/A _6352_/B VGND VGND VPWR VPWR _4019_/S sky130_fd_sc_hd__and2_4
XFILLER_38_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5965_ _5980_/A _5965_/B VGND VGND VPWR VPWR _5971_/B sky130_fd_sc_hd__nor2_8
X_4916_ _4515_/B _5026_/A _4962_/C _4972_/A _4818_/B VGND VGND VPWR VPWR _4991_/A
+ sky130_fd_sc_hd__o221ai_1
X_5896_ _6698_/Q _5626_/X _5647_/X _6458_/Q VGND VGND VPWR VPWR _5896_/X sky130_fd_sc_hd__a22o_1
XFILLER_32_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_178_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4847_ _4581_/A _4831_/X _4845_/X _4846_/X VGND VGND VPWR VPWR _4847_/X sky130_fd_sc_hd__o211a_1
XFILLER_138_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4778_ _4799_/A _4778_/B _4778_/C VGND VGND VPWR VPWR _4935_/A sky130_fd_sc_hd__nand3_1
XFILLER_165_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3729_ _7027_/Q _5478_/A _4020_/A _6466_/Q VGND VGND VPWR VPWR _3729_/X sky130_fd_sc_hd__a22o_1
X_6517_ _7022_/CLK _6517_/D fanout517/X VGND VGND VPWR VPWR _6517_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_174_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6448_ _7050_/CLK _6448_/D fanout515/X VGND VGND VPWR VPWR _6448_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_134_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_164_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6379_ _6400_/A _6399_/B VGND VGND VPWR VPWR _6379_/X sky130_fd_sc_hd__and2_1
XFILLER_121_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_169_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_386 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_654 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_94_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5750_ _6926_/Q _5633_/X _5646_/X _6998_/Q VGND VGND VPWR VPWR _5750_/X sky130_fd_sc_hd__a22o_1
XFILLER_97_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4701_ _4701_/A _5005_/B VGND VGND VPWR VPWR _4711_/A sky130_fd_sc_hd__nor2_1
X_5681_ _6811_/Q _5627_/X _5636_/X _6819_/Q VGND VGND VPWR VPWR _5681_/X sky130_fd_sc_hd__a22o_1
XFILLER_148_626 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4632_ _4632_/A _4632_/B VGND VGND VPWR VPWR _4799_/B sky130_fd_sc_hd__nand2_1
XFILLER_8_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_175_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_163_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4563_ _4574_/A _4563_/B VGND VGND VPWR VPWR _5088_/B sky130_fd_sc_hd__nand2_1
XFILLER_156_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold603 _4036_/X VGND VGND VPWR VPWR _6478_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_190_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold614 _7174_/A VGND VGND VPWR VPWR hold614/X sky130_fd_sc_hd__dlygate4sd3_1
X_6302_ _6302_/A _6302_/B _6302_/C _6004_/B VGND VGND VPWR VPWR _6302_/X sky130_fd_sc_hd__or4b_1
X_3514_ _7083_/Q _5538_/A _5502_/A _7051_/Q VGND VGND VPWR VPWR _3514_/X sky130_fd_sc_hd__a22o_1
Xhold625 _4265_/X VGND VGND VPWR VPWR _6668_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_155_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold636 _6448_/Q VGND VGND VPWR VPWR hold636/X sky130_fd_sc_hd__dlygate4sd3_1
X_4494_ _4549_/B _4586_/B VGND VGND VPWR VPWR _4911_/A sky130_fd_sc_hd__nor2_1
Xhold647 _4155_/X VGND VGND VPWR VPWR _6568_/D sky130_fd_sc_hd__dlygate4sd3_1
Xmax_cap355 _3533_/A VGND VGND VPWR VPWR _3531_/A sky130_fd_sc_hd__buf_12
Xmax_cap366 _5947_/Y VGND VGND VPWR VPWR _6291_/A2 sky130_fd_sc_hd__buf_12
Xhold658 _6809_/Q VGND VGND VPWR VPWR hold658/X sky130_fd_sc_hd__dlygate4sd3_1
X_6233_ _6662_/Q _6294_/A2 _6294_/B1 _6712_/Q VGND VGND VPWR VPWR _6233_/X sky130_fd_sc_hd__a22o_1
XFILLER_171_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmax_cap377 _5969_/C VGND VGND VPWR VPWR _6294_/B1 sky130_fd_sc_hd__buf_12
XFILLER_116_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3445_ _6895_/Q _5325_/A _5244_/A _6823_/Q _3442_/X VGND VGND VPWR VPWR _3471_/A
+ sky130_fd_sc_hd__a221o_1
Xhold669 _6871_/Q VGND VGND VPWR VPWR hold669/X sky130_fd_sc_hd__dlygate4sd3_1
Xmax_cap388 _5963_/X VGND VGND VPWR VPWR _5974_/B sky130_fd_sc_hd__buf_12
Xmax_cap399 _5649_/X VGND VGND VPWR VPWR _5807_/B1 sky130_fd_sc_hd__buf_12
XTAP_930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6164_ _6969_/Q _5955_/X _6294_/B1 _7046_/Q _6163_/X VGND VGND VPWR VPWR _6167_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_131_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3376_ _6857_/Q _3374_/Y _4077_/S _3953_/B _3373_/X VGND VGND VPWR VPWR _3395_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_134_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5115_ _4551_/B _4615_/X _4631_/X _4973_/B VGND VGND VPWR VPWR _5116_/C sky130_fd_sc_hd__o22a_1
XTAP_974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1303 _6910_/Q VGND VGND VPWR VPWR _5348_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1314 hold1314/A VGND VGND VPWR VPWR wb_dat_o[19] sky130_fd_sc_hd__buf_12
X_6095_ _7006_/Q _6290_/A2 wire390/X _6854_/Q _6094_/X VGND VGND VPWR VPWR _6102_/A
+ sky130_fd_sc_hd__a221o_1
XTAP_996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1325 _4175_/A1 VGND VGND VPWR VPWR hold1325/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_57_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1336 hold1336/A VGND VGND VPWR VPWR wb_dat_o[16] sky130_fd_sc_hd__buf_12
XFILLER_57_359 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1347 _6316_/A1 VGND VGND VPWR VPWR hold1347/X sky130_fd_sc_hd__dlygate4sd3_1
X_5046_ _4576_/X _4686_/B _4977_/B VGND VGND VPWR VPWR _5046_/X sky130_fd_sc_hd__a21o_1
XFILLER_27_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1358 hold1358/A VGND VGND VPWR VPWR wb_dat_o[20] sky130_fd_sc_hd__buf_12
Xhold1369 hold1506/X VGND VGND VPWR VPWR hold1369/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_84_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_234 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6997_ _7083_/CLK _6997_/D fanout518/X VGND VGND VPWR VPWR _6997_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_43_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5948_ _5977_/A _5963_/C _5981_/C VGND VGND VPWR VPWR _5948_/X sky130_fd_sc_hd__and3_4
XFILLER_139_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_178_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_626 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5879_ _6657_/Q _5923_/B VGND VGND VPWR VPWR _5879_/X sky130_fd_sc_hd__and2b_1
XFILLER_126_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_331 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_161_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_191_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_307 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_746 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_157_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_129_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_144_106 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_144_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_334 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3230_ _6417_/Q _6416_/Q _6415_/Q _6485_/Q VGND VGND VPWR VPWR _3231_/S sky130_fd_sc_hd__or4bb_1
XFILLER_113_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_592 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6920_ _7017_/CLK _6920_/D fanout515/X VGND VGND VPWR VPWR _6920_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_62_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6851_ _7056_/CLK _6851_/D fanout504/X VGND VGND VPWR VPWR _6851_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_90_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_671 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5802_ _3224_/Y _5646_/A _5667_/B VGND VGND VPWR VPWR _5802_/Y sky130_fd_sc_hd__a21oi_2
X_3994_ _3994_/A0 _5530_/A1 _4001_/S VGND VGND VPWR VPWR _3994_/X sky130_fd_sc_hd__mux2_1
X_6782_ _7069_/CLK _6782_/D fanout516/X VGND VGND VPWR VPWR _6782_/Q sky130_fd_sc_hd__dfrtp_1
X_5733_ _6789_/Q _5667_/X _5723_/X _5732_/X _3174_/Y VGND VGND VPWR VPWR _5733_/X
+ sky130_fd_sc_hd__o221a_2
XFILLER_31_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_175_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5664_ _6874_/Q _5914_/A2 _5919_/B1 _6890_/Q VGND VGND VPWR VPWR _5664_/X sky130_fd_sc_hd__a22o_1
XFILLER_148_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_163_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_54_csclk _7000_/CLK VGND VGND VPWR VPWR _7032_/CLK sky130_fd_sc_hd__clkbuf_16
X_4615_ _4631_/A _4615_/B VGND VGND VPWR VPWR _4615_/X sky130_fd_sc_hd__or2_2
X_5595_ _5595_/A1 _5571_/Y _5596_/B _5594_/X VGND VGND VPWR VPWR _7100_/D sky130_fd_sc_hd__a31o_1
XFILLER_135_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold400 _4282_/X VGND VGND VPWR VPWR _6682_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold411 _6948_/Q VGND VGND VPWR VPWR hold411/X sky130_fd_sc_hd__dlygate4sd3_1
X_4546_ _4721_/B _4649_/A _4788_/A _4921_/A _4581_/A VGND VGND VPWR VPWR _4546_/X
+ sky130_fd_sc_hd__o32a_1
Xhold422 _5341_/X VGND VGND VPWR VPWR _6904_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold433 _6932_/Q VGND VGND VPWR VPWR hold433/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold444 _5360_/X VGND VGND VPWR VPWR _6921_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold455 _7057_/Q VGND VGND VPWR VPWR hold455/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_190_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold466 _5449_/X VGND VGND VPWR VPWR _7000_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4477_ _4692_/A _4479_/A VGND VGND VPWR VPWR _4506_/A sky130_fd_sc_hd__or2_1
Xhold477 _6425_/Q VGND VGND VPWR VPWR hold477/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold488 _5214_/X VGND VGND VPWR VPWR _6791_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6216_ _6661_/Q _6294_/A2 _5975_/C _6701_/Q _6215_/X VGND VGND VPWR VPWR _6217_/B
+ sky130_fd_sc_hd__a221o_1
Xhold499 _6437_/Q VGND VGND VPWR VPWR hold499/X sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_69_csclk _7000_/CLK VGND VGND VPWR VPWR _7071_/CLK sky130_fd_sc_hd__clkbuf_16
X_3428_ input41/X _4092_/S _5271_/A _6848_/Q VGND VGND VPWR VPWR _3428_/X sky130_fd_sc_hd__a22o_1
X_7196_ _7196_/A VGND VGND VPWR VPWR _7196_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_38_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6147_ _6816_/Q _5936_/X _5947_/Y _7032_/Q _6146_/X VGND VGND VPWR VPWR _6152_/B
+ sky130_fd_sc_hd__a221o_1
X_3359_ _7054_/Q _5502_/A _5478_/A _7033_/Q VGND VGND VPWR VPWR _3359_/X sky130_fd_sc_hd__a22o_1
Xhold1100 _5169_/X VGND VGND VPWR VPWR _6755_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1111 _6625_/Q VGND VGND VPWR VPWR _4226_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1122 _4262_/X VGND VGND VPWR VPWR _6665_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1133 _7067_/Q VGND VGND VPWR VPWR _5525_/A0 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1144 _4322_/X VGND VGND VPWR VPWR _6715_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6078_ _6789_/Q _5975_/X _6068_/X _6077_/X _3174_/Y VGND VGND VPWR VPWR _6078_/X
+ sky130_fd_sc_hd__o221a_2
Xhold1155 _7039_/Q VGND VGND VPWR VPWR _5494_/A0 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1166 _5530_/X VGND VGND VPWR VPWR _7071_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1177 _7034_/Q VGND VGND VPWR VPWR _5488_/A0 sky130_fd_sc_hd__dlygate4sd3_1
X_5029_ _4515_/B _5026_/B _4581_/X _4774_/A _4833_/X VGND VGND VPWR VPWR _5038_/B
+ sky130_fd_sc_hd__o2111a_1
XTAP_2605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1188 _5285_/X VGND VGND VPWR VPWR _6854_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1199 _6914_/Q VGND VGND VPWR VPWR _5353_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_66_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_392 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_167_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_166_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_182_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_166_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_182_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_134_150 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_134_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_178 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_151_71 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_189_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4400_ _4737_/B _4892_/A VGND VGND VPWR VPWR _4401_/B sky130_fd_sc_hd__or2_1
XFILLER_173_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5380_ _5380_/A0 _5488_/A1 _5387_/S VGND VGND VPWR VPWR _5380_/X sky130_fd_sc_hd__mux2_1
X_4331_ _4679_/A _4542_/A VGND VGND VPWR VPWR _4746_/B sky130_fd_sc_hd__nand2b_1
XFILLER_99_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_323 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7050_ _7050_/CLK _7050_/D fanout516/X VGND VGND VPWR VPWR _7050_/Q sky130_fd_sc_hd__dfrtp_4
X_4262_ _4262_/A0 _6353_/A1 _4266_/S VGND VGND VPWR VPWR _4262_/X sky130_fd_sc_hd__mux2_1
XFILLER_141_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6001_ _6906_/Q _5972_/A _5949_/X _7063_/Q _6000_/X VGND VGND VPWR VPWR _6001_/Y
+ sky130_fd_sc_hd__a221oi_1
X_3213_ _6853_/Q VGND VGND VPWR VPWR _3213_/Y sky130_fd_sc_hd__inv_2
XFILLER_101_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4193_ hold827/X _5505_/A1 _4195_/S VGND VGND VPWR VPWR _4193_/X sky130_fd_sc_hd__mux2_1
XFILLER_79_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_435 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6903_ _6999_/CLK _6903_/D fanout523/X VGND VGND VPWR VPWR _6903_/Q sky130_fd_sc_hd__dfrtp_2
X_6834_ _7071_/CLK _6834_/D fanout504/X VGND VGND VPWR VPWR _6834_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_50_332 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6765_ _6965_/CLK _6765_/D fanout514/X VGND VGND VPWR VPWR _6765_/Q sky130_fd_sc_hd__dfrtp_4
X_3977_ hold990/X _6354_/A1 _3983_/S VGND VGND VPWR VPWR _3977_/X sky130_fd_sc_hd__mux2_1
X_5716_ _6845_/Q _5922_/B1 _5926_/A2 _6805_/Q VGND VGND VPWR VPWR _5716_/X sky130_fd_sc_hd__a22o_1
XFILLER_148_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6696_ _6696_/CLK _6696_/D fanout495/X VGND VGND VPWR VPWR _6696_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_148_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5647_ _5667_/A _5649_/C _5650_/B VGND VGND VPWR VPWR _5647_/X sky130_fd_sc_hd__and3_4
XFILLER_148_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_459 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_191_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5578_ _5578_/A1 _5571_/Y _5577_/B _5579_/B VGND VGND VPWR VPWR _7095_/D sky130_fd_sc_hd__a31o_1
XFILLER_151_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold230 _5167_/X VGND VGND VPWR VPWR _6754_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold241 _6912_/Q VGND VGND VPWR VPWR hold241/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold252 _5177_/X VGND VGND VPWR VPWR _6761_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_117_695 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4529_ _4481_/Y _4492_/Y _4527_/X _4755_/A _4883_/A VGND VGND VPWR VPWR _4529_/X
+ sky130_fd_sc_hd__o41a_1
XFILLER_6_8 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold263 _6683_/Q VGND VGND VPWR VPWR hold263/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold274 _5368_/X VGND VGND VPWR VPWR _6928_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold285 _6516_/Q VGND VGND VPWR VPWR hold285/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold296 _4089_/X VGND VGND VPWR VPWR _6514_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_172_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_172_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7179_ _7179_/A VGND VGND VPWR VPWR _7179_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_131_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_103 _3943_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_114 _3951_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_125 _3894_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_164_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_136 _6294_/B1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_147 _5534_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_158 _3931_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_169 hold588/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_146_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_8 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_164 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput9 mask_rev_in[14] VGND VGND VPWR VPWR input9/X sky130_fd_sc_hd__clkbuf_2
XFILLER_92_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3900_ _4335_/C _3900_/B _3900_/C _3900_/D VGND VGND VPWR VPWR _3901_/D sky130_fd_sc_hd__nor4_1
X_4880_ _5087_/B _4879_/X _4960_/B VGND VGND VPWR VPWR _4881_/D sky130_fd_sc_hd__a21bo_1
XFILLER_189_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3831_ hold37/A hold71/A hold78/A VGND VGND VPWR VPWR _3847_/B sky130_fd_sc_hd__and3_1
XFILLER_32_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6550_ _6769_/CLK _6550_/D _6399_/A VGND VGND VPWR VPWR _6550_/Q sky130_fd_sc_hd__dfrtp_4
X_3762_ _6786_/Q _5208_/A _5181_/A _6764_/Q VGND VGND VPWR VPWR _3762_/X sky130_fd_sc_hd__a22o_1
X_5501_ hold467/X _5519_/A1 _5501_/S VGND VGND VPWR VPWR _5501_/X sky130_fd_sc_hd__mux2_1
XFILLER_9_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_146_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3693_ _6787_/Q _5208_/A _4002_/A _6451_/Q VGND VGND VPWR VPWR _3693_/X sky130_fd_sc_hd__a22o_1
X_6481_ _6686_/CLK _6481_/D fanout492/X VGND VGND VPWR VPWR _6481_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_146_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5432_ hold533/X _5519_/A1 _5432_/S VGND VGND VPWR VPWR _5432_/X sky130_fd_sc_hd__mux2_1
XFILLER_145_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput302 _3950_/X VGND VGND VPWR VPWR ser_rx sky130_fd_sc_hd__buf_12
XFILLER_145_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_161_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput313 hold1369/X VGND VGND VPWR VPWR wb_ack_o sky130_fd_sc_hd__buf_12
XFILLER_133_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5363_ _5363_/A0 _5495_/A1 _5369_/S VGND VGND VPWR VPWR _5363_/X sky130_fd_sc_hd__mux2_1
XFILLER_99_310 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput324 hold1313/X VGND VGND VPWR VPWR hold1314/A sky130_fd_sc_hd__buf_12
Xoutput335 hold1315/X VGND VGND VPWR VPWR hold1316/A sky130_fd_sc_hd__buf_12
XFILLER_114_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7102_ _7124_/CLK _7102_/D fanout503/X VGND VGND VPWR VPWR _7102_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_99_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4314_ hold459/X _5534_/A1 _4314_/S VGND VGND VPWR VPWR _4314_/X sky130_fd_sc_hd__mux2_1
XFILLER_87_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5294_ _5294_/A0 _5465_/A1 _5297_/S VGND VGND VPWR VPWR _5294_/X sky130_fd_sc_hd__mux2_1
XFILLER_113_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_141_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4245_ hold901/X _5189_/A1 hold63/X VGND VGND VPWR VPWR _4245_/X sky130_fd_sc_hd__mux2_1
X_7033_ _7033_/CLK _7033_/D fanout507/X VGND VGND VPWR VPWR _7033_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_101_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4176_ _3625_/X _4176_/A1 _4180_/S VGND VGND VPWR VPWR _6586_/D sky130_fd_sc_hd__mux2_1
XFILLER_142_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6817_ _6969_/CLK _6817_/D fanout507/X VGND VGND VPWR VPWR _6817_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_11_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6748_ _7010_/CLK _6748_/D fanout498/X VGND VGND VPWR VPWR _6748_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_7_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6679_ _7155_/CLK _6679_/D _6370_/A VGND VGND VPWR VPWR _6679_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_176_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_191_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_191_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_516 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_104_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_116_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_120_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xmgmt_gpio_14_buff_inst _3931_/X VGND VGND VPWR VPWR mgmt_gpio_out[14] sky130_fd_sc_hd__clkbuf_8
XFILLER_58_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_427 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_186_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_157_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_173_80 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4030_ hold640/X _4289_/A1 _4031_/S VGND VGND VPWR VPWR _4030_/X sky130_fd_sc_hd__mux2_1
XFILLER_111_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_711 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5981_ _5981_/A _5981_/B _5981_/C VGND VGND VPWR VPWR _5981_/X sky130_fd_sc_hd__and3_4
XFILLER_80_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4932_ _5112_/A _4932_/B _4932_/C VGND VGND VPWR VPWR _4940_/C sky130_fd_sc_hd__and3_1
X_4863_ _4594_/X _4620_/B _5088_/C _4933_/C _4862_/X VGND VGND VPWR VPWR _4879_/C
+ sky130_fd_sc_hd__o2111a_1
X_6602_ _6683_/CLK _6602_/D fanout509/X VGND VGND VPWR VPWR _6602_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA_14 _5478_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3814_ _3814_/A _3814_/B _3814_/C _3814_/D VGND VGND VPWR VPWR _3815_/D sky130_fd_sc_hd__nor4_1
XANTENNA_25 _3433_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_36 _4321_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4794_ _4479_/A _4921_/A _5043_/B _4676_/B VGND VGND VPWR VPWR _4813_/B sky130_fd_sc_hd__o22a_1
XFILLER_177_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_47 _3816_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_192_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_58 _5937_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_146_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6533_ _6711_/CLK _6533_/D fanout486/X VGND VGND VPWR VPWR _6533_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA_69 _6467_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3745_ _3745_/A _3745_/B _3745_/C _3745_/D VGND VGND VPWR VPWR _3746_/D sky130_fd_sc_hd__nor4_1
XFILLER_118_234 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6464_ _6559_/CLK _6464_/D _3264_/A VGND VGND VPWR VPWR _6464_/Q sky130_fd_sc_hd__dfrtp_1
X_3676_ _6627_/Q _4225_/A _4214_/A _6621_/Q _3675_/X VGND VGND VPWR VPWR _3683_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_161_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5415_ _5415_/A _5529_/B VGND VGND VPWR VPWR _5423_/S sky130_fd_sc_hd__and2_4
XFILLER_173_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6395_ _6396_/A _6396_/B VGND VGND VPWR VPWR _6395_/X sky130_fd_sc_hd__and2_1
XFILLER_133_248 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5346_ hold355/X _5523_/A1 _5351_/S VGND VGND VPWR VPWR _5346_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput176 _3211_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[10] sky130_fd_sc_hd__buf_12
XFILLER_102_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput187 _3200_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[20] sky130_fd_sc_hd__buf_12
Xoutput198 _3190_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[30] sky130_fd_sc_hd__buf_12
XFILLER_141_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5277_ hold673/X _5544_/A1 _5279_/S VGND VGND VPWR VPWR _5277_/X sky130_fd_sc_hd__mux2_1
X_7016_ _7017_/CLK _7016_/D fanout515/X VGND VGND VPWR VPWR _7016_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_101_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4228_ hold819/X _5505_/A1 _4230_/S VGND VGND VPWR VPWR _4228_/X sky130_fd_sc_hd__mux2_1
XFILLER_46_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4159_ _3747_/Y _4159_/A1 _4165_/S VGND VGND VPWR VPWR _6571_/D sky130_fd_sc_hd__mux2_1
XFILLER_28_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_471 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_532 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_340 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_192_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_424 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_174_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput12 mask_rev_in[17] VGND VGND VPWR VPWR input12/X sky130_fd_sc_hd__clkbuf_2
Xinput23 mask_rev_in[27] VGND VGND VPWR VPWR input23/X sky130_fd_sc_hd__buf_2
Xinput34 mask_rev_in[8] VGND VGND VPWR VPWR input34/X sky130_fd_sc_hd__clkbuf_1
Xinput45 mgmt_gpio_in[18] VGND VGND VPWR VPWR input45/X sky130_fd_sc_hd__clkbuf_4
X_3530_ _7006_/Q _5451_/A _4151_/A _6569_/Q _3528_/X VGND VGND VPWR VPWR _3535_/C
+ sky130_fd_sc_hd__a221o_1
Xinput56 mgmt_gpio_in[28] VGND VGND VPWR VPWR input56/X sky130_fd_sc_hd__dlymetal6s2s_1
Xinput67 mgmt_gpio_in[3] VGND VGND VPWR VPWR _3263_/C sky130_fd_sc_hd__buf_6
Xhold807 _6428_/Q VGND VGND VPWR VPWR hold807/X sky130_fd_sc_hd__dlygate4sd3_1
Xinput78 spi_csb VGND VGND VPWR VPWR input78/X sky130_fd_sc_hd__clkbuf_1
XFILLER_128_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold818 _3964_/X VGND VGND VPWR VPWR _6420_/D sky130_fd_sc_hd__dlygate4sd3_1
Xinput89 spimemio_flash_io2_do VGND VGND VPWR VPWR input89/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold829 _6621_/Q VGND VGND VPWR VPWR hold829/X sky130_fd_sc_hd__dlygate4sd3_1
X_3461_ _3461_/A _3461_/B _3461_/C _3460_/Y VGND VGND VPWR VPWR _3471_/C sky130_fd_sc_hd__or4b_1
XFILLER_143_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5200_ _5200_/A0 hold588/X _5207_/S VGND VGND VPWR VPWR _5200_/X sky130_fd_sc_hd__mux2_1
XFILLER_42_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6180_ _6180_/A1 _5612_/Y _6178_/X _6179_/X VGND VGND VPWR VPWR _7126_/D sky130_fd_sc_hd__o22a_1
X_3392_ _3557_/A _3487_/A VGND VGND VPWR VPWR _5511_/A sky130_fd_sc_hd__nor2_8
XFILLER_170_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5131_ _5131_/A _5131_/B _5131_/C _5130_/X VGND VGND VPWR VPWR _5131_/X sky130_fd_sc_hd__or4b_1
XFILLER_69_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5062_ _5062_/A _5062_/B _5062_/C VGND VGND VPWR VPWR _5112_/B sky130_fd_sc_hd__and3_1
Xhold1507 _6640_/Q VGND VGND VPWR VPWR _3948_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1518 hold37/A VGND VGND VPWR VPWR _3852_/A1 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1529 _7099_/Q VGND VGND VPWR VPWR _5591_/A1 sky130_fd_sc_hd__dlygate4sd3_1
X_4013_ hold515/X _5534_/A1 _4013_/S VGND VGND VPWR VPWR _4013_/X sky130_fd_sc_hd__mux2_1
XFILLER_37_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_224 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5964_ _5964_/A _5965_/B VGND VGND VPWR VPWR _5973_/C sky130_fd_sc_hd__nor2_8
X_4915_ _4915_/A _4915_/B _4960_/C VGND VGND VPWR VPWR _5062_/A sky130_fd_sc_hd__and3_1
XFILLER_178_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5895_ _5895_/A _5895_/B VGND VGND VPWR VPWR _5895_/X sky130_fd_sc_hd__or2_1
XFILLER_178_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4846_ _4721_/B _5026_/A _4788_/A _5106_/A VGND VGND VPWR VPWR _4846_/X sky130_fd_sc_hd__o31a_1
XFILLER_21_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4777_ _4883_/C _5020_/A _4776_/X _4363_/Y VGND VGND VPWR VPWR _4881_/B sky130_fd_sc_hd__a31o_1
XFILLER_193_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6516_ _7060_/CLK _6516_/D fanout521/X VGND VGND VPWR VPWR _6516_/Q sky130_fd_sc_hd__dfrtp_1
X_3728_ input72/X hold76/A _4139_/A _6556_/Q _3727_/X VGND VGND VPWR VPWR _3736_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_4_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6447_ _6881_/CLK _6447_/D fanout523/X VGND VGND VPWR VPWR _6447_/Q sky130_fd_sc_hd__dfrtp_2
X_3659_ _6844_/Q _5271_/A _4139_/A _6557_/Q VGND VGND VPWR VPWR _3659_/X sky130_fd_sc_hd__a22o_1
XFILLER_161_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6378_ _6399_/A _6399_/B VGND VGND VPWR VPWR _6378_/X sky130_fd_sc_hd__and2_1
XFILLER_121_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_611 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5329_ hold557/X _5515_/A1 _5333_/S VGND VGND VPWR VPWR _5329_/X sky130_fd_sc_hd__mux2_1
XFILLER_102_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_730 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_180_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_189_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_113_708 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_94_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4700_ _4701_/A _4717_/B VGND VGND VPWR VPWR _4767_/B sky130_fd_sc_hd__nor2_1
XTAP_1191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5680_ _6963_/Q _5648_/X _5919_/B1 _6891_/Q VGND VGND VPWR VPWR _5680_/X sky130_fd_sc_hd__a22o_1
XFILLER_148_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_435 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4631_ _4631_/A _4672_/B VGND VGND VPWR VPWR _4631_/X sky130_fd_sc_hd__or2_2
XFILLER_147_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4562_ _4943_/A _4565_/B VGND VGND VPWR VPWR _4563_/B sky130_fd_sc_hd__nor2_1
XFILLER_162_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6301_ _6669_/Q _5977_/X _6298_/X _6300_/X VGND VGND VPWR VPWR _6302_/C sky130_fd_sc_hd__a211o_1
XFILLER_143_310 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold604 _7184_/A VGND VGND VPWR VPWR hold604/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold615 _4068_/X VGND VGND VPWR VPWR _6500_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3513_ _6446_/Q _3361_/Y _4096_/A _7199_/A _3512_/X VGND VGND VPWR VPWR _3518_/C
+ sky130_fd_sc_hd__a221o_1
Xhold626 _6673_/Q VGND VGND VPWR VPWR hold626/X sky130_fd_sc_hd__dlygate4sd3_1
X_4493_ _5043_/A _4748_/A VGND VGND VPWR VPWR _5074_/A sky130_fd_sc_hd__or2_1
Xhold637 _4000_/X VGND VGND VPWR VPWR _6448_/D sky130_fd_sc_hd__dlygate4sd3_1
Xmax_cap356 _3706_/B VGND VGND VPWR VPWR _5168_/A sky130_fd_sc_hd__buf_12
Xhold648 _6558_/Q VGND VGND VPWR VPWR hold648/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmax_cap367 _5601_/Y VGND VGND VPWR VPWR _6295_/A2 sky130_fd_sc_hd__buf_8
X_6232_ _6647_/Q _5950_/X _5952_/Y _7153_/Q _6231_/X VGND VGND VPWR VPWR _6232_/X
+ sky130_fd_sc_hd__a221o_1
Xhold659 _5234_/X VGND VGND VPWR VPWR _6809_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_131_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3444_ _6431_/Q _3975_/A _5415_/A _6975_/Q VGND VGND VPWR VPWR _3444_/X sky130_fd_sc_hd__a22o_1
Xmax_cap378 _5972_/C VGND VGND VPWR VPWR _6294_/A2 sky130_fd_sc_hd__buf_12
Xmax_cap389 _5962_/X VGND VGND VPWR VPWR _6285_/A2 sky130_fd_sc_hd__buf_12
XFILLER_131_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6163_ _6849_/Q _5939_/X _5942_/X _6945_/Q VGND VGND VPWR VPWR _6163_/X sky130_fd_sc_hd__a22o_1
X_3375_ _3571_/A _3560_/B VGND VGND VPWR VPWR _4077_/S sky130_fd_sc_hd__nor2_8
XFILLER_170_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5114_ _4695_/B _5043_/X _5052_/X _5082_/X VGND VGND VPWR VPWR _5114_/X sky130_fd_sc_hd__o211a_1
Xhold1304 _5348_/X VGND VGND VPWR VPWR _6910_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6094_ _6982_/Q _6176_/A2 _6282_/A2 _6998_/Q VGND VGND VPWR VPWR _6094_/X sky130_fd_sc_hd__a22o_1
XTAP_986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1315 _6314_/A1 VGND VGND VPWR VPWR hold1315/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1326 hold1326/A VGND VGND VPWR VPWR wb_dat_o[10] sky130_fd_sc_hd__buf_12
Xhold1337 _4159_/A1 VGND VGND VPWR VPWR hold1337/X sky130_fd_sc_hd__dlygate4sd3_1
X_5045_ _4703_/B _5043_/X _5044_/X _4995_/X VGND VGND VPWR VPWR _5085_/B sky130_fd_sc_hd__o211ai_1
Xhold1348 hold1348/A VGND VGND VPWR VPWR wb_dat_o[31] sky130_fd_sc_hd__buf_12
Xhold1359 _6315_/A1 VGND VGND VPWR VPWR hold1359/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_27_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_246 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6996_ _7039_/CLK _6996_/D fanout498/X VGND VGND VPWR VPWR _6996_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_80_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5947_ _5959_/A _5980_/B VGND VGND VPWR VPWR _5947_/Y sky130_fd_sc_hd__nor2_8
XFILLER_178_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5878_ _6697_/Q _5626_/X _5629_/X _6467_/Q _5877_/X VGND VGND VPWR VPWR _5886_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_139_638 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4829_ _4943_/A _4943_/B _4565_/B VGND VGND VPWR VPWR _4829_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_193_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_660 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_181_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_343 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_124_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_758 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_189_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_190 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_363 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_144_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_172_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_346 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1 hold1/A VGND VGND VPWR VPWR hold1/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_94_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_179 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6850_ _7063_/CLK _6850_/D fanout504/X VGND VGND VPWR VPWR _6850_/Q sky130_fd_sc_hd__dfstp_1
X_5801_ _5801_/A1 _6305_/A2 _5799_/X _5800_/X VGND VGND VPWR VPWR _7112_/D sky130_fd_sc_hd__o22a_1
XFILLER_90_683 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6781_ _7017_/CLK _6781_/D fanout515/X VGND VGND VPWR VPWR _6781_/Q sky130_fd_sc_hd__dfrtp_1
X_3993_ _3993_/A _5511_/B VGND VGND VPWR VPWR _4001_/S sky130_fd_sc_hd__and2_4
X_5732_ _6973_/Q _5644_/X _5724_/X _5726_/X _5731_/X VGND VGND VPWR VPWR _5732_/X
+ sky130_fd_sc_hd__a2111o_2
XFILLER_31_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5663_ _6834_/Q _5617_/X _5920_/A2 _6826_/Q VGND VGND VPWR VPWR _5663_/X sky130_fd_sc_hd__a22o_1
XFILLER_148_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4614_ _4614_/A _4630_/B VGND VGND VPWR VPWR _4615_/B sky130_fd_sc_hd__or2_4
XFILLER_135_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5594_ _6508_/Q _5979_/A _5979_/B VGND VGND VPWR VPWR _5594_/X sky130_fd_sc_hd__and3_1
XFILLER_129_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_191_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold401 _6894_/Q VGND VGND VPWR VPWR hold401/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_163_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4545_ _4545_/A _4632_/B VGND VGND VPWR VPWR _4788_/A sky130_fd_sc_hd__nand2_8
Xhold412 _5391_/X VGND VGND VPWR VPWR _6948_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold423 _7038_/Q VGND VGND VPWR VPWR hold423/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold434 _5373_/X VGND VGND VPWR VPWR _6932_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold445 _6714_/Q VGND VGND VPWR VPWR hold445/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold456 _5514_/X VGND VGND VPWR VPWR _7057_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_171_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4476_ _4554_/A _4629_/B VGND VGND VPWR VPWR _4943_/C sky130_fd_sc_hd__or2_1
Xhold467 _7046_/Q VGND VGND VPWR VPWR hold467/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_387 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold478 _3974_/X VGND VGND VPWR VPWR _6425_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6215_ _6605_/Q wire390/X _5978_/X _6696_/Q VGND VGND VPWR VPWR _6215_/X sky130_fd_sc_hd__a22o_1
Xhold489 _6935_/Q VGND VGND VPWR VPWR hold489/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_131_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3427_ _6800_/Q _5217_/A _5415_/A _6976_/Q _3426_/X VGND VGND VPWR VPWR _3432_/C
+ sky130_fd_sc_hd__a221o_1
X_7195_ _7195_/A VGND VGND VPWR VPWR _7195_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_131_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_131_368 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6146_ _6856_/Q _5975_/A _5975_/C _7053_/Q VGND VGND VPWR VPWR _6146_/X sky130_fd_sc_hd__a22o_1
XFILLER_38_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3358_ _3797_/A _3563_/A VGND VGND VPWR VPWR _5478_/A sky130_fd_sc_hd__nor2_8
XTAP_772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1101 _6694_/Q VGND VGND VPWR VPWR _4296_/A0 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1112 _4226_/X VGND VGND VPWR VPWR _6625_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1123 _6751_/Q VGND VGND VPWR VPWR _5164_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_57_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6077_ _6077_/A _6077_/B _6077_/C _5975_/X VGND VGND VPWR VPWR _6077_/X sky130_fd_sc_hd__or4b_1
Xhold1134 _5525_/X VGND VGND VPWR VPWR _7067_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1145 _6650_/Q VGND VGND VPWR VPWR _4244_/A0 sky130_fd_sc_hd__dlygate4sd3_1
X_3289_ hold81/X _3440_/A VGND VGND VPWR VPWR _3797_/A sky130_fd_sc_hd__or2_4
Xhold1156 _5494_/X VGND VGND VPWR VPWR _7039_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1167 _6970_/Q VGND VGND VPWR VPWR _5416_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_73_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1178 _5488_/X VGND VGND VPWR VPWR _7034_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_57_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5028_ _4587_/A _5025_/Y _5027_/Y _4828_/A VGND VGND VPWR VPWR _5037_/A sky130_fd_sc_hd__o22a_1
XTAP_2606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1189 _6555_/Q VGND VGND VPWR VPWR _4140_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_650 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_717 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_683 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_599 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6979_ _7011_/CLK _6979_/D fanout500/X VGND VGND VPWR VPWR _6979_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_110_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_179_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_154_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_182_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_162 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold990 _6427_/Q VGND VGND VPWR VPWR hold990/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_135_73 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_135_95 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_330 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_352 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_158_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_185_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_172_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4330_ _4679_/A _4542_/A VGND VGND VPWR VPWR _4448_/A sky130_fd_sc_hd__and2b_1
XFILLER_141_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4261_ _4261_/A _5187_/B VGND VGND VPWR VPWR _4266_/S sky130_fd_sc_hd__and2_2
X_6000_ _6978_/Q _5943_/Y _5953_/Y _6994_/Q VGND VGND VPWR VPWR _6000_/X sky130_fd_sc_hd__a22o_1
XFILLER_140_154 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3212_ _6861_/Q VGND VGND VPWR VPWR _3212_/Y sky130_fd_sc_hd__inv_2
X_4192_ hold937/X _5189_/A1 _4195_/S VGND VGND VPWR VPWR _4192_/X sky130_fd_sc_hd__mux2_1
XFILLER_39_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6902_ _7082_/CLK hold24/X fanout519/X VGND VGND VPWR VPWR _6902_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_23_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6833_ _6887_/CLK _6833_/D fanout524/X VGND VGND VPWR VPWR _6833_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_24_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_519 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6764_ _7071_/CLK _6764_/D fanout504/X VGND VGND VPWR VPWR _6764_/Q sky130_fd_sc_hd__dfrtp_1
X_3976_ _3976_/A0 _5488_/A1 _3983_/S VGND VGND VPWR VPWR _3976_/X sky130_fd_sc_hd__mux2_1
X_5715_ _6989_/Q _5622_/X _5624_/X _6829_/Q VGND VGND VPWR VPWR _5715_/X sky130_fd_sc_hd__a22o_1
X_6695_ _6695_/CLK _6695_/D fanout490/X VGND VGND VPWR VPWR _6695_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_176_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5646_ _5646_/A _5646_/B _5649_/C VGND VGND VPWR VPWR _5646_/X sky130_fd_sc_hd__and3_4
XFILLER_40_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_164_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_191_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5577_ _7095_/Q _5577_/B VGND VGND VPWR VPWR _5579_/B sky130_fd_sc_hd__nor2_1
XFILLER_117_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_163_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold220 _5450_/X VGND VGND VPWR VPWR _7001_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_2_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold231 _6517_/Q VGND VGND VPWR VPWR hold231/X sky130_fd_sc_hd__dlygate4sd3_1
X_4528_ _4977_/B _4692_/C _4965_/B VGND VGND VPWR VPWR _4755_/A sky130_fd_sc_hd__nor3_1
XFILLER_191_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold242 _5350_/X VGND VGND VPWR VPWR _6912_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_132_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold253 _7074_/Q VGND VGND VPWR VPWR hold253/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold264 _4283_/X VGND VGND VPWR VPWR _6683_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_131_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold275 hold275/A VGND VGND VPWR VPWR hold275/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_132_655 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4459_ _4943_/A _4828_/A VGND VGND VPWR VPWR _4505_/D sky130_fd_sc_hd__or2_1
Xhold286 _4093_/X VGND VGND VPWR VPWR _6516_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold297 _7075_/Q VGND VGND VPWR VPWR hold297/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_131_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7178_ _7178_/A VGND VGND VPWR VPWR _7178_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_105_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6129_ _6129_/A1 _5612_/A _5612_/B VGND VGND VPWR VPWR _6129_/X sky130_fd_sc_hd__o21a_1
XTAP_580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_403 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_104 _3943_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_115 _3247_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_126 _3894_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_137 _6285_/A2 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_148 _5533_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_159 _3939_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_179_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_182_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_674 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_162_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_91_200 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_53_csclk _7000_/CLK VGND VGND VPWR VPWR _7033_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_92_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_189_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3830_ _6485_/Q _3830_/B VGND VGND VPWR VPWR _3857_/S sky130_fd_sc_hd__nand2b_4
Xclkbuf_leaf_68_csclk _7000_/CLK VGND VGND VPWR VPWR _7055_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_32_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_686 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3761_ _3761_/A _3761_/B VGND VGND VPWR VPWR _5181_/A sky130_fd_sc_hd__nor2_1
XFILLER_13_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5500_ hold211/X hold114/X _5501_/S VGND VGND VPWR VPWR _5500_/X sky130_fd_sc_hd__mux2_1
XFILLER_192_319 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6480_ _6769_/CLK _6480_/D fanout492/X VGND VGND VPWR VPWR _6480_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_72_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3692_ _6923_/Q _5361_/A _5460_/A _7011_/Q _3691_/X VGND VGND VPWR VPWR _3713_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_146_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_187_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5431_ hold257/X hold114/X _5432_/S VGND VGND VPWR VPWR _5431_/X sky130_fd_sc_hd__mux2_1
Xoutput303 _5605_/A VGND VGND VPWR VPWR serial_clock sky130_fd_sc_hd__buf_12
Xoutput314 hold1349/X VGND VGND VPWR VPWR hold1350/A sky130_fd_sc_hd__buf_12
X_5362_ _5362_/A0 _5530_/A1 _5369_/S VGND VGND VPWR VPWR _5362_/X sky130_fd_sc_hd__mux2_1
Xoutput325 hold1343/X VGND VGND VPWR VPWR hold1344/A sky130_fd_sc_hd__buf_12
Xoutput336 hold1351/X VGND VGND VPWR VPWR hold1352/A sky130_fd_sc_hd__buf_12
XFILLER_99_322 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7101_ _7124_/CLK _7101_/D fanout502/X VGND VGND VPWR VPWR _7101_/Q sky130_fd_sc_hd__dfstp_1
X_4313_ hold561/X _5491_/A1 _4314_/S VGND VGND VPWR VPWR _4313_/X sky130_fd_sc_hd__mux2_1
X_5293_ hold523/X _5515_/A1 _5297_/S VGND VGND VPWR VPWR _5293_/X sky130_fd_sc_hd__mux2_1
X_7032_ _7032_/CLK _7032_/D fanout507/X VGND VGND VPWR VPWR _7032_/Q sky130_fd_sc_hd__dfrtp_2
X_4244_ _4244_/A0 _5308_/A1 hold63/X VGND VGND VPWR VPWR _4244_/X sky130_fd_sc_hd__mux2_1
XFILLER_114_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4175_ _3684_/X _4175_/A1 _4180_/S VGND VGND VPWR VPWR _6585_/D sky130_fd_sc_hd__mux2_1
XFILLER_67_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6816_ _6969_/CLK _6816_/D fanout506/X VGND VGND VPWR VPWR _6816_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_50_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6747_ _7034_/CLK _6747_/D fanout488/X VGND VGND VPWR VPWR _6747_/Q sky130_fd_sc_hd__dfrtp_2
X_3959_ _3247_/A hold587/X _3959_/S VGND VGND VPWR VPWR _3959_/X sky130_fd_sc_hd__mux2_8
XFILLER_183_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6678_ _6718_/CLK _6678_/D _6401_/A VGND VGND VPWR VPWR _6678_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_136_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5629_ _5667_/A _5650_/B _5651_/C VGND VGND VPWR VPWR _5629_/X sky130_fd_sc_hd__and3_4
XFILLER_164_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout530 _4746_/A VGND VGND VPWR VPWR _4554_/A sky130_fd_sc_hd__buf_8
XFILLER_120_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_285 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_179 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_360 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_170_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_173_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5980_ _5980_/A _5980_/B VGND VGND VPWR VPWR _5980_/Y sky130_fd_sc_hd__nor2_8
XFILLER_92_564 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4931_ _4931_/A VGND VGND VPWR VPWR _4932_/C sky130_fd_sc_hd__clkinv_2
XFILLER_178_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4862_ _4862_/A _4862_/B VGND VGND VPWR VPWR _4862_/X sky130_fd_sc_hd__or2_1
XFILLER_177_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6601_ _6689_/CLK _6601_/D fanout509/X VGND VGND VPWR VPWR _6601_/Q sky130_fd_sc_hd__dfstp_1
X_3813_ _3813_/A _3813_/B VGND VGND VPWR VPWR _3814_/D sky130_fd_sc_hd__or2_1
XANTENNA_15 _5478_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_26 _3461_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4793_ _4793_/A _4793_/B VGND VGND VPWR VPWR _4793_/Y sky130_fd_sc_hd__nand2_1
XANTENNA_37 _4225_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_193_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_48 _5351_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6532_ _6707_/CLK _6532_/D fanout486/X VGND VGND VPWR VPWR _6532_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA_59 _5941_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3744_ _6427_/Q _3975_/A _4133_/A _6551_/Q _3743_/X VGND VGND VPWR VPWR _3745_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_192_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_192_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_146_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6463_ _6683_/CLK _6463_/D fanout509/X VGND VGND VPWR VPWR _6463_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_118_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3675_ _6567_/Q _4151_/A _4133_/A _6552_/Q VGND VGND VPWR VPWR _3675_/X sky130_fd_sc_hd__a22o_1
XFILLER_106_408 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5414_ hold847/X _5537_/A1 _5414_/S VGND VGND VPWR VPWR _5414_/X sky130_fd_sc_hd__mux2_1
X_6394_ _6396_/A _6396_/B VGND VGND VPWR VPWR _6394_/X sky130_fd_sc_hd__and2_1
X_5345_ hold963/X _5495_/A1 _5351_/S VGND VGND VPWR VPWR _5345_/X sky130_fd_sc_hd__mux2_1
Xoutput177 _3210_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[11] sky130_fd_sc_hd__buf_12
Xoutput188 _3199_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[21] sky130_fd_sc_hd__buf_12
X_5276_ _5276_/A0 _5465_/A1 _5279_/S VGND VGND VPWR VPWR _5276_/X sky130_fd_sc_hd__mux2_1
Xoutput199 _3189_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[31] sky130_fd_sc_hd__buf_12
XFILLER_101_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_135 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7015_ _7060_/CLK _7015_/D fanout522/X VGND VGND VPWR VPWR _7015_/Q sky130_fd_sc_hd__dfrtp_2
X_4227_ _4227_/A0 _5189_/A1 _4230_/S VGND VGND VPWR VPWR _4227_/X sky130_fd_sc_hd__mux2_1
XFILLER_56_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4158_ _3816_/X _4158_/A1 _4165_/S VGND VGND VPWR VPWR _6570_/D sky130_fd_sc_hd__mux2_1
XFILLER_28_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4089_ hold295/X _4088_/X _4095_/S VGND VGND VPWR VPWR _4089_/X sky130_fd_sc_hd__mux2_1
XFILLER_43_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_178_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_168_157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_544 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_514 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_474 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_400 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_436 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_175_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_174_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput13 mask_rev_in[18] VGND VGND VPWR VPWR input13/X sky130_fd_sc_hd__clkbuf_1
XFILLER_128_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput24 mask_rev_in[28] VGND VGND VPWR VPWR input24/X sky130_fd_sc_hd__clkbuf_2
Xinput35 mask_rev_in[9] VGND VGND VPWR VPWR input35/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_155_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput46 mgmt_gpio_in[19] VGND VGND VPWR VPWR input46/X sky130_fd_sc_hd__buf_2
Xinput57 mgmt_gpio_in[29] VGND VGND VPWR VPWR input57/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_6_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput68 mgmt_gpio_in[5] VGND VGND VPWR VPWR _3950_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_143_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold808 _3978_/X VGND VGND VPWR VPWR _6428_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_6_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput79 spi_enabled VGND VGND VPWR VPWR _3951_/B sky130_fd_sc_hd__clkbuf_4
Xhold819 _6627_/Q VGND VGND VPWR VPWR hold819/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_183_683 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3460_ _3460_/A _3460_/B _3460_/C VGND VGND VPWR VPWR _3460_/Y sky130_fd_sc_hd__nor3_1
XFILLER_155_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_131_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3391_ _3761_/A _3391_/B VGND VGND VPWR VPWR _5520_/A sky130_fd_sc_hd__nor2_8
XFILLER_130_208 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5130_ _4748_/B _4745_/B _4940_/B _5129_/X VGND VGND VPWR VPWR _5130_/X sky130_fd_sc_hd__o211a_1
XFILLER_35_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1508 _6489_/Q VGND VGND VPWR VPWR _3905_/B1 sky130_fd_sc_hd__dlygate4sd3_1
X_5061_ _5061_/A _5100_/B _5061_/C _5061_/D VGND VGND VPWR VPWR _5062_/C sky130_fd_sc_hd__and4_1
XFILLER_96_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1519 hold29/A VGND VGND VPWR VPWR _3846_/A1 sky130_fd_sc_hd__dlygate4sd3_1
X_4012_ hold581/X _5491_/A1 _4013_/S VGND VGND VPWR VPWR _4012_/X sky130_fd_sc_hd__mux2_1
XFILLER_92_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_383 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5963_ _5979_/A _5977_/A _5963_/C VGND VGND VPWR VPWR _5963_/X sky130_fd_sc_hd__and3_4
XFILLER_52_236 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_opt_4_0_csclk clkbuf_3_6_0_csclk/X VGND VGND VPWR VPWR clkbuf_opt_4_0_csclk/X
+ sky130_fd_sc_hd__clkbuf_16
X_4914_ _4914_/A _4914_/B VGND VGND VPWR VPWR _4914_/Y sky130_fd_sc_hd__nand2_1
XFILLER_80_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5894_ _6708_/Q _5630_/X _5634_/X _6688_/Q VGND VGND VPWR VPWR _5895_/B sky130_fd_sc_hd__a22o_1
XFILLER_178_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_280 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4845_ _4515_/B _4831_/X _4833_/X _4844_/X VGND VGND VPWR VPWR _4845_/X sky130_fd_sc_hd__o211a_1
XFILLER_32_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4776_ _5022_/B _4703_/A _4898_/B _4746_/X _4775_/X VGND VGND VPWR VPWR _4776_/X
+ sky130_fd_sc_hd__o2111a_1
XFILLER_165_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6515_ _7022_/CLK _6515_/D fanout517/X VGND VGND VPWR VPWR _6515_/Q sky130_fd_sc_hd__dfrtp_1
X_3727_ _7019_/Q hold18/A _5397_/A _6955_/Q VGND VGND VPWR VPWR _3727_/X sky130_fd_sc_hd__a22o_1
XFILLER_146_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6446_ _7041_/CLK _6446_/D fanout518/X VGND VGND VPWR VPWR _6446_/Q sky130_fd_sc_hd__dfrtp_4
X_3658_ _6900_/Q _5334_/A _5289_/A _6860_/Q _3657_/X VGND VGND VPWR VPWR _3661_/C
+ sky130_fd_sc_hd__a221o_1
X_6377_ _6400_/A _6399_/B VGND VGND VPWR VPWR _6377_/X sky130_fd_sc_hd__and2_1
X_3589_ _6797_/Q _5217_/A _4133_/A _6553_/Q VGND VGND VPWR VPWR _3589_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_623 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5328_ hold337/X _5541_/A1 _5333_/S VGND VGND VPWR VPWR _5328_/X sky130_fd_sc_hd__mux2_1
XFILLER_88_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5259_ hold743/X _5457_/A1 _5261_/S VGND VGND VPWR VPWR _5259_/X sky130_fd_sc_hd__mux2_1
XFILLER_87_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_575 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_149_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_171_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_374 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_154_61 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_179_80 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4630_ _4630_/A _4630_/B VGND VGND VPWR VPWR _4672_/B sky130_fd_sc_hd__or2_2
XFILLER_8_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4561_ _4561_/A _4561_/B VGND VGND VPWR VPWR _4565_/B sky130_fd_sc_hd__or2_1
X_6300_ _6464_/Q _5943_/Y _6300_/B1 _6623_/Q _6299_/X VGND VGND VPWR VPWR _6300_/X
+ sky130_fd_sc_hd__a221o_1
X_3512_ _6934_/Q hold41/A _4038_/A _6484_/Q VGND VGND VPWR VPWR _3512_/X sky130_fd_sc_hd__a22o_1
XFILLER_116_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold605 _4053_/X VGND VGND VPWR VPWR _6493_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_7_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold616 _6717_/Q VGND VGND VPWR VPWR hold616/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_143_322 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4492_ _4622_/A _4703_/A VGND VGND VPWR VPWR _4492_/Y sky130_fd_sc_hd__nor2_1
Xhold627 _4271_/X VGND VGND VPWR VPWR _6673_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold638 _7186_/A VGND VGND VPWR VPWR hold638/X sky130_fd_sc_hd__dlygate4sd3_1
X_6231_ _6657_/Q _6288_/A2 _5977_/X _6667_/Q VGND VGND VPWR VPWR _6231_/X sky130_fd_sc_hd__a22o_1
Xhold649 _4143_/X VGND VGND VPWR VPWR _6558_/D sky130_fd_sc_hd__dlygate4sd3_1
Xmax_cap357 hold76/X VGND VGND VPWR VPWR _4092_/S sky130_fd_sc_hd__buf_6
X_3443_ _7044_/Q _5493_/A _3355_/Y input17/X VGND VGND VPWR VPWR _3443_/X sky130_fd_sc_hd__a22o_2
XFILLER_170_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_cap368 hold52/X VGND VGND VPWR VPWR hold53/A sky130_fd_sc_hd__buf_12
Xmax_cap379 _5953_/Y VGND VGND VPWR VPWR _6282_/A2 sky130_fd_sc_hd__buf_8
XFILLER_131_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6162_ _6817_/Q _5936_/X _5972_/B _7062_/Q _6161_/X VGND VGND VPWR VPWR _6168_/C
+ sky130_fd_sc_hd__a221o_1
XTAP_921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3374_ _3374_/A _3390_/B VGND VGND VPWR VPWR _3374_/Y sky130_fd_sc_hd__nor2_8
XTAP_932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5113_ _4994_/A _5065_/Y _5108_/Y _5131_/C _5112_/X VGND VGND VPWR VPWR _5113_/X
+ sky130_fd_sc_hd__o41a_1
XTAP_954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6093_ _6093_/A _6093_/B _6093_/C _6092_/Y VGND VGND VPWR VPWR _6093_/X sky130_fd_sc_hd__or4b_1
XTAP_976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1305 hold1395/X VGND VGND VPWR VPWR hold1305/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1316 hold1316/A VGND VGND VPWR VPWR wb_dat_o[29] sky130_fd_sc_hd__buf_12
Xhold1327 _4188_/A1 VGND VGND VPWR VPWR hold1327/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5044_ _4901_/B _4962_/X _4615_/B _4678_/A VGND VGND VPWR VPWR _5044_/X sky130_fd_sc_hd__a211o_1
Xhold1338 hold1338/A VGND VGND VPWR VPWR wb_dat_o[17] sky130_fd_sc_hd__buf_12
XFILLER_38_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1349 _4182_/A1 VGND VGND VPWR VPWR hold1349/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_72_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6995_ _7046_/CLK _6995_/D fanout500/X VGND VGND VPWR VPWR _6995_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_25_258 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5946_ _5981_/A _5979_/A _5963_/C VGND VGND VPWR VPWR _5946_/X sky130_fd_sc_hd__and3_4
XFILLER_41_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5877_ _6552_/Q _5639_/X _5649_/X _6677_/Q VGND VGND VPWR VPWR _5877_/X sky130_fd_sc_hd__a22o_1
XFILLER_179_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4828_ _4828_/A _5026_/A VGND VGND VPWR VPWR _4828_/X sky130_fd_sc_hd__or2_1
XFILLER_138_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4759_ _4965_/A _4703_/B _4505_/D VGND VGND VPWR VPWR _5007_/B sky130_fd_sc_hd__o21a_1
XFILLER_107_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_193_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_161_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6429_ _7034_/CLK _6429_/D fanout489/X VGND VGND VPWR VPWR _6429_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_134_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_187_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_375 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_165_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_152_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_99_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_180_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_228 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_140_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold2 hold2/A VGND VGND VPWR VPWR hold2/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_181_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_456 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5800_ _7111_/Q _5612_/A _5612_/B VGND VGND VPWR VPWR _5800_/X sky130_fd_sc_hd__o21a_1
XFILLER_23_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6780_ _7069_/CLK _6780_/D fanout521/X VGND VGND VPWR VPWR _6780_/Q sky130_fd_sc_hd__dfrtp_1
X_3992_ hold491/X _5519_/A1 _3992_/S VGND VGND VPWR VPWR _3992_/X sky130_fd_sc_hd__mux2_1
XFILLER_90_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5731_ _6837_/Q _5928_/A2 _5727_/X _5728_/X _5730_/X VGND VGND VPWR VPWR _5731_/X
+ sky130_fd_sc_hd__a2111o_1
XFILLER_176_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_176_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_188_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5662_ _7010_/Q _5620_/X _5629_/X _7018_/Q _5635_/X VGND VGND VPWR VPWR _5662_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_175_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_176_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4613_ _4617_/B _4888_/A _4613_/C VGND VGND VPWR VPWR _4630_/B sky130_fd_sc_hd__nand3b_4
X_5593_ _5593_/A _5962_/B VGND VGND VPWR VPWR _5596_/B sky130_fd_sc_hd__nand2_1
XFILLER_191_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_163_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4544_ _4544_/A _4544_/B VGND VGND VPWR VPWR _4632_/B sky130_fd_sc_hd__xnor2_4
Xhold402 _5330_/X VGND VGND VPWR VPWR _6894_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_144_631 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold413 _6741_/Q VGND VGND VPWR VPWR hold413/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold424 _5492_/X VGND VGND VPWR VPWR _7038_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold435 _6793_/Q VGND VGND VPWR VPWR hold435/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold446 _4320_/X VGND VGND VPWR VPWR _6714_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4475_ _4554_/A _4629_/B VGND VGND VPWR VPWR _4793_/A sky130_fd_sc_hd__nor2_4
XFILLER_116_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold457 _6554_/Q VGND VGND VPWR VPWR hold457/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold468 _5501_/X VGND VGND VPWR VPWR _7046_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6214_ _6691_/Q _5972_/B _5976_/Y _6476_/Q _6213_/X VGND VGND VPWR VPWR _6217_/A
+ sky130_fd_sc_hd__a221o_1
Xhold479 _7037_/Q VGND VGND VPWR VPWR hold479/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_399 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3426_ _6992_/Q hold34/A hold41/A _6936_/Q VGND VGND VPWR VPWR _3426_/X sky130_fd_sc_hd__a22o_1
X_7194_ _7194_/A VGND VGND VPWR VPWR _7194_/X sky130_fd_sc_hd__clkbuf_1
XTAP_740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6145_ _6984_/Q _6176_/A2 _6299_/A2 _6800_/Q _6144_/X VGND VGND VPWR VPWR _6152_/A
+ sky130_fd_sc_hd__a221o_1
XTAP_751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3357_ _3557_/A _3719_/A VGND VGND VPWR VPWR _5502_/A sky130_fd_sc_hd__nor2_8
XFILLER_100_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1102 _4296_/X VGND VGND VPWR VPWR _6694_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1113 _6609_/Q VGND VGND VPWR VPWR _4203_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1124 _5164_/X VGND VGND VPWR VPWR _6751_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6076_ _7029_/Q _5947_/Y _6073_/X _6075_/X VGND VGND VPWR VPWR _6077_/C sky130_fd_sc_hd__a211o_1
Xhold1135 _6786_/Q VGND VGND VPWR VPWR _5209_/A0 sky130_fd_sc_hd__dlygate4sd3_1
X_3288_ hold39/X hold51/X VGND VGND VPWR VPWR _3440_/A sky130_fd_sc_hd__or2_1
Xhold1146 _4244_/X VGND VGND VPWR VPWR _6650_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_57_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5027_ _5027_/A VGND VGND VPWR VPWR _5027_/Y sky130_fd_sc_hd__inv_2
Xhold1157 _7059_/Q VGND VGND VPWR VPWR _5516_/A0 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1168 _5416_/X VGND VGND VPWR VPWR _6970_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_73_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1179 _7026_/Q VGND VGND VPWR VPWR _5479_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_26_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_191 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6978_ _6978_/CLK _6978_/D fanout490/X VGND VGND VPWR VPWR _6978_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_81_695 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5929_ _6474_/Q _5622_/X _5929_/B1 _6469_/Q _5928_/X VGND VGND VPWR VPWR _5929_/Y
+ sky130_fd_sc_hd__a221oi_1
XFILLER_179_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_403 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_186_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_147_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_135_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_135_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold980 _6915_/Q VGND VGND VPWR VPWR hold980/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold991 _3977_/X VGND VGND VPWR VPWR _6427_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_189_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_189_347 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_126_620 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4260_ hold579/X _6357_/A1 _4260_/S VGND VGND VPWR VPWR _4260_/X sky130_fd_sc_hd__mux2_1
XFILLER_5_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_347 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3211_ _6869_/Q VGND VGND VPWR VPWR _3211_/Y sky130_fd_sc_hd__inv_2
X_4191_ _4191_/A0 _5308_/A1 _4195_/S VGND VGND VPWR VPWR _4191_/X sky130_fd_sc_hd__mux2_1
XFILLER_140_166 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_94_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6901_ _7058_/CLK _6901_/D fanout521/X VGND VGND VPWR VPWR _6901_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_47_191 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6832_ _6887_/CLK _6832_/D fanout524/X VGND VGND VPWR VPWR _6832_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_35_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3975_ _3975_/A _6352_/B VGND VGND VPWR VPWR _3983_/S sky130_fd_sc_hd__and2_2
X_6763_ _7039_/CLK _6763_/D fanout498/X VGND VGND VPWR VPWR _6763_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_149_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_149_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5714_ _3204_/Y _5923_/B _5667_/B VGND VGND VPWR VPWR _5714_/Y sky130_fd_sc_hd__a21oi_1
X_6694_ _7067_/CLK _6694_/D _3264_/A VGND VGND VPWR VPWR _6694_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_109_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5645_ _5667_/A _5645_/B _5650_/B VGND VGND VPWR VPWR _5645_/X sky130_fd_sc_hd__and3_4
XFILLER_191_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_163_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5576_ _7095_/Q _7094_/Q VGND VGND VPWR VPWR _5651_/B sky130_fd_sc_hd__nor2_4
XFILLER_156_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold210 _5242_/X VGND VGND VPWR VPWR _6816_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4527_ _4596_/B _4448_/A _4557_/B _4959_/A _4526_/X VGND VGND VPWR VPWR _4527_/X
+ sky130_fd_sc_hd__a311o_1
Xhold221 _6530_/Q VGND VGND VPWR VPWR hold221/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold232 _4095_/X VGND VGND VPWR VPWR _6517_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold243 _6766_/Q VGND VGND VPWR VPWR hold243/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold254 _5533_/X VGND VGND VPWR VPWR _7074_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold265 _6463_/Q VGND VGND VPWR VPWR hold265/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_131_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4458_ _4570_/B _4554_/A _4596_/B VGND VGND VPWR VPWR _4549_/B sky130_fd_sc_hd__or3b_4
Xhold276 _4049_/X VGND VGND VPWR VPWR _6491_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_49_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold287 hold287/A VGND VGND VPWR VPWR hold287/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_132_667 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold298 _5534_/X VGND VGND VPWR VPWR _7075_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3409_ _6904_/Q _5334_/A _5289_/A _6864_/Q VGND VGND VPWR VPWR _3409_/X sky130_fd_sc_hd__a22o_1
X_7177_ _7177_/A VGND VGND VPWR VPWR _7177_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_58_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_131_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4389_ _4592_/A _4409_/B _4617_/B VGND VGND VPWR VPWR _4390_/B sky130_fd_sc_hd__a21oi_1
XTAP_570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6128_ _6791_/Q _5975_/X _6118_/X _6127_/X _3174_/Y VGND VGND VPWR VPWR _6128_/X
+ sky130_fd_sc_hd__o221a_4
XFILLER_100_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6059_ _6845_/Q _5939_/X _6299_/A2 _6797_/Q VGND VGND VPWR VPWR _6059_/X sky130_fd_sc_hd__a22o_1
XFILLER_73_415 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_105 _7198_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_116 _3247_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_127 _3894_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_138 _5919_/B1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_149 _5515_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_139_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_154_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_182_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_686 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_150_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_162_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_212 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3760_ _6882_/Q hold83/A _4273_/A _6675_/Q _3759_/X VGND VGND VPWR VPWR _3778_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_158_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_192_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3691_ _6661_/Q _4255_/A _6352_/A _7152_/Q VGND VGND VPWR VPWR _3691_/X sky130_fd_sc_hd__a22o_1
XFILLER_173_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_145_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5430_ hold155/X hold142/X _5432_/S VGND VGND VPWR VPWR _5430_/X sky130_fd_sc_hd__mux2_1
XFILLER_145_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5361_ _5361_/A _5529_/B VGND VGND VPWR VPWR _5369_/S sky130_fd_sc_hd__and2_4
Xoutput304 _3439_/X VGND VGND VPWR VPWR serial_data_1 sky130_fd_sc_hd__buf_12
XFILLER_161_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_173_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput315 hold1325/X VGND VGND VPWR VPWR hold1326/A sky130_fd_sc_hd__buf_12
XFILLER_114_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput326 hold1357/X VGND VGND VPWR VPWR hold1358/A sky130_fd_sc_hd__buf_12
Xoutput337 hold1359/X VGND VGND VPWR VPWR hold1360/A sky130_fd_sc_hd__buf_12
X_4312_ hold801/X _6355_/A1 _4314_/S VGND VGND VPWR VPWR _4312_/X sky130_fd_sc_hd__mux2_1
X_7100_ _7131_/CLK _7100_/D fanout502/X VGND VGND VPWR VPWR _7100_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_99_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5292_ hold323/X _5523_/A1 _5297_/S VGND VGND VPWR VPWR _5292_/X sky130_fd_sc_hd__mux2_1
XFILLER_113_133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7031_ _7031_/CLK _7031_/D fanout522/X VGND VGND VPWR VPWR _7031_/Q sky130_fd_sc_hd__dfrtp_1
X_4243_ hold62/X _5187_/B VGND VGND VPWR VPWR hold63/A sky130_fd_sc_hd__and2_2
XFILLER_141_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4174_ _3747_/Y _4174_/A1 _4180_/S VGND VGND VPWR VPWR _6584_/D sky130_fd_sc_hd__mux2_1
XFILLER_67_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_234 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6815_ _7060_/CLK _6815_/D fanout521/X VGND VGND VPWR VPWR _6815_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_168_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6746_ _6746_/CLK _6746_/D fanout488/X VGND VGND VPWR VPWR _6746_/Q sky130_fd_sc_hd__dfstp_4
X_3958_ _3958_/A _5529_/B VGND VGND VPWR VPWR _3974_/S sky130_fd_sc_hd__and2_2
XFILLER_50_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6677_ _6711_/CLK _6677_/D fanout486/X VGND VGND VPWR VPWR _6677_/Q sky130_fd_sc_hd__dfstp_2
X_3889_ _6507_/Q _3887_/B _3886_/X _3876_/B _3889_/B2 VGND VGND VPWR VPWR _6509_/D
+ sky130_fd_sc_hd__a32o_1
XFILLER_137_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_149_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5628_ _5667_/A _5645_/B _5650_/B VGND VGND VPWR VPWR _5628_/X sky130_fd_sc_hd__and3b_4
XFILLER_136_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5559_ _5559_/A VGND VGND VPWR VPWR _5561_/B sky130_fd_sc_hd__clkinv_2
XFILLER_183_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_116_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout520 fanout525/X VGND VGND VPWR VPWR fanout520/X sky130_fd_sc_hd__buf_8
XFILLER_116_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_404 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_3_1_0_wb_clk_i clkbuf_3_1_0_wb_clk_i/A VGND VGND VPWR VPWR _7130_/CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_27_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_187_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_127_203 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_108_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_291 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_584 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_576 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4930_ _4959_/A _4999_/B _4930_/C _5087_/B VGND VGND VPWR VPWR _4931_/A sky130_fd_sc_hd__or4b_2
XFILLER_80_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4861_ _5005_/A _4861_/B VGND VGND VPWR VPWR _4933_/C sky130_fd_sc_hd__or2_1
XTAP_2790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6600_ _6630_/CLK _6600_/D fanout495/X VGND VGND VPWR VPWR _6600_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_82_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3812_ _6625_/Q _4225_/A _5142_/A _6735_/Q _3811_/X VGND VGND VPWR VPWR _3813_/B
+ sky130_fd_sc_hd__a221o_1
XANTENNA_16 _3360_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4792_ _4587_/A _4921_/A _5043_/B _4703_/B VGND VGND VPWR VPWR _4933_/B sky130_fd_sc_hd__o22a_1
XFILLER_177_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_27 _3461_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_38 _3502_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_177_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_49 _5369_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3743_ input44/X _3343_/Y _4145_/A _6561_/Q VGND VGND VPWR VPWR _3743_/X sky130_fd_sc_hd__a22o_1
X_6531_ _7082_/CLK hold28/X fanout520/X VGND VGND VPWR VPWR _6531_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_9_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_146_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3674_ _3674_/A _3674_/B _3674_/C _3673_/Y VGND VGND VPWR VPWR _3684_/C sky130_fd_sc_hd__or4b_2
X_6462_ _6699_/CLK _6462_/D fanout509/X VGND VGND VPWR VPWR _6462_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_134_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5413_ hold205/X hold114/X _5414_/S VGND VGND VPWR VPWR _5413_/X sky130_fd_sc_hd__mux2_1
XFILLER_146_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_161_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6393_ _6396_/A _6396_/B VGND VGND VPWR VPWR _6393_/X sky130_fd_sc_hd__and2_1
X_5344_ _5344_/A0 _5530_/A1 _5351_/S VGND VGND VPWR VPWR _5344_/X sky130_fd_sc_hd__mux2_1
XFILLER_161_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput178 _3209_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[12] sky130_fd_sc_hd__buf_12
XFILLER_114_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5275_ hold511/X _5515_/A1 _5279_/S VGND VGND VPWR VPWR _5275_/X sky130_fd_sc_hd__mux2_1
Xoutput189 _3198_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[22] sky130_fd_sc_hd__buf_12
XFILLER_102_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4226_ _4226_/A0 _6353_/A1 _4230_/S VGND VGND VPWR VPWR _4226_/X sky130_fd_sc_hd__mux2_1
XFILLER_87_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7014_ _7083_/CLK _7014_/D fanout518/X VGND VGND VPWR VPWR _7014_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_68_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4157_ _6639_/Q _4181_/B VGND VGND VPWR VPWR _4165_/S sky130_fd_sc_hd__nand2_8
XFILLER_110_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4088_ hold173/X hold23/X _4092_/S VGND VGND VPWR VPWR _4088_/X sky130_fd_sc_hd__mux2_1
XFILLER_71_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6729_ _3939_/A1 _6729_/D _6381_/X VGND VGND VPWR VPWR _6729_/Q sky130_fd_sc_hd__dfrtn_1
XFILLER_137_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_149_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_52_csclk _7000_/CLK VGND VGND VPWR VPWR _6969_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_152_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_191_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_486 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_67_csclk _7000_/CLK VGND VGND VPWR VPWR _7056_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_59_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_407 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_159_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_174_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput14 mask_rev_in[19] VGND VGND VPWR VPWR input14/X sky130_fd_sc_hd__clkbuf_2
Xinput25 mask_rev_in[29] VGND VGND VPWR VPWR input25/X sky130_fd_sc_hd__clkbuf_1
XFILLER_174_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput36 mgmt_gpio_in[0] VGND VGND VPWR VPWR _3952_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_128_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_167_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput47 mgmt_gpio_in[1] VGND VGND VPWR VPWR input47/X sky130_fd_sc_hd__clkbuf_2
Xinput58 mgmt_gpio_in[2] VGND VGND VPWR VPWR _3247_/A sky130_fd_sc_hd__buf_12
XFILLER_10_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput69 mgmt_gpio_in[6] VGND VGND VPWR VPWR input69/X sky130_fd_sc_hd__clkbuf_1
XFILLER_183_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold809 _6452_/Q VGND VGND VPWR VPWR hold809/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_183_695 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_537 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3390_ _3706_/A _3390_/B VGND VGND VPWR VPWR _5253_/A sky130_fd_sc_hd__nor2_8
XFILLER_184_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5060_ _5019_/Y _5102_/A _5059_/X _5003_/X VGND VGND VPWR VPWR _6723_/D sky130_fd_sc_hd__a211o_1
XFILLER_28_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1509 hold14/A VGND VGND VPWR VPWR _3839_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_96_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4011_ hold811/X _6355_/A1 _4013_/S VGND VGND VPWR VPWR _4011_/X sky130_fd_sc_hd__mux2_1
XFILLER_96_178 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_234 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5962_ _5977_/A _5962_/B _5963_/C VGND VGND VPWR VPWR _5962_/X sky130_fd_sc_hd__and3_4
XFILLER_92_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4913_ _5010_/B _4913_/B _4913_/C _4913_/D VGND VGND VPWR VPWR _4914_/B sky130_fd_sc_hd__and4b_1
X_5893_ _7154_/Q _5614_/X _5914_/A2 hold65/A VGND VGND VPWR VPWR _5895_/A sky130_fd_sc_hd__a22o_1
XFILLER_61_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4844_ _4513_/A _4831_/X _4834_/X _4842_/X _4843_/X VGND VGND VPWR VPWR _4844_/X
+ sky130_fd_sc_hd__o2111a_1
XFILLER_60_292 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4775_ _4751_/Y _5074_/A _4902_/B _4775_/D VGND VGND VPWR VPWR _4775_/X sky130_fd_sc_hd__and4b_1
XFILLER_119_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6514_ _7069_/CLK _6514_/D fanout515/X VGND VGND VPWR VPWR _7180_/A sky130_fd_sc_hd__dfrtp_1
X_3726_ _3726_/A _3726_/B _3726_/C _3726_/D VGND VGND VPWR VPWR _3746_/B sky130_fd_sc_hd__nor4_1
XFILLER_107_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6445_ _7082_/CLK _6445_/D fanout519/X VGND VGND VPWR VPWR _6445_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_106_217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3657_ _6804_/Q _5226_/A _4231_/A _6632_/Q VGND VGND VPWR VPWR _3657_/X sky130_fd_sc_hd__a22o_1
XFILLER_173_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_164_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6376_ _6400_/A _6399_/B VGND VGND VPWR VPWR _6376_/X sky130_fd_sc_hd__and2_1
X_3588_ _3588_/A _3588_/B _3588_/C _3587_/Y VGND VGND VPWR VPWR _3625_/B sky130_fd_sc_hd__or4b_1
XFILLER_115_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5327_ hold996/X _5495_/A1 _5333_/S VGND VGND VPWR VPWR _5327_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_114_272 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5258_ _5258_/A0 _5465_/A1 _5261_/S VGND VGND VPWR VPWR _5258_/X sky130_fd_sc_hd__mux2_1
XFILLER_87_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4209_ _4209_/A0 _5308_/A1 _4213_/S VGND VGND VPWR VPWR _4209_/X sky130_fd_sc_hd__mux2_1
XFILLER_102_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5189_ hold895/X _5189_/A1 _5189_/S VGND VGND VPWR VPWR _5189_/X sky130_fd_sc_hd__mux2_1
XFILLER_113_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_113_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_189_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_132_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_164_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_180_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_120_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_370 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_188_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_92 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_128_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4560_ _4513_/A _4515_/B _4629_/B VGND VGND VPWR VPWR _4579_/A sky130_fd_sc_hd__a21o_1
XFILLER_155_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3511_ _3554_/A _3628_/B VGND VGND VPWR VPWR _4038_/A sky130_fd_sc_hd__nor2_8
Xhold606 _6581_/Q VGND VGND VPWR VPWR hold606/X sky130_fd_sc_hd__dlygate4sd3_1
X_4491_ _4943_/A _4586_/B VGND VGND VPWR VPWR _4514_/B sky130_fd_sc_hd__or2_1
Xhold617 _4324_/X VGND VGND VPWR VPWR _6717_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold628 _7049_/Q VGND VGND VPWR VPWR hold628/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_143_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6230_ _6230_/A1 _6305_/A2 _6228_/X _6229_/X VGND VGND VPWR VPWR _7128_/D sky130_fd_sc_hd__o22a_1
X_3442_ _6799_/Q _5217_/A hold41/A _6935_/Q VGND VGND VPWR VPWR _3442_/X sky130_fd_sc_hd__a22o_1
Xhold639 _4057_/X VGND VGND VPWR VPWR _6495_/D sky130_fd_sc_hd__dlygate4sd3_1
Xmax_cap369 hold40/X VGND VGND VPWR VPWR _3487_/A sky130_fd_sc_hd__buf_12
XTAP_900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6161_ _6889_/Q _6296_/A2 _6284_/B1 _6865_/Q VGND VGND VPWR VPWR _6161_/X sky130_fd_sc_hd__a22o_1
X_3373_ _7001_/Q _5442_/A _5190_/A input60/X VGND VGND VPWR VPWR _3373_/X sky130_fd_sc_hd__a22o_1
XTAP_911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5112_ _5112_/A _5112_/B _5112_/C VGND VGND VPWR VPWR _5112_/X sky130_fd_sc_hd__and3_1
XTAP_955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6092_ _6092_/A _6092_/B VGND VGND VPWR VPWR _6092_/Y sky130_fd_sc_hd__nor2_1
XTAP_966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_264 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1306 hold1306/A VGND VGND VPWR VPWR wb_dat_o[18] sky130_fd_sc_hd__buf_12
XTAP_988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1317 _4176_/A1 VGND VGND VPWR VPWR hold1317/X sky130_fd_sc_hd__dlygate4sd3_1
X_5043_ _5043_/A _5043_/B VGND VGND VPWR VPWR _5043_/X sky130_fd_sc_hd__and2_2
XTAP_999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1328 hold1328/A VGND VGND VPWR VPWR wb_dat_o[6] sky130_fd_sc_hd__buf_12
XFILLER_84_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1339 _4177_/A1 VGND VGND VPWR VPWR hold1339/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_93_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_0_wbbd_sck _7149_/Q VGND VGND VPWR VPWR clkbuf_0_wbbd_sck/X sky130_fd_sc_hd__clkbuf_16
X_6994_ _6994_/CLK _6994_/D fanout490/X VGND VGND VPWR VPWR _6994_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_80_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5945_ _5978_/B _5962_/B _5963_/C VGND VGND VPWR VPWR _5973_/A sky130_fd_sc_hd__and3_4
XFILLER_80_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5876_ _6601_/Q _5632_/X _5872_/X _5873_/X _5875_/X VGND VGND VPWR VPWR _5876_/X
+ sky130_fd_sc_hd__a2111o_2
XFILLER_178_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4827_ _4943_/B _4921_/A _4622_/A VGND VGND VPWR VPWR _4942_/C sky130_fd_sc_hd__a21o_1
XFILLER_21_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4758_ _4587_/A _4549_/B _4703_/Y VGND VGND VPWR VPWR _4763_/A sky130_fd_sc_hd__o21ba_1
XFILLER_147_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_153_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_193_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_515 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3709_ _6435_/Q _3984_/A _5253_/A _6827_/Q VGND VGND VPWR VPWR _3709_/X sky130_fd_sc_hd__a22o_1
XFILLER_134_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4689_ _5043_/A _4695_/B VGND VGND VPWR VPWR _4689_/Y sky130_fd_sc_hd__nor2_1
XFILLER_162_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6428_ _6994_/CLK _6428_/D fanout489/X VGND VGND VPWR VPWR _6428_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_122_507 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_570 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6359_ _6399_/A _6399_/B VGND VGND VPWR VPWR _6359_/X sky130_fd_sc_hd__and2_1
XFILLER_88_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_140_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_702 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_152_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_487 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold3 hold3/A VGND VGND VPWR VPWR hold3/X sky130_fd_sc_hd__buf_6
XFILLER_181_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3991_ hold267/X hold114/X _3992_/S VGND VGND VPWR VPWR _3991_/X sky130_fd_sc_hd__mux2_1
X_5730_ _7013_/Q _5921_/A2 _5729_/X VGND VGND VPWR VPWR _5730_/X sky130_fd_sc_hd__a21o_1
XFILLER_95_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_188_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5661_ _7002_/Q _5614_/X _5657_/X _5658_/X _5660_/X VGND VGND VPWR VPWR _5661_/X
+ sky130_fd_sc_hd__a2111o_1
XFILLER_30_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4612_ _4671_/B _4861_/B VGND VGND VPWR VPWR _4612_/X sky130_fd_sc_hd__or2_1
X_5592_ _7100_/Q _7099_/Q VGND VGND VPWR VPWR _5962_/B sky130_fd_sc_hd__and2_2
XFILLER_191_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4543_ _4394_/Y _5026_/A input99/X _4390_/A VGND VGND VPWR VPWR _4799_/A sky130_fd_sc_hd__o211ai_4
Xhold403 _6712_/Q VGND VGND VPWR VPWR hold403/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold414 _5150_/X VGND VGND VPWR VPWR _6741_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_128_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_144_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold425 _6940_/Q VGND VGND VPWR VPWR hold425/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold436 _5216_/X VGND VGND VPWR VPWR _6793_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4474_ _4977_/B _4692_/C VGND VGND VPWR VPWR _4556_/A sky130_fd_sc_hd__or2_1
Xhold447 _6864_/Q VGND VGND VPWR VPWR hold447/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold458 _4138_/X VGND VGND VPWR VPWR _6554_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_143_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold469 _6746_/Q VGND VGND VPWR VPWR hold469/X sky130_fd_sc_hd__dlygate4sd3_1
X_6213_ _6561_/Q _5969_/A _5973_/C _6620_/Q VGND VGND VPWR VPWR _6213_/X sky130_fd_sc_hd__a22o_1
XFILLER_143_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3425_ _6920_/Q _5352_/A _5244_/A _6824_/Q _3424_/X VGND VGND VPWR VPWR _3432_/B
+ sky130_fd_sc_hd__a221o_1
X_7193_ _7193_/A VGND VGND VPWR VPWR _7193_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_131_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3356_ _7009_/Q _5451_/A _3355_/Y input19/X VGND VGND VPWR VPWR _3356_/X sky130_fd_sc_hd__a22o_1
X_6144_ _6888_/Q _6296_/A2 _5946_/X _6840_/Q VGND VGND VPWR VPWR _6144_/X sky130_fd_sc_hd__a22o_1
XTAP_741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1103 _6550_/Q VGND VGND VPWR VPWR _4134_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_85_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1114 _4203_/X VGND VGND VPWR VPWR _6609_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3287_ hold50/X VGND VGND VPWR VPWR hold51/A sky130_fd_sc_hd__inv_2
X_6075_ _6965_/Q _5955_/X _6294_/A2 _7082_/Q _6074_/X VGND VGND VPWR VPWR _6075_/X
+ sky130_fd_sc_hd__a221o_1
Xhold1125 _6695_/Q VGND VGND VPWR VPWR _4298_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1136 _5209_/X VGND VGND VPWR VPWR _6786_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_100_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1147 _6735_/Q VGND VGND VPWR VPWR _5143_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_38_340 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5026_ _5026_/A _5026_/B VGND VGND VPWR VPWR _5027_/A sky130_fd_sc_hd__nand2_1
Xhold1158 _5516_/X VGND VGND VPWR VPWR _7059_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1169 _6675_/Q VGND VGND VPWR VPWR _4274_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_9 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6977_ _7080_/CLK _6977_/D fanout515/X VGND VGND VPWR VPWR _6977_/Q sky130_fd_sc_hd__dfrtp_1
X_5928_ _6582_/Q _5928_/A2 _5928_/B1 _6618_/Q VGND VGND VPWR VPWR _5928_/X sky130_fd_sc_hd__a22o_1
XFILLER_139_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5859_ _6466_/Q _5629_/X _5644_/X _6451_/Q _5858_/X VGND VGND VPWR VPWR _5864_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_186_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_135_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_182_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_356 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_624 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold970 _5522_/X VGND VGND VPWR VPWR _7064_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold981 _5354_/X VGND VGND VPWR VPWR _6915_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_122_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold992 _6843_/Q VGND VGND VPWR VPWR hold992/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_273 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_189_359 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_158_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_407 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_632 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_176_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3210_ _6877_/Q VGND VGND VPWR VPWR _3210_/Y sky130_fd_sc_hd__inv_2
XFILLER_113_359 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4190_ _4190_/A hold7/X VGND VGND VPWR VPWR _4195_/S sky130_fd_sc_hd__and2_4
XFILLER_79_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_140_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_192_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6900_ _7022_/CLK hold13/X fanout517/X VGND VGND VPWR VPWR _6900_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_48_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6831_ _7042_/CLK _6831_/D fanout523/X VGND VGND VPWR VPWR _6831_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_23_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6762_ _6976_/CLK _6762_/D fanout497/X VGND VGND VPWR VPWR _6762_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_62_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3974_ hold477/X _5519_/A1 _3974_/S VGND VGND VPWR VPWR _3974_/X sky130_fd_sc_hd__mux2_1
X_5713_ _5713_/A1 _6305_/A2 _5711_/X _5712_/X VGND VGND VPWR VPWR _7108_/D sky130_fd_sc_hd__o22a_1
X_6693_ _7067_/CLK _6693_/D _3264_/A VGND VGND VPWR VPWR _6693_/Q sky130_fd_sc_hd__dfrtp_4
X_5644_ _5667_/A _5645_/B _5648_/C VGND VGND VPWR VPWR _5644_/X sky130_fd_sc_hd__and3_4
XFILLER_176_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5575_ _5575_/A1 _5573_/B _5571_/Y _5574_/Y VGND VGND VPWR VPWR _7094_/D sky130_fd_sc_hd__a31o_1
Xhold200 _5176_/X VGND VGND VPWR VPWR _6760_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold211 _7045_/Q VGND VGND VPWR VPWR hold211/X sky130_fd_sc_hd__dlygate4sd3_1
X_4526_ _4922_/B _4526_/B _4526_/C _4898_/A VGND VGND VPWR VPWR _4526_/X sky130_fd_sc_hd__or4b_1
XFILLER_191_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold222 _4110_/X VGND VGND VPWR VPWR _6530_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold233 _6896_/Q VGND VGND VPWR VPWR hold233/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold244 _5185_/X VGND VGND VPWR VPWR _6766_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold255 _7080_/Q VGND VGND VPWR VPWR hold255/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_132_624 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold266 _4018_/X VGND VGND VPWR VPWR _6463_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4457_ _4554_/A _4691_/A _4570_/B VGND VGND VPWR VPWR _5025_/B sky130_fd_sc_hd__nor3_4
XFILLER_171_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold277 _7081_/Q VGND VGND VPWR VPWR hold277/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_49_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold288 _4055_/X VGND VGND VPWR VPWR _6494_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold299 _7155_/Q VGND VGND VPWR VPWR hold299/X sky130_fd_sc_hd__dlygate4sd3_1
X_3408_ _6840_/Q _5262_/A _3405_/X _3407_/X VGND VGND VPWR VPWR _3433_/B sky130_fd_sc_hd__a211o_1
XFILLER_132_679 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7176_ _7176_/A VGND VGND VPWR VPWR _7176_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_172_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4388_ _4545_/A _4530_/B VGND VGND VPWR VPWR _4403_/A sky130_fd_sc_hd__nand2_1
XFILLER_58_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6127_ _6127_/A _6127_/B _6127_/C _6004_/B VGND VGND VPWR VPWR _6127_/X sky130_fd_sc_hd__or4b_1
XTAP_571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3339_ _3706_/B _3554_/B VGND VGND VPWR VPWR _3339_/Y sky130_fd_sc_hd__nor2_8
XTAP_582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6058_ _6813_/Q _5936_/X _6289_/A2 _7074_/Q _6057_/X VGND VGND VPWR VPWR _6068_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_73_427 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5009_ _4692_/A _4495_/X _4597_/Y _4965_/B VGND VGND VPWR VPWR _5016_/C sky130_fd_sc_hd__o22a_1
XTAP_2405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_106 _7198_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_117 _3247_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_128 _3894_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_139 _5925_/B1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_726 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_610 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_654 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_146_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_711 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3690_ _6811_/Q _5235_/A _4008_/A _6456_/Q _3689_/X VGND VGND VPWR VPWR _3713_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_118_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5360_ hold443/X _5519_/A1 _5360_/S VGND VGND VPWR VPWR _5360_/X sky130_fd_sc_hd__mux2_1
Xoutput305 _3403_/X VGND VGND VPWR VPWR serial_data_2 sky130_fd_sc_hd__buf_12
XFILLER_58_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput316 hold1317/X VGND VGND VPWR VPWR hold1318/A sky130_fd_sc_hd__buf_12
XFILLER_5_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput327 hold1307/X VGND VGND VPWR VPWR hold1308/A sky130_fd_sc_hd__buf_12
XFILLER_126_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4311_ hold887/X _5189_/A1 _4314_/S VGND VGND VPWR VPWR _4311_/X sky130_fd_sc_hd__mux2_1
Xoutput338 hold1347/X VGND VGND VPWR VPWR hold1348/A sky130_fd_sc_hd__buf_12
XFILLER_126_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5291_ hold917/X _5531_/A1 _5297_/S VGND VGND VPWR VPWR _5291_/X sky130_fd_sc_hd__mux2_1
XFILLER_153_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7030_ _7083_/CLK _7030_/D fanout517/X VGND VGND VPWR VPWR _7030_/Q sky130_fd_sc_hd__dfrtp_1
X_4242_ hold385/X _5534_/A1 _4242_/S VGND VGND VPWR VPWR _4242_/X sky130_fd_sc_hd__mux2_1
XFILLER_113_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4173_ _3816_/X _4173_/A1 _4180_/S VGND VGND VPWR VPWR _6583_/D sky130_fd_sc_hd__mux2_1
XFILLER_95_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_622 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6814_ _6990_/CLK _6814_/D _6396_/A VGND VGND VPWR VPWR _6814_/Q sky130_fd_sc_hd__dfrtp_1
X_6745_ _6746_/CLK _6745_/D fanout488/X VGND VGND VPWR VPWR _6745_/Q sky130_fd_sc_hd__dfrtp_4
X_3957_ hold5/X _6351_/A2 _6624_/Q VGND VGND VPWR VPWR hold6/A sky130_fd_sc_hd__mux2_8
XFILLER_31_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6676_ _6769_/CLK _6676_/D fanout492/X VGND VGND VPWR VPWR _6676_/Q sky130_fd_sc_hd__dfrtp_4
X_3888_ _3886_/X _3887_/Y _6506_/Q _6763_/Q VGND VGND VPWR VPWR _6508_/D sky130_fd_sc_hd__a2bb2o_1
X_5627_ _5646_/A _5645_/B _5651_/B VGND VGND VPWR VPWR _5627_/X sky130_fd_sc_hd__and3b_4
X_5558_ _7088_/Q _7089_/Q _7090_/Q _5558_/D VGND VGND VPWR VPWR _5559_/A sky130_fd_sc_hd__and4_1
XFILLER_3_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4509_ _4692_/A _4943_/B _4549_/B _4495_/X VGND VGND VPWR VPWR _4510_/C sky130_fd_sc_hd__a31o_1
XFILLER_132_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5489_ hold943/X _6354_/A1 _5492_/S VGND VGND VPWR VPWR _5489_/X sky130_fd_sc_hd__mux2_1
Xfanout510 fanout526/X VGND VGND VPWR VPWR fanout510/X sky130_fd_sc_hd__buf_4
Xfanout521 fanout522/X VGND VGND VPWR VPWR fanout521/X sky130_fd_sc_hd__buf_8
X_7159_ _3939_/A1 _7159_/D _6389_/X VGND VGND VPWR VPWR _7159_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_58_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_318 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_186_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_128_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_182_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_135_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_151_752 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_544 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4860_ _4542_/A _5048_/A _5068_/A VGND VGND VPWR VPWR _5088_/C sky130_fd_sc_hd__a21oi_1
XTAP_2780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_154 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3811_ input20/X _3384_/Y _5487_/A _7034_/Q VGND VGND VPWR VPWR _3811_/X sky130_fd_sc_hd__a22o_1
XFILLER_60_463 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4791_ _4921_/A _4791_/B VGND VGND VPWR VPWR _4821_/C sky130_fd_sc_hd__or2_1
XANTENNA_17 _3361_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_28 _3461_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_39 _4255_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6530_ _7041_/CLK _6530_/D fanout519/X VGND VGND VPWR VPWR _6530_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_13_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3742_ _6867_/Q _5298_/A _4112_/B input47/X _3741_/X VGND VGND VPWR VPWR _3745_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_158_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_192_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_186_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6461_ _7038_/CLK _6461_/D fanout490/X VGND VGND VPWR VPWR _6461_/Q sky130_fd_sc_hd__dfrtp_2
X_3673_ _6744_/Q _5151_/A _3629_/Y _6765_/Q _3672_/X VGND VGND VPWR VPWR _3673_/Y
+ sky130_fd_sc_hd__a221oi_1
X_5412_ hold681/X _5544_/A1 _5414_/S VGND VGND VPWR VPWR _5412_/X sky130_fd_sc_hd__mux2_1
XFILLER_161_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6392_ _6396_/A _6396_/B VGND VGND VPWR VPWR _6392_/X sky130_fd_sc_hd__and2_1
XFILLER_161_527 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5343_ _5343_/A _5511_/B VGND VGND VPWR VPWR _5351_/S sky130_fd_sc_hd__and2_4
XFILLER_114_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput179 _3208_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[13] sky130_fd_sc_hd__buf_12
XFILLER_87_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5274_ hold311/X _5523_/A1 _5279_/S VGND VGND VPWR VPWR _5274_/X sky130_fd_sc_hd__mux2_1
XFILLER_114_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7013_ _7042_/CLK _7013_/D fanout520/X VGND VGND VPWR VPWR _7013_/Q sky130_fd_sc_hd__dfrtp_4
X_4225_ _4225_/A hold7/X VGND VGND VPWR VPWR _4230_/S sky130_fd_sc_hd__and2_4
X_4156_ hold885/X _4236_/A1 _4156_/S VGND VGND VPWR VPWR _4156_/X sky130_fd_sc_hd__mux2_1
XFILLER_56_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4087_ hold697/X _4086_/X _4095_/S VGND VGND VPWR VPWR _4087_/X sky130_fd_sc_hd__mux2_1
XFILLER_24_600 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4989_ _4748_/B _4719_/B _4725_/B _4972_/A VGND VGND VPWR VPWR _4989_/X sky130_fd_sc_hd__o22a_1
X_6728_ _3939_/A1 _6728_/D _6380_/X VGND VGND VPWR VPWR _6728_/Q sky130_fd_sc_hd__dfrtn_1
XFILLER_149_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6659_ _6699_/CLK _6659_/D fanout509/X VGND VGND VPWR VPWR _6659_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_109_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_192_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_192_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_191_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout351 _5612_/Y VGND VGND VPWR VPWR _6305_/A2 sky130_fd_sc_hd__buf_6
XFILLER_59_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput15 mask_rev_in[1] VGND VGND VPWR VPWR input15/X sky130_fd_sc_hd__clkbuf_1
Xinput26 mask_rev_in[2] VGND VGND VPWR VPWR input26/X sky130_fd_sc_hd__clkbuf_1
XFILLER_167_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_168_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput37 mgmt_gpio_in[10] VGND VGND VPWR VPWR input37/X sky130_fd_sc_hd__clkbuf_1
XFILLER_168_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput48 mgmt_gpio_in[20] VGND VGND VPWR VPWR input48/X sky130_fd_sc_hd__clkbuf_2
Xinput59 mgmt_gpio_in[30] VGND VGND VPWR VPWR input59/X sky130_fd_sc_hd__clkbuf_4
XFILLER_116_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_184_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_413 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4010_ hold565/X _4299_/A1 _4013_/S VGND VGND VPWR VPWR _4010_/X sky130_fd_sc_hd__mux2_1
XFILLER_84_319 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5961_ _5976_/A _5965_/B VGND VGND VPWR VPWR _5975_/A sky130_fd_sc_hd__nor2_4
XFILLER_80_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4912_ _4912_/A _4912_/B _4912_/C _5017_/D VGND VGND VPWR VPWR _4913_/D sky130_fd_sc_hd__and4_1
XFILLER_33_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5892_ _6602_/Q _5632_/X _5926_/B1 _6548_/Q _5890_/X VGND VGND VPWR VPWR _5892_/X
+ sky130_fd_sc_hd__a221o_1
X_4843_ _4586_/B _4831_/X _4585_/X _5017_/A VGND VGND VPWR VPWR _4843_/X sky130_fd_sc_hd__o211a_1
XFILLER_119_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4774_ _4774_/A _4774_/B _4774_/C _4774_/D VGND VGND VPWR VPWR _4775_/D sky130_fd_sc_hd__and4_1
XFILLER_193_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6513_ _7069_/CLK _6513_/D fanout515/X VGND VGND VPWR VPWR _7179_/A sky130_fd_sc_hd__dfrtp_1
XFILLER_193_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3725_ _6819_/Q _5244_/A _4096_/A input62/X _3724_/X VGND VGND VPWR VPWR _3726_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_119_546 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6444_ _7082_/CLK _6444_/D fanout519/X VGND VGND VPWR VPWR _6444_/Q sky130_fd_sc_hd__dfrtp_4
X_3656_ _6717_/Q _4321_/A _5145_/A _6739_/Q _3655_/X VGND VGND VPWR VPWR _3661_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_146_387 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6375_ _6399_/A _6401_/B VGND VGND VPWR VPWR _6375_/X sky130_fd_sc_hd__and2_1
X_3587_ _6805_/Q _5226_/A _4139_/A _6558_/Q _3586_/X VGND VGND VPWR VPWR _3587_/Y
+ sky130_fd_sc_hd__a221oi_1
X_5326_ _5326_/A0 _5530_/A1 _5333_/S VGND VGND VPWR VPWR _5326_/X sky130_fd_sc_hd__mux2_1
XFILLER_114_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5257_ hold305/X _5515_/A1 _5261_/S VGND VGND VPWR VPWR _5257_/X sky130_fd_sc_hd__mux2_1
XFILLER_88_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4208_ _4208_/A hold7/X VGND VGND VPWR VPWR _4213_/S sky130_fd_sc_hd__and2_2
XFILLER_180_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5188_ _5188_/A0 _5308_/A1 _5189_/S VGND VGND VPWR VPWR _5188_/X sky130_fd_sc_hd__mux2_1
XFILLER_29_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4139_ _4139_/A hold7/X VGND VGND VPWR VPWR _4144_/S sky130_fd_sc_hd__and2_2
XFILLER_43_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_192_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_162 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_330 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_175_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_332 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3510_ _6798_/Q _5217_/A _4249_/A _6659_/Q _3508_/X VGND VGND VPWR VPWR _3518_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_7_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4490_ _4495_/A _4490_/B VGND VGND VPWR VPWR _4586_/B sky130_fd_sc_hd__or2_4
Xhold607 _4170_/X VGND VGND VPWR VPWR _6581_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_155_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold618 _6652_/Q VGND VGND VPWR VPWR hold618/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold629 _5505_/X VGND VGND VPWR VPWR _7049_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3441_ _3761_/A _5161_/B VGND VGND VPWR VPWR _4096_/A sky130_fd_sc_hd__nor2_8
XFILLER_6_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_171_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6160_ _7033_/Q _5947_/Y _6296_/B1 _6905_/Q _6159_/X VGND VGND VPWR VPWR _6168_/B
+ sky130_fd_sc_hd__a221o_1
XTAP_901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3372_ _3797_/A _3761_/A VGND VGND VPWR VPWR _5190_/A sky130_fd_sc_hd__nor2_8
XTAP_912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5111_ _4594_/X _4615_/B _4936_/X _5110_/X VGND VGND VPWR VPWR _5131_/C sky130_fd_sc_hd__o211ai_4
XTAP_934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6091_ _7059_/Q _5972_/B _6284_/B1 _6862_/Q _6090_/X VGND VGND VPWR VPWR _6092_/B
+ sky130_fd_sc_hd__a221o_1
XTAP_956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1307 hold1393/X VGND VGND VPWR VPWR hold1307/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_69_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_628 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1318 hold1318/A VGND VGND VPWR VPWR wb_dat_o[11] sky130_fd_sc_hd__buf_12
X_5042_ _4707_/B _5041_/Y _4971_/C VGND VGND VPWR VPWR _5058_/B sky130_fd_sc_hd__a21o_1
XTAP_989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_511 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1329 _4179_/A1 VGND VGND VPWR VPWR hold1329/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_38_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6993_ _7029_/CLK hold36/X fanout519/X VGND VGND VPWR VPWR _6993_/Q sky130_fd_sc_hd__dfrtp_4
Xclkbuf_leaf_51_csclk clkbuf_opt_4_0_csclk/X VGND VGND VPWR VPWR _7078_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_80_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5944_ _5979_/B _5962_/B _5963_/C VGND VGND VPWR VPWR _5972_/A sky130_fd_sc_hd__and3_4
XFILLER_80_399 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5875_ _6472_/Q _5622_/X _5642_/X _6462_/Q _5874_/X VGND VGND VPWR VPWR _5875_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_33_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4826_ _4455_/Y _4566_/B _4574_/A VGND VGND VPWR VPWR _4839_/B sky130_fd_sc_hd__o21ai_1
Xclkbuf_leaf_66_csclk _7000_/CLK VGND VGND VPWR VPWR _6984_/CLK sky130_fd_sc_hd__clkbuf_16
X_4757_ _4549_/B _4495_/X _4717_/B _4394_/Y VGND VGND VPWR VPWR _4766_/B sky130_fd_sc_hd__o22a_1
X_3708_ _7040_/Q _5493_/A _4237_/A _6646_/Q _3707_/X VGND VGND VPWR VPWR _3711_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_107_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_527 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4688_ _4901_/B _4719_/B VGND VGND VPWR VPWR _4720_/A sky130_fd_sc_hd__nor2_1
X_6427_ _7034_/CLK _6427_/D fanout489/X VGND VGND VPWR VPWR _6427_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_161_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3639_ _6996_/Q _5442_/A _5179_/B _6759_/Q VGND VGND VPWR VPWR _3639_/X sky130_fd_sc_hd__a22o_1
XFILLER_122_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6358_ _6400_/A _6399_/B VGND VGND VPWR VPWR _6358_/X sky130_fd_sc_hd__and2_1
XFILLER_161_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_582 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5309_ hold973/X _5531_/A1 _5315_/S VGND VGND VPWR VPWR _5309_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_130_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6289_ _6674_/Q _6289_/A2 _5957_/X _6709_/Q _6288_/X VGND VGND VPWR VPWR _6292_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_76_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_19_csclk clkbuf_3_5_0_csclk/X VGND VGND VPWR VPWR _6998_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_140_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_714 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_138_630 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_652 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_313 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold4 hold4/A VGND VGND VPWR VPWR hold4/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_66_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_171 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3990_ _3990_/A0 hold142/X _3992_/S VGND VGND VPWR VPWR _3990_/X sky130_fd_sc_hd__mux2_1
XFILLER_22_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_148_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5660_ _6970_/Q _5644_/X _5649_/X _6930_/Q _5659_/X VGND VGND VPWR VPWR _5660_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_88_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4611_ _4678_/A _4962_/C VGND VGND VPWR VPWR _4861_/B sky130_fd_sc_hd__or2_4
X_5591_ _5591_/A1 _5593_/A _5590_/Y VGND VGND VPWR VPWR _7099_/D sky130_fd_sc_hd__a21oi_1
XFILLER_129_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4542_ _4542_/A _4613_/C _4542_/C VGND VGND VPWR VPWR _4634_/A sky130_fd_sc_hd__and3_1
XFILLER_129_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold404 _4318_/X VGND VGND VPWR VPWR _6712_/D sky130_fd_sc_hd__dlygate4sd3_1
Xwire390 _5975_/A VGND VGND VPWR VPWR wire390/X sky130_fd_sc_hd__buf_8
XFILLER_143_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold415 _6657_/Q VGND VGND VPWR VPWR hold415/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold426 _5382_/X VGND VGND VPWR VPWR _6940_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_144_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4473_ _4554_/A _4691_/A _4448_/A VGND VGND VPWR VPWR _4965_/B sky130_fd_sc_hd__or3b_4
Xhold437 _6422_/Q VGND VGND VPWR VPWR hold437/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold448 _5296_/X VGND VGND VPWR VPWR _6864_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6212_ _7035_/Q _6295_/A2 _5943_/Y _6461_/Q _6211_/X VGND VGND VPWR VPWR _6218_/C
+ sky130_fd_sc_hd__a221o_1
Xhold459 _6709_/Q VGND VGND VPWR VPWR hold459/X sky130_fd_sc_hd__dlygate4sd3_1
X_3424_ _6896_/Q _5325_/A _5520_/A _7069_/Q VGND VGND VPWR VPWR _3424_/X sky130_fd_sc_hd__a22o_1
X_7192_ _7192_/A VGND VGND VPWR VPWR _7192_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_98_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_131_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6143_ _6143_/A _6143_/B _6143_/C _6142_/Y VGND VGND VPWR VPWR _6143_/X sky130_fd_sc_hd__or4b_2
XTAP_731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3355_ _5168_/A _3538_/B VGND VGND VPWR VPWR _3355_/Y sky130_fd_sc_hd__nor2_8
XTAP_742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1104 _4134_/X VGND VGND VPWR VPWR _6550_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_100_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6074_ _6957_/Q _5957_/X _5978_/X _6949_/Q VGND VGND VPWR VPWR _6074_/X sky130_fd_sc_hd__a22o_1
XTAP_786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3286_ hold49/X _3286_/A1 _6624_/Q VGND VGND VPWR VPWR hold50/A sky130_fd_sc_hd__mux2_2
Xhold1115 _7083_/Q VGND VGND VPWR VPWR _5543_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1126 _4298_/X VGND VGND VPWR VPWR _6695_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1137 _6898_/Q VGND VGND VPWR VPWR _5335_/A0 sky130_fd_sc_hd__dlygate4sd3_1
X_5025_ _5025_/A _5025_/B VGND VGND VPWR VPWR _5025_/Y sky130_fd_sc_hd__nor2_2
Xhold1148 _5143_/X VGND VGND VPWR VPWR _6735_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_85_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1159 _6926_/Q VGND VGND VPWR VPWR _5366_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_38_352 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6976_ _6976_/CLK _6976_/D fanout501/X VGND VGND VPWR VPWR _6976_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_80_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_159_9 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5927_ _6564_/Q _5927_/A2 _5646_/X _6484_/Q _5926_/X VGND VGND VPWR VPWR _5930_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_22_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5858_ _5667_/B _5857_/X _6620_/Q _5914_/A2 VGND VGND VPWR VPWR _5858_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_22_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4809_ _4921_/A _4788_/A _4636_/B _4665_/C VGND VGND VPWR VPWR _4812_/C sky130_fd_sc_hd__o31a_1
X_5789_ _6448_/Q _5917_/B1 _5786_/X _5788_/X VGND VGND VPWR VPWR _5789_/X sky130_fd_sc_hd__a211o_1
XFILLER_119_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_181_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_99 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold960 _4269_/X VGND VGND VPWR VPWR _6671_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_150_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold971 _7048_/Q VGND VGND VPWR VPWR hold971/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_135_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold982 _6995_/Q VGND VGND VPWR VPWR hold982/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold993 _5273_/X VGND VGND VPWR VPWR _6843_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_122_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_285 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_419 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_192_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_642 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6830_ _6988_/CLK _6830_/D _6396_/A VGND VGND VPWR VPWR _6830_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_62_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_163 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6761_ _6976_/CLK _6761_/D fanout497/X VGND VGND VPWR VPWR _6761_/Q sky130_fd_sc_hd__dfrtp_1
X_3973_ hold25/X hold96/X _6624_/Q VGND VGND VPWR VPWR hold97/A sky130_fd_sc_hd__mux2_2
X_5712_ _7107_/Q _5612_/A _5612_/B VGND VGND VPWR VPWR _5712_/X sky130_fd_sc_hd__o21a_1
X_6692_ _7067_/CLK _6692_/D _3264_/A VGND VGND VPWR VPWR _6692_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_176_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_176_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5643_ _5646_/A _5643_/B _5650_/B VGND VGND VPWR VPWR _5643_/X sky130_fd_sc_hd__and3b_4
XFILLER_148_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5574_ _5577_/B VGND VGND VPWR VPWR _5574_/Y sky130_fd_sc_hd__inv_2
Xhold201 _6792_/Q VGND VGND VPWR VPWR hold201/X sky130_fd_sc_hd__dlygate4sd3_1
X_4525_ _4525_/A _4732_/A _4525_/C _4523_/X VGND VGND VPWR VPWR _4526_/B sky130_fd_sc_hd__or4b_1
Xhold212 _5500_/X VGND VGND VPWR VPWR _7045_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold223 _7086_/Q VGND VGND VPWR VPWR hold223/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold234 _5332_/X VGND VGND VPWR VPWR _6896_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold245 _6633_/Q VGND VGND VPWR VPWR hold245/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold256 _5540_/X VGND VGND VPWR VPWR _7080_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4456_ _4884_/A _4947_/B VGND VGND VPWR VPWR _4456_/Y sky130_fd_sc_hd__nand2_2
Xhold267 _6440_/Q VGND VGND VPWR VPWR hold267/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_131_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold278 _5541_/X VGND VGND VPWR VPWR _7081_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3407_ _6440_/Q _3984_/A _5379_/A _6944_/Q _3406_/X VGND VGND VPWR VPWR _3407_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_131_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold289 _7191_/A VGND VGND VPWR VPWR hold289/X sky130_fd_sc_hd__dlygate4sd3_1
X_7175_ _7175_/A VGND VGND VPWR VPWR _7175_/X sky130_fd_sc_hd__clkbuf_1
X_4387_ _4545_/A _4564_/A _4564_/B VGND VGND VPWR VPWR _4574_/A sky130_fd_sc_hd__and3_2
XFILLER_86_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_723 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6126_ _7031_/Q _5947_/Y _6123_/X _6125_/X VGND VGND VPWR VPWR _6127_/C sky130_fd_sc_hd__a211o_1
XTAP_561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3338_ _3354_/A _3401_/B VGND VGND VPWR VPWR _3554_/B sky130_fd_sc_hd__or2_4
XFILLER_100_511 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6057_ _7066_/Q _6283_/A2 wire390/X _6853_/Q _6056_/X VGND VGND VPWR VPWR _6057_/X
+ sky130_fd_sc_hd__a221o_1
X_3269_ hold56/X hold29/X _3856_/S VGND VGND VPWR VPWR hold30/A sky130_fd_sc_hd__mux2_1
X_5008_ _5008_/A _5008_/B _5008_/C _5008_/D VGND VGND VPWR VPWR _5018_/A sky130_fd_sc_hd__and4_1
XFILLER_73_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_631 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_107 _7198_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_118 input50/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_129 _3894_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_121_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_164_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_152 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6959_ _6999_/CLK _6959_/D fanout523/X VGND VGND VPWR VPWR _6959_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_179_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_179_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_738 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_622 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_182_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_146_42 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_64 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_146_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold790 _4258_/X VGND VGND VPWR VPWR _6662_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_162_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_91_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1490 _7164_/Q VGND VGND VPWR VPWR _3252_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_55_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_163 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_2_0__f_mgmt_gpio_in[4] clkbuf_0_mgmt_gpio_in[4]/X VGND VGND VPWR VPWR _7171_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_158_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_158_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput306 _3934_/X VGND VGND VPWR VPWR serial_load sky130_fd_sc_hd__buf_12
Xoutput317 hold1339/X VGND VGND VPWR VPWR hold1340/A sky130_fd_sc_hd__buf_12
XFILLER_160_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4310_ _4310_/A0 _6353_/A1 _4314_/S VGND VGND VPWR VPWR _4310_/X sky130_fd_sc_hd__mux2_1
Xoutput328 hold1311/X VGND VGND VPWR VPWR hold1312/A sky130_fd_sc_hd__buf_12
XFILLER_114_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5290_ _5290_/A0 _5530_/A1 _5297_/S VGND VGND VPWR VPWR _5290_/X sky130_fd_sc_hd__mux2_1
Xoutput339 hold1341/X VGND VGND VPWR VPWR hold1342/A sky130_fd_sc_hd__buf_12
XFILLER_113_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4241_ hold485/X _5491_/A1 _4242_/S VGND VGND VPWR VPWR _4241_/X sky130_fd_sc_hd__mux2_1
XFILLER_114_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_179 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4172_ _6637_/Q _6308_/B VGND VGND VPWR VPWR _4180_/S sky130_fd_sc_hd__nand2_8
XFILLER_28_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_586 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6813_ _7054_/CLK _6813_/D fanout503/X VGND VGND VPWR VPWR _6813_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_51_634 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6744_ _6746_/CLK _6744_/D fanout484/X VGND VGND VPWR VPWR _6744_/Q sky130_fd_sc_hd__dfrtp_4
X_3956_ _6642_/Q _3956_/B VGND VGND VPWR VPWR _6639_/D sky130_fd_sc_hd__and2_1
X_6675_ _6711_/CLK _6675_/D fanout486/X VGND VGND VPWR VPWR _6675_/Q sky130_fd_sc_hd__dfrtp_4
X_3887_ _6507_/Q _3887_/B VGND VGND VPWR VPWR _3887_/Y sky130_fd_sc_hd__nand2_1
XFILLER_137_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5626_ _5667_/A _5643_/B _5648_/C VGND VGND VPWR VPWR _5626_/X sky130_fd_sc_hd__and3_4
XFILLER_176_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5557_ _5557_/A1 _5550_/Y _5555_/Y _5556_/X VGND VGND VPWR VPWR _7089_/D sky130_fd_sc_hd__a22o_1
XFILLER_117_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4508_ _4943_/A _4943_/B _4479_/A VGND VGND VPWR VPWR _4510_/B sky130_fd_sc_hd__a21o_1
XFILLER_117_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5488_ _5488_/A0 _5488_/A1 _5492_/S VGND VGND VPWR VPWR _5488_/X sky130_fd_sc_hd__mux2_1
XFILLER_104_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_9 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_444 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4439_ _4977_/B _4680_/A VGND VGND VPWR VPWR _4439_/Y sky130_fd_sc_hd__nor2_1
Xfanout500 fanout526/X VGND VGND VPWR VPWR fanout500/X sky130_fd_sc_hd__buf_8
XFILLER_160_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout511 fanout513/X VGND VGND VPWR VPWR _3264_/A sky130_fd_sc_hd__buf_8
XFILLER_59_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout522 fanout525/X VGND VGND VPWR VPWR fanout522/X sky130_fd_sc_hd__buf_4
X_7158_ _7171_/CLK _7158_/D _6388_/X VGND VGND VPWR VPWR _7158_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_76_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6109_ _6943_/Q _5942_/X _5981_/X _6935_/Q VGND VGND VPWR VPWR _6109_/X sky130_fd_sc_hd__a22o_1
X_7089_ _7131_/CLK _7089_/D fanout502/X VGND VGND VPWR VPWR _7089_/Q sky130_fd_sc_hd__dfrtp_2
XTAP_391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_236 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_186_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_179_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_488 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_211 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3810_ _7087_/Q _5179_/B _4261_/A _6665_/Q _3809_/X VGND VGND VPWR VPWR _3813_/A
+ sky130_fd_sc_hd__a221o_1
X_4790_ _4985_/A _4924_/B _4785_/B VGND VGND VPWR VPWR _4791_/B sky130_fd_sc_hd__or3b_1
XFILLER_32_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_18 _3984_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_158_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_29 _3461_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3741_ _6676_/Q _4273_/A _4151_/A _6566_/Q VGND VGND VPWR VPWR _3741_/X sky130_fd_sc_hd__a22o_1
XFILLER_13_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_192_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_374 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6460_ _7038_/CLK _6460_/D fanout490/X VGND VGND VPWR VPWR _6460_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_70_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3672_ _7049_/Q _5502_/A _4273_/A _6677_/Q VGND VGND VPWR VPWR _3672_/X sky130_fd_sc_hd__a22o_1
X_5411_ hold86/X hold23/X _5414_/S VGND VGND VPWR VPWR hold87/A sky130_fd_sc_hd__mux2_1
X_6391_ _6396_/A _6396_/B VGND VGND VPWR VPWR _6391_/X sky130_fd_sc_hd__and2_1
X_5342_ hold915/X _5537_/A1 _5342_/S VGND VGND VPWR VPWR _5342_/X sky130_fd_sc_hd__mux2_1
XFILLER_161_539 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_142_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5273_ hold992/X _5495_/A1 _5279_/S VGND VGND VPWR VPWR _5273_/X sky130_fd_sc_hd__mux2_1
XFILLER_99_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7012_ _7051_/CLK _7012_/D fanout514/X VGND VGND VPWR VPWR _7012_/Q sky130_fd_sc_hd__dfrtp_1
X_4224_ _6624_/Q _6306_/B _4221_/X _5040_/B _3168_/A VGND VGND VPWR VPWR _4224_/X
+ sky130_fd_sc_hd__a2111o_1
X_4155_ hold646/X _4289_/A1 _4156_/S VGND VGND VPWR VPWR _4155_/X sky130_fd_sc_hd__mux2_1
XFILLER_28_406 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4086_ hold519/X _5515_/A1 _4092_/S VGND VGND VPWR VPWR _4086_/X sky130_fd_sc_hd__mux2_1
XFILLER_71_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_612 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_639 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4988_ _4988_/A _4988_/B VGND VGND VPWR VPWR _4999_/C sky130_fd_sc_hd__nor2_1
X_6727_ _3939_/A1 _6727_/D _6379_/X VGND VGND VPWR VPWR _6727_/Q sky130_fd_sc_hd__dfrtn_1
X_3939_ input83/X _3939_/A1 _6403_/Q VGND VGND VPWR VPWR _3939_/X sky130_fd_sc_hd__mux2_1
XFILLER_183_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6658_ _6683_/CLK _6658_/D fanout509/X VGND VGND VPWR VPWR _6658_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_125_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5609_ _6507_/Q _5609_/B VGND VGND VPWR VPWR _5609_/Y sky130_fd_sc_hd__nor2_1
XFILLER_3_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6589_ _7137_/CLK _6589_/D VGND VGND VPWR VPWR _6589_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_124_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_105_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_263 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_328 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_32 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_718 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput16 mask_rev_in[20] VGND VGND VPWR VPWR input16/X sky130_fd_sc_hd__buf_2
Xinput27 mask_rev_in[30] VGND VGND VPWR VPWR input27/X sky130_fd_sc_hd__clkbuf_1
Xinput38 mgmt_gpio_in[11] VGND VGND VPWR VPWR input38/X sky130_fd_sc_hd__clkbuf_4
Xinput49 mgmt_gpio_in[21] VGND VGND VPWR VPWR input49/X sky130_fd_sc_hd__clkbuf_1
XFILLER_128_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_143_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_151_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_425 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_296 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5960_ _5968_/A _5979_/A _5977_/A VGND VGND VPWR VPWR _5972_/C sky130_fd_sc_hd__and3_1
XFILLER_53_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4911_ _4911_/A _4911_/B _4911_/C VGND VGND VPWR VPWR _5017_/D sky130_fd_sc_hd__nor3_2
X_5891_ _3205_/Y _5923_/B _5667_/B VGND VGND VPWR VPWR _5891_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_45_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4842_ _4495_/X _4831_/X _5132_/C _4840_/X _4841_/X VGND VGND VPWR VPWR _4842_/X
+ sky130_fd_sc_hd__o2111a_1
XFILLER_20_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4773_ _5043_/A _4901_/B _4899_/B VGND VGND VPWR VPWR _4774_/D sky130_fd_sc_hd__a21o_1
XFILLER_165_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3724_ _6995_/Q _5442_/A _5163_/A _6752_/Q VGND VGND VPWR VPWR _3724_/X sky130_fd_sc_hd__a22o_1
X_6512_ _7060_/CLK _6512_/D fanout521/X VGND VGND VPWR VPWR _6512_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_174_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6443_ _7046_/CLK _6443_/D fanout500/X VGND VGND VPWR VPWR _6443_/Q sky130_fd_sc_hd__dfstp_1
X_3655_ input37/X _4092_/S _5388_/A _6948_/Q VGND VGND VPWR VPWR _3655_/X sky130_fd_sc_hd__a22o_1
XFILLER_146_399 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6374_ _6400_/A _6399_/B VGND VGND VPWR VPWR _6374_/X sky130_fd_sc_hd__and2_1
X_3586_ _6813_/Q _5235_/A _4151_/A _6568_/Q VGND VGND VPWR VPWR _3586_/X sky130_fd_sc_hd__a22o_1
X_5325_ _5325_/A _5529_/B VGND VGND VPWR VPWR _5333_/S sky130_fd_sc_hd__and2_4
XFILLER_130_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_142_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5256_ hold325/X _5541_/A1 _5261_/S VGND VGND VPWR VPWR _5256_/X sky130_fd_sc_hd__mux2_1
X_4207_ hold907/X _4236_/A1 _4207_/S VGND VGND VPWR VPWR _4207_/X sky130_fd_sc_hd__mux2_1
XFILLER_87_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5187_ _5187_/A _5187_/B VGND VGND VPWR VPWR _5189_/S sky130_fd_sc_hd__and2_1
XFILLER_29_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4138_ hold457/X _6357_/A1 _4138_/S VGND VGND VPWR VPWR _4138_/X sky130_fd_sc_hd__mux2_1
XFILLER_113_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4069_ hold180/X _5533_/A1 _4077_/S VGND VGND VPWR VPWR _4069_/X sky130_fd_sc_hd__mux2_1
XFILLER_56_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_169_436 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_149_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_152_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_192_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_174 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_180_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_120_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_342 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_344 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold608 _7069_/Q VGND VGND VPWR VPWR hold608/X sky130_fd_sc_hd__dlygate4sd3_1
X_3440_ _3440_/A _3440_/B VGND VGND VPWR VPWR _5161_/B sky130_fd_sc_hd__or2_4
Xhold619 _4246_/X VGND VGND VPWR VPWR _6652_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_171_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3371_ _3554_/A _3487_/A VGND VGND VPWR VPWR _5442_/A sky130_fd_sc_hd__nor2_8
XFILLER_112_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5110_ _5110_/A _5110_/B _5110_/C VGND VGND VPWR VPWR _5110_/X sky130_fd_sc_hd__and3_1
XTAP_924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6090_ _6806_/Q _5973_/B _6285_/A2 _6894_/Q VGND VGND VPWR VPWR _6090_/X sky130_fd_sc_hd__a22o_1
XTAP_946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5041_ _5043_/B _4672_/B _4686_/B _5021_/B VGND VGND VPWR VPWR _5041_/Y sky130_fd_sc_hd__o211ai_1
XTAP_979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1308 hold1308/A VGND VGND VPWR VPWR wb_dat_o[21] sky130_fd_sc_hd__buf_12
Xhold1319 _4189_/A1 VGND VGND VPWR VPWR hold1319/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_38_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_0_wb_clk_i wb_clk_i VGND VGND VPWR VPWR clkbuf_0_wb_clk_i/X sky130_fd_sc_hd__clkbuf_16
XFILLER_93_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6992_ _7029_/CLK _6992_/D fanout523/X VGND VGND VPWR VPWR _6992_/Q sky130_fd_sc_hd__dfrtp_4
X_5943_ _5976_/A _5953_/B VGND VGND VPWR VPWR _5943_/Y sky130_fd_sc_hd__nor2_8
XFILLER_53_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5874_ _6482_/Q _5646_/X _5919_/B1 _6632_/Q VGND VGND VPWR VPWR _5874_/X sky130_fd_sc_hd__a22o_1
XFILLER_139_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4825_ _4946_/A _4944_/A _4946_/C VGND VGND VPWR VPWR _5089_/A sky130_fd_sc_hd__nand3_1
XFILLER_193_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_193_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4756_ _4965_/A _4695_/B _4520_/X VGND VGND VPWR VPWR _4774_/B sky130_fd_sc_hd__o21a_1
X_3707_ _6947_/Q _5388_/A _5142_/A _6736_/Q VGND VGND VPWR VPWR _3707_/X sky130_fd_sc_hd__a22o_1
XFILLER_146_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4687_ _4692_/C _4687_/B VGND VGND VPWR VPWR _5081_/A sky130_fd_sc_hd__or2_1
XFILLER_162_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_19 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_539 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6426_ _7034_/CLK _6426_/D fanout489/X VGND VGND VPWR VPWR _6426_/Q sky130_fd_sc_hd__dfstp_1
X_3638_ _6812_/Q _5235_/A _4196_/A _6606_/Q VGND VGND VPWR VPWR _3638_/X sky130_fd_sc_hd__a22o_1
XFILLER_162_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3569_ _3568_/X _6731_/Q _3749_/S VGND VGND VPWR VPWR _6731_/D sky130_fd_sc_hd__mux2_1
X_6357_ hold299/X _6357_/A1 hold54/X VGND VGND VPWR VPWR _6357_/X sky130_fd_sc_hd__mux2_1
XFILLER_115_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5308_ _5308_/A0 _5308_/A1 _5315_/S VGND VGND VPWR VPWR _5308_/X sky130_fd_sc_hd__mux2_1
XFILLER_88_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6288_ _6659_/Q _6288_/A2 _5969_/A _6564_/Q VGND VGND VPWR VPWR _6288_/X sky130_fd_sc_hd__a22o_1
XFILLER_48_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5239_ hold193/X _5533_/A1 _5243_/S VGND VGND VPWR VPWR _5239_/X sky130_fd_sc_hd__mux2_1
XFILLER_29_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_124_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_375 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_20 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_152_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_137_185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_140_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold5 hold5/A VGND VGND VPWR VPWR hold5/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_181_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_183 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_740 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4610_ _4678_/A _4701_/A VGND VGND VPWR VPWR _4745_/B sky130_fd_sc_hd__or2_4
XFILLER_175_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5590_ _7099_/Q _5571_/Y _5593_/A VGND VGND VPWR VPWR _5590_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_175_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4541_ _4542_/A _4541_/B _4541_/C VGND VGND VPWR VPWR _4544_/B sky130_fd_sc_hd__and3_1
XFILLER_191_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_174 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold405 _6608_/Q VGND VGND VPWR VPWR hold405/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold416 _4252_/X VGND VGND VPWR VPWR _6657_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_144_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4472_ _4472_/A _4561_/A VGND VGND VPWR VPWR _4515_/B sky130_fd_sc_hd__or2_4
Xhold427 _6872_/Q VGND VGND VPWR VPWR hold427/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_183_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold438 _3968_/X VGND VGND VPWR VPWR _6422_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_144_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold449 _6469_/Q VGND VGND VPWR VPWR hold449/X sky130_fd_sc_hd__dlygate4sd3_1
X_6211_ _6556_/Q _6259_/A2 _5963_/X _6566_/Q VGND VGND VPWR VPWR _6211_/X sky130_fd_sc_hd__a22o_1
X_3423_ _6816_/Q _5235_/A _5307_/A _6880_/Q _3422_/X VGND VGND VPWR VPWR _3432_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_89_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7191_ _7191_/A VGND VGND VPWR VPWR _7191_/X sky130_fd_sc_hd__clkbuf_1
XTAP_710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6142_ _6142_/A _6142_/B VGND VGND VPWR VPWR _6142_/Y sky130_fd_sc_hd__nor2_1
X_3354_ _3354_/A _3440_/B VGND VGND VPWR VPWR _3538_/B sky130_fd_sc_hd__or2_4
XTAP_721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6073_ _6821_/Q _5969_/A _6294_/B1 _7042_/Q VGND VGND VPWR VPWR _6073_/X sky130_fd_sc_hd__a22o_1
Xhold1105 _6480_/Q VGND VGND VPWR VPWR _4039_/A0 sky130_fd_sc_hd__dlygate4sd3_1
X_3285_ hold48/X hold37/X _3856_/S VGND VGND VPWR VPWR hold49/A sky130_fd_sc_hd__mux2_1
XTAP_776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1116 _5543_/X VGND VGND VPWR VPWR _7083_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5024_ _4479_/A _5026_/B _5023_/X _4836_/X VGND VGND VPWR VPWR _5038_/A sky130_fd_sc_hd__o211a_1
Xhold1127 _6950_/Q VGND VGND VPWR VPWR _5393_/A0 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1138 _5335_/X VGND VGND VPWR VPWR _6898_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1149 _6862_/Q VGND VGND VPWR VPWR _5294_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_1909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6975_ _6976_/CLK _6975_/D fanout497/X VGND VGND VPWR VPWR _6975_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5926_ _6554_/Q _5926_/A2 _5926_/B1 _6549_/Q VGND VGND VPWR VPWR _5926_/X sky130_fd_sc_hd__a22o_1
XFILLER_22_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_167_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5857_ _6656_/Q _5923_/B VGND VGND VPWR VPWR _5857_/X sky130_fd_sc_hd__and2b_1
XFILLER_70_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4808_ _4725_/B _4972_/A _4581_/X VGND VGND VPWR VPWR _4818_/C sky130_fd_sc_hd__o21a_1
XFILLER_186_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5788_ _6928_/Q _5633_/X _5646_/X _7000_/Q _5787_/X VGND VGND VPWR VPWR _5788_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_119_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4739_ _4739_/A VGND VGND VPWR VPWR _4739_/Y sky130_fd_sc_hd__inv_2
XFILLER_147_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6409_ _3500_/A1 _6409_/D _6365_/X VGND VGND VPWR VPWR hold37/A sky130_fd_sc_hd__dfrtp_1
Xhold950 _4305_/X VGND VGND VPWR VPWR _6701_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_1_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold961 _6579_/Q VGND VGND VPWR VPWR hold961/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold972 _5504_/X VGND VGND VPWR VPWR _7048_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold983 _5444_/X VGND VGND VPWR VPWR _6995_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_135_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold994 _6464_/Q VGND VGND VPWR VPWR hold994/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_103_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_448 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_640 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_676 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_100_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_678 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_50_csclk clkbuf_opt_1_0_csclk/X VGND VGND VPWR VPWR _7070_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_125_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_65_csclk clkbuf_3_2_0_csclk/X VGND VGND VPWR VPWR _7011_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_94_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_654 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6760_ _6789_/CLK _6760_/D fanout497/X VGND VGND VPWR VPWR _6760_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_62_175 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3972_ hold237/X hold114/X _3974_/S VGND VGND VPWR VPWR _3972_/X sky130_fd_sc_hd__mux2_1
XFILLER_62_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5711_ _6788_/Q _5667_/X _5703_/X _5710_/X _5610_/A VGND VGND VPWR VPWR _5711_/X
+ sky130_fd_sc_hd__o221a_2
X_6691_ _7067_/CLK _6691_/D _3264_/A VGND VGND VPWR VPWR _6691_/Q sky130_fd_sc_hd__dfrtp_4
X_5642_ _5667_/A _5643_/B _5646_/B VGND VGND VPWR VPWR _5642_/X sky130_fd_sc_hd__and3_4
XFILLER_176_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5573_ _7094_/Q _5573_/B VGND VGND VPWR VPWR _5577_/B sky130_fd_sc_hd__or2_1
XFILLER_129_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold202 _5215_/X VGND VGND VPWR VPWR _6792_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_144_431 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4524_ _5043_/A _4789_/B VGND VGND VPWR VPWR _4525_/C sky130_fd_sc_hd__nor2_1
XFILLER_191_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold213 _6944_/Q VGND VGND VPWR VPWR hold213/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold224 _5546_/X VGND VGND VPWR VPWR _7086_/D sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_18_csclk clkbuf_3_5_0_csclk/X VGND VGND VPWR VPWR _7059_/CLK sky130_fd_sc_hd__clkbuf_16
Xhold235 _7032_/Q VGND VGND VPWR VPWR hold235/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold246 _4235_/X VGND VGND VPWR VPWR _6633_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4455_ _5021_/A VGND VGND VPWR VPWR _4455_/Y sky130_fd_sc_hd__inv_2
Xhold257 _6984_/Q VGND VGND VPWR VPWR hold257/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold268 _3991_/X VGND VGND VPWR VPWR _6440_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold279 _6444_/Q VGND VGND VPWR VPWR hold279/X sky130_fd_sc_hd__dlygate4sd3_1
X_3406_ _7045_/Q _5493_/A _5538_/A _7085_/Q VGND VGND VPWR VPWR _3406_/X sky130_fd_sc_hd__a22o_1
X_7174_ _7174_/A VGND VGND VPWR VPWR _7174_/X sky130_fd_sc_hd__clkbuf_1
X_4386_ _4564_/A _4564_/B VGND VGND VPWR VPWR _4530_/B sky130_fd_sc_hd__and2_1
XFILLER_131_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3337_ _5168_/A _3761_/B VGND VGND VPWR VPWR _3958_/A sky130_fd_sc_hd__nor2_8
X_6125_ _6959_/Q _5957_/X _6284_/B1 _6863_/Q _6124_/X VGND VGND VPWR VPWR _6125_/X
+ sky130_fd_sc_hd__a221o_1
XTAP_551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_735 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3268_ hold106/X _6724_/Q _6624_/Q VGND VGND VPWR VPWR _3268_/X sky130_fd_sc_hd__mux2_8
X_6056_ _6981_/Q _6176_/A2 _6290_/A2 _7005_/Q VGND VGND VPWR VPWR _6056_/X sky130_fd_sc_hd__a22o_1
XFILLER_45_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5007_ _5007_/A _5007_/B _5007_/C VGND VGND VPWR VPWR _5073_/B sky130_fd_sc_hd__and3_1
XTAP_2407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3199_ _6957_/Q VGND VGND VPWR VPWR _3199_/Y sky130_fd_sc_hd__inv_2
XFILLER_54_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_108 _7198_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_119 input38/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_687 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6958_ _6988_/CLK _6958_/D fanout518/X VGND VGND VPWR VPWR _6958_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_41_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5909_ _6543_/Q _5667_/X _5902_/X _5908_/X _5610_/A VGND VGND VPWR VPWR _5909_/X
+ sky130_fd_sc_hd__o221a_2
X_6889_ _7058_/CLK hold85/X fanout524/X VGND VGND VPWR VPWR _6889_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_139_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_155_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_108_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_100_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_146_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_162_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold780 _5490_/X VGND VGND VPWR VPWR _7036_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold791 _6661_/Q VGND VGND VPWR VPWR hold791/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_150_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_459 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1480 hold88/A VGND VGND VPWR VPWR _3256_/A1 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1491 _7111_/Q VGND VGND VPWR VPWR _5779_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_17_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_189_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_187_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_173_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput307 _3933_/X VGND VGND VPWR VPWR serial_resetn sky130_fd_sc_hd__buf_12
Xoutput318 hold1321/X VGND VGND VPWR VPWR hold1322/A sky130_fd_sc_hd__buf_12
Xoutput329 hold1309/X VGND VGND VPWR VPWR hold1310/A sky130_fd_sc_hd__buf_12
XFILLER_114_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_99_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4240_ hold775/X _6355_/A1 _4242_/S VGND VGND VPWR VPWR _4240_/X sky130_fd_sc_hd__mux2_1
XFILLER_113_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4171_ hold543/X _6357_/A1 _4171_/S VGND VGND VPWR VPWR _4171_/X sky130_fd_sc_hd__mux2_1
XFILLER_67_212 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_96_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_598 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6812_ _6998_/CLK _6812_/D _3264_/A VGND VGND VPWR VPWR _6812_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_36_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_646 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6743_ _6746_/CLK _6743_/D fanout484/X VGND VGND VPWR VPWR _6743_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_189_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3955_ _6644_/Q _3956_/B VGND VGND VPWR VPWR _6636_/D sky130_fd_sc_hd__and2_1
XFILLER_189_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_370 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6674_ _6689_/CLK _6674_/D fanout510/X VGND VGND VPWR VPWR _6674_/Q sky130_fd_sc_hd__dfstp_1
X_3886_ _5968_/A _5981_/A _5979_/A VGND VGND VPWR VPWR _3886_/X sky130_fd_sc_hd__and3_1
X_5625_ _5646_/A _5646_/B _5649_/C VGND VGND VPWR VPWR _5625_/X sky130_fd_sc_hd__and3b_4
XFILLER_137_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5556_ _7088_/Q _7089_/Q _6509_/Q _6507_/Q _5612_/A VGND VGND VPWR VPWR _5556_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_145_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4507_ _4554_/A _4570_/B _4587_/A _4505_/X _4506_/X VGND VGND VPWR VPWR _4510_/A
+ sky130_fd_sc_hd__o311a_1
X_5487_ _5487_/A _6352_/B VGND VGND VPWR VPWR _5492_/S sky130_fd_sc_hd__and2_2
XFILLER_160_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4438_ _4613_/C _4630_/A _4592_/B VGND VGND VPWR VPWR _4680_/A sky130_fd_sc_hd__or3b_1
Xfanout501 fanout502/X VGND VGND VPWR VPWR fanout501/X sky130_fd_sc_hd__buf_8
XFILLER_132_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout512 fanout513/X VGND VGND VPWR VPWR _6396_/A sky130_fd_sc_hd__buf_6
Xfanout523 fanout524/X VGND VGND VPWR VPWR fanout523/X sky130_fd_sc_hd__buf_8
XFILLER_59_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7157_ _7157_/CLK _7157_/D _3264_/X VGND VGND VPWR VPWR _7157_/Q sky130_fd_sc_hd__dfstp_2
X_4369_ _4499_/B _4449_/C VGND VGND VPWR VPWR _4707_/B sky130_fd_sc_hd__nor2_8
XFILLER_59_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6108_ _6855_/Q wire390/X _6282_/B1 _6975_/Q _6107_/X VGND VGND VPWR VPWR _6118_/A
+ sky130_fd_sc_hd__a221o_1
XTAP_392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7088_ _7131_/CLK _7088_/D fanout502/X VGND VGND VPWR VPWR _7088_/Q sky130_fd_sc_hd__dfrtp_2
X_6039_ _7081_/Q _6294_/A2 _5975_/C _7049_/Q _6038_/X VGND VGND VPWR VPWR _6042_/A
+ sky130_fd_sc_hd__a221o_1
XTAP_2204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_148_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_186_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_128_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_191 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_19 _5388_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3740_ _6883_/Q hold83/A hold34/A _6987_/Q _3739_/X VGND VGND VPWR VPWR _3745_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_119_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3671_ _6972_/Q _5415_/A _4032_/A _6477_/Q _3631_/X VGND VGND VPWR VPWR _3674_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_158_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5410_ hold569/X _5515_/A1 _5414_/S VGND VGND VPWR VPWR _5410_/X sky130_fd_sc_hd__mux2_1
XFILLER_173_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6390_ _6396_/A _6396_/B VGND VGND VPWR VPWR _6390_/X sky130_fd_sc_hd__and2_1
XFILLER_126_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5341_ hold421/X _5545_/A1 _5342_/S VGND VGND VPWR VPWR _5341_/X sky130_fd_sc_hd__mux2_1
XFILLER_142_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5272_ _5272_/A0 _5521_/A1 _5279_/S VGND VGND VPWR VPWR _5272_/X sky130_fd_sc_hd__mux2_1
X_7011_ _7011_/CLK _7011_/D fanout500/X VGND VGND VPWR VPWR _7011_/Q sky130_fd_sc_hd__dfstp_1
X_4223_ _6640_/Q _4223_/B VGND VGND VPWR VPWR _5040_/B sky130_fd_sc_hd__nand2b_4
X_4154_ hold813/X _5505_/A1 _4156_/S VGND VGND VPWR VPWR _4154_/X sky130_fd_sc_hd__mux2_1
XFILLER_68_554 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4085_ hold481/X _4084_/X _4095_/S VGND VGND VPWR VPWR _4085_/X sky130_fd_sc_hd__mux2_1
XFILLER_55_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_207 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_624 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4987_ _4988_/A _4791_/B _4793_/Y VGND VGND VPWR VPWR _5062_/B sky130_fd_sc_hd__o21a_1
X_6726_ _7140_/CLK _6726_/D _4181_/B VGND VGND VPWR VPWR _6726_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_177_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3938_ _6404_/Q _3940_/B VGND VGND VPWR VPWR _3938_/Y sky130_fd_sc_hd__nor2_1
XFILLER_177_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_206 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6657_ _6699_/CLK _6657_/D fanout509/X VGND VGND VPWR VPWR _6657_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_177_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3869_ hold5/A _6402_/Q _6396_/B VGND VGND VPWR VPWR _3869_/X sky130_fd_sc_hd__o21a_1
XFILLER_176_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5608_ _5608_/A1 _5605_/B _5607_/X VGND VGND VPWR VPWR _7105_/D sky130_fd_sc_hd__a21o_1
X_6588_ _7137_/CLK _6588_/D VGND VGND VPWR VPWR _6588_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_191_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5539_ hold652/X hold588/X _5546_/S VGND VGND VPWR VPWR _5539_/X sky130_fd_sc_hd__mux2_1
XFILLER_105_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_132_286 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_44 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_568 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_443 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput17 mask_rev_in[21] VGND VGND VPWR VPWR input17/X sky130_fd_sc_hd__clkbuf_1
Xinput28 mask_rev_in[31] VGND VGND VPWR VPWR input28/X sky130_fd_sc_hd__clkbuf_2
XFILLER_168_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput39 mgmt_gpio_in[12] VGND VGND VPWR VPWR _3954_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_109_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_170_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_182_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_546 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_708 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4910_ _4430_/C _4892_/B _5073_/A _5100_/C _4741_/X VGND VGND VPWR VPWR _4913_/C
+ sky130_fd_sc_hd__o2111a_1
XFILLER_80_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_590 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5890_ _6473_/Q _5622_/X _5920_/A2 _6568_/Q VGND VGND VPWR VPWR _5890_/X sky130_fd_sc_hd__a22o_1
XFILLER_61_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4841_ _4479_/A _4831_/X _4836_/X _4506_/A _4933_/A VGND VGND VPWR VPWR _4841_/X
+ sky130_fd_sc_hd__o2111a_1
XTAP_2590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_487 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4772_ _4720_/A _4772_/B _4772_/C VGND VGND VPWR VPWR _4774_/C sky130_fd_sc_hd__and3b_1
XFILLER_20_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_159_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6511_ _7017_/CLK _6511_/D fanout515/X VGND VGND VPWR VPWR _6511_/Q sky130_fd_sc_hd__dfrtp_1
X_3723_ _6851_/Q _3374_/Y _4279_/A _6681_/Q _3722_/X VGND VGND VPWR VPWR _3726_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_158_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6442_ _7039_/CLK _6442_/D fanout498/X VGND VGND VPWR VPWR _6442_/Q sky130_fd_sc_hd__dfstp_1
X_3654_ input54/X _5190_/A _4127_/A _6547_/Q _3653_/X VGND VGND VPWR VPWR _3661_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_134_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_146_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6373_ _6399_/A _6399_/B VGND VGND VPWR VPWR _6373_/X sky130_fd_sc_hd__and2_1
Xclkbuf_3_0_0_wb_clk_i clkbuf_3_1_0_wb_clk_i/A VGND VGND VPWR VPWR _7123_/CLK sky130_fd_sc_hd__clkbuf_8
X_3585_ _6917_/Q _5352_/A _5244_/A _6821_/Q _3584_/X VGND VGND VPWR VPWR _3588_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_161_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_359 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5324_ _5324_/A0 hold27/X hold84/X VGND VGND VPWR VPWR hold85/A sky130_fd_sc_hd__mux2_1
XFILLER_114_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5255_ hold975/X _5495_/A1 _5261_/S VGND VGND VPWR VPWR _5255_/X sky130_fd_sc_hd__mux2_1
XFILLER_57_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4206_ _4206_/A0 hold46/X _4207_/S VGND VGND VPWR VPWR hold47/A sky130_fd_sc_hd__mux2_1
X_5186_ hold650/X hold588/X _5186_/S VGND VGND VPWR VPWR _5186_/X sky130_fd_sc_hd__mux2_1
XFILLER_56_502 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4137_ hold622/X _4289_/A1 _4138_/S VGND VGND VPWR VPWR _4137_/X sky130_fd_sc_hd__mux2_1
X_4068_ hold614/X _4067_/X _4078_/S VGND VGND VPWR VPWR _4068_/X sky130_fd_sc_hd__mux2_1
XFILLER_71_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6709_ _6718_/CLK _6709_/D fanout496/X VGND VGND VPWR VPWR _6709_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_184_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_164_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_164_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_192_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_118_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_164_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_152_348 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_668 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_568 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_398 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_187_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold609 _5527_/X VGND VGND VPWR VPWR _7069_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_128_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3370_ _6905_/Q _5334_/A _3356_/X _3362_/X _3369_/X VGND VGND VPWR VPWR _3396_/B
+ sky130_fd_sc_hd__a2111o_1
XTAP_903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5040_ _4960_/Y _5040_/B _5087_/B _5061_/C VGND VGND VPWR VPWR _5119_/A sky130_fd_sc_hd__and4b_1
XTAP_969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1309 hold1394/X VGND VGND VPWR VPWR hold1309/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_93_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6991_ _7029_/CLK _6991_/D fanout519/X VGND VGND VPWR VPWR _6991_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_93_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5942_ _5979_/B _5981_/B _5981_/C VGND VGND VPWR VPWR _5942_/X sky130_fd_sc_hd__and3_4
XFILLER_92_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5873_ _6567_/Q _5920_/A2 _5926_/B1 _6547_/Q VGND VGND VPWR VPWR _5873_/X sky130_fd_sc_hd__a22o_1
XFILLER_179_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4824_ _4915_/A _4823_/X _4915_/B VGND VGND VPWR VPWR _4881_/C sky130_fd_sc_hd__a21bo_1
XFILLER_138_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_159_470 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4755_ _4755_/A _4959_/C VGND VGND VPWR VPWR _5020_/A sky130_fd_sc_hd__nor2_1
X_3706_ _3706_/A _3706_/B VGND VGND VPWR VPWR _5142_/A sky130_fd_sc_hd__nor2_4
X_4686_ _4691_/C _4686_/B VGND VGND VPWR VPWR _4686_/X sky130_fd_sc_hd__or2_1
XFILLER_162_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_164 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6425_ _7073_/CLK _6425_/D fanout497/X VGND VGND VPWR VPWR _6425_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_161_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3637_ _6884_/Q hold83/A _5325_/A _6892_/Q VGND VGND VPWR VPWR _3637_/X sky130_fd_sc_hd__a22o_1
XFILLER_146_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6356_ _6356_/A0 hold46/X hold54/X VGND VGND VPWR VPWR hold55/A sky130_fd_sc_hd__mux2_1
X_3568_ _3627_/A1 _4186_/A0 _3685_/S VGND VGND VPWR VPWR _3568_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5307_ _5307_/A _5511_/B VGND VGND VPWR VPWR _5315_/S sky130_fd_sc_hd__and2_4
XFILLER_161_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6287_ _6694_/Q _5972_/B _5973_/B _6554_/Q _6286_/X VGND VGND VPWR VPWR _6293_/C
+ sky130_fd_sc_hd__a221o_1
X_3499_ _3557_/A _3554_/B VGND VGND VPWR VPWR _4255_/A sky130_fd_sc_hd__nor2_4
XFILLER_88_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5238_ hold381/X _5523_/A1 _5243_/S VGND VGND VPWR VPWR _5238_/X sky130_fd_sc_hd__mux2_1
XFILLER_69_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5169_ _5308_/A1 _5169_/A1 _5169_/S VGND VGND VPWR VPWR _5169_/X sky130_fd_sc_hd__mux2_1
XFILLER_56_343 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_387 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_32 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_149_21 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_130_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_137_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_180_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold6 hold6/A VGND VGND VPWR VPWR hold6/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_75_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_188_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_276 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_129_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4540_ _4793_/A _4623_/B VGND VGND VPWR VPWR _4540_/Y sky130_fd_sc_hd__nor2_1
XFILLER_128_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_143_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire392 _5956_/X VGND VGND VPWR VPWR _5973_/B sky130_fd_sc_hd__buf_12
Xhold406 _4201_/X VGND VGND VPWR VPWR _6608_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_128_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4471_ _4471_/A _4471_/B VGND VGND VPWR VPWR _4899_/B sky130_fd_sc_hd__or2_2
XFILLER_183_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold417 _6888_/Q VGND VGND VPWR VPWR hold417/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold428 _5305_/X VGND VGND VPWR VPWR _6872_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6210_ _6681_/Q _5949_/X _5973_/B _6551_/Q _6209_/X VGND VGND VPWR VPWR _6218_/B
+ sky130_fd_sc_hd__a221o_1
Xhold439 _7052_/Q VGND VGND VPWR VPWR hold439/X sky130_fd_sc_hd__dlygate4sd3_1
X_3422_ _6912_/Q _5343_/A _3419_/X _3421_/X VGND VGND VPWR VPWR _3422_/X sky130_fd_sc_hd__a211o_1
X_7190_ _7190_/A VGND VGND VPWR VPWR _7190_/X sky130_fd_sc_hd__clkbuf_1
XTAP_700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6141_ _6920_/Q _5937_/X _6285_/B1 _7016_/Q _6140_/X VGND VGND VPWR VPWR _6142_/B
+ sky130_fd_sc_hd__a221o_1
XTAP_711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_744 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3353_ hold73/X hold80/X VGND VGND VPWR VPWR _3440_/B sky130_fd_sc_hd__nand2b_1
XFILLER_112_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_243 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6072_ _7050_/Q _5975_/C _6290_/B1 _7021_/Q _6071_/X VGND VGND VPWR VPWR _6077_/B
+ sky130_fd_sc_hd__a221o_1
XTAP_766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3284_ hold38/X _4983_/A1 _6624_/Q VGND VGND VPWR VPWR hold39/A sky130_fd_sc_hd__mux2_2
XTAP_777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1106 _4039_/X VGND VGND VPWR VPWR _6480_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_97_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1117 _6450_/Q VGND VGND VPWR VPWR _4003_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_100_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5023_ _4549_/B _4640_/B _4495_/X VGND VGND VPWR VPWR _5023_/X sky130_fd_sc_hd__a21o_1
Xhold1128 _5393_/X VGND VGND VPWR VPWR _6950_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1139 _6858_/Q VGND VGND VPWR VPWR _5290_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_38_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6974_ _6990_/CLK _6974_/D fanout513/X VGND VGND VPWR VPWR _6974_/Q sky130_fd_sc_hd__dfrtp_2
X_5925_ _6669_/Q _5633_/X _5925_/B1 _6719_/Q _5924_/X VGND VGND VPWR VPWR _5930_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_179_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5856_ _6561_/Q _5636_/X _5919_/B1 _6631_/Q _5855_/X VGND VGND VPWR VPWR _5864_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_167_716 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4807_ _4640_/B _4588_/B _4671_/B _4687_/B VGND VGND VPWR VPWR _5108_/A sky130_fd_sc_hd__o22a_1
X_5787_ _6912_/Q _5628_/X _5927_/A2 _6824_/Q VGND VGND VPWR VPWR _5787_/X sky130_fd_sc_hd__a22o_1
XFILLER_119_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4738_ _4672_/X _5021_/C _4885_/A VGND VGND VPWR VPWR _4739_/A sky130_fd_sc_hd__a21oi_1
XFILLER_119_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_175 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_635 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_107_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4669_ _4644_/X _4666_/X _4915_/B VGND VGND VPWR VPWR _4669_/Y sky130_fd_sc_hd__a21boi_1
X_6408_ _3500_/A1 _6408_/D _6364_/X VGND VGND VPWR VPWR hold71/A sky130_fd_sc_hd__dfrtp_2
Xhold940 _5282_/X VGND VGND VPWR VPWR _6851_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold951 _6646_/Q VGND VGND VPWR VPWR hold951/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold962 _4168_/X VGND VGND VPWR VPWR _6579_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold973 _6875_/Q VGND VGND VPWR VPWR hold973/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold984 hold984/A VGND VGND VPWR VPWR hold984/X sky130_fd_sc_hd__dlygate4sd3_1
X_6339_ _6642_/Q _6339_/A2 _6339_/B1 _4222_/B _6338_/X VGND VGND VPWR VPWR _6339_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_89_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold995 _4019_/X VGND VGND VPWR VPWR _6464_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_49_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_652 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_688 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_552 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_138_462 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_134 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3971_ hold112/X _3971_/A1 _6624_/Q VGND VGND VPWR VPWR _3971_/X sky130_fd_sc_hd__mux2_8
XFILLER_62_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5710_ _6804_/Q _5926_/A2 _5704_/X _5707_/X _5709_/X VGND VGND VPWR VPWR _5710_/X
+ sky130_fd_sc_hd__a2111o_1
XFILLER_93_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6690_ _7067_/CLK _6690_/D _3264_/A VGND VGND VPWR VPWR _6690_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_188_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_149_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5641_ _3180_/Y _5923_/B _5667_/B VGND VGND VPWR VPWR _5641_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_191_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5572_ _5609_/B _5643_/B _5645_/B _5572_/B1 _5565_/X VGND VGND VPWR VPWR _7093_/D
+ sky130_fd_sc_hd__o32a_1
Xclkbuf_1_0_1_csclk clkbuf_1_0_1_csclk/A VGND VGND VPWR VPWR clkbuf_2_1_0_csclk/A
+ sky130_fd_sc_hd__clkbuf_8
X_4523_ _4523_/A _5074_/A _4523_/C _4523_/D VGND VGND VPWR VPWR _4523_/X sky130_fd_sc_hd__and4_1
XFILLER_116_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold203 _7053_/Q VGND VGND VPWR VPWR hold203/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold214 _5386_/X VGND VGND VPWR VPWR _6944_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_144_443 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold225 _6790_/Q VGND VGND VPWR VPWR hold225/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold236 _5485_/X VGND VGND VPWR VPWR _7032_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4454_ _4789_/A _4692_/C VGND VGND VPWR VPWR _5021_/A sky130_fd_sc_hd__or2_1
Xhold247 _6976_/Q VGND VGND VPWR VPWR hold247/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold258 _5431_/X VGND VGND VPWR VPWR _6984_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold269 _6432_/Q VGND VGND VPWR VPWR hold269/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3405_ _6808_/Q _5226_/A _5511_/A _7061_/Q VGND VGND VPWR VPWR _3405_/X sky130_fd_sc_hd__a22o_1
X_7173_ _7173_/A VGND VGND VPWR VPWR _7173_/X sky130_fd_sc_hd__clkbuf_1
X_4385_ _4436_/A _4541_/B _4541_/C VGND VGND VPWR VPWR _4564_/B sky130_fd_sc_hd__nand3_1
XTAP_530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6124_ _6807_/Q _5973_/B _6300_/B1 _6879_/Q VGND VGND VPWR VPWR _6124_/X sky130_fd_sc_hd__a22o_1
XTAP_541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3336_ _3366_/A _3401_/B VGND VGND VPWR VPWR _3761_/B sky130_fd_sc_hd__or2_4
XTAP_552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6055_ _6079_/A2 _6305_/A2 _6053_/X _6054_/X VGND VGND VPWR VPWR _7121_/D sky130_fd_sc_hd__o22a_1
XTAP_585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3267_ hold48/X hold105/X _3266_/Y VGND VGND VPWR VPWR _3267_/X sky130_fd_sc_hd__a21bo_1
XFILLER_100_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5006_ _4401_/X _4885_/B _5005_/X _4736_/X VGND VGND VPWR VPWR _5007_/C sky130_fd_sc_hd__o211a_1
X_3198_ _6965_/Q VGND VGND VPWR VPWR _3198_/Y sky130_fd_sc_hd__inv_2
XTAP_2408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_109 _3953_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_666 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6957_ _7082_/CLK _6957_/D fanout519/X VGND VGND VPWR VPWR _6957_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_54_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5908_ _6678_/Q _5649_/X _5903_/X _5905_/X _5907_/X VGND VGND VPWR VPWR _5908_/X
+ sky130_fd_sc_hd__a2111o_1
XFILLER_167_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6888_ _6999_/CLK _6888_/D fanout523/X VGND VGND VPWR VPWR _6888_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_179_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5839_ _7034_/Q _5645_/X _5648_/X _6715_/Q _5838_/X VGND VGND VPWR VPWR _5842_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_22_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_139_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_139_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_163_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold770 _4107_/X VGND VGND VPWR VPWR _6527_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold781 _6764_/Q VGND VGND VPWR VPWR hold781/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold792 _4257_/X VGND VGND VPWR VPWR _6661_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_39_20 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1470 _7171_/Q VGND VGND VPWR VPWR _3229_/A1 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1481 _7124_/Q VGND VGND VPWR VPWR _6154_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_29_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1492 _7122_/Q VGND VGND VPWR VPWR _6080_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_91_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_189_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_185_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_185_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput308 _3951_/X VGND VGND VPWR VPWR spi_sdi sky130_fd_sc_hd__buf_12
Xoutput319 hold1329/X VGND VGND VPWR VPWR hold1330/A sky130_fd_sc_hd__buf_12
XFILLER_4_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4170_ hold606/X _4289_/A1 _4171_/S VGND VGND VPWR VPWR _4170_/X sky130_fd_sc_hd__mux2_1
XFILLER_95_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6811_ _7046_/CLK _6811_/D fanout497/X VGND VGND VPWR VPWR _6811_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_23_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6742_ _6746_/CLK _6742_/D fanout484/X VGND VGND VPWR VPWR _6742_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_51_658 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3954_ _6769_/Q _3954_/B VGND VGND VPWR VPWR _3954_/X sky130_fd_sc_hd__and2_2
XFILLER_50_168 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6673_ _6708_/CLK _6673_/D _6400_/A VGND VGND VPWR VPWR _6673_/Q sky130_fd_sc_hd__dfstp_1
X_3885_ _7100_/Q _7099_/Q VGND VGND VPWR VPWR _5979_/A sky130_fd_sc_hd__and2b_4
XFILLER_31_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5624_ _5646_/A _5648_/C _5651_/C VGND VGND VPWR VPWR _5624_/X sky130_fd_sc_hd__and3b_4
XFILLER_31_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_136_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5555_ _7088_/Q _7089_/Q VGND VGND VPWR VPWR _5555_/Y sky130_fd_sc_hd__nand2_1
XFILLER_129_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4506_ _4506_/A _4506_/B _4506_/C VGND VGND VPWR VPWR _4506_/X sky130_fd_sc_hd__and3_1
XFILLER_144_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5486_ hold967/X _5537_/A1 _5486_/S VGND VGND VPWR VPWR _5486_/X sky130_fd_sc_hd__mux2_1
XFILLER_172_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_160_744 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4437_ _4617_/B _4888_/A VGND VGND VPWR VPWR _4592_/B sky130_fd_sc_hd__nor2_1
Xfanout502 fanout503/X VGND VGND VPWR VPWR fanout502/X sky130_fd_sc_hd__buf_8
Xfanout513 fanout526/X VGND VGND VPWR VPWR fanout513/X sky130_fd_sc_hd__buf_6
X_7156_ _7171_/CLK _7156_/D _6387_/X VGND VGND VPWR VPWR hold5/A sky130_fd_sc_hd__dfrtn_1
Xfanout524 fanout525/X VGND VGND VPWR VPWR fanout524/X sky130_fd_sc_hd__buf_8
X_4368_ _4368_/A _4544_/A VGND VGND VPWR VPWR _4449_/C sky130_fd_sc_hd__or2_2
XFILLER_86_511 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6107_ _6927_/Q _5977_/X _6290_/B1 _7023_/Q _6106_/X VGND VGND VPWR VPWR _6107_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_58_235 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3319_ _3328_/A hold60/X VGND VGND VPWR VPWR _3533_/A sky130_fd_sc_hd__or2_4
X_7087_ _7131_/CLK _7087_/D fanout501/X VGND VGND VPWR VPWR _7087_/Q sky130_fd_sc_hd__dfrtp_2
X_4299_ hold567/X _4299_/A1 _4302_/S VGND VGND VPWR VPWR _4299_/X sky130_fd_sc_hd__mux2_1
XTAP_393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_566 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6038_ _6836_/Q _5946_/X wire390/X _6852_/Q VGND VGND VPWR VPWR _6038_/X sky130_fd_sc_hd__a22o_1
XTAP_2205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_260 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_179 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_64_csclk clkbuf_3_2_0_csclk/X VGND VGND VPWR VPWR _7027_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_10_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_108_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_79_csclk _6661_/CLK VGND VGND VPWR VPWR _6697_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_2_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_17_csclk clkbuf_3_5_0_csclk/X VGND VGND VPWR VPWR _6988_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_2761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_186_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_158_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_158_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_186_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3670_ _6988_/Q hold34/A _6352_/A _7153_/Q _3630_/X VGND VGND VPWR VPWR _3674_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_9_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5340_ hold731/X _5457_/A1 _5342_/S VGND VGND VPWR VPWR _5340_/X sky130_fd_sc_hd__mux2_1
XFILLER_56_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5271_ _5271_/A _5511_/B VGND VGND VPWR VPWR _5279_/S sky130_fd_sc_hd__and2_4
XFILLER_99_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7010_ _7010_/CLK _7010_/D fanout498/X VGND VGND VPWR VPWR _7010_/Q sky130_fd_sc_hd__dfstp_1
X_4222_ _6640_/Q _4222_/B VGND VGND VPWR VPWR _4222_/X sky130_fd_sc_hd__and2b_4
XFILLER_68_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4153_ hold921/X _5189_/A1 _4156_/S VGND VGND VPWR VPWR _4153_/X sky130_fd_sc_hd__mux2_1
XFILLER_68_566 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_374 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4084_ hold369/X _5541_/A1 _4092_/S VGND VGND VPWR VPWR _4084_/X sky130_fd_sc_hd__mux2_1
XFILLER_55_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_411 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4986_ _4977_/B _4640_/X _4902_/B _5112_/A _5061_/D VGND VGND VPWR VPWR _5001_/A
+ sky130_fd_sc_hd__o2111a_1
X_3937_ input84/X _3263_/C _6404_/Q VGND VGND VPWR VPWR _3937_/X sky130_fd_sc_hd__mux2_2
XFILLER_51_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6725_ _7137_/CLK _6725_/D _4181_/B VGND VGND VPWR VPWR _6725_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_137_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6656_ _6696_/CLK _6656_/D fanout495/X VGND VGND VPWR VPWR _6656_/Q sky130_fd_sc_hd__dfrtp_1
X_3868_ _6485_/Q _3867_/A _3867_/Y _6487_/Q VGND VGND VPWR VPWR _6485_/D sky130_fd_sc_hd__a22o_1
XFILLER_176_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5607_ _7089_/Q _6509_/Q _5607_/C _7088_/Q VGND VGND VPWR VPWR _5607_/X sky130_fd_sc_hd__and4b_1
X_6587_ _7137_/CLK _6587_/D VGND VGND VPWR VPWR _6587_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_118_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3799_ _6954_/Q _5397_/A _4002_/A _6450_/Q _3798_/X VGND VGND VPWR VPWR _3802_/C
+ sky130_fd_sc_hd__a221o_1
X_5538_ _5538_/A _5538_/B VGND VGND VPWR VPWR _5546_/S sky130_fd_sc_hd__and2_4
XFILLER_11_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5469_ hold18/X _5538_/B VGND VGND VPWR VPWR hold19/A sky130_fd_sc_hd__and2_4
XFILLER_132_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7139_ _7140_/CLK _7139_/D VGND VGND VPWR VPWR _7139_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_47_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_187_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_455 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_42 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_168_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput18 mask_rev_in[22] VGND VGND VPWR VPWR input18/X sky130_fd_sc_hd__clkbuf_1
XFILLER_128_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput29 mask_rev_in[3] VGND VGND VPWR VPWR input29/X sky130_fd_sc_hd__clkbuf_1
XFILLER_182_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_240 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_151_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_184_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4840_ _4587_/A _4831_/X _4839_/X _5007_/A _4828_/X VGND VGND VPWR VPWR _4840_/X
+ sky130_fd_sc_hd__o2111a_1
XTAP_2580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4771_ _4549_/B _4515_/B _4717_/A _4717_/B _4770_/X VGND VGND VPWR VPWR _4772_/C
+ sky130_fd_sc_hd__o221a_1
XFILLER_159_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6510_ _7069_/CLK _6510_/D fanout515/X VGND VGND VPWR VPWR _6510_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_20_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3722_ _7072_/Q _5529_/A _5190_/A input53/X VGND VGND VPWR VPWR _3722_/X sky130_fd_sc_hd__a22o_1
XFILLER_119_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_159_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6441_ _7034_/CLK _6441_/D fanout488/X VGND VGND VPWR VPWR _6441_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_146_335 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3653_ _6980_/Q _5424_/A _5511_/A _7057_/Q VGND VGND VPWR VPWR _3653_/X sky130_fd_sc_hd__a22o_1
XFILLER_173_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6372_ _6399_/A _6399_/B VGND VGND VPWR VPWR _6372_/X sky130_fd_sc_hd__and2_1
XFILLER_115_711 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3584_ _7082_/Q _5538_/A _5502_/A _7050_/Q VGND VGND VPWR VPWR _3584_/X sky130_fd_sc_hd__a22o_1
X_5323_ hold417/X _5545_/A1 hold84/X VGND VGND VPWR VPWR _5323_/X sky130_fd_sc_hd__mux2_1
XFILLER_115_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5254_ _5254_/A0 _5488_/A1 _5261_/S VGND VGND VPWR VPWR _5254_/X sky130_fd_sc_hd__mux2_1
X_4205_ hold797/X _6355_/A1 _4207_/S VGND VGND VPWR VPWR _4205_/X sky130_fd_sc_hd__mux2_1
XFILLER_87_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5185_ hold243/X hold90/X _5186_/S VGND VGND VPWR VPWR _5185_/X sky130_fd_sc_hd__mux2_1
Xclkbuf_3_6_0_csclk clkbuf_3_7_0_csclk/A VGND VGND VPWR VPWR clkbuf_3_6_0_csclk/X
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_68_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4136_ hold821/X _5505_/A1 _4138_/S VGND VGND VPWR VPWR _4136_/X sky130_fd_sc_hd__mux2_1
XFILLER_68_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4067_ hold363/X _5532_/A1 _4077_/S VGND VGND VPWR VPWR _4067_/X sky130_fd_sc_hd__mux2_1
XFILLER_37_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_731 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4969_ _4977_/B _4965_/C _4671_/B _4679_/Y VGND VGND VPWR VPWR _5081_/C sky130_fd_sc_hd__o31a_1
XFILLER_149_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6708_ _6708_/CLK _6708_/D _6401_/A VGND VGND VPWR VPWR _6708_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_177_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6639_ _7150_/CLK _6639_/D _6308_/B VGND VGND VPWR VPWR _6639_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_98_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_187_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_458 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_143_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6990_ _6990_/CLK _6990_/D fanout513/X VGND VGND VPWR VPWR _6990_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_53_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5941_ _5980_/A _5953_/B VGND VGND VPWR VPWR _5941_/Y sky130_fd_sc_hd__nor2_8
XFILLER_34_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5872_ _5872_/A _5872_/B VGND VGND VPWR VPWR _5872_/X sky130_fd_sc_hd__or2_1
XFILLER_34_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4823_ _4977_/B _4692_/C _4962_/C _5100_/B _4822_/X VGND VGND VPWR VPWR _4823_/X
+ sky130_fd_sc_hd__o311a_1
XFILLER_21_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4754_ _4713_/A _4715_/B _4514_/B VGND VGND VPWR VPWR _5017_/C sky130_fd_sc_hd__o21a_1
XFILLER_159_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3705_ _6835_/Q _5262_/A _4026_/A _6471_/Q _3704_/X VGND VGND VPWR VPWR _3711_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_119_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4685_ _4884_/A _4619_/Y _4683_/Y _4684_/Y VGND VGND VPWR VPWR _5085_/A sky130_fd_sc_hd__a211o_1
XFILLER_174_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6424_ _7073_/CLK _6424_/D fanout497/X VGND VGND VPWR VPWR _6424_/Q sky130_fd_sc_hd__dfstp_2
X_3636_ _7012_/Q _5460_/A _4285_/A _6687_/Q VGND VGND VPWR VPWR _3636_/X sky130_fd_sc_hd__a22o_1
XFILLER_162_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_176 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6355_ hold863/X _6355_/A1 hold54/A VGND VGND VPWR VPWR _6355_/X sky130_fd_sc_hd__mux2_1
XFILLER_127_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_162_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3567_ _3567_/A _3567_/B _3567_/C VGND VGND VPWR VPWR _3567_/Y sky130_fd_sc_hd__nand3_2
XFILLER_108_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_703 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5306_ hold841/X _5537_/A1 _5306_/S VGND VGND VPWR VPWR _5306_/X sky130_fd_sc_hd__mux2_1
X_6286_ _6603_/Q _5939_/X _6286_/B1 _6474_/Q VGND VGND VPWR VPWR _6286_/X sky130_fd_sc_hd__a22o_1
X_3498_ _7075_/Q _5529_/A _3355_/Y input16/X _3497_/X VGND VGND VPWR VPWR _3502_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_130_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5237_ hold957/X _5495_/A1 _5243_/S VGND VGND VPWR VPWR _5237_/X sky130_fd_sc_hd__mux2_1
XFILLER_88_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5168_ _5168_/A _5183_/B _5187_/B VGND VGND VPWR VPWR _5169_/S sky130_fd_sc_hd__or3b_2
XFILLER_84_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4119_ hold271/X hold114/X _4120_/S VGND VGND VPWR VPWR _4119_/X sky130_fd_sc_hd__mux2_1
XFILLER_56_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5099_ _5102_/A _5079_/Y _5098_/X _5071_/X VGND VGND VPWR VPWR _6724_/D sky130_fd_sc_hd__a211o_1
XFILLER_83_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_314 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_140_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_68 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_44 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_149_33 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_149_99 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_180_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_180_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_133_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_181_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_181_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_94_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold7 hold7/A VGND VGND VPWR VPWR hold7/X sky130_fd_sc_hd__buf_8
XFILLER_75_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_129_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4470_ _4470_/A _4640_/B VGND VGND VPWR VPWR _4922_/B sky130_fd_sc_hd__nor2_1
Xhold407 hold407/A VGND VGND VPWR VPWR hold407/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_143_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold418 _5323_/X VGND VGND VPWR VPWR _6888_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3421_ _6424_/Q _3958_/A _5442_/A _7000_/Q _3420_/X VGND VGND VPWR VPWR _3421_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_99_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold429 _6765_/Q VGND VGND VPWR VPWR hold429/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_143_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_98_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_171_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6140_ _7061_/Q _5972_/B _6284_/B1 _6864_/Q VGND VGND VPWR VPWR _6140_/X sky130_fd_sc_hd__a22o_1
XFILLER_131_319 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3352_ hold33/X _3391_/B VGND VGND VPWR VPWR _5451_/A sky130_fd_sc_hd__nor2_8
XTAP_712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_112_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6071_ _7058_/Q _5972_/B _5973_/B _6805_/Q VGND VGND VPWR VPWR _6071_/X sky130_fd_sc_hd__a22o_1
XTAP_756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_255 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3283_ hold37/X hold71/A _3856_/S VGND VGND VPWR VPWR hold38/A sky130_fd_sc_hd__mux2_1
XTAP_767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1107 _6475_/Q VGND VGND VPWR VPWR _4033_/A0 sky130_fd_sc_hd__dlygate4sd3_1
X_5022_ _5022_/A _5022_/B VGND VGND VPWR VPWR _5089_/B sky130_fd_sc_hd__or2_1
XTAP_789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1118 _4003_/X VGND VGND VPWR VPWR _6450_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_112_599 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1129 _6982_/Q VGND VGND VPWR VPWR _5429_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_93_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6973_ _7082_/CLK _6973_/D fanout520/X VGND VGND VPWR VPWR _6973_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_53_347 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5924_ _5667_/B _5923_/X _6699_/Q _5924_/B2 VGND VGND VPWR VPWR _5924_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_179_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_166 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5855_ _6556_/Q _5627_/X _5630_/X _6706_/Q VGND VGND VPWR VPWR _5855_/X sky130_fd_sc_hd__a22o_1
XFILLER_21_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4806_ _4640_/B _4495_/X _4725_/B _4676_/B VGND VGND VPWR VPWR _4806_/X sky130_fd_sc_hd__o22a_1
XFILLER_167_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5786_ _6816_/Q _5913_/A2 _5785_/X VGND VGND VPWR VPWR _5786_/X sky130_fd_sc_hd__a21o_1
XFILLER_119_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4737_ _4894_/B _4737_/B _5025_/B VGND VGND VPWR VPWR _5021_/C sky130_fd_sc_hd__or3b_1
XFILLER_135_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_135_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_174_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4668_ _4965_/C _4703_/B VGND VGND VPWR VPWR _4668_/X sky130_fd_sc_hd__or2_1
XFILLER_119_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_647 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6407_ _3939_/A1 _6407_/D _6363_/X VGND VGND VPWR VPWR hold78/A sky130_fd_sc_hd__dfrtp_2
X_3619_ _6957_/Q _5397_/A _4002_/A _6453_/Q _3618_/X VGND VGND VPWR VPWR _3623_/C
+ sky130_fd_sc_hd__a221o_1
Xhold930 _5147_/X VGND VGND VPWR VPWR _6738_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold941 _6736_/Q VGND VGND VPWR VPWR hold941/X sky130_fd_sc_hd__dlygate4sd3_1
X_4599_ _4631_/A _5005_/A VGND VGND VPWR VPWR _4703_/B sky130_fd_sc_hd__or2_4
XFILLER_190_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold952 _4239_/X VGND VGND VPWR VPWR _6646_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_162_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold963 _6907_/Q VGND VGND VPWR VPWR hold963/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_162_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold974 _5309_/X VGND VGND VPWR VPWR _6875_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_115_371 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6338_ _6644_/Q _6338_/A2 _6338_/B1 _6643_/Q VGND VGND VPWR VPWR _6338_/X sky130_fd_sc_hd__a22o_1
Xhold985 _4114_/X VGND VGND VPWR VPWR _6533_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold996 _6891_/Q VGND VGND VPWR VPWR hold996/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_115_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6269_ _6648_/Q _5950_/X _6294_/A2 _6663_/Q VGND VGND VPWR VPWR _6269_/X sky130_fd_sc_hd__a22o_1
XFILLER_130_341 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_2_3_0_csclk clkbuf_2_3_0_csclk/A VGND VGND VPWR VPWR clkbuf_3_7_0_csclk/A
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_57_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_623 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_564 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_176_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_176_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_146 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_179 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_127 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_192_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_192_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3970_ hold153/X hold142/X _3974_/S VGND VGND VPWR VPWR _3970_/X sky130_fd_sc_hd__mux2_1
XFILLER_188_330 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5640_ _5643_/B _5651_/B VGND VGND VPWR VPWR _5667_/B sky130_fd_sc_hd__nand2_8
XFILLER_86_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5571_ _6506_/Q _5609_/B VGND VGND VPWR VPWR _5571_/Y sky130_fd_sc_hd__nand2_1
X_4522_ _4901_/B _4899_/B _4588_/B _4943_/B VGND VGND VPWR VPWR _4523_/D sky130_fd_sc_hd__o22a_1
Xhold204 _5509_/X VGND VGND VPWR VPWR _7053_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_7_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold215 _7188_/A VGND VGND VPWR VPWR hold215/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_7_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold226 _5213_/X VGND VGND VPWR VPWR _6790_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_144_455 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4453_ _4613_/C _4614_/A _4592_/B VGND VGND VPWR VPWR _4692_/C sky130_fd_sc_hd__or3b_4
Xhold237 _6424_/Q VGND VGND VPWR VPWR hold237/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_172_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold248 _5422_/X VGND VGND VPWR VPWR _6976_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_144_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold259 _6658_/Q VGND VGND VPWR VPWR hold259/X sky130_fd_sc_hd__dlygate4sd3_1
X_3404_ _7024_/Q hold18/A _5388_/A _6952_/Q VGND VGND VPWR VPWR _3404_/X sky130_fd_sc_hd__a22o_1
X_4384_ _4541_/B _4541_/C _4436_/A VGND VGND VPWR VPWR _4564_/A sky130_fd_sc_hd__a21o_1
XTAP_520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6123_ _6991_/Q _6286_/B1 _6282_/A2 _6999_/Q VGND VGND VPWR VPWR _6123_/X sky130_fd_sc_hd__a22o_1
X_3335_ hold73/X hold80/X VGND VGND VPWR VPWR _3401_/B sky130_fd_sc_hd__nand2_1
XTAP_531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6054_ _6507_/Q _6054_/A2 _5611_/X VGND VGND VPWR VPWR _6054_/X sky130_fd_sc_hd__a21o_1
XTAP_575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3266_ hold105/X hold29/X VGND VGND VPWR VPWR _3266_/Y sky130_fd_sc_hd__nand2b_1
XTAP_586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5005_ _5005_/A _5005_/B VGND VGND VPWR VPWR _5005_/X sky130_fd_sc_hd__or2_1
XFILLER_39_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3197_ _6973_/Q VGND VGND VPWR VPWR _3197_/Y sky130_fd_sc_hd__inv_2
XTAP_2409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6956_ _7083_/CLK _6956_/D fanout517/X VGND VGND VPWR VPWR _6956_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_41_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5907_ _6581_/Q _5617_/X _5639_/X _6553_/Q _5906_/X VGND VGND VPWR VPWR _5907_/X
+ sky130_fd_sc_hd__a221o_1
X_6887_ _6887_/CLK _6887_/D fanout524/X VGND VGND VPWR VPWR _6887_/Q sky130_fd_sc_hd__dfrtp_2
X_5838_ _6650_/Q _5922_/A2 _5632_/X _6599_/Q VGND VGND VPWR VPWR _5838_/X sky130_fd_sc_hd__a22o_1
X_5769_ _6871_/Q _5625_/X _5643_/X _6887_/Q _5768_/X VGND VGND VPWR VPWR _5769_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_148_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_175_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_135_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_680 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold760 _5194_/X VGND VGND VPWR VPWR _6773_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold771 _6510_/Q VGND VGND VPWR VPWR hold771/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold782 _5182_/X VGND VGND VPWR VPWR _6764_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold793 _7189_/A VGND VGND VPWR VPWR hold793/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_39_32 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1460 _7119_/Q VGND VGND VPWR VPWR _6029_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_17_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1471 _7141_/Q VGND VGND VPWR VPWR _6325_/A1 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1482 _6778_/Q VGND VGND VPWR VPWR hold1482/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1493 hold21/A VGND VGND VPWR VPWR _3252_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput309 _3946_/X VGND VGND VPWR VPWR spimemio_flash_io0_di sky130_fd_sc_hd__buf_12
XFILLER_154_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_141_403 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6810_ _7073_/CLK _6810_/D fanout498/X VGND VGND VPWR VPWR _6810_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_91_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6741_ _7037_/CLK _6741_/D fanout484/X VGND VGND VPWR VPWR _6741_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_189_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3953_ _6768_/Q _3953_/B VGND VGND VPWR VPWR _3953_/X sky130_fd_sc_hd__and2_2
XFILLER_50_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3884_ _7097_/Q _7098_/Q VGND VGND VPWR VPWR _5959_/A sky130_fd_sc_hd__nand2b_4
X_6672_ _6689_/CLK _6672_/D fanout510/X VGND VGND VPWR VPWR _6672_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_188_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5623_ _5667_/A _5649_/C _5650_/B VGND VGND VPWR VPWR _5623_/X sky130_fd_sc_hd__and3b_4
X_5554_ _5554_/A _5561_/A _5554_/C VGND VGND VPWR VPWR _7088_/D sky130_fd_sc_hd__and3_1
XFILLER_129_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4505_ _4503_/Y _4505_/B _5007_/A _4505_/D VGND VGND VPWR VPWR _4505_/X sky130_fd_sc_hd__and4b_1
X_5485_ hold235/X hold114/X _5486_/S VGND VGND VPWR VPWR _5485_/X sky130_fd_sc_hd__mux2_1
XFILLER_145_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_160_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4436_ _4436_/A _4590_/A VGND VGND VPWR VPWR _4977_/B sky130_fd_sc_hd__or2_4
XFILLER_132_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_160_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout503 fanout526/X VGND VGND VPWR VPWR fanout503/X sky130_fd_sc_hd__buf_8
Xfanout514 fanout525/X VGND VGND VPWR VPWR fanout514/X sky130_fd_sc_hd__clkbuf_16
X_7155_ _7155_/CLK _7155_/D fanout510/X VGND VGND VPWR VPWR _7155_/Q sky130_fd_sc_hd__dfrtp_2
X_4367_ _4613_/C _4367_/B VGND VGND VPWR VPWR _4894_/B sky130_fd_sc_hd__nand2_2
Xfanout525 fanout526/X VGND VGND VPWR VPWR fanout525/X sky130_fd_sc_hd__buf_8
X_3318_ _3571_/B _5168_/A VGND VGND VPWR VPWR _3975_/A sky130_fd_sc_hd__nor2_8
XFILLER_86_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_98_383 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6106_ _7007_/Q _6290_/A2 _6294_/A2 _7084_/Q VGND VGND VPWR VPWR _6106_/X sky130_fd_sc_hd__a22o_1
XFILLER_112_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7086_ _7086_/CLK _7086_/D fanout515/X VGND VGND VPWR VPWR _7086_/Q sky130_fd_sc_hd__dfrtp_1
X_4298_ _4298_/A0 _6353_/A1 _4302_/S VGND VGND VPWR VPWR _4298_/X sky130_fd_sc_hd__mux2_1
XFILLER_86_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3249_ _3248_/Y _3242_/A _3249_/S VGND VGND VPWR VPWR _7167_/D sky130_fd_sc_hd__mux2_1
XFILLER_86_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6037_ _6820_/Q _5969_/A _5957_/X _6956_/Q _6036_/X VGND VGND VPWR VPWR _6043_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_86_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6939_ _6945_/CLK _6939_/D fanout506/X VGND VGND VPWR VPWR _6939_/Q sky130_fd_sc_hd__dfstp_1
XPHY_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_44 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_0_csclk _3936_/X VGND VGND VPWR VPWR clkbuf_0_csclk/X sky130_fd_sc_hd__clkbuf_16
XFILLER_135_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_163_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold590 _6617_/Q VGND VGND VPWR VPWR hold590/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_96_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_173_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_173_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_1_0_0_csclk clkbuf_0_csclk/X VGND VGND VPWR VPWR clkbuf_1_0_1_csclk/A sky130_fd_sc_hd__clkbuf_8
XFILLER_18_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1290 _5231_/X VGND VGND VPWR VPWR _6806_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_45_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_272 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5270_ _5270_/A0 _5537_/A1 _5270_/S VGND VGND VPWR VPWR _5270_/X sky130_fd_sc_hd__mux2_1
XFILLER_114_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4221_ _6636_/Q _6637_/Q _6639_/Q _3167_/Y VGND VGND VPWR VPWR _4221_/X sky130_fd_sc_hd__or4b_1
XFILLER_99_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4152_ _4152_/A0 _5308_/A1 _4156_/S VGND VGND VPWR VPWR _4152_/X sky130_fd_sc_hd__mux2_1
XFILLER_110_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4083_ hold315/X _4082_/X _4095_/S VGND VGND VPWR VPWR _4083_/X sky130_fd_sc_hd__mux2_1
XFILLER_83_515 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_548 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_291 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_423 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4985_ _4985_/A _4985_/B VGND VGND VPWR VPWR _5061_/D sky130_fd_sc_hd__or2_1
XFILLER_23_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6724_ _7137_/CLK _6724_/D _4181_/B VGND VGND VPWR VPWR _6724_/Q sky130_fd_sc_hd__dfrtp_1
X_3936_ _6624_/Q _3936_/A2 _6396_/B _3935_/Y VGND VGND VPWR VPWR _3936_/X sky130_fd_sc_hd__a22o_2
XFILLER_189_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_3_2_0_csclk clkbuf_3_3_0_csclk/A VGND VGND VPWR VPWR clkbuf_3_2_0_csclk/X
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_176_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6655_ _6696_/CLK _6655_/D fanout495/X VGND VGND VPWR VPWR _6655_/Q sky130_fd_sc_hd__dfrtp_1
X_3867_ _3867_/A _3867_/B VGND VGND VPWR VPWR _3867_/Y sky130_fd_sc_hd__nor2_1
X_5606_ _5606_/A1 _5605_/B _5605_/Y _6507_/Q VGND VGND VPWR VPWR _7104_/D sky130_fd_sc_hd__a22o_1
XFILLER_164_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_192_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6586_ _7137_/CLK _6586_/D VGND VGND VPWR VPWR _6586_/Q sky130_fd_sc_hd__dfxtp_1
X_3798_ _6742_/Q _5151_/A _5170_/B _7173_/A VGND VGND VPWR VPWR _3798_/X sky130_fd_sc_hd__a22o_1
X_5537_ hold679/X _5537_/A1 _5537_/S VGND VGND VPWR VPWR _5537_/X sky130_fd_sc_hd__mux2_1
XFILLER_118_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_191_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5468_ hold195/X hold27/X _5468_/S VGND VGND VPWR VPWR _5468_/X sky130_fd_sc_hd__mux2_1
XFILLER_127_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4419_ _4613_/C _4419_/B VGND VGND VPWR VPWR _4944_/B sky130_fd_sc_hd__and2_1
XFILLER_160_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5399_ hold182/X hold90/X _5399_/S VGND VGND VPWR VPWR _5399_/X sky130_fd_sc_hd__mux2_1
X_7138_ _7140_/CLK _7138_/D VGND VGND VPWR VPWR _7138_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_143_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7069_ _7069_/CLK _7069_/D fanout516/X VGND VGND VPWR VPWR _7069_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_100_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_626 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_506 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput19 mask_rev_in[23] VGND VGND VPWR VPWR input19/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_168_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_109_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_170_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_97_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4770_ _4770_/A _4770_/B _5008_/C VGND VGND VPWR VPWR _4770_/X sky130_fd_sc_hd__and3_1
XTAP_1891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3721_ input21/X _3384_/Y _4225_/A _6626_/Q _3720_/X VGND VGND VPWR VPWR _3726_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_158_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_159_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6440_ _7034_/CLK _6440_/D fanout488/X VGND VGND VPWR VPWR _6440_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_146_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3652_ _3951_/A _4096_/A _3636_/X _3650_/X _3651_/X VGND VGND VPWR VPWR _3667_/B
+ sky130_fd_sc_hd__a2111o_1
XFILLER_174_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6371_ _6399_/A _6399_/B VGND VGND VPWR VPWR _6371_/X sky130_fd_sc_hd__and2_1
X_3583_ _6893_/Q _5325_/A _5163_/A _6754_/Q _3576_/X VGND VGND VPWR VPWR _3588_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_127_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5322_ hold767/X _5457_/A1 hold84/A VGND VGND VPWR VPWR _5322_/X sky130_fd_sc_hd__mux2_1
XFILLER_142_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5253_ _5253_/A _5511_/B VGND VGND VPWR VPWR _5261_/S sky130_fd_sc_hd__and2_4
X_4204_ hold903/X _5189_/A1 _4207_/S VGND VGND VPWR VPWR _4204_/X sky130_fd_sc_hd__mux2_1
X_5184_ hold429/X _5541_/A1 _5186_/S VGND VGND VPWR VPWR _5184_/X sky130_fd_sc_hd__mux2_1
XFILLER_68_331 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4135_ hold867/X _5189_/A1 _4138_/S VGND VGND VPWR VPWR _4135_/X sky130_fd_sc_hd__mux2_1
XFILLER_29_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_63_csclk clkbuf_3_2_0_csclk/X VGND VGND VPWR VPWR _7039_/CLK sky130_fd_sc_hd__clkbuf_16
X_4066_ _4066_/A0 _4065_/X _4078_/S VGND VGND VPWR VPWR _4066_/X sky130_fd_sc_hd__mux2_1
XFILLER_83_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_743 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_78_csclk _6661_/CLK VGND VGND VPWR VPWR _6695_/CLK sky130_fd_sc_hd__clkbuf_16
X_4968_ _4745_/B _4973_/B _4966_/X _4967_/X VGND VGND VPWR VPWR _4979_/B sky130_fd_sc_hd__o211a_1
X_6707_ _6707_/CLK _6707_/D fanout486/X VGND VGND VPWR VPWR _6707_/Q sky130_fd_sc_hd__dfstp_1
X_3919_ _6521_/Q input81/X _3951_/B VGND VGND VPWR VPWR _3919_/X sky130_fd_sc_hd__mux2_8
XFILLER_149_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4899_ _4965_/A _4899_/B VGND VGND VPWR VPWR _4899_/Y sky130_fd_sc_hd__nor2_1
XFILLER_177_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_164_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6638_ _7150_/CLK _6638_/D _6308_/B VGND VGND VPWR VPWR _6638_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_106_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6569_ _6632_/CLK _6569_/D _3264_/A VGND VGND VPWR VPWR _6569_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_3_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_152_328 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_145_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_16_csclk clkbuf_3_5_0_csclk/X VGND VGND VPWR VPWR _7043_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_105_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_275 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5940_ _7099_/Q _5940_/B _7102_/Q _7100_/Q VGND VGND VPWR VPWR _5953_/B sky130_fd_sc_hd__or4b_4
XFILLER_53_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5871_ _6562_/Q _5636_/X _5913_/B1 _6627_/Q _5870_/X VGND VGND VPWR VPWR _5872_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_179_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4822_ _4679_/A _4575_/A _4862_/A _4793_/Y _4821_/X VGND VGND VPWR VPWR _4822_/X
+ sky130_fd_sc_hd__o311a_1
XFILLER_166_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4753_ _4943_/A _4495_/X _4701_/A _4715_/B VGND VGND VPWR VPWR _5136_/B sky130_fd_sc_hd__o22a_1
X_3704_ input15/X _3339_/Y _5145_/A _6738_/Q VGND VGND VPWR VPWR _3704_/X sky130_fd_sc_hd__a22o_1
XFILLER_159_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4684_ _5005_/A _4717_/B VGND VGND VPWR VPWR _4684_/Y sky130_fd_sc_hd__nor2_1
XFILLER_146_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6423_ _7073_/CLK _6423_/D fanout497/X VGND VGND VPWR VPWR _6423_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_174_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3635_ _6924_/Q _5361_/A _3958_/A _6420_/Q VGND VGND VPWR VPWR _3635_/X sky130_fd_sc_hd__a22o_1
XFILLER_147_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_162_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6354_ _6354_/A0 _6354_/A1 hold54/A VGND VGND VPWR VPWR _6354_/X sky130_fd_sc_hd__mux2_1
X_3566_ _3566_/A _3566_/B _3566_/C _3566_/D VGND VGND VPWR VPWR _3567_/C sky130_fd_sc_hd__and4_1
XFILLER_161_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5305_ hold427/X _5545_/A1 _5306_/S VGND VGND VPWR VPWR _5305_/X sky130_fd_sc_hd__mux2_1
XFILLER_103_715 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_170_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3497_ _6862_/Q _5289_/A _4315_/A _6714_/Q VGND VGND VPWR VPWR _3497_/X sky130_fd_sc_hd__a22o_1
X_6285_ _6634_/Q _6285_/A2 _6285_/B1 _6479_/Q _6284_/X VGND VGND VPWR VPWR _6293_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_103_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_748 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5236_ _5236_/A0 _5530_/A1 _5243_/S VGND VGND VPWR VPWR _5236_/X sky130_fd_sc_hd__mux2_1
XFILLER_130_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5167_ hold229/X _5533_/A1 _5167_/S VGND VGND VPWR VPWR _5167_/X sky130_fd_sc_hd__mux2_1
XFILLER_56_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4118_ _4118_/A0 hold142/X _4120_/S VGND VGND VPWR VPWR _4118_/X sky130_fd_sc_hd__mux2_1
XFILLER_68_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5098_ _6724_/Q _4222_/X _5086_/X _5097_/X VGND VGND VPWR VPWR _5098_/X sky130_fd_sc_hd__a211o_1
XFILLER_37_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4049_ hold275/X _4048_/X _4061_/S VGND VGND VPWR VPWR _4049_/X sky130_fd_sc_hd__mux2_1
XFILLER_37_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_149_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_153_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_180_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_140_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_407 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_470 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold8 hold8/A VGND VGND VPWR VPWR hold8/X sky130_fd_sc_hd__buf_6
XFILLER_75_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_188_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_190_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_171_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_328 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold408 _4102_/X VGND VGND VPWR VPWR _6523_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold419 _6936_/Q VGND VGND VPWR VPWR hold419/X sky130_fd_sc_hd__dlygate4sd3_1
X_3420_ input32/X _3339_/Y _5424_/A _6984_/Q VGND VGND VPWR VPWR _3420_/X sky130_fd_sc_hd__a22o_1
XFILLER_99_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_131_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_143_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3351_ _3354_/A hold74/X VGND VGND VPWR VPWR _3391_/B sky130_fd_sc_hd__or2_4
XFILLER_112_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3282_ hold80/X hold73/X VGND VGND VPWR VPWR hold81/A sky130_fd_sc_hd__nand2b_1
XFILLER_98_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_112_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6070_ _6829_/Q _5974_/B _5977_/X _6925_/Q _6069_/X VGND VGND VPWR VPWR _6077_/A
+ sky130_fd_sc_hd__a221o_1
XTAP_746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1108 _4033_/X VGND VGND VPWR VPWR _6475_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5021_ _5021_/A _5021_/B _5021_/C VGND VGND VPWR VPWR _5021_/X sky130_fd_sc_hd__and3_1
XFILLER_112_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1119 _7030_/Q VGND VGND VPWR VPWR _5483_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_78_492 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_93_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6972_ _7075_/CLK _6972_/D fanout514/X VGND VGND VPWR VPWR _6972_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_53_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_359 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5923_ _6659_/Q _5923_/B VGND VGND VPWR VPWR _5923_/X sky130_fd_sc_hd__and2b_1
XFILLER_80_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5854_ _6615_/Q _5928_/B1 _5850_/X _5851_/X _5853_/X VGND VGND VPWR VPWR _5854_/X
+ sky130_fd_sc_hd__a2111o_1
XFILLER_22_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4805_ _4921_/A _4495_/X _5043_/B _4597_/Y VGND VGND VPWR VPWR _4805_/X sky130_fd_sc_hd__o22a_1
XFILLER_167_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5785_ _6968_/Q _5925_/B1 _5650_/X _6896_/Q VGND VGND VPWR VPWR _5785_/X sky130_fd_sc_hd__a22o_1
XFILLER_166_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4736_ _4885_/A _4736_/B VGND VGND VPWR VPWR _4736_/X sky130_fd_sc_hd__or2_1
XFILLER_174_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4667_ _5043_/B _4725_/B _4672_/B _4788_/A VGND VGND VPWR VPWR _4812_/A sky130_fd_sc_hd__a211o_1
X_6406_ _3939_/A1 _6406_/D _6362_/X VGND VGND VPWR VPWR _6406_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_135_659 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold920 _5279_/X VGND VGND VPWR VPWR _6849_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3618_ _6925_/Q _5361_/A _5415_/A _6973_/Q VGND VGND VPWR VPWR _3618_/X sky130_fd_sc_hd__a22o_1
XFILLER_190_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold931 _6466_/Q VGND VGND VPWR VPWR hold931/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_162_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4598_ _4617_/B _4613_/C _4630_/A _4888_/A VGND VGND VPWR VPWR _5005_/A sky130_fd_sc_hd__or4b_4
Xhold942 _5144_/X VGND VGND VPWR VPWR _6736_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_122_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold953 _7040_/Q VGND VGND VPWR VPWR hold953/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold964 _5345_/X VGND VGND VPWR VPWR _6907_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_1_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6337_ _6336_/X _6337_/A1 _6346_/S VGND VGND VPWR VPWR _7145_/D sky130_fd_sc_hd__mux2_1
X_3549_ _3563_/A _5161_/B VGND VGND VPWR VPWR _4008_/A sky130_fd_sc_hd__nor2_4
Xhold975 _6827_/Q VGND VGND VPWR VPWR hold975/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold986 _6605_/Q VGND VGND VPWR VPWR hold986/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_1_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold997 _5327_/X VGND VGND VPWR VPWR _6891_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_88_234 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6268_ _6268_/A _6268_/B _6268_/C _6267_/Y VGND VGND VPWR VPWR _6268_/X sky130_fd_sc_hd__or4b_2
XFILLER_142_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5219_ hold923/X _5531_/A1 _5225_/S VGND VGND VPWR VPWR _5219_/X sky130_fd_sc_hd__mux2_1
XFILLER_103_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6199_ _6599_/Q _5939_/X _5953_/Y _6480_/Q _6198_/X VGND VGND VPWR VPWR _6200_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_84_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_462 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_185_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_181_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_497 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_180_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_180_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_140_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_353 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_418 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_188_342 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_206 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5570_ _5570_/A _6508_/Q VGND VGND VPWR VPWR _5597_/B sky130_fd_sc_hd__nor2_1
XFILLER_79_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4521_ _4943_/B _4581_/A _5106_/A _4519_/X _4520_/X VGND VGND VPWR VPWR _4523_/C
+ sky130_fd_sc_hd__o2111a_1
XFILLER_156_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_144_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold205 _6968_/Q VGND VGND VPWR VPWR hold205/X sky130_fd_sc_hd__dlygate4sd3_1
X_4452_ _4613_/C _4630_/A _4592_/B VGND VGND VPWR VPWR _4947_/B sky130_fd_sc_hd__and3b_2
Xhold216 _4061_/X VGND VGND VPWR VPWR _6497_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold227 _6977_/Q VGND VGND VPWR VPWR hold227/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold238 _3972_/X VGND VGND VPWR VPWR _6424_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold249 _6563_/Q VGND VGND VPWR VPWR hold249/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3403_ _7131_/Q _6761_/Q _6762_/Q VGND VGND VPWR VPWR _3403_/X sky130_fd_sc_hd__mux2_2
XFILLER_144_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7171_ _7171_/CLK _7171_/D _6401_/X VGND VGND VPWR VPWR _7171_/Q sky130_fd_sc_hd__dfrtp_1
X_4383_ _4888_/A _4542_/C _4383_/C VGND VGND VPWR VPWR _4541_/C sky130_fd_sc_hd__and3_1
XFILLER_131_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6122_ _6911_/Q _5972_/A _6285_/B1 _7015_/Q _6121_/X VGND VGND VPWR VPWR _6127_/B
+ sky130_fd_sc_hd__a221o_1
XTAP_521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3334_ _7086_/Q _5538_/A _5298_/A _6873_/Q VGND VGND VPWR VPWR _3334_/X sky130_fd_sc_hd__a22o_2
XFILLER_124_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6053_ _6788_/Q _5975_/X _6043_/X _6052_/X _3174_/Y VGND VGND VPWR VPWR _6053_/X
+ sky130_fd_sc_hd__o221a_2
XTAP_576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3265_ _7171_/Q hold5/A _6487_/Q _3858_/B VGND VGND VPWR VPWR _7156_/D sky130_fd_sc_hd__o211a_1
XTAP_587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5004_ _4965_/B _4973_/A _4743_/Y _5017_/A VGND VGND VPWR VPWR _5004_/X sky130_fd_sc_hd__o211a_1
X_3196_ _6981_/Q VGND VGND VPWR VPWR _3196_/Y sky130_fd_sc_hd__inv_2
XFILLER_38_164 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6955_ _7083_/CLK _6955_/D fanout519/X VGND VGND VPWR VPWR _6955_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_81_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5906_ _6468_/Q _5629_/X _5631_/X _6612_/Q VGND VGND VPWR VPWR _5906_/X sky130_fd_sc_hd__a22o_1
X_6886_ _7043_/CLK _6886_/D fanout518/X VGND VGND VPWR VPWR _6886_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_179_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5837_ _6470_/Q _5622_/X _5626_/X _6695_/Q _5836_/X VGND VGND VPWR VPWR _5842_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_167_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5768_ _6903_/Q _5623_/X _5637_/X _6855_/Q VGND VGND VPWR VPWR _5768_/X sky130_fd_sc_hd__a22o_1
XFILLER_5_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4719_ _4965_/A _4719_/B VGND VGND VPWR VPWR _4720_/C sky130_fd_sc_hd__nor2_1
X_5699_ _6924_/Q _5633_/X _5646_/X _6996_/Q VGND VGND VPWR VPWR _5699_/X sky130_fd_sc_hd__a22o_1
XFILLER_107_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_135_478 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_190_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold750 _5544_/X VGND VGND VPWR VPWR _7084_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold761 _6837_/Q VGND VGND VPWR VPWR hold761/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold772 _4081_/X VGND VGND VPWR VPWR _6510_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold783 _6557_/Q VGND VGND VPWR VPWR hold783/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_1_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold794 _5191_/X VGND VGND VPWR VPWR _6770_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_39_44 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1450 _7106_/Q VGND VGND VPWR VPWR _5690_/A1 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1461 _7158_/Q VGND VGND VPWR VPWR _3904_/A2 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1472 _7104_/Q VGND VGND VPWR VPWR _5606_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_29_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1483 hold10/A VGND VGND VPWR VPWR _6331_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_72_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1494 _7108_/Q VGND VGND VPWR VPWR _5713_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_185_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_187_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_185_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_138_294 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_415 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6740_ _7037_/CLK _6740_/D fanout484/X VGND VGND VPWR VPWR _6740_/Q sky130_fd_sc_hd__dfrtp_4
X_3952_ _3952_/A input1/X VGND VGND VPWR VPWR _3952_/X sky130_fd_sc_hd__and2_1
XFILLER_189_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6671_ _6708_/CLK _6671_/D _6400_/A VGND VGND VPWR VPWR _6671_/Q sky130_fd_sc_hd__dfrtp_1
X_3883_ _7097_/Q _7098_/Q VGND VGND VPWR VPWR _5981_/A sky130_fd_sc_hd__and2b_2
X_5622_ _5667_/A _5646_/B _5651_/C VGND VGND VPWR VPWR _5622_/X sky130_fd_sc_hd__and3_4
X_5553_ _7088_/Q _5558_/D VGND VGND VPWR VPWR _5554_/C sky130_fd_sc_hd__nand2_1
XFILLER_191_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_191_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4504_ _5043_/A _4885_/A _4692_/C _4640_/B _4748_/A VGND VGND VPWR VPWR _4505_/B
+ sky130_fd_sc_hd__o32a_1
X_5484_ hold727/X _5544_/A1 _5486_/S VGND VGND VPWR VPWR _5484_/X sky130_fd_sc_hd__mux2_1
XFILLER_144_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4435_ _4542_/A _4435_/B VGND VGND VPWR VPWR _4435_/Y sky130_fd_sc_hd__nor2_1
XFILLER_144_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout504 fanout526/X VGND VGND VPWR VPWR fanout504/X sky130_fd_sc_hd__buf_8
X_7154_ _7155_/CLK hold55/X _6370_/A VGND VGND VPWR VPWR _7154_/Q sky130_fd_sc_hd__dfrtp_1
Xfanout515 fanout525/X VGND VGND VPWR VPWR fanout515/X sky130_fd_sc_hd__buf_8
X_4366_ _4554_/A _4570_/B VGND VGND VPWR VPWR _4417_/B sky130_fd_sc_hd__or2_1
Xfanout526 input75/X VGND VGND VPWR VPWR fanout526/X sky130_fd_sc_hd__buf_12
X_6105_ _6129_/A1 _5612_/Y _6103_/X _6104_/X VGND VGND VPWR VPWR _6105_/X sky130_fd_sc_hd__o22a_1
XFILLER_113_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3317_ _5168_/A VGND VGND VPWR VPWR _3317_/Y sky130_fd_sc_hd__inv_2
XFILLER_113_684 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7085_ _7086_/CLK _7085_/D fanout525/X VGND VGND VPWR VPWR _7085_/Q sky130_fd_sc_hd__dfrtp_2
X_4297_ _4297_/A hold7/X VGND VGND VPWR VPWR _4302_/S sky130_fd_sc_hd__and2_4
XFILLER_112_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6036_ _6812_/Q _5936_/X _6286_/B1 _6988_/Q VGND VGND VPWR VPWR _6036_/X sky130_fd_sc_hd__a22o_1
X_3248_ _7167_/Q _6485_/Q _3247_/Y VGND VGND VPWR VPWR _3248_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_67_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3179_ _6489_/Q VGND VGND VPWR VPWR _3179_/Y sky130_fd_sc_hd__inv_2
XTAP_2207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6938_ _6978_/CLK _6938_/D fanout500/X VGND VGND VPWR VPWR _6938_/Q sky130_fd_sc_hd__dfstp_1
XPHY_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6869_ _6999_/CLK _6869_/D fanout524/X VGND VGND VPWR VPWR _6869_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_155_518 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_151_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_459 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold580 _4260_/X VGND VGND VPWR VPWR _6664_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold591 _4212_/X VGND VGND VPWR VPWR _6617_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_173_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1280 _5303_/X VGND VGND VPWR VPWR _6870_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1291 _6446_/Q VGND VGND VPWR VPWR _3998_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_186_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_173_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_185_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_173_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_126_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4220_ _6643_/Q _6642_/Q _6644_/Q VGND VGND VPWR VPWR _4223_/B sky130_fd_sc_hd__nor3_2
X_4151_ _4151_/A hold7/X VGND VGND VPWR VPWR _4156_/S sky130_fd_sc_hd__and2_2
XFILLER_83_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4082_ hold207/X hold90/X _4092_/S VGND VGND VPWR VPWR _4082_/X sky130_fd_sc_hd__mux2_1
XFILLER_83_527 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_435 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4984_ _4984_/A _4984_/B _4984_/C VGND VGND VPWR VPWR _5067_/B sky130_fd_sc_hd__nand3_2
X_6723_ _7140_/CLK _6723_/D _4181_/B VGND VGND VPWR VPWR _6723_/Q sky130_fd_sc_hd__dfrtp_1
X_3935_ _6624_/Q _3935_/B VGND VGND VPWR VPWR _3935_/Y sky130_fd_sc_hd__nor2_2
X_6654_ _7155_/CLK _6654_/D _6370_/A VGND VGND VPWR VPWR _6654_/Q sky130_fd_sc_hd__dfrtp_2
X_3866_ _7104_/Q _6757_/Q _6762_/Q VGND VGND VPWR VPWR _5605_/A sky130_fd_sc_hd__mux2_2
XFILLER_176_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5605_ _5605_/A _5605_/B VGND VGND VPWR VPWR _5605_/Y sky130_fd_sc_hd__nor2_1
XFILLER_164_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6585_ _7137_/CLK _6585_/D VGND VGND VPWR VPWR _6585_/Q sky130_fd_sc_hd__dfxtp_1
X_3797_ _3797_/A _5168_/A VGND VGND VPWR VPWR _5170_/B sky130_fd_sc_hd__nor2_1
XFILLER_176_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5536_ _5536_/A0 hold114/X _5537_/S VGND VGND VPWR VPWR _5536_/X sky130_fd_sc_hd__mux2_1
X_5467_ hold620/X _5545_/A1 _5468_/S VGND VGND VPWR VPWR _5467_/X sky130_fd_sc_hd__mux2_1
XFILLER_160_543 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4418_ _4691_/A _4418_/B VGND VGND VPWR VPWR _4943_/B sky130_fd_sc_hd__nand2_8
X_5398_ _5398_/A0 _5521_/A1 _5405_/S VGND VGND VPWR VPWR _5398_/X sky130_fd_sc_hd__mux2_1
XFILLER_99_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_682 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7137_ _7137_/CLK _7137_/D VGND VGND VPWR VPWR _7137_/Q sky130_fd_sc_hd__dfxtp_1
X_4349_ _4356_/B _4592_/A _4617_/B VGND VGND VPWR VPWR _4350_/B sky130_fd_sc_hd__a21oi_1
XFILLER_86_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_654 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7068_ _7084_/CLK _7068_/D fanout514/X VGND VGND VPWR VPWR _7068_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_86_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_207 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6019_ _6803_/Q _5973_/B _5974_/B _6827_/Q VGND VGND VPWR VPWR _6019_/X sky130_fd_sc_hd__a22o_1
XFILLER_39_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_638 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_146_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_182_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_167 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_124_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_124_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_151_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_719 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3720_ _6875_/Q _5307_/A _5158_/A _6749_/Q VGND VGND VPWR VPWR _3720_/X sky130_fd_sc_hd__a22o_1
XFILLER_159_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_490 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_158_175 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3651_ _6796_/Q _5217_/A _4249_/A _6657_/Q _3638_/X VGND VGND VPWR VPWR _3651_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_158_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_173_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6370_ _6370_/A _6401_/B VGND VGND VPWR VPWR _6370_/X sky130_fd_sc_hd__and2_1
X_3582_ _6683_/Q _4279_/A _4261_/A _6668_/Q _3581_/X VGND VGND VPWR VPWR _3588_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_127_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5321_ _5321_/A0 _5465_/A1 hold84/A VGND VGND VPWR VPWR _5321_/X sky130_fd_sc_hd__mux2_1
XFILLER_5_380 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5252_ hold185/X hold27/X _5252_/S VGND VGND VPWR VPWR _5252_/X sky130_fd_sc_hd__mux2_1
X_4203_ _4203_/A0 _5308_/A1 _4207_/S VGND VGND VPWR VPWR _4203_/X sky130_fd_sc_hd__mux2_1
X_5183_ _5183_/A _5183_/B _5511_/B VGND VGND VPWR VPWR _5186_/S sky130_fd_sc_hd__nor3b_4
XFILLER_68_343 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4134_ _4134_/A0 _5308_/A1 _4138_/S VGND VGND VPWR VPWR _4134_/X sky130_fd_sc_hd__mux2_1
XFILLER_3_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_462 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_313 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4065_ hold984/X _6354_/A1 _4112_/B VGND VGND VPWR VPWR _4065_/X sky130_fd_sc_hd__mux2_1
XFILLER_83_357 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4967_ _4501_/B _4748_/B _4695_/B _4962_/X VGND VGND VPWR VPWR _4967_/X sky130_fd_sc_hd__o22a_1
X_3918_ _6519_/Q input78/X _3951_/B VGND VGND VPWR VPWR _3918_/X sky130_fd_sc_hd__mux2_8
X_6706_ _6769_/CLK _6706_/D fanout492/X VGND VGND VPWR VPWR _6706_/Q sky130_fd_sc_hd__dfrtp_1
X_4898_ _4898_/A _4898_/B VGND VGND VPWR VPWR _5100_/C sky130_fd_sc_hd__and2_1
XFILLER_149_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6637_ _7150_/CLK _6637_/D _6308_/B VGND VGND VPWR VPWR _6637_/Q sky130_fd_sc_hd__dfrtp_2
X_3849_ _3848_/X _3849_/A1 _3857_/S VGND VGND VPWR VPWR _6410_/D sky130_fd_sc_hd__mux2_1
XFILLER_192_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_137_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6568_ _6683_/CLK _6568_/D fanout496/X VGND VGND VPWR VPWR _6568_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_152_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_106_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5519_ hold301/X _5519_/A1 _5519_/S VGND VGND VPWR VPWR _5519_/X sky130_fd_sc_hd__mux2_1
X_6499_ _6711_/CLK _6499_/D fanout486/X VGND VGND VPWR VPWR _6499_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_106_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_700 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_413 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_435 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_179_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_552 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_287 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_187_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_168_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_156_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_183_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_170_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_112_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_111_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5870_ _6616_/Q _5928_/B1 _5634_/X _6687_/Q VGND VGND VPWR VPWR _5870_/X sky130_fd_sc_hd__a22o_1
XFILLER_179_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4821_ _4525_/C _4724_/B _4821_/C _4821_/D VGND VGND VPWR VPWR _4821_/X sky130_fd_sc_hd__and4bb_1
XFILLER_178_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4752_ _4703_/A _4676_/B _4506_/C VGND VGND VPWR VPWR _4752_/X sky130_fd_sc_hd__o21a_1
X_3703_ _6843_/Q _5271_/A _5379_/A _6939_/Q _3702_/X VGND VGND VPWR VPWR _3711_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_174_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4683_ _4703_/B _4683_/B VGND VGND VPWR VPWR _4683_/Y sky130_fd_sc_hd__nor2_1
X_6422_ _7010_/CLK _6422_/D fanout498/X VGND VGND VPWR VPWR _6422_/Q sky130_fd_sc_hd__dfstp_1
X_3634_ _6436_/Q _3984_/A _4315_/A _6712_/Q VGND VGND VPWR VPWR _3634_/X sky130_fd_sc_hd__a22o_1
XFILLER_134_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6353_ _6353_/A0 _6353_/A1 hold54/A VGND VGND VPWR VPWR _6353_/X sky130_fd_sc_hd__mux2_1
XFILLER_127_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3565_ _3565_/A _3565_/B _3565_/C _3565_/D VGND VGND VPWR VPWR _3566_/D sky130_fd_sc_hd__nor4_1
X_5304_ hold669/X _5544_/A1 _5306_/S VGND VGND VPWR VPWR _5304_/X sky130_fd_sc_hd__mux2_1
X_6284_ _6618_/Q _5971_/A _6284_/B1 _6613_/Q VGND VGND VPWR VPWR _6284_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3496_ _3554_/A _3560_/B VGND VGND VPWR VPWR _4315_/A sky130_fd_sc_hd__nor2_8
XFILLER_103_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5235_ _5235_/A _5529_/B VGND VGND VPWR VPWR _5243_/S sky130_fd_sc_hd__and2_4
XFILLER_69_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5166_ hold397/X _5532_/A1 _5167_/S VGND VGND VPWR VPWR _5166_/X sky130_fd_sc_hd__mux2_1
XFILLER_69_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4117_ hold379/X _5534_/A1 _4120_/S VGND VGND VPWR VPWR _4117_/X sky130_fd_sc_hd__mux2_1
X_5097_ _5091_/A _5124_/B _5134_/A _5121_/B VGND VGND VPWR VPWR _5097_/X sky130_fd_sc_hd__o31a_1
XFILLER_84_666 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4048_ hold126/X hold90/X _4103_/B VGND VGND VPWR VPWR _4048_/X sky130_fd_sc_hd__mux2_1
XFILLER_17_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5999_ _6818_/Q _5969_/A _5951_/X _7071_/Q _5998_/X VGND VGND VPWR VPWR _6003_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_52_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_602 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_177_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_177_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_177_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_137_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_627 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_660 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput290 _6437_/Q VGND VGND VPWR VPWR pll_trim[3] sky130_fd_sc_hd__buf_12
XFILLER_181_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold9 hold9/A VGND VGND VPWR VPWR hold9/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_87_482 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_235 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_62_csclk clkbuf_3_2_0_csclk/X VGND VGND VPWR VPWR _7073_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_116_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold409 _6667_/Q VGND VGND VPWR VPWR hold409/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_7_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3350_ _3797_/A _3525_/A VGND VGND VPWR VPWR _5334_/A sky130_fd_sc_hd__nor2_8
XTAP_703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_77_csclk _6661_/CLK VGND VGND VPWR VPWR _7038_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3281_ hold79/X _6720_/Q _6624_/Q VGND VGND VPWR VPWR hold80/A sky130_fd_sc_hd__mux2_1
XFILLER_151_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5020_ _5020_/A _5020_/B VGND VGND VPWR VPWR _5102_/A sky130_fd_sc_hd__and2_1
XTAP_769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1109 _6599_/Q VGND VGND VPWR VPWR _4191_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_66_600 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6971_ _7073_/CLK _6971_/D fanout497/X VGND VGND VPWR VPWR _6971_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_93_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5922_ _6654_/Q _5922_/A2 _5922_/B1 _6603_/Q _5921_/X VGND VGND VPWR VPWR _5930_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_22_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5853_ _6579_/Q _5617_/X _5920_/A2 _6566_/Q _5852_/X VGND VGND VPWR VPWR _5853_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_110_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_15_csclk clkbuf_3_5_0_csclk/X VGND VGND VPWR VPWR _6990_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_61_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4804_ _4921_/A _4588_/B _5043_/B _4695_/B VGND VGND VPWR VPWR _4819_/A sky130_fd_sc_hd__o22a_1
X_5784_ _6952_/Q _5924_/B2 _5912_/B1 _7032_/Q _5783_/X VGND VGND VPWR VPWR _5784_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_9_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4735_ _4401_/B _4549_/B _4703_/A _4615_/B VGND VGND VPWR VPWR _4736_/B sky130_fd_sc_hd__o22a_1
XFILLER_159_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4666_ _4666_/A _4666_/B _4666_/C VGND VGND VPWR VPWR _4666_/X sky130_fd_sc_hd__and3_1
XFILLER_135_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6405_ _3939_/A1 _6405_/D _6361_/X VGND VGND VPWR VPWR _6405_/Q sky130_fd_sc_hd__dfrtp_4
X_3617_ input14/X _3355_/Y _5379_/A _6941_/Q _3570_/X VGND VGND VPWR VPWR _3623_/B
+ sky130_fd_sc_hd__a221o_1
Xhold910 _5387_/X VGND VGND VPWR VPWR _6945_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_134_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold921 _6566_/Q VGND VGND VPWR VPWR hold921/X sky130_fd_sc_hd__dlygate4sd3_1
X_4597_ _4707_/B _4707_/C VGND VGND VPWR VPWR _4597_/Y sky130_fd_sc_hd__nand2_8
Xhold932 _4022_/X VGND VGND VPWR VPWR _6466_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold943 _7035_/Q VGND VGND VPWR VPWR hold943/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_162_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold954 _5495_/X VGND VGND VPWR VPWR _7040_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6336_ _6644_/Q _6336_/A2 _6336_/B1 _6643_/Q _6335_/X VGND VGND VPWR VPWR _6336_/X
+ sky130_fd_sc_hd__a221o_1
X_3548_ _3548_/A _3548_/B _3548_/C VGND VGND VPWR VPWR _3566_/C sky130_fd_sc_hd__nor3_1
Xhold965 _7009_/Q VGND VGND VPWR VPWR hold965/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_143_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold976 _5255_/X VGND VGND VPWR VPWR _6827_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold987 _4198_/X VGND VGND VPWR VPWR _6605_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold998 _6686_/Q VGND VGND VPWR VPWR hold998/X sky130_fd_sc_hd__dlygate4sd3_1
X_6267_ _6267_/A _6267_/B VGND VGND VPWR VPWR _6267_/Y sky130_fd_sc_hd__nor2_1
X_3479_ _3552_/A _3538_/B VGND VGND VPWR VPWR _4297_/A sky130_fd_sc_hd__nor2_4
XFILLER_88_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5218_ _5218_/A0 _5530_/A1 _5225_/S VGND VGND VPWR VPWR _5218_/X sky130_fd_sc_hd__mux2_1
XFILLER_76_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6198_ _6555_/Q _6259_/A2 _5972_/A _6650_/Q VGND VGND VPWR VPWR _6198_/X sky130_fd_sc_hd__a22o_1
X_5149_ hold497/X _5491_/A1 _5150_/S VGND VGND VPWR VPWR _5149_/X sky130_fd_sc_hd__mux2_1
XFILLER_72_603 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_179 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_599 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_176_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_671 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_706 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_400 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_176_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_188_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_148_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_148_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4520_ _4943_/A _4581_/A VGND VGND VPWR VPWR _4520_/X sky130_fd_sc_hd__or2_1
XFILLER_172_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold206 _5413_/X VGND VGND VPWR VPWR _6968_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4451_ _4613_/C _4614_/A VGND VGND VPWR VPWR _4617_/A sky130_fd_sc_hd__or2_1
Xhold217 _6758_/Q VGND VGND VPWR VPWR hold217/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_172_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold228 _5423_/X VGND VGND VPWR VPWR _6977_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold239 _6789_/Q VGND VGND VPWR VPWR hold239/X sky130_fd_sc_hd__dlygate4sd3_1
X_3402_ _5183_/A hold53/X VGND VGND VPWR VPWR _5179_/B sky130_fd_sc_hd__nor2_8
XFILLER_171_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7170_ _3939_/A1 _7170_/D _6400_/X VGND VGND VPWR VPWR _7170_/Q sky130_fd_sc_hd__dfrtp_1
X_4382_ _4542_/C _4383_/C VGND VGND VPWR VPWR _4390_/A sky130_fd_sc_hd__and2_1
XFILLER_125_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6121_ _6447_/Q _5601_/Y _6176_/A2 _6983_/Q VGND VGND VPWR VPWR _6121_/X sky130_fd_sc_hd__a22o_1
XTAP_511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3333_ _3525_/A _3487_/A VGND VGND VPWR VPWR _5298_/A sky130_fd_sc_hd__nor2_8
XFILLER_112_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6052_ _6052_/A _6052_/B _6052_/C _6004_/B VGND VGND VPWR VPWR _6052_/X sky130_fd_sc_hd__or4b_1
XTAP_566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3264_ _3264_/A _6396_/B VGND VGND VPWR VPWR _3264_/X sky130_fd_sc_hd__and2_1
XFILLER_98_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5003_ _5062_/A _5003_/B VGND VGND VPWR VPWR _5003_/X sky130_fd_sc_hd__and2_1
XTAP_599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3195_ _6989_/Q VGND VGND VPWR VPWR _3195_/Y sky130_fd_sc_hd__inv_2
XFILLER_38_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_422 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6954_ _7083_/CLK _6954_/D fanout518/X VGND VGND VPWR VPWR _6954_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_179_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5905_ _6648_/Q _5918_/A2 _5918_/B1 _6607_/Q _5904_/X VGND VGND VPWR VPWR _5905_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_81_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_179_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6885_ _7058_/CLK _6885_/D fanout524/X VGND VGND VPWR VPWR _6885_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_22_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5836_ _5667_/B _5835_/X _6614_/Q _5928_/B1 VGND VGND VPWR VPWR _5836_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_167_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5767_ _6927_/Q _5633_/X _5646_/X _6999_/Q VGND VGND VPWR VPWR _5767_/X sky130_fd_sc_hd__a22o_1
X_4718_ _4718_/A _4718_/B _4718_/C _4697_/X VGND VGND VPWR VPWR _4720_/B sky130_fd_sc_hd__or4b_1
X_5698_ _6972_/Q _5644_/X _5807_/B1 _6932_/Q _5697_/X VGND VGND VPWR VPWR _5698_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_147_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4649_ _4649_/A _4649_/B VGND VGND VPWR VPWR _4985_/B sky130_fd_sc_hd__or2_1
XFILLER_190_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold740 _5311_/X VGND VGND VPWR VPWR _6877_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold751 _7042_/Q VGND VGND VPWR VPWR hold751/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_190_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold762 _5266_/X VGND VGND VPWR VPWR _6837_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold773 _6702_/Q VGND VGND VPWR VPWR hold773/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold784 _4142_/X VGND VGND VPWR VPWR _6557_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_143_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6319_ _6320_/B _6348_/B1 _6643_/Q VGND VGND VPWR VPWR _6322_/B sky130_fd_sc_hd__a21boi_1
Xhold795 _6436_/Q VGND VGND VPWR VPWR hold795/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_131_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1440 _6729_/Q VGND VGND VPWR VPWR _3686_/A1 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1451 _6637_/Q VGND VGND VPWR VPWR _3871_/B1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_29_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1462 _7105_/Q VGND VGND VPWR VPWR _5608_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_45_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1473 hold96/A VGND VGND VPWR VPWR _6346_/A1 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1484 _7121_/Q VGND VGND VPWR VPWR _6079_/A2 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_176_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1495 _7131_/Q VGND VGND VPWR VPWR _6305_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_647 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_187_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_187_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_153_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_427 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3951_ _3951_/A _3951_/B VGND VGND VPWR VPWR _3951_/X sky130_fd_sc_hd__and2_1
XFILLER_44_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_190 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6670_ _6708_/CLK _6670_/D _6400_/A VGND VGND VPWR VPWR _6670_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_91_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3882_ _5940_/B _7102_/Q VGND VGND VPWR VPWR _5968_/A sky130_fd_sc_hd__and2_2
XFILLER_149_538 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5621_ _7093_/Q _7092_/Q VGND VGND VPWR VPWR _5651_/C sky130_fd_sc_hd__and2b_2
XFILLER_188_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5552_ _6507_/Q _3880_/B _5550_/Y _6509_/Q VGND VGND VPWR VPWR _5561_/A sky130_fd_sc_hd__a211o_1
XFILLER_145_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_191_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4503_ _4425_/X _4503_/B _4503_/C _4503_/D VGND VGND VPWR VPWR _4503_/Y sky130_fd_sc_hd__nand4b_1
XFILLER_191_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5483_ _5483_/A0 _5543_/A1 _5486_/S VGND VGND VPWR VPWR _5483_/X sky130_fd_sc_hd__mux2_1
X_4434_ _4557_/B _4677_/B VGND VGND VPWR VPWR _4898_/A sky130_fd_sc_hd__nand2_1
XFILLER_6_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7153_ _7153_/CLK _7153_/D _3940_/B VGND VGND VPWR VPWR _7153_/Q sky130_fd_sc_hd__dfstp_2
X_4365_ _4554_/A _4570_/B VGND VGND VPWR VPWR _4418_/B sky130_fd_sc_hd__nor2_2
Xfanout505 fanout526/X VGND VGND VPWR VPWR fanout505/X sky130_fd_sc_hd__buf_4
XFILLER_98_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout516 fanout525/X VGND VGND VPWR VPWR fanout516/X sky130_fd_sc_hd__buf_6
X_6104_ _6507_/Q _7122_/Q _5611_/X VGND VGND VPWR VPWR _6104_/X sky130_fd_sc_hd__a21o_1
Xfanout527 _4181_/B VGND VGND VPWR VPWR _6308_/B sky130_fd_sc_hd__buf_12
X_3316_ _3328_/A _3328_/B VGND VGND VPWR VPWR _3706_/B sky130_fd_sc_hd__nand2b_4
XFILLER_112_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7084_ _7084_/CLK _7084_/D fanout522/X VGND VGND VPWR VPWR _7084_/Q sky130_fd_sc_hd__dfrtp_1
X_4296_ _4296_/A0 _5543_/A1 _4296_/S VGND VGND VPWR VPWR _4296_/X sky130_fd_sc_hd__mux2_1
XFILLER_58_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_696 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6035_ _6884_/Q _6296_/A2 _6290_/B1 _7020_/Q _6034_/X VGND VGND VPWR VPWR _6043_/B
+ sky130_fd_sc_hd__a221o_1
X_3247_ _3247_/A _6485_/Q VGND VGND VPWR VPWR _3247_/Y sky130_fd_sc_hd__nand2_1
XTAP_396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3178_ _4544_/A VGND VGND VPWR VPWR _4436_/A sky130_fd_sc_hd__inv_2
XTAP_2208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6937_ _7029_/CLK hold43/X fanout523/X VGND VGND VPWR VPWR _6937_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6868_ _7083_/CLK _6868_/D fanout518/X VGND VGND VPWR VPWR _6868_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_22_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5819_ _6817_/Q _5913_/A2 _5628_/X _6913_/Q VGND VGND VPWR VPWR _5819_/X sky130_fd_sc_hd__a22o_1
XFILLER_22_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6799_ _7042_/CLK _6799_/D fanout519/X VGND VGND VPWR VPWR _6799_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_10_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_175_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_163_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_190_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold570 _5410_/X VGND VGND VPWR VPWR _6965_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_2_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold581 _6458_/Q VGND VGND VPWR VPWR hold581/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold592 _7061_/Q VGND VGND VPWR VPWR hold592/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_150_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1270 _5438_/X VGND VGND VPWR VPWR _6990_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_17_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1281 hold1541/X VGND VGND VPWR VPWR _4064_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_57_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1292 _3998_/X VGND VGND VPWR VPWR _6446_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_186_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_186_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_186_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_276 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_202 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_438 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_141_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4150_ hold531/X _6357_/A1 _4150_/S VGND VGND VPWR VPWR _4150_/X sky130_fd_sc_hd__mux2_1
XFILLER_95_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4081_ hold771/X _4080_/X _4095_/S VGND VGND VPWR VPWR _4081_/X sky130_fd_sc_hd__mux2_1
XFILLER_49_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4983_ _4983_/A1 _5040_/B _4941_/Y _4982_/X VGND VGND VPWR VPWR _6722_/D sky130_fd_sc_hd__o22a_1
XFILLER_51_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6722_ _7150_/CLK _6722_/D _4181_/B VGND VGND VPWR VPWR _6722_/Q sky130_fd_sc_hd__dfrtp_1
X_3934_ _7105_/Q _6758_/Q _6762_/Q VGND VGND VPWR VPWR _3934_/X sky130_fd_sc_hd__mux2_1
X_3865_ _3259_/B _3826_/A _3864_/X _3825_/B _6402_/Q VGND VGND VPWR VPWR _6402_/D
+ sky130_fd_sc_hd__a32o_1
X_6653_ _7155_/CLK hold64/X _6370_/A VGND VGND VPWR VPWR _6653_/Q sky130_fd_sc_hd__dfrtp_4
X_5604_ _3876_/A _5610_/A _5564_/Y _5603_/Y VGND VGND VPWR VPWR _5605_/B sky130_fd_sc_hd__a31o_1
XFILLER_118_711 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3796_ _6898_/Q _5334_/A _4214_/A _6619_/Q _3795_/X VGND VGND VPWR VPWR _3802_/B
+ sky130_fd_sc_hd__a221o_1
X_6584_ _7137_/CLK _6584_/D VGND VGND VPWR VPWR _6584_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_191_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5535_ hold189/X hold142/X _5537_/S VGND VGND VPWR VPWR _5535_/X sky130_fd_sc_hd__mux2_1
XFILLER_11_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_703 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5466_ hold687/X _5544_/A1 _5468_/S VGND VGND VPWR VPWR _5466_/X sky130_fd_sc_hd__mux2_1
XFILLER_160_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_172_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4417_ _4596_/B _4417_/B VGND VGND VPWR VPWR _4944_/A sky130_fd_sc_hd__nor2_2
XFILLER_160_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5397_ _5397_/A _5538_/B VGND VGND VPWR VPWR _5405_/S sky130_fd_sc_hd__and2_4
XFILLER_59_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7136_ _7140_/CLK _7136_/D VGND VGND VPWR VPWR _7136_/Q sky130_fd_sc_hd__dfxtp_1
X_4348_ _4450_/A _4590_/A VGND VGND VPWR VPWR _4901_/A sky130_fd_sc_hd__or2_4
XFILLER_99_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7067_ _7067_/CLK _7067_/D fanout513/X VGND VGND VPWR VPWR _7067_/Q sky130_fd_sc_hd__dfrtp_1
X_4279_ _4279_/A _5187_/B VGND VGND VPWR VPWR _4284_/S sky130_fd_sc_hd__and2_4
XFILLER_101_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_219 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6018_ _6883_/Q _5973_/A _5971_/B _6859_/Q _6017_/X VGND VGND VPWR VPWR _6026_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_39_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_655 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_167_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_109_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_163_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_235 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_408 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_159_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_174_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3650_ _6908_/Q _5343_/A _4038_/A _6482_/Q _3637_/X VGND VGND VPWR VPWR _3650_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_158_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_173_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3581_ input46/X _4103_/B _5520_/A _7066_/Q VGND VGND VPWR VPWR _3581_/X sky130_fd_sc_hd__a22o_1
X_5320_ hold349/X _5515_/A1 hold84/X VGND VGND VPWR VPWR _5320_/X sky130_fd_sc_hd__mux2_1
XFILLER_54_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_680 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5251_ hold632/X _5545_/A1 _5252_/S VGND VGND VPWR VPWR _5251_/X sky130_fd_sc_hd__mux2_1
XFILLER_114_235 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4202_ _4202_/A hold7/X VGND VGND VPWR VPWR _4207_/S sky130_fd_sc_hd__and2_4
X_5182_ _5530_/A1 hold781/X _5182_/S VGND VGND VPWR VPWR _5182_/X sky130_fd_sc_hd__mux2_1
XFILLER_96_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4133_ _4133_/A hold7/X VGND VGND VPWR VPWR _4138_/S sky130_fd_sc_hd__and2_4
XFILLER_68_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4064_ _4064_/A0 _4063_/X _4078_/S VGND VGND VPWR VPWR _4064_/X sky130_fd_sc_hd__mux2_1
XFILLER_83_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_211 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4966_ _4719_/B _4676_/B _4973_/B VGND VGND VPWR VPWR _4966_/X sky130_fd_sc_hd__a21o_1
X_6705_ _6707_/CLK _6705_/D fanout486/X VGND VGND VPWR VPWR _6705_/Q sky130_fd_sc_hd__dfrtp_1
X_3917_ _6518_/Q input80/X _3951_/B VGND VGND VPWR VPWR _3917_/X sky130_fd_sc_hd__mux2_8
X_4897_ _4894_/B _4885_/A _4737_/B _4885_/B _4739_/Y VGND VGND VPWR VPWR _5105_/A
+ sky130_fd_sc_hd__o41a_1
XFILLER_165_603 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6636_ _7150_/CLK _6636_/D _6308_/B VGND VGND VPWR VPWR _6636_/Q sky130_fd_sc_hd__dfrtp_4
X_3848_ hold37/A _6488_/Q _3841_/B _3847_/X VGND VGND VPWR VPWR _3848_/X sky130_fd_sc_hd__a22o_1
XFILLER_177_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_164_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3779_ _6555_/Q _4139_/A _4151_/A _6565_/Q VGND VGND VPWR VPWR _3779_/X sky130_fd_sc_hd__a22o_1
X_6567_ _6633_/CLK _6567_/D fanout509/X VGND VGND VPWR VPWR _6567_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_138_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_192_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5518_ hold592/X _5545_/A1 _5519_/S VGND VGND VPWR VPWR _5518_/X sky130_fd_sc_hd__mux2_1
X_6498_ _6707_/CLK _6498_/D fanout486/X VGND VGND VPWR VPWR _6498_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_145_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5449_ hold465/X hold114/X _5450_/S VGND VGND VPWR VPWR _5449_/X sky130_fd_sc_hd__mux2_1
XFILLER_78_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_120_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7119_ _7123_/CLK _7119_/D fanout499/X VGND VGND VPWR VPWR _7119_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_87_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_1__f_wbbd_sck clkbuf_0_wbbd_sck/X VGND VGND VPWR VPWR _3936_/A2 sky130_fd_sc_hd__clkbuf_16
XFILLER_179_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_188_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_491 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_127 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_8 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_151_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4820_ _5067_/A _4820_/B _4984_/B _4984_/A VGND VGND VPWR VPWR _4821_/D sky130_fd_sc_hd__and4b_1
XTAP_2391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4751_ _4885_/A _4465_/B _4901_/B _4523_/A VGND VGND VPWR VPWR _4751_/Y sky130_fd_sc_hd__o31ai_1
XFILLER_193_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3702_ _6686_/Q _4285_/A _4121_/A _6541_/Q VGND VGND VPWR VPWR _3702_/X sky130_fd_sc_hd__a22o_1
X_4682_ _4965_/A _4965_/B VGND VGND VPWR VPWR _4683_/B sky130_fd_sc_hd__and2_1
XFILLER_119_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3633_ input26/X _3339_/Y _4121_/A _6542_/Q VGND VGND VPWR VPWR _3633_/X sky130_fd_sc_hd__a22o_1
X_6421_ _6994_/CLK _6421_/D fanout489/X VGND VGND VPWR VPWR _6421_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_146_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_319 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6352_ _6352_/A _6352_/B VGND VGND VPWR VPWR hold54/A sky130_fd_sc_hd__and2_2
X_3564_ _6438_/Q _3984_/A _4303_/A _6704_/Q _3562_/X VGND VGND VPWR VPWR _3565_/D
+ sky130_fd_sc_hd__a221o_2
XFILLER_108_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_161_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5303_ _5303_/A0 _5465_/A1 _5306_/S VGND VGND VPWR VPWR _5303_/X sky130_fd_sc_hd__mux2_1
X_6283_ _6684_/Q _6283_/A2 _5981_/X _6679_/Q _6282_/X VGND VGND VPWR VPWR _6293_/A
+ sky130_fd_sc_hd__a221o_1
X_3495_ _6422_/Q _3958_/A _3360_/Y input7/X _3494_/X VGND VGND VPWR VPWR _3502_/B
+ sky130_fd_sc_hd__a221o_4
XFILLER_170_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5234_ hold658/X _5537_/A1 _5234_/S VGND VGND VPWR VPWR _5234_/X sky130_fd_sc_hd__mux2_1
XFILLER_69_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5165_ _5165_/A0 _5495_/A1 _5167_/S VGND VGND VPWR VPWR _5165_/X sky130_fd_sc_hd__mux2_1
XFILLER_130_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4116_ hold180/X _5533_/A1 _4120_/S VGND VGND VPWR VPWR _4116_/X sky130_fd_sc_hd__mux2_1
XFILLER_69_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5096_ _4587_/A _5026_/B _5037_/A _5095_/X VGND VGND VPWR VPWR _5134_/A sky130_fd_sc_hd__o211ai_1
XFILLER_84_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_678 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4047_ _4047_/A0 _4046_/X _4061_/S VGND VGND VPWR VPWR _4047_/X sky130_fd_sc_hd__mux2_1
XFILLER_37_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_553 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5998_ _6938_/Q _5942_/X _5973_/C _6874_/Q _5984_/X VGND VGND VPWR VPWR _5998_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_24_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4949_ _5025_/A _4947_/B _4566_/B VGND VGND VPWR VPWR _4949_/X sky130_fd_sc_hd__a21o_1
XFILLER_33_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_137_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6619_ _6686_/CLK _6619_/D fanout492/X VGND VGND VPWR VPWR _6619_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_193_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_192_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput280 _6420_/Q VGND VGND VPWR VPWR pll_trim[18] sky130_fd_sc_hd__buf_12
Xoutput291 _6438_/Q VGND VGND VPWR VPWR pll_trim[4] sky130_fd_sc_hd__buf_12
XFILLER_121_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_604 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_188_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_169_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_400 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_444 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_171_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3280_ hold78/X _3247_/A _3856_/S VGND VGND VPWR VPWR hold79/A sky130_fd_sc_hd__mux2_1
XTAP_726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_612 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6970_ _7010_/CLK _6970_/D fanout498/X VGND VGND VPWR VPWR _6970_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_19_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_626 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5921_ _6479_/Q _5921_/A2 _5644_/X _6454_/Q VGND VGND VPWR VPWR _5921_/X sky130_fd_sc_hd__a22o_1
XFILLER_179_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5852_ _7035_/Q _5645_/X _5649_/X _6676_/Q VGND VGND VPWR VPWR _5852_/X sky130_fd_sc_hd__a22o_1
XFILLER_34_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4803_ _4513_/A _4921_/A _5043_/B _4973_/A VGND VGND VPWR VPWR _4817_/C sky130_fd_sc_hd__o22a_1
XFILLER_21_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5783_ _7016_/Q _5921_/A2 _5915_/A2 _6960_/Q _5781_/X VGND VGND VPWR VPWR _5783_/X
+ sky130_fd_sc_hd__a221o_1
X_4734_ _4721_/B _4715_/B _4520_/X VGND VGND VPWR VPWR _4734_/X sky130_fd_sc_hd__o21a_1
XFILLER_119_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4665_ _4732_/A _5061_/A _4665_/C _4665_/D VGND VGND VPWR VPWR _4666_/C sky130_fd_sc_hd__and4b_1
XFILLER_190_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_162_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6404_ _7171_/CLK _6404_/D _6360_/X VGND VGND VPWR VPWR _6404_/Q sky130_fd_sc_hd__dfrtp_4
Xhold900 _4323_/X VGND VGND VPWR VPWR _6716_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3616_ _6789_/Q _5208_/A _4038_/A _6483_/Q _3615_/X VGND VGND VPWR VPWR _3623_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_174_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_190_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold911 _6897_/Q VGND VGND VPWR VPWR hold911/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold922 _4153_/X VGND VGND VPWR VPWR _6566_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4596_ _4746_/A _4596_/B _4595_/B VGND VGND VPWR VPWR _4725_/B sky130_fd_sc_hd__or3b_4
Xhold933 _6620_/Q VGND VGND VPWR VPWR hold933/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold944 _5489_/X VGND VGND VPWR VPWR _7035_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6335_ _6642_/Q _6335_/A2 _6335_/B1 _4222_/B VGND VGND VPWR VPWR _6335_/X sky130_fd_sc_hd__a22o_1
X_3547_ _6757_/Q _5179_/B _4237_/A _6649_/Q _3546_/X VGND VGND VPWR VPWR _3548_/C
+ sky130_fd_sc_hd__a221o_4
Xhold955 _6971_/Q VGND VGND VPWR VPWR hold955/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold966 _5459_/X VGND VGND VPWR VPWR _7009_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_103_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold977 _6711_/Q VGND VGND VPWR VPWR hold977/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold988 _6939_/Q VGND VGND VPWR VPWR hold988/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_88_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3478_ hold61/X _5183_/B VGND VGND VPWR VPWR hold62/A sky130_fd_sc_hd__nor2_8
Xhold999 _4287_/X VGND VGND VPWR VPWR _6686_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6266_ _6693_/Q _5972_/B _5959_/Y _6617_/Q _6265_/X VGND VGND VPWR VPWR _6267_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_170_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5217_ _5217_/A _5511_/B VGND VGND VPWR VPWR _5225_/S sky130_fd_sc_hd__and2_4
X_6197_ _7034_/Q _6295_/A2 _5973_/C _6619_/Q _6196_/X VGND VGND VPWR VPWR _6200_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_69_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5148_ hold785/X _6355_/A1 _5150_/S VGND VGND VPWR VPWR _5148_/X sky130_fd_sc_hd__mux2_1
XFILLER_151_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5079_ _5079_/A _5106_/B VGND VGND VPWR VPWR _5079_/Y sky130_fd_sc_hd__nand2_1
XFILLER_44_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_704 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_193_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_403 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_436 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_180_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_82 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_604 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_534 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_144_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_172_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4450_ _4450_/A _4632_/A VGND VGND VPWR VPWR _4471_/B sky130_fd_sc_hd__nand2_1
Xhold207 _6779_/Q VGND VGND VPWR VPWR hold207/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_156_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold218 _5174_/X VGND VGND VPWR VPWR _6758_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_171_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold229 _6754_/Q VGND VGND VPWR VPWR hold229/X sky130_fd_sc_hd__dlygate4sd3_1
X_3401_ hold39/X _3401_/B hold51/X VGND VGND VPWR VPWR hold52/A sky130_fd_sc_hd__or3b_4
X_4381_ _4617_/B _4613_/C VGND VGND VPWR VPWR _4383_/C sky130_fd_sc_hd__and2_1
X_3332_ _3571_/A _3706_/A VGND VGND VPWR VPWR _5538_/A sky130_fd_sc_hd__nor2_8
X_6120_ _6903_/Q _6296_/B1 _5978_/X _6951_/Q _6119_/X VGND VGND VPWR VPWR _6127_/A
+ sky130_fd_sc_hd__a221o_1
XTAP_501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3263_ _6764_/Q _6813_/Q _3263_/C VGND VGND VPWR VPWR _3263_/Y sky130_fd_sc_hd__nor3_2
X_6051_ _6972_/Q _6282_/B1 _6048_/X _6050_/X VGND VGND VPWR VPWR _6052_/C sky130_fd_sc_hd__a211o_1
XTAP_556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_206 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5002_ _5067_/B _5002_/B _5131_/A _5001_/X VGND VGND VPWR VPWR _5003_/B sky130_fd_sc_hd__or4b_1
X_3194_ _6997_/Q VGND VGND VPWR VPWR _3194_/Y sky130_fd_sc_hd__inv_2
XFILLER_78_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_434 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6953_ _7078_/CLK _6953_/D fanout507/X VGND VGND VPWR VPWR _6953_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_53_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5904_ _6617_/Q _5928_/B1 _5913_/B1 _6628_/Q VGND VGND VPWR VPWR _5904_/X sky130_fd_sc_hd__a22o_1
X_6884_ _7083_/CLK _6884_/D fanout518/X VGND VGND VPWR VPWR _6884_/Q sky130_fd_sc_hd__dfrtp_2
X_5835_ _6655_/Q _5923_/B VGND VGND VPWR VPWR _5835_/X sky130_fd_sc_hd__and2b_1
XFILLER_14_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_528 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5766_ _6983_/Q _5642_/X _5807_/B1 _6935_/Q _5758_/Y VGND VGND VPWR VPWR _5766_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_148_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4717_ _4717_/A _4717_/B VGND VGND VPWR VPWR _4718_/C sky130_fd_sc_hd__nor2_1
XFILLER_175_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5697_ _5667_/B _5693_/X _5642_/X _6980_/Q VGND VGND VPWR VPWR _5697_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_175_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4648_ _4922_/B _4915_/A _4648_/C _4648_/D VGND VGND VPWR VPWR _4666_/B sky130_fd_sc_hd__and4b_1
XFILLER_135_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold730 _5403_/X VGND VGND VPWR VPWR _6959_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold741 _6941_/Q VGND VGND VPWR VPWR hold741/X sky130_fd_sc_hd__dlygate4sd3_1
X_4579_ _4579_/A _4579_/B _4579_/C _5110_/A VGND VGND VPWR VPWR _4579_/X sky130_fd_sc_hd__and4_1
Xhold752 _5497_/X VGND VGND VPWR VPWR _7042_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold763 _6853_/Q VGND VGND VPWR VPWR hold763/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold774 _4306_/X VGND VGND VPWR VPWR _6702_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6318_ _6320_/B _6318_/B VGND VGND VPWR VPWR _6318_/Y sky130_fd_sc_hd__nand2_1
Xhold785 _6739_/Q VGND VGND VPWR VPWR hold785/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_1_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold796 _3987_/X VGND VGND VPWR VPWR _6436_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_131_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6249_ _6601_/Q _5939_/X _5953_/Y _6482_/Q _6248_/X VGND VGND VPWR VPWR _6250_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_39_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1430 _6722_/Q VGND VGND VPWR VPWR _4983_/A1 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1441 _6732_/Q VGND VGND VPWR VPWR _3473_/A1 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1452 _6575_/Q VGND VGND VPWR VPWR _4163_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_57_464 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1463 _7144_/Q VGND VGND VPWR VPWR _6334_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_45_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1474 _7120_/Q VGND VGND VPWR VPWR _6054_/A2 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_72_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_61_csclk clkbuf_3_2_0_csclk/X VGND VGND VPWR VPWR _6976_/CLK sky130_fd_sc_hd__clkbuf_16
Xhold1485 hold44/A VGND VGND VPWR VPWR _3254_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1496 _7125_/Q VGND VGND VPWR VPWR _6179_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_84_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_659 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_76_csclk _6661_/CLK VGND VGND VPWR VPWR _7034_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_9_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_139_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_141_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_14_csclk clkbuf_3_5_0_csclk/X VGND VGND VPWR VPWR _7067_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_96_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold90 hold90/A VGND VGND VPWR VPWR hold90/X sky130_fd_sc_hd__clkbuf_16
Xclkbuf_leaf_29_csclk clkbuf_3_7_0_csclk/X VGND VGND VPWR VPWR _7082_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_91_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3950_ _3950_/A _3950_/B VGND VGND VPWR VPWR _3950_/X sky130_fd_sc_hd__and2_1
XFILLER_50_128 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3881_ _5610_/A _3887_/B _5609_/B VGND VGND VPWR VPWR _6507_/D sky130_fd_sc_hd__o21ai_1
XFILLER_149_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5620_ _5667_/A _5643_/B _5650_/B VGND VGND VPWR VPWR _5620_/X sky130_fd_sc_hd__and3_4
XFILLER_84_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5551_ _7088_/Q _5558_/D VGND VGND VPWR VPWR _5554_/A sky130_fd_sc_hd__or2_1
XFILLER_157_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4502_ _4471_/A _4885_/A _4965_/A _4501_/X VGND VGND VPWR VPWR _4503_/B sky130_fd_sc_hd__o31a_1
X_5482_ hold745/X _5542_/A1 _5486_/S VGND VGND VPWR VPWR _5482_/X sky130_fd_sc_hd__mux2_1
XFILLER_117_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4433_ _4596_/B _4746_/B _4554_/A VGND VGND VPWR VPWR _4965_/A sky130_fd_sc_hd__or3b_4
XFILLER_172_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7152_ _7153_/CLK _7152_/D _3940_/B VGND VGND VPWR VPWR _7152_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_116_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4364_ _4542_/A _4679_/A VGND VGND VPWR VPWR _4570_/B sky130_fd_sc_hd__nand2b_4
Xfanout506 fanout507/X VGND VGND VPWR VPWR fanout506/X sky130_fd_sc_hd__buf_8
X_6103_ _6790_/Q _6004_/B _6093_/X _6102_/X _3174_/Y VGND VGND VPWR VPWR _6103_/X
+ sky130_fd_sc_hd__o221a_4
Xfanout517 fanout525/X VGND VGND VPWR VPWR fanout517/X sky130_fd_sc_hd__buf_8
X_3315_ hold31/X hold59/X VGND VGND VPWR VPWR _3328_/B sky130_fd_sc_hd__nor2_2
Xfanout528 input164/X VGND VGND VPWR VPWR _4181_/B sky130_fd_sc_hd__clkbuf_16
XFILLER_112_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4295_ hold171/X hold46/X _4296_/S VGND VGND VPWR VPWR _4295_/X sky130_fd_sc_hd__mux2_1
X_7083_ _7083_/CLK _7083_/D fanout517/X VGND VGND VPWR VPWR _7083_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_112_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3246_ _3246_/A _3246_/B VGND VGND VPWR VPWR _7168_/D sky130_fd_sc_hd__xnor2_1
X_6034_ _7065_/Q _6283_/A2 _6296_/B1 _6900_/Q VGND VGND VPWR VPWR _6034_/X sky130_fd_sc_hd__a22o_1
XTAP_397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3177_ _4334_/B VGND VGND VPWR VPWR _3177_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_54_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6936_ _7042_/CLK _6936_/D fanout523/X VGND VGND VPWR VPWR _6936_/Q sky130_fd_sc_hd__dfrtp_2
XPHY_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_139 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_180 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6867_ _7074_/CLK _6867_/D fanout505/X VGND VGND VPWR VPWR _6867_/Q sky130_fd_sc_hd__dfstp_1
X_5818_ _6969_/Q _5925_/B1 _5650_/X _6897_/Q VGND VGND VPWR VPWR _5818_/X sky130_fd_sc_hd__a22o_1
X_6798_ _6988_/CLK _6798_/D _6396_/A VGND VGND VPWR VPWR _6798_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_10_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5749_ _6902_/Q _5623_/X _5625_/X _6870_/Q _5748_/X VGND VGND VPWR VPWR _5754_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_182_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_182_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold560 _4281_/X VGND VGND VPWR VPWR _6681_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold571 _6659_/Q VGND VGND VPWR VPWR hold571/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold582 _4012_/X VGND VGND VPWR VPWR _6458_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold593 _5518_/X VGND VGND VPWR VPWR _7061_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_173_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1260 _4256_/X VGND VGND VPWR VPWR _6660_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_18_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1271 _6518_/Q VGND VGND VPWR VPWR _4097_/A0 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1282 _4064_/X VGND VGND VPWR VPWR _6498_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_85_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1293 _6846_/Q VGND VGND VPWR VPWR _5276_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_122 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_186_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_185_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_99_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_288 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_141_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4080_ _5200_/A0 hold588/X _4092_/S VGND VGND VPWR VPWR _4080_/X sky130_fd_sc_hd__mux2_1
XFILLER_64_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4982_ _5020_/B _4914_/Y _4981_/X VGND VGND VPWR VPWR _4982_/X sky130_fd_sc_hd__a21o_1
X_6721_ _3931_/A1 _6721_/D _4181_/B VGND VGND VPWR VPWR _6721_/Q sky130_fd_sc_hd__dfrtp_1
X_3933_ _7103_/Q _6759_/Q _6762_/Q VGND VGND VPWR VPWR _3933_/X sky130_fd_sc_hd__mux2_1
XFILLER_51_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6652_ _7155_/CLK _6652_/D _6370_/A VGND VGND VPWR VPWR _6652_/Q sky130_fd_sc_hd__dfstp_1
X_3864_ _7170_/Q _6402_/Q _6485_/Q VGND VGND VPWR VPWR _3864_/X sky130_fd_sc_hd__o21ba_1
X_5603_ _5607_/C _5555_/Y _3876_/A VGND VGND VPWR VPWR _5603_/Y sky130_fd_sc_hd__a21oi_1
X_6583_ _7137_/CLK _6583_/D VGND VGND VPWR VPWR _6583_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_118_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3795_ _6874_/Q _5307_/A _4249_/A _6655_/Q VGND VGND VPWR VPWR _3795_/X sky130_fd_sc_hd__a22o_1
XFILLER_118_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5534_ hold297/X _5534_/A1 _5537_/S VGND VGND VPWR VPWR _5534_/X sky130_fd_sc_hd__mux2_1
XFILLER_8_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_191_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_715 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5465_ _5465_/A0 _5465_/A1 _5468_/S VGND VGND VPWR VPWR _5465_/X sky130_fd_sc_hd__mux2_1
X_4416_ _4419_/B _4416_/B _4535_/A VGND VGND VPWR VPWR _4479_/A sky130_fd_sc_hd__or3b_4
X_5396_ hold677/X _5537_/A1 _5396_/S VGND VGND VPWR VPWR _5396_/X sky130_fd_sc_hd__mux2_1
XFILLER_132_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7135_ _7140_/CLK _7135_/D VGND VGND VPWR VPWR _7135_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_113_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_160_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4347_ _4368_/A _4499_/B VGND VGND VPWR VPWR _4590_/A sky130_fd_sc_hd__or2_2
XFILLER_86_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7066_ _7067_/CLK _7066_/D _3264_/A VGND VGND VPWR VPWR _7066_/Q sky130_fd_sc_hd__dfrtp_2
X_4278_ hold303/X _6357_/A1 _4278_/S VGND VGND VPWR VPWR _4278_/X sky130_fd_sc_hd__mux2_1
X_6017_ _6835_/Q _5946_/X _5971_/A _6867_/Q VGND VGND VPWR VPWR _6017_/X sky130_fd_sc_hd__a22o_1
X_3229_ _3247_/A _3229_/A1 _3229_/S VGND VGND VPWR VPWR _7171_/D sky130_fd_sc_hd__mux2_1
XFILLER_100_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_0__f_wbbd_sck clkbuf_0_wbbd_sck/X VGND VGND VPWR VPWR _6347_/A1 sky130_fd_sc_hd__clkbuf_16
XTAP_1327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6919_ _7046_/CLK _6919_/D fanout503/X VGND VGND VPWR VPWR _6919_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_23_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_155_306 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_108_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_247 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold390 _3989_/X VGND VGND VPWR VPWR _6438_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_37_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_378 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1090 _4280_/X VGND VGND VPWR VPWR _6680_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_93_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_93_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_155 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3580_ _6869_/Q _5298_/A hold62/A _6653_/Q _3579_/X VGND VGND VPWR VPWR _3625_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_173_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_173_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_173_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_142_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5250_ hold683/X _5544_/A1 _5252_/S VGND VGND VPWR VPWR _5250_/X sky130_fd_sc_hd__mux2_1
XFILLER_47_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4201_ hold405/X _5534_/A1 _4201_/S VGND VGND VPWR VPWR _4201_/X sky130_fd_sc_hd__mux2_1
XFILLER_130_718 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5181_ _5181_/A _5529_/B VGND VGND VPWR VPWR _5182_/S sky130_fd_sc_hd__nand2_1
XFILLER_96_610 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4132_ hold431/X _5534_/A1 _4132_/S VGND VGND VPWR VPWR _4132_/X sky130_fd_sc_hd__mux2_1
XFILLER_110_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4063_ _4113_/A0 _6353_/A1 _4112_/B VGND VGND VPWR VPWR _4063_/X sky130_fd_sc_hd__mux2_1
XFILLER_110_486 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4965_ _4965_/A _4965_/B _4965_/C VGND VGND VPWR VPWR _4973_/B sky130_fd_sc_hd__and3_2
X_6704_ _7034_/CLK _6704_/D fanout488/X VGND VGND VPWR VPWR _6704_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_51_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_149_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3916_ _3185_/Y input82/X _3951_/B VGND VGND VPWR VPWR _3916_/X sky130_fd_sc_hd__mux2_8
XFILLER_177_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4896_ _4901_/B _4719_/B _4895_/Y _4774_/A VGND VGND VPWR VPWR _4906_/A sky130_fd_sc_hd__o211a_1
XFILLER_149_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6635_ _7150_/CLK _6635_/D _6308_/B VGND VGND VPWR VPWR _6635_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_22_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3847_ hold48/A _3847_/B VGND VGND VPWR VPWR _3847_/X sky130_fd_sc_hd__or2_1
XFILLER_165_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_165_637 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6566_ _6630_/CLK _6566_/D fanout496/X VGND VGND VPWR VPWR _6566_/Q sky130_fd_sc_hd__dfrtp_1
X_3778_ _3778_/A _3778_/B _3778_/C wire347/X VGND VGND VPWR VPWR _3816_/B sky130_fd_sc_hd__or4b_1
XFILLER_164_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5517_ hold693/X _5544_/A1 _5519_/S VGND VGND VPWR VPWR _5517_/X sky130_fd_sc_hd__mux2_1
XFILLER_145_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6497_ _7082_/CLK _6497_/D fanout519/X VGND VGND VPWR VPWR _7188_/A sky130_fd_sc_hd__dfrtp_1
XFILLER_105_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_160_320 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5448_ hold671/X _5544_/A1 _5450_/S VGND VGND VPWR VPWR _5448_/X sky130_fd_sc_hd__mux2_1
XFILLER_105_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_154_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5379_ _5379_/A _5529_/B VGND VGND VPWR VPWR _5387_/S sky130_fd_sc_hd__and2_4
XFILLER_160_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7118_ _7130_/CLK _7118_/D fanout488/X VGND VGND VPWR VPWR _7118_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_87_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7049_ _7075_/CLK _7049_/D fanout514/X VGND VGND VPWR VPWR _7049_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_47_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_155_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_179_707 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_256 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_239 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4750_ _4977_/B _4692_/C _4965_/B _4549_/B _4622_/A VGND VGND VPWR VPWR _4912_/A
+ sky130_fd_sc_hd__o32a_1
XTAP_1691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3701_ _6915_/Q _5352_/A _5226_/A _6803_/Q _3700_/X VGND VGND VPWR VPWR _3712_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_186_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4681_ _4965_/B _4630_/B _4576_/X _5021_/B VGND VGND VPWR VPWR _4681_/X sky130_fd_sc_hd__o211a_1
X_6420_ _6994_/CLK _6420_/D fanout489/X VGND VGND VPWR VPWR _6420_/Q sky130_fd_sc_hd__dfstp_1
X_3632_ _6788_/Q _5208_/A _3384_/Y input22/X VGND VGND VPWR VPWR _3632_/X sky130_fd_sc_hd__a22o_1
XFILLER_174_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_134_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6351_ _3168_/A _6351_/A2 _5040_/B _6350_/X VGND VGND VPWR VPWR _7150_/D sky130_fd_sc_hd__o31a_1
X_3563_ _3563_/A _3761_/B VGND VGND VPWR VPWR _4303_/A sky130_fd_sc_hd__nor2_4
XFILLER_127_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5302_ hold343/X _5515_/A1 _5306_/S VGND VGND VPWR VPWR _5302_/X sky130_fd_sc_hd__mux2_1
X_6282_ _6484_/Q _6282_/A2 _6282_/B1 _6454_/Q _6281_/X VGND VGND VPWR VPWR _6282_/X
+ sky130_fd_sc_hd__a221o_1
X_3494_ _6902_/Q _5334_/A _3433_/A _3493_/Y VGND VGND VPWR VPWR _3494_/X sky130_fd_sc_hd__a211o_2
XFILLER_142_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5233_ hold473/X _5545_/A1 _5234_/S VGND VGND VPWR VPWR _5233_/X sky130_fd_sc_hd__mux2_1
Xclkbuf_opt_3_0_csclk _6684_/CLK VGND VGND VPWR VPWR clkbuf_opt_3_0_csclk/X sky130_fd_sc_hd__clkbuf_16
X_5164_ _5164_/A0 _5530_/A1 _5167_/S VGND VGND VPWR VPWR _5164_/X sky130_fd_sc_hd__mux2_1
XFILLER_124_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4115_ hold363/X _5532_/A1 _4120_/S VGND VGND VPWR VPWR _4115_/X sky130_fd_sc_hd__mux2_1
XFILLER_84_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5095_ _5022_/A _4479_/A _4506_/C _4933_/A VGND VGND VPWR VPWR _5095_/X sky130_fd_sc_hd__o211a_1
XFILLER_68_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4046_ hold893/X _5521_/A1 _4103_/B VGND VGND VPWR VPWR _4046_/X sky130_fd_sc_hd__mux2_1
XFILLER_17_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5997_ _7039_/Q _5969_/C _5983_/X _5992_/X _5996_/X VGND VGND VPWR VPWR _6003_/A
+ sky130_fd_sc_hd__a2111o_1
XFILLER_52_565 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4948_ _5025_/A _4557_/B _4851_/B VGND VGND VPWR VPWR _5121_/A sky130_fd_sc_hd__a21oi_2
XFILLER_178_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4879_ _5058_/A _4879_/B _4879_/C _4879_/D VGND VGND VPWR VPWR _4879_/X sky130_fd_sc_hd__and4b_1
XFILLER_20_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6618_ _6632_/CLK _6618_/D _3264_/A VGND VGND VPWR VPWR _6618_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_165_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_192_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6549_ _6746_/CLK _6549_/D fanout489/X VGND VGND VPWR VPWR _6549_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_106_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_161_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput270 _6744_/Q VGND VGND VPWR VPWR pll_sel[2] sky130_fd_sc_hd__buf_12
Xoutput281 _6421_/Q VGND VGND VPWR VPWR pll_trim[19] sky130_fd_sc_hd__buf_12
Xoutput292 _6439_/Q VGND VGND VPWR VPWR pll_trim[5] sky130_fd_sc_hd__buf_12
XFILLER_121_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_521 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_169_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_456 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_607 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_171_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_139_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_624 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_171_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5920_ _6569_/Q _5920_/A2 _5916_/X _5917_/X _5919_/X VGND VGND VPWR VPWR _5920_/X
+ sky130_fd_sc_hd__a2111o_1
XFILLER_81_638 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5851_ _6461_/Q _5642_/X _5648_/X _6716_/Q VGND VGND VPWR VPWR _5851_/X sky130_fd_sc_hd__a22o_1
XFILLER_34_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_548 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4802_ _4513_/A _4640_/B _4725_/B _4745_/B VGND VGND VPWR VPWR _4817_/B sky130_fd_sc_hd__o22a_1
X_5782_ _3223_/Y _5923_/B _5667_/B VGND VGND VPWR VPWR _5782_/Y sky130_fd_sc_hd__a21oi_1
X_4733_ _4733_/A VGND VGND VPWR VPWR _4902_/B sky130_fd_sc_hd__clkinv_2
X_4664_ _4664_/A _4664_/B _4664_/C _4664_/D VGND VGND VPWR VPWR _4665_/D sky130_fd_sc_hd__and4_1
XFILLER_119_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6403_ _7171_/CLK _6403_/D _6359_/X VGND VGND VPWR VPWR _6403_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_119_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3615_ _7005_/Q _5451_/A _5487_/A _7037_/Q VGND VGND VPWR VPWR _3615_/X sky130_fd_sc_hd__a22o_1
XFILLER_128_670 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold901 _6651_/Q VGND VGND VPWR VPWR hold901/X sky130_fd_sc_hd__dlygate4sd3_1
X_4595_ _4691_/A _4595_/B VGND VGND VPWR VPWR _4595_/Y sky130_fd_sc_hd__nand2_1
Xhold912 _5333_/X VGND VGND VPWR VPWR _6897_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold923 _6795_/Q VGND VGND VPWR VPWR hold923/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_190_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold934 _4216_/X VGND VGND VPWR VPWR _6620_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6334_ _6333_/X _6334_/A1 _6346_/S VGND VGND VPWR VPWR _7144_/D sky130_fd_sc_hd__mux2_1
X_3546_ input24/X _3384_/Y _4127_/A _6549_/Q VGND VGND VPWR VPWR _3546_/X sky130_fd_sc_hd__a22o_1
Xhold945 _7056_/Q VGND VGND VPWR VPWR hold945/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_127_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold956 _5417_/X VGND VGND VPWR VPWR _6971_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold967 _7033_/Q VGND VGND VPWR VPWR hold967/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold978 _4317_/X VGND VGND VPWR VPWR _6711_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold989 _5381_/X VGND VGND VPWR VPWR _6939_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6265_ _6628_/Q _5973_/A _5946_/X _6581_/Q VGND VGND VPWR VPWR _6265_/X sky130_fd_sc_hd__a22o_1
X_3477_ _6854_/Q _3374_/Y _4166_/A _6582_/Q _3476_/X VGND VGND VPWR VPWR _3489_/A
+ sky130_fd_sc_hd__a221o_1
X_5216_ hold435/X _5519_/A1 _5216_/S VGND VGND VPWR VPWR _5216_/X sky130_fd_sc_hd__mux2_1
XFILLER_103_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6196_ _6460_/Q _5943_/Y _5948_/X _6545_/Q VGND VGND VPWR VPWR _6196_/X sky130_fd_sc_hd__a22o_1
XFILLER_28_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5147_ hold929/X _6354_/A1 _5150_/S VGND VGND VPWR VPWR _5147_/X sky130_fd_sc_hd__mux2_1
XFILLER_29_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5078_ _4430_/C _4892_/B _4893_/Y _5077_/X _4741_/X VGND VGND VPWR VPWR _5106_/B
+ sky130_fd_sc_hd__o2111a_1
XFILLER_44_318 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4029_ hold845/X _5505_/A1 _4031_/S VGND VGND VPWR VPWR _4029_/X sky130_fd_sc_hd__mux2_1
XFILLER_13_716 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_161_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_87_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_307 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_156_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_172_735 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold208 _5201_/X VGND VGND VPWR VPWR _6779_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold219 _7001_/Q VGND VGND VPWR VPWR hold219/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_172_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3400_ _3706_/B _3487_/A VGND VGND VPWR VPWR _3433_/A sky130_fd_sc_hd__nor2_4
XFILLER_125_651 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4380_ _4592_/A _4409_/B VGND VGND VPWR VPWR _4435_/B sky130_fd_sc_hd__nand2_1
XFILLER_125_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3331_ _6793_/Q _5208_/A hold83/A _6889_/Q _3327_/X VGND VGND VPWR VPWR _3349_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_112_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6050_ _6444_/Q _5601_/Y _5978_/X _6948_/Q _6049_/X VGND VGND VPWR VPWR _6050_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_112_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3262_ _3904_/A2 _3260_/X _3862_/S _3247_/A VGND VGND VPWR VPWR _7158_/D sky130_fd_sc_hd__a22o_1
XTAP_557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5001_ _5001_/A _5062_/B _5070_/B _5110_/B VGND VGND VPWR VPWR _5001_/X sky130_fd_sc_hd__and4_1
XTAP_579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3193_ _7005_/Q VGND VGND VPWR VPWR _3193_/Y sky130_fd_sc_hd__inv_2
XFILLER_66_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6952_ _7017_/CLK _6952_/D fanout515/X VGND VGND VPWR VPWR _6952_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_81_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5903_ _6463_/Q _5642_/X _5644_/X _6453_/Q _5891_/Y VGND VGND VPWR VPWR _5903_/X
+ sky130_fd_sc_hd__a221o_1
X_6883_ _7029_/CLK _6883_/D fanout519/X VGND VGND VPWR VPWR _6883_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_179_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5834_ _6450_/Q _5644_/X _5919_/B1 _6630_/Q _5833_/X VGND VGND VPWR VPWR _5842_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_61_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5765_ _7015_/Q _5921_/A2 _5760_/X _5763_/X _5764_/X VGND VGND VPWR VPWR _5765_/X
+ sky130_fd_sc_hd__a2111o_1
X_4716_ _4606_/Y _4673_/Y _4714_/X _4715_/Y VGND VGND VPWR VPWR _4718_/B sky130_fd_sc_hd__a211o_1
X_5696_ _6948_/Q _5924_/B2 _5912_/B1 _7028_/Q _5695_/X VGND VGND VPWR VPWR _5696_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_148_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4647_ _4575_/X _4745_/B _4676_/B _4725_/B _4646_/X VGND VGND VPWR VPWR _4648_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_162_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_190_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold720 _5367_/X VGND VGND VPWR VPWR _6927_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4578_ _4828_/A _4640_/B VGND VGND VPWR VPWR _5110_/A sky130_fd_sc_hd__or2_1
Xhold731 _6903_/Q VGND VGND VPWR VPWR hold731/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_162_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold742 _5383_/X VGND VGND VPWR VPWR _6941_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_122_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold753 _6482_/Q VGND VGND VPWR VPWR hold753/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold764 _5284_/X VGND VGND VPWR VPWR _6853_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6317_ _6320_/B _6317_/A2 _6640_/Q VGND VGND VPWR VPWR _6317_/X sky130_fd_sc_hd__a21bo_1
XFILLER_103_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3529_ _3531_/A _3554_/B VGND VGND VPWR VPWR _4151_/A sky130_fd_sc_hd__nor2_8
XFILLER_143_470 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold775 _6647_/Q VGND VGND VPWR VPWR hold775/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold786 _5148_/X VGND VGND VPWR VPWR _6739_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold797 _6611_/Q VGND VGND VPWR VPWR hold797/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_103_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6248_ _6557_/Q _6259_/A2 _5972_/A _6652_/Q VGND VGND VPWR VPWR _6248_/X sky130_fd_sc_hd__a22o_1
XFILLER_131_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6179_ _6179_/A1 _3878_/Y _5610_/Y VGND VGND VPWR VPWR _6179_/X sky130_fd_sc_hd__o21a_1
XFILLER_162_59 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1420 _6571_/Q VGND VGND VPWR VPWR _4159_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_130_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1431 _5405_/S VGND VGND VPWR VPWR _5399_/S sky130_fd_sc_hd__dlygate4sd3_1
Xhold1442 _3473_/X VGND VGND VPWR VPWR _6732_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1453 _6572_/Q VGND VGND VPWR VPWR _4160_/A1 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1464 _6624_/Q VGND VGND VPWR VPWR _3959_/S sky130_fd_sc_hd__dlygate4sd3_1
Xhold1475 _7109_/Q VGND VGND VPWR VPWR _5756_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_57_476 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1486 _3253_/X VGND VGND VPWR VPWR _7163_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1497 _7112_/Q VGND VGND VPWR VPWR _5801_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_187_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_187_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_187_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_154_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_71 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_131 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold80 hold80/A VGND VGND VPWR VPWR hold80/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_75_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold91 hold91/A VGND VGND VPWR VPWR hold91/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_152_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3880_ _5605_/A _3880_/B VGND VGND VPWR VPWR _3887_/B sky130_fd_sc_hd__nor2_1
XFILLER_189_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_188_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5550_ _5558_/D VGND VGND VPWR VPWR _5550_/Y sky130_fd_sc_hd__inv_2
XFILLER_77_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4501_ _5043_/A _4501_/B VGND VGND VPWR VPWR _4501_/X sky130_fd_sc_hd__or2_1
XFILLER_157_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5481_ hold100/X hold3/X _5486_/S VGND VGND VPWR VPWR _5481_/X sky130_fd_sc_hd__mux2_1
XFILLER_172_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4432_ _4554_/A _4691_/A _4448_/A VGND VGND VPWR VPWR _4677_/B sky130_fd_sc_hd__and3_2
XFILLER_144_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7151_ _7153_/CLK _7151_/D _3940_/B VGND VGND VPWR VPWR _7151_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_125_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4363_ _4883_/A VGND VGND VPWR VPWR _4363_/Y sky130_fd_sc_hd__inv_2
Xfanout507 fanout526/X VGND VGND VPWR VPWR fanout507/X sky130_fd_sc_hd__buf_8
X_6102_ _6102_/A _6102_/B _6102_/C _6004_/B VGND VGND VPWR VPWR _6102_/X sky130_fd_sc_hd__or4b_1
X_3314_ _3571_/B hold61/X VGND VGND VPWR VPWR _5352_/A sky130_fd_sc_hd__nor2_8
Xfanout518 fanout520/X VGND VGND VPWR VPWR fanout518/X sky130_fd_sc_hd__buf_8
X_7082_ _7082_/CLK _7082_/D fanout520/X VGND VGND VPWR VPWR _7082_/Q sky130_fd_sc_hd__dfrtp_4
Xfanout529 _4779_/A VGND VGND VPWR VPWR _4613_/C sky130_fd_sc_hd__clkbuf_8
XFILLER_98_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4294_ hold341/X _5523_/A1 _4296_/S VGND VGND VPWR VPWR _4294_/X sky130_fd_sc_hd__mux2_1
X_6033_ _6908_/Q _5972_/A _6282_/A2 _6996_/Q _6032_/X VGND VGND VPWR VPWR _6043_/A
+ sky130_fd_sc_hd__a221o_1
X_3245_ _3245_/A _3245_/B VGND VGND VPWR VPWR _3246_/B sky130_fd_sc_hd__nor2_1
XFILLER_112_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3176_ _7101_/Q VGND VGND VPWR VPWR _5940_/B sky130_fd_sc_hd__clkinv_2
XFILLER_132_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6935_ _7086_/CLK _6935_/D fanout516/X VGND VGND VPWR VPWR _6935_/Q sky130_fd_sc_hd__dfrtp_1
XPHY_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6866_ _7075_/CLK _6866_/D fanout505/X VGND VGND VPWR VPWR _6866_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_34_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5817_ _5817_/A _5817_/B VGND VGND VPWR VPWR _5817_/X sky130_fd_sc_hd__or2_1
X_6797_ _7046_/CLK _6797_/D fanout500/X VGND VGND VPWR VPWR _6797_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_167_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5748_ _5667_/B _5747_/X _5644_/X _6974_/Q VGND VGND VPWR VPWR _5748_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_157_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5679_ _6923_/Q _5633_/X _5646_/X _6995_/Q VGND VGND VPWR VPWR _5679_/X sky130_fd_sc_hd__a22o_1
XFILLER_136_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold550 _4125_/X VGND VGND VPWR VPWR _6543_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_173_14 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold561 _6708_/Q VGND VGND VPWR VPWR hold561/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_1_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold572 _4254_/X VGND VGND VPWR VPWR _6659_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold583 _6698_/Q VGND VGND VPWR VPWR hold583/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold594 _7008_/Q VGND VGND VPWR VPWR hold594/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_77_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_181_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1250 _5503_/X VGND VGND VPWR VPWR _7047_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1261 _6974_/Q VGND VGND VPWR VPWR _5420_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_57_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1272 _4097_/X VGND VGND VPWR VPWR _6518_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1283 _6958_/Q VGND VGND VPWR VPWR _5402_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1294 _5276_/X VGND VGND VPWR VPWR _6846_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_118 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_185_134 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_540 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_154_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_302 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput170 wb_we_i VGND VGND VPWR VPWR _6320_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_36_402 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4981_ _5087_/C _4959_/X _4980_/Y _4222_/X VGND VGND VPWR VPWR _4981_/X sky130_fd_sc_hd__a211o_1
XFILLER_91_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3932_ _6515_/Q input93/X _6767_/Q VGND VGND VPWR VPWR _3932_/X sky130_fd_sc_hd__mux2_2
X_6720_ _7150_/CLK _6720_/D _6308_/B VGND VGND VPWR VPWR _6720_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_149_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6651_ _6769_/CLK _6651_/D _6399_/A VGND VGND VPWR VPWR _6651_/Q sky130_fd_sc_hd__dfrtp_1
X_3863_ _3905_/B1 _3825_/B _3863_/B1 VGND VGND VPWR VPWR _6403_/D sky130_fd_sc_hd__a21o_1
XFILLER_32_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5602_ _7102_/Q _5571_/Y _5598_/A _5601_/Y _6508_/Q VGND VGND VPWR VPWR _7102_/D
+ sky130_fd_sc_hd__a32o_1
X_6582_ _6689_/CLK _6582_/D fanout509/X VGND VGND VPWR VPWR _6582_/Q sky130_fd_sc_hd__dfrtp_2
X_3794_ input4/X _3339_/Y _5415_/A _6970_/Q _3793_/X VGND VGND VPWR VPWR _3802_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_176_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_192_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5533_ hold253/X _5533_/A1 _5537_/S VGND VGND VPWR VPWR _5533_/X sky130_fd_sc_hd__mux2_1
XFILLER_185_690 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_60_csclk clkbuf_3_2_0_csclk/X VGND VGND VPWR VPWR _6789_/CLK sky130_fd_sc_hd__clkbuf_16
X_5464_ hold755/X _5542_/A1 _5468_/S VGND VGND VPWR VPWR _5464_/X sky130_fd_sc_hd__mux2_1
XFILLER_133_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4415_ _4419_/B _4416_/B VGND VGND VPWR VPWR _4561_/A sky130_fd_sc_hd__or2_1
X_5395_ hold612/X _5545_/A1 _5396_/S VGND VGND VPWR VPWR _5395_/X sky130_fd_sc_hd__mux2_1
XFILLER_99_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7134_ _7140_/CLK _7134_/D VGND VGND VPWR VPWR _7134_/Q sky130_fd_sc_hd__dfxtp_1
X_4346_ _4346_/A _4346_/B VGND VGND VPWR VPWR _4450_/A sky130_fd_sc_hd__or2_1
XFILLER_59_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_75_csclk _6661_/CLK VGND VGND VPWR VPWR _6994_/CLK sky130_fd_sc_hd__clkbuf_16
X_7065_ _7067_/CLK _7065_/D fanout513/X VGND VGND VPWR VPWR _7065_/Q sky130_fd_sc_hd__dfrtp_4
Xfanout359 _3878_/Y VGND VGND VPWR VPWR _5612_/A sky130_fd_sc_hd__buf_6
X_4277_ hold596/X _4289_/A1 _4278_/S VGND VGND VPWR VPWR _4277_/X sky130_fd_sc_hd__mux2_1
XFILLER_100_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6016_ _6939_/Q _5942_/X _5972_/B _7056_/Q _6009_/X VGND VGND VPWR VPWR _6026_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_39_240 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3228_ _6485_/Q _3685_/S VGND VGND VPWR VPWR _3229_/S sky130_fd_sc_hd__nand2_1
XFILLER_55_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_276 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6918_ _6988_/CLK _6918_/D _6396_/A VGND VGND VPWR VPWR _6918_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_23_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_13_csclk clkbuf_3_5_0_csclk/X VGND VGND VPWR VPWR _6632_/CLK sky130_fd_sc_hd__clkbuf_16
X_6849_ _6945_/CLK _6849_/D fanout506/X VGND VGND VPWR VPWR _6849_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_50_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_155_318 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_148_381 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_28_csclk clkbuf_3_5_0_csclk/X VGND VGND VPWR VPWR _7041_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_184_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold380 _4117_/X VGND VGND VPWR VPWR _6536_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold391 _6704_/Q VGND VGND VPWR VPWR hold391/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_2_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1080 _4047_/X VGND VGND VPWR VPWR _6490_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1091 _6499_/Q VGND VGND VPWR VPWR _4066_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_18_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_220 hold90/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_268 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_186_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_158_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_174_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_146_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_142_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4200_ hold507/X _5491_/A1 _4201_/S VGND VGND VPWR VPWR _4200_/X sky130_fd_sc_hd__mux2_1
X_5180_ _5180_/A1 hold53/X _5530_/A1 hold663/X _5529_/B VGND VGND VPWR VPWR _5180_/X
+ sky130_fd_sc_hd__o311a_1
XFILLER_96_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4131_ hold529/X _5491_/A1 _4132_/S VGND VGND VPWR VPWR _4131_/X sky130_fd_sc_hd__mux2_1
XFILLER_95_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_655 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4062_ _6396_/B _3560_/B _4077_/S _4044_/X _5511_/B VGND VGND VPWR VPWR _4078_/S
+ sky130_fd_sc_hd__o221a_4
XFILLER_96_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_198 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_498 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4964_ _4615_/X _4962_/X _4963_/X _4961_/X VGND VGND VPWR VPWR _4979_/A sky130_fd_sc_hd__o211a_1
XFILLER_51_246 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6703_ _7034_/CLK _6703_/D fanout488/X VGND VGND VPWR VPWR _6703_/Q sky130_fd_sc_hd__dfrtp_2
X_3915_ _3184_/Y input90/X _3915_/S VGND VGND VPWR VPWR _3915_/X sky130_fd_sc_hd__mux2_2
XFILLER_189_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4895_ _4895_/A _4895_/B VGND VGND VPWR VPWR _4895_/Y sky130_fd_sc_hd__nand2_1
XFILLER_177_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3846_ _3845_/X _3846_/A1 _3857_/S VGND VGND VPWR VPWR _6411_/D sky130_fd_sc_hd__mux2_1
X_6634_ _7067_/CLK _6634_/D _3264_/A VGND VGND VPWR VPWR _6634_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_20_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_192_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_649 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3777_ _3777_/A _3777_/B _3777_/C _3777_/D VGND VGND VPWR VPWR _3777_/Y sky130_fd_sc_hd__nor4_1
X_6565_ _6565_/CLK _6565_/D fanout495/X VGND VGND VPWR VPWR _6565_/Q sky130_fd_sc_hd__dfrtp_2
X_5516_ _5516_/A0 _5543_/A1 _5519_/S VGND VGND VPWR VPWR _5516_/X sky130_fd_sc_hd__mux2_1
XFILLER_133_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6496_ _7041_/CLK _6496_/D fanout519/X VGND VGND VPWR VPWR _7187_/A sky130_fd_sc_hd__dfrtp_1
XFILLER_118_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5447_ _5447_/A0 _5543_/A1 _5450_/S VGND VGND VPWR VPWR _5447_/X sky130_fd_sc_hd__mux2_1
XFILLER_133_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_160_332 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5378_ _5378_/A0 hold27/X hold42/X VGND VGND VPWR VPWR hold43/A sky130_fd_sc_hd__mux2_1
XFILLER_59_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7117_ _7130_/CLK _7117_/D fanout484/X VGND VGND VPWR VPWR _7117_/Q sky130_fd_sc_hd__dfrtp_1
X_4329_ _4679_/A _4575_/A VGND VGND VPWR VPWR _4789_/A sky130_fd_sc_hd__or2_1
XFILLER_101_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_346 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7048_ _7071_/CLK _7048_/D fanout505/X VGND VGND VPWR VPWR _7048_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_101_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_408 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_168_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_144_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_502 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_144_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_202 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_371 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_268 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_159_410 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3700_ _6979_/Q _5424_/A _5343_/A _6907_/Q VGND VGND VPWR VPWR _3700_/X sky130_fd_sc_hd__a22o_1
XFILLER_53_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4680_ _4680_/A _4725_/B VGND VGND VPWR VPWR _4686_/B sky130_fd_sc_hd__or2_1
XFILLER_147_627 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3631_ input5/X _3360_/Y _4303_/A _6702_/Q VGND VGND VPWR VPWR _3631_/X sky130_fd_sc_hd__a22o_1
XFILLER_147_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6350_ _3903_/A _4222_/B _6317_/X _6349_/X _6320_/B VGND VGND VPWR VPWR _6350_/X
+ sky130_fd_sc_hd__a32o_1
X_3562_ _6544_/Q _4121_/A _4261_/A _6669_/Q VGND VGND VPWR VPWR _3562_/X sky130_fd_sc_hd__a22o_1
XFILLER_155_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_161_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5301_ hold329/X _5541_/A1 _5306_/S VGND VGND VPWR VPWR _5301_/X sky130_fd_sc_hd__mux2_1
X_6281_ _6559_/Q _5936_/X _5942_/X _6689_/Q VGND VGND VPWR VPWR _6281_/X sky130_fd_sc_hd__a22o_1
XFILLER_142_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3493_ _5168_/A hold53/A VGND VGND VPWR VPWR _3493_/Y sky130_fd_sc_hd__nor2_1
XFILLER_115_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5232_ hold689/X _5544_/A1 _5234_/S VGND VGND VPWR VPWR _5232_/X sky130_fd_sc_hd__mux2_1
XFILLER_142_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_376 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5163_ _5163_/A _5529_/B VGND VGND VPWR VPWR _5167_/S sky130_fd_sc_hd__and2_1
X_4114_ hold984/X _6354_/A1 _4120_/S VGND VGND VPWR VPWR _4114_/X sky130_fd_sc_hd__mux2_1
XFILLER_96_463 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5094_ _5094_/A _5094_/B VGND VGND VPWR VPWR _5124_/B sky130_fd_sc_hd__nand2_1
XFILLER_84_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4045_ _6396_/B _5183_/B _4103_/B _4044_/X _5511_/B VGND VGND VPWR VPWR _4061_/S
+ sky130_fd_sc_hd__o221a_4
XFILLER_17_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5996_ _5996_/A _5996_/B VGND VGND VPWR VPWR _5996_/X sky130_fd_sc_hd__or2_1
XPHY_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4947_ _4947_/A _4947_/B _4947_/C VGND VGND VPWR VPWR _4947_/X sky130_fd_sc_hd__and3_1
X_4878_ _4878_/A _4878_/B _4878_/C VGND VGND VPWR VPWR _4879_/D sky130_fd_sc_hd__and3_1
XFILLER_165_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6617_ _6698_/CLK _6617_/D _6401_/A VGND VGND VPWR VPWR _6617_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_193_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3829_ _6487_/Q _3858_/B _3867_/B _3856_/S VGND VGND VPWR VPWR _3830_/B sky130_fd_sc_hd__a31o_1
XFILLER_165_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_165_479 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6548_ _7038_/CLK _6548_/D fanout489/X VGND VGND VPWR VPWR _6548_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_192_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_180_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6479_ _6632_/CLK _6479_/D _3264_/A VGND VGND VPWR VPWR _6479_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_121_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput260 _6750_/Q VGND VGND VPWR VPWR pll_bypass sky130_fd_sc_hd__buf_12
Xoutput271 _6434_/Q VGND VGND VPWR VPWR pll_trim[0] sky130_fd_sc_hd__buf_12
Xoutput282 _6435_/Q VGND VGND VPWR VPWR pll_trim[1] sky130_fd_sc_hd__buf_12
Xoutput293 _6440_/Q VGND VGND VPWR VPWR pll_trim[6] sky130_fd_sc_hd__buf_12
XFILLER_59_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_198 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_385 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_156_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_144_619 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_171_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_124_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_179 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_179_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5850_ _5850_/A _5850_/B VGND VGND VPWR VPWR _5850_/X sky130_fd_sc_hd__or2_1
XFILLER_61_352 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4801_ _4640_/B _4515_/B _4725_/B _4973_/A VGND VGND VPWR VPWR _5065_/A sky130_fd_sc_hd__o22a_1
XTAP_2190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5781_ _7008_/Q _5912_/A2 _5618_/X _6880_/Q VGND VGND VPWR VPWR _5781_/X sky130_fd_sc_hd__a22o_1
XFILLER_21_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4732_ _4732_/A _4732_/B VGND VGND VPWR VPWR _4733_/A sky130_fd_sc_hd__or2_1
XFILLER_147_435 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4663_ _4713_/A _4861_/B _4658_/X _4662_/X VGND VGND VPWR VPWR _4664_/D sky130_fd_sc_hd__o211a_1
X_6402_ _3939_/A1 _6402_/D _6358_/X VGND VGND VPWR VPWR _6402_/Q sky130_fd_sc_hd__dfrtp_4
X_3614_ _3614_/A _3614_/B _3614_/C _3614_/D VGND VGND VPWR VPWR _3624_/B sky130_fd_sc_hd__nor4_1
X_4594_ _4678_/A _4748_/B VGND VGND VPWR VPWR _4594_/X sky130_fd_sc_hd__or2_4
XFILLER_190_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold902 _4245_/X VGND VGND VPWR VPWR _6651_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_128_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold913 _6449_/Q VGND VGND VPWR VPWR hold913/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_134_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold924 _5219_/X VGND VGND VPWR VPWR _6795_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3545_ _5183_/A _3761_/B VGND VGND VPWR VPWR _4127_/A sky130_fd_sc_hd__nor2_8
XFILLER_155_490 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6333_ _6642_/Q _6333_/A2 _6333_/B1 _4222_/B _6332_/X VGND VGND VPWR VPWR _6333_/X
+ sky130_fd_sc_hd__a221o_1
Xhold935 _6556_/Q VGND VGND VPWR VPWR hold935/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_143_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold946 _5513_/X VGND VGND VPWR VPWR _7056_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold957 _6811_/Q VGND VGND VPWR VPWR hold957/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold968 _5486_/X VGND VGND VPWR VPWR _7033_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6264_ _7037_/Q _6295_/A2 _5951_/X _6673_/Q _6263_/X VGND VGND VPWR VPWR _6267_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_103_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold979 hold979/A VGND VGND VPWR VPWR hold979/X sky130_fd_sc_hd__dlygate4sd3_1
X_3476_ _6942_/Q _5379_/A _4014_/A _6464_/Q VGND VGND VPWR VPWR _3476_/X sky130_fd_sc_hd__a22o_1
XFILLER_143_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5215_ hold201/X hold114/X _5216_/S VGND VGND VPWR VPWR _5215_/X sky130_fd_sc_hd__mux2_1
XFILLER_142_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6195_ _6470_/Q _5941_/Y _6285_/A2 _6630_/Q _6194_/X VGND VGND VPWR VPWR _6201_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_97_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5146_ _5146_/A0 _6353_/A1 _5150_/S VGND VGND VPWR VPWR _5146_/X sky130_fd_sc_hd__mux2_1
XFILLER_28_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5077_ _4965_/B _4972_/A _4772_/B _5004_/X _4515_/X VGND VGND VPWR VPWR _5077_/X
+ sky130_fd_sc_hd__o2111a_1
XFILLER_151_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4028_ hold577/X _4299_/A1 _4031_/S VGND VGND VPWR VPWR _4028_/X sky130_fd_sc_hd__mux2_1
XFILLER_84_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_371 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_522 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_59 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5979_ _5979_/A _5979_/B _5981_/B VGND VGND VPWR VPWR _5979_/X sky130_fd_sc_hd__and3_4
XFILLER_100_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_166_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_178_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_422 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_179 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_319 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_276 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold209 _6816_/Q VGND VGND VPWR VPWR hold209/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_172_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3330_ hold82/X _3525_/A VGND VGND VPWR VPWR hold83/A sky130_fd_sc_hd__nor2_8
XFILLER_125_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3261_ _6415_/Q _3261_/B VGND VGND VPWR VPWR _3862_/S sky130_fd_sc_hd__nor2_1
XFILLER_124_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5000_ _5000_/A VGND VGND VPWR VPWR _5110_/B sky130_fd_sc_hd__inv_2
XTAP_569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3192_ _7013_/Q VGND VGND VPWR VPWR _3192_/Y sky130_fd_sc_hd__inv_2
XFILLER_66_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_94_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6951_ _7031_/CLK _6951_/D fanout522/X VGND VGND VPWR VPWR _6951_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_53_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5902_ _6558_/Q _5627_/X _5897_/X _5898_/X _5901_/X VGND VGND VPWR VPWR _5902_/X
+ sky130_fd_sc_hd__a2111o_1
XFILLER_34_330 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6882_ _7083_/CLK _6882_/D fanout518/X VGND VGND VPWR VPWR _6882_/Q sky130_fd_sc_hd__dfstp_4
X_5833_ _7151_/Q _5614_/X _5647_/X _6455_/Q VGND VGND VPWR VPWR _5833_/X sky130_fd_sc_hd__a22o_1
XFILLER_34_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5764_ _6951_/Q _5924_/B2 _5912_/B1 _7031_/Q VGND VGND VPWR VPWR _5764_/X sky130_fd_sc_hd__a22o_1
X_4715_ _4717_/A _4715_/B VGND VGND VPWR VPWR _4715_/Y sky130_fd_sc_hd__nor2_1
XFILLER_175_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5695_ _7012_/Q _5921_/A2 _5915_/A2 _6956_/Q _5694_/X VGND VGND VPWR VPWR _5695_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_135_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4646_ _4725_/B _4597_/Y _4745_/B _4595_/Y _4645_/X VGND VGND VPWR VPWR _4646_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_175_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_162_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_163_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold710 _5374_/X VGND VGND VPWR VPWR _6933_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold721 _7007_/Q VGND VGND VPWR VPWR hold721/X sky130_fd_sc_hd__dlygate4sd3_1
X_4577_ _4943_/A _4692_/A _4748_/B _4574_/Y _4692_/C VGND VGND VPWR VPWR _4579_/C
+ sky130_fd_sc_hd__a311o_1
XFILLER_190_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_162_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold732 _5340_/X VGND VGND VPWR VPWR _6903_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold743 _6831_/Q VGND VGND VPWR VPWR hold743/X sky130_fd_sc_hd__dlygate4sd3_1
X_6316_ _3396_/X _6316_/A1 _6316_/S VGND VGND VPWR VPWR _7140_/D sky130_fd_sc_hd__mux2_1
Xhold754 _4041_/X VGND VGND VPWR VPWR _6482_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_131_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3528_ _6990_/Q hold34/A _4032_/A _6479_/Q VGND VGND VPWR VPWR _3528_/X sky130_fd_sc_hd__a22o_1
Xhold765 _7194_/A VGND VGND VPWR VPWR hold765/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_190_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold776 _4240_/X VGND VGND VPWR VPWR _6647_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold787 _6672_/Q VGND VGND VPWR VPWR hold787/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_143_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold798 _4205_/X VGND VGND VPWR VPWR _6611_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6247_ _7036_/Q _6295_/A2 _5973_/C _6621_/Q _6246_/X VGND VGND VPWR VPWR _6250_/A
+ sky130_fd_sc_hd__a221o_1
X_3459_ _6791_/Q _5208_/A _5502_/A _7052_/Q _3458_/X VGND VGND VPWR VPWR _3460_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_162_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1410 _6592_/Q VGND VGND VPWR VPWR _4183_/A1 sky130_fd_sc_hd__dlygate4sd3_1
X_6178_ _6793_/Q _6004_/B _6168_/X _6177_/X _5610_/A VGND VGND VPWR VPWR _6178_/X
+ sky130_fd_sc_hd__o221a_2
XFILLER_29_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1421 _6725_/Q VGND VGND VPWR VPWR _3270_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_111_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1432 _5399_/X VGND VGND VPWR VPWR _6955_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_84_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1443 _6730_/Q VGND VGND VPWR VPWR _3627_/A1 sky130_fd_sc_hd__dlygate4sd3_1
X_5129_ _4988_/A _4586_/B _4725_/B _4597_/Y _5132_/B VGND VGND VPWR VPWR _5129_/X
+ sky130_fd_sc_hd__o221a_1
Xhold1454 _6723_/Q VGND VGND VPWR VPWR _3286_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_29_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1465 _7146_/Q VGND VGND VPWR VPWR _6340_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_45_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1476 _5735_/X VGND VGND VPWR VPWR _7109_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_57_488 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1487 hold1/A VGND VGND VPWR VPWR _3255_/A1 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1498 _7168_/Q VGND VGND VPWR VPWR _3245_/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_344 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_187_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_187_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_187_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_181_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_746 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_611 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold70 hold70/A VGND VGND VPWR VPWR hold70/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_48_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold81 hold81/A VGND VGND VPWR VPWR hold81/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold92 hold92/A VGND VGND VPWR VPWR hold92/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_29_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_480 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_189_699 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4500_ _4692_/C _4691_/C VGND VGND VPWR VPWR _4501_/B sky130_fd_sc_hd__or2_2
X_5480_ _5480_/A0 _5495_/A1 _5486_/S VGND VGND VPWR VPWR _5480_/X sky130_fd_sc_hd__mux2_1
XFILLER_172_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_144_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_172_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_1 _5406_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4431_ _4557_/B VGND VGND VPWR VPWR _4470_/A sky130_fd_sc_hd__inv_2
XFILLER_172_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_144_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4362_ _5043_/A _4622_/A _6644_/Q VGND VGND VPWR VPWR _4883_/A sky130_fd_sc_hd__o21a_1
X_7150_ _7150_/CLK _7150_/D _4181_/B VGND VGND VPWR VPWR _7150_/Q sky130_fd_sc_hd__dfrtp_1
X_3313_ _3328_/A _3313_/B VGND VGND VPWR VPWR hold61/A sky130_fd_sc_hd__nand2_8
XFILLER_112_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6101_ _7075_/Q _6289_/A2 _6098_/X _6100_/X VGND VGND VPWR VPWR _6102_/C sky130_fd_sc_hd__a211o_1
Xfanout508 fanout510/X VGND VGND VPWR VPWR _6370_/A sky130_fd_sc_hd__buf_6
X_7081_ _7082_/CLK _7081_/D fanout519/X VGND VGND VPWR VPWR _7081_/Q sky130_fd_sc_hd__dfrtp_2
X_4293_ hold165/X hold90/X _4296_/S VGND VGND VPWR VPWR _4293_/X sky130_fd_sc_hd__mux2_1
Xfanout519 fanout520/X VGND VGND VPWR VPWR fanout519/X sky130_fd_sc_hd__buf_8
X_3244_ _7169_/Q _3245_/B _3243_/Y _3245_/A VGND VGND VPWR VPWR _3244_/X sky130_fd_sc_hd__o22a_1
X_6032_ _7028_/Q _5947_/Y _5973_/B _6804_/Q _6031_/X VGND VGND VPWR VPWR _6032_/X
+ sky130_fd_sc_hd__a221o_1
XTAP_388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3175_ _6508_/Q VGND VGND VPWR VPWR _5609_/B sky130_fd_sc_hd__clkinv_2
XFILLER_94_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6934_ _6998_/CLK _6934_/D fanout513/X VGND VGND VPWR VPWR _6934_/Q sky130_fd_sc_hd__dfrtp_1
XPHY_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6865_ _7078_/CLK _6865_/D fanout507/X VGND VGND VPWR VPWR _6865_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_22_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5816_ _7009_/Q _5912_/A2 _5816_/B1 _6945_/Q _5815_/X VGND VGND VPWR VPWR _5817_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_22_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6796_ _6988_/CLK _6796_/D _6396_/A VGND VGND VPWR VPWR _6796_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_22_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_179_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5747_ _6918_/Q _5923_/B VGND VGND VPWR VPWR _5747_/X sky130_fd_sc_hd__and2b_1
XFILLER_157_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_182_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5678_ _6931_/Q _5807_/B1 _5674_/X _5675_/X _5677_/X VGND VGND VPWR VPWR _5678_/X
+ sky130_fd_sc_hd__a2111o_1
XFILLER_175_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4629_ _4691_/A _4629_/B _4793_/B VGND VGND VPWR VPWR _4666_/A sky130_fd_sc_hd__or3b_1
XFILLER_135_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold540 _4219_/X VGND VGND VPWR VPWR _6623_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold551 _6674_/Q VGND VGND VPWR VPWR hold551/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold562 _4313_/X VGND VGND VPWR VPWR _6708_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_173_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold573 _6474_/Q VGND VGND VPWR VPWR hold573/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold584 _4301_/X VGND VGND VPWR VPWR _6698_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold595 _5458_/X VGND VGND VPWR VPWR _7008_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_77_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1240 _5254_/X VGND VGND VPWR VPWR _6826_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_18_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1251 _6794_/Q VGND VGND VPWR VPWR _5218_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_85_572 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1262 _5420_/X VGND VGND VPWR VPWR _6974_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1273 _6918_/Q VGND VGND VPWR VPWR _5357_/A0 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1284 _5402_/X VGND VGND VPWR VPWR _6958_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1295 _7014_/Q VGND VGND VPWR VPWR _5465_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_146 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_139_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_99_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput160 wb_dat_i[6] VGND VGND VPWR VPWR _6342_/B1 sky130_fd_sc_hd__clkbuf_1
XFILLER_36_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4980_ _5087_/B _4979_/X _4960_/Y VGND VGND VPWR VPWR _4980_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_17_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3931_ _6516_/Q _3931_/A1 _6765_/Q VGND VGND VPWR VPWR _3931_/X sky130_fd_sc_hd__mux2_1
XFILLER_32_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_177_603 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6650_ _6711_/CLK _6650_/D fanout486/X VGND VGND VPWR VPWR _6650_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_149_316 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3862_ _6404_/Q _7159_/Q _3862_/S VGND VGND VPWR VPWR _6404_/D sky130_fd_sc_hd__mux2_1
X_5601_ _5964_/A _5980_/B VGND VGND VPWR VPWR _5601_/Y sky130_fd_sc_hd__nor2_8
XFILLER_149_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6581_ _6718_/CLK _6581_/D _6401_/A VGND VGND VPWR VPWR _6581_/Q sky130_fd_sc_hd__dfrtp_2
X_3793_ input71/X hold76/A _4038_/A _6480_/Q VGND VGND VPWR VPWR _3793_/X sky130_fd_sc_hd__a22o_1
X_5532_ hold367/X _5532_/A1 _5537_/S VGND VGND VPWR VPWR _5532_/X sky130_fd_sc_hd__mux2_1
XFILLER_157_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_9_csclk _6684_/CLK VGND VGND VPWR VPWR _6699_/CLK sky130_fd_sc_hd__clkbuf_16
X_5463_ hold905/X _5505_/A1 _5468_/S VGND VGND VPWR VPWR _5463_/X sky130_fd_sc_hd__mux2_1
XFILLER_117_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4414_ _4542_/A _5022_/A VGND VGND VPWR VPWR _4692_/A sky130_fd_sc_hd__or2_4
X_5394_ hold725/X _5544_/A1 _5396_/S VGND VGND VPWR VPWR _5394_/X sky130_fd_sc_hd__mux2_1
XFILLER_99_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7133_ _7137_/CLK _7133_/D VGND VGND VPWR VPWR _7133_/Q sky130_fd_sc_hd__dfxtp_1
X_4345_ _4544_/A _4541_/B _4345_/C VGND VGND VPWR VPWR _4346_/B sky130_fd_sc_hd__and3_1
XFILLER_98_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4276_ hold799/X _6355_/A1 _4278_/S VGND VGND VPWR VPWR _4276_/X sky130_fd_sc_hd__mux2_1
Xfanout349 _5975_/X VGND VGND VPWR VPWR _6004_/B sky130_fd_sc_hd__buf_12
X_7064_ _7071_/CLK _7064_/D fanout504/X VGND VGND VPWR VPWR _7064_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_100_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6015_ _7027_/Q _6291_/A2 _6007_/X _6012_/X _6014_/X VGND VGND VPWR VPWR _6027_/B
+ sky130_fd_sc_hd__a2111o_1
X_3227_ _6417_/Q _6416_/Q _6415_/Q VGND VGND VPWR VPWR _3817_/C sky130_fd_sc_hd__nor3_2
XFILLER_86_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_252 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_288 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6917_ _7029_/CLK _6917_/D fanout519/X VGND VGND VPWR VPWR _6917_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_52_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6848_ _6961_/CLK _6848_/D fanout521/X VGND VGND VPWR VPWR _6848_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_167_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6779_ _7017_/CLK _6779_/D fanout515/X VGND VGND VPWR VPWR _6779_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_183_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_108_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_151_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_190_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold370 _5202_/X VGND VGND VPWR VPWR _6780_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_2_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold381 _6812_/Q VGND VGND VPWR VPWR hold381/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold392 _4308_/X VGND VGND VPWR VPWR _6704_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_77_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1070 _7173_/A VGND VGND VPWR VPWR _5170_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1081 _7178_/A VGND VGND VPWR VPWR _4078_/A0 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1092 _4066_/X VGND VGND VPWR VPWR _6499_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_210 hold114/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_221 hold142/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_631 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_102 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_686 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_139_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_130_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4130_ hold823/X _6355_/A1 _4132_/S VGND VGND VPWR VPWR _4130_/X sky130_fd_sc_hd__mux2_1
XFILLER_96_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_667 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4061_ hold215/X _4060_/X _4061_/S VGND VGND VPWR VPWR _4061_/X sky130_fd_sc_hd__mux2_1
XFILLER_49_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_572 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4963_ _4687_/B _4615_/B _4683_/B _4703_/B VGND VGND VPWR VPWR _4963_/X sky130_fd_sc_hd__o22a_1
X_6702_ _7034_/CLK _6702_/D fanout490/X VGND VGND VPWR VPWR _6702_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_51_258 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3914_ _3183_/Y input92/X _3915_/S VGND VGND VPWR VPWR _3914_/X sky130_fd_sc_hd__mux2_2
XFILLER_32_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4894_ _4894_/A _4894_/B VGND VGND VPWR VPWR _4895_/B sky130_fd_sc_hd__nor2_1
XFILLER_149_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6633_ _6633_/CLK _6633_/D fanout509/X VGND VGND VPWR VPWR _6633_/Q sky130_fd_sc_hd__dfrtp_1
X_3845_ _3267_/X _3266_/Y _3845_/S VGND VGND VPWR VPWR _3845_/X sky130_fd_sc_hd__mux2_1
XFILLER_20_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6564_ _6689_/CLK _6564_/D fanout510/X VGND VGND VPWR VPWR _6564_/Q sky130_fd_sc_hd__dfrtp_2
X_3776_ _6810_/Q _5235_/A _5379_/A _6938_/Q _3775_/X VGND VGND VPWR VPWR _3777_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_138_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5515_ hold359/X _5515_/A1 _5519_/S VGND VGND VPWR VPWR _5515_/X sky130_fd_sc_hd__mux2_1
X_6495_ _7041_/CLK _6495_/D fanout518/X VGND VGND VPWR VPWR _7186_/A sky130_fd_sc_hd__dfrtp_1
XFILLER_145_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5446_ hold857/X _5542_/A1 _5450_/S VGND VGND VPWR VPWR _5446_/X sky130_fd_sc_hd__mux2_1
XFILLER_160_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5377_ hold419/X _5545_/A1 hold42/X VGND VGND VPWR VPWR _5377_/X sky130_fd_sc_hd__mux2_1
XFILLER_160_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7116_ _7130_/CLK _7116_/D fanout484/X VGND VGND VPWR VPWR _7116_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_59_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4328_ _4575_/A VGND VGND VPWR VPWR _4328_/Y sky130_fd_sc_hd__inv_2
XFILLER_101_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_358 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7047_ _7055_/CLK _7047_/D fanout500/X VGND VGND VPWR VPWR _7047_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_74_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4259_ hold654/X _4289_/A1 _4260_/S VGND VGND VPWR VPWR _4259_/X sky130_fd_sc_hd__mux2_1
XFILLER_28_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_380 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_514 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_147_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_187_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_74_csclk clkbuf_3_2_0_csclk/X VGND VGND VPWR VPWR _7010_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_147_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3630_ _6428_/Q _3975_/A _3572_/Y input97/X VGND VGND VPWR VPWR _3630_/X sky130_fd_sc_hd__a22o_1
XFILLER_147_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_146_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3561_ hold61/X _3761_/B VGND VGND VPWR VPWR _4261_/A sky130_fd_sc_hd__nor2_4
X_5300_ _5300_/A0 _5531_/A1 _5306_/S VGND VGND VPWR VPWR _5300_/X sky130_fd_sc_hd__mux2_1
XFILLER_142_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6280_ _7130_/Q _6305_/A2 _6278_/X _6279_/X VGND VGND VPWR VPWR _7130_/D sky130_fd_sc_hd__o22a_1
X_3492_ _6870_/Q _5298_/A _5151_/A _6746_/Q _3491_/X VGND VGND VPWR VPWR _3502_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_142_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5231_ _5231_/A0 _5465_/A1 _5234_/S VGND VGND VPWR VPWR _5231_/X sky130_fd_sc_hd__mux2_1
XFILLER_102_219 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_388 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5162_ _5488_/A1 _5162_/A1 _5162_/S VGND VGND VPWR VPWR _5162_/X sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_12_csclk clkbuf_opt_2_0_csclk/X VGND VGND VPWR VPWR _7155_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_111_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4113_ _4113_/A0 _6353_/A1 _4120_/S VGND VGND VPWR VPWR _4113_/X sky130_fd_sc_hd__mux2_1
X_5093_ _4549_/B _4515_/B _4834_/X _5037_/D VGND VGND VPWR VPWR _5094_/B sky130_fd_sc_hd__o211a_1
XFILLER_96_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4044_ _6396_/B _5190_/A VGND VGND VPWR VPWR _4044_/X sky130_fd_sc_hd__and2b_1
XFILLER_37_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_27_csclk clkbuf_3_5_0_csclk/X VGND VGND VPWR VPWR _7083_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_64_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_92_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5995_ _6986_/Q _5941_/Y wire390/X _6850_/Q _5994_/X VGND VGND VPWR VPWR _5996_/B
+ sky130_fd_sc_hd__a221o_1
XPHY_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4946_ _4946_/A _5025_/B _4946_/C VGND VGND VPWR VPWR _4958_/C sky130_fd_sc_hd__and3_1
XFILLER_178_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_193_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4877_ _4877_/A _4877_/B _4877_/C _4877_/D VGND VGND VPWR VPWR _4878_/C sky130_fd_sc_hd__and4_1
XFILLER_193_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6616_ _6633_/CLK _6616_/D _6370_/A VGND VGND VPWR VPWR _6616_/Q sky130_fd_sc_hd__dfstp_1
X_3828_ _7167_/Q _3828_/B VGND VGND VPWR VPWR _3867_/B sky130_fd_sc_hd__nand2_1
XFILLER_165_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6547_ _6697_/CLK _6547_/D fanout489/X VGND VGND VPWR VPWR _6547_/Q sky130_fd_sc_hd__dfrtp_4
X_3759_ _6645_/Q _4237_/A _4008_/A _6455_/Q VGND VGND VPWR VPWR _3759_/X sky130_fd_sc_hd__a22o_1
XFILLER_152_119 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6478_ _6718_/CLK _6478_/D _6401_/A VGND VGND VPWR VPWR _6478_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_106_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5429_ _5429_/A0 _5543_/A1 _5432_/S VGND VGND VPWR VPWR _5429_/X sky130_fd_sc_hd__mux2_1
Xoutput250 _3938_/Y VGND VGND VPWR VPWR pad_flash_csb_oeb sky130_fd_sc_hd__buf_12
Xoutput261 _6736_/Q VGND VGND VPWR VPWR pll_dco_ena sky130_fd_sc_hd__buf_12
XFILLER_121_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput272 _6428_/Q VGND VGND VPWR VPWR pll_trim[10] sky130_fd_sc_hd__buf_12
Xoutput283 _6422_/Q VGND VGND VPWR VPWR pll_trim[20] sky130_fd_sc_hd__buf_12
Xoutput294 _6441_/Q VGND VGND VPWR VPWR pll_trim[7] sky130_fd_sc_hd__buf_12
XFILLER_181_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_188_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_397 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_424 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_99_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_164_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_1_1_1_wb_clk_i clkbuf_1_1_1_wb_clk_i/A VGND VGND VPWR VPWR clkbuf_2_3_0_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_8
XTAP_707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_180 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4800_ _4921_/A _4586_/B _5043_/B _4745_/B VGND VGND VPWR VPWR _4816_/A sky130_fd_sc_hd__o22a_1
XTAP_2180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5780_ _6992_/Q _5622_/X _5624_/X _6832_/Q VGND VGND VPWR VPWR _5780_/X sky130_fd_sc_hd__a22o_1
XFILLER_14_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4731_ _4535_/A _4435_/Y _4715_/B _4394_/Y VGND VGND VPWR VPWR _5016_/A sky130_fd_sc_hd__o2bb2a_1
XFILLER_187_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_159_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4662_ _4662_/A _4662_/B _4662_/C VGND VGND VPWR VPWR _4662_/X sky130_fd_sc_hd__and3_1
XFILLER_147_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6401_ _6401_/A _6401_/B VGND VGND VPWR VPWR _6401_/X sky130_fd_sc_hd__and2_1
X_3613_ input29/X _3339_/Y _3360_/Y input6/X _3612_/X VGND VGND VPWR VPWR _3614_/D
+ sky130_fd_sc_hd__a221o_2
X_4593_ _4678_/A _4671_/B VGND VGND VPWR VPWR _4719_/B sky130_fd_sc_hd__or2_4
Xhold903 _6610_/Q VGND VGND VPWR VPWR hold903/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold914 _4001_/X VGND VGND VPWR VPWR _6449_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6332_ _6644_/Q _6332_/A2 _6332_/B1 _6643_/Q VGND VGND VPWR VPWR _6332_/X sky130_fd_sc_hd__a22o_1
X_3544_ hold61/X _5161_/B VGND VGND VPWR VPWR _4237_/A sky130_fd_sc_hd__nor2_4
Xhold925 _6561_/Q VGND VGND VPWR VPWR hold925/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold936 _4141_/X VGND VGND VPWR VPWR _6556_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold947 _6899_/Q VGND VGND VPWR VPWR hold947/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_142_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold958 _5237_/X VGND VGND VPWR VPWR _6811_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold969 _7064_/Q VGND VGND VPWR VPWR hold969/X sky130_fd_sc_hd__dlygate4sd3_1
X_6263_ _6473_/Q _5941_/Y _5978_/X _6698_/Q VGND VGND VPWR VPWR _6263_/X sky130_fd_sc_hd__a22o_1
XFILLER_89_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3475_ _3552_/A _3560_/B VGND VGND VPWR VPWR _4014_/A sky130_fd_sc_hd__nor2_4
XFILLER_103_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_143_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5214_ hold487/X _5526_/A1 _5216_/S VGND VGND VPWR VPWR _5214_/X sky130_fd_sc_hd__mux2_1
X_6194_ _6550_/Q _5973_/B _5963_/X _6565_/Q VGND VGND VPWR VPWR _6194_/X sky130_fd_sc_hd__a22o_1
X_5145_ _5145_/A _6352_/B VGND VGND VPWR VPWR _5150_/S sky130_fd_sc_hd__and2_2
XFILLER_29_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5076_ _5100_/A _5136_/C _5102_/B _5101_/B VGND VGND VPWR VPWR _5079_/A sky130_fd_sc_hd__and4_1
XFILLER_44_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4027_ _4027_/A0 _5308_/A1 _4031_/S VGND VGND VPWR VPWR _4027_/X sky130_fd_sc_hd__mux2_1
XFILLER_37_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5978_ _5979_/A _5978_/B _5981_/B VGND VGND VPWR VPWR _5978_/X sky130_fd_sc_hd__and3_4
XFILLER_12_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4929_ _4929_/A _4929_/B VGND VGND VPWR VPWR _4999_/B sky130_fd_sc_hd__or2_1
XFILLER_166_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_176_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmgmt_gpio_9_buff_inst _3921_/X VGND VGND VPWR VPWR mgmt_gpio_out[9] sky130_fd_sc_hd__clkbuf_8
XFILLER_118_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_134_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_161_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_180 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_711 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_184_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_171_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_166_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_124_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3260_ _7159_/Q _6415_/Q _3261_/B VGND VGND VPWR VPWR _3260_/X sky130_fd_sc_hd__a21o_1
XFILLER_140_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_667 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3191_ _7021_/Q VGND VGND VPWR VPWR _3191_/Y sky130_fd_sc_hd__inv_2
XFILLER_182_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6950_ _6988_/CLK _6950_/D fanout517/X VGND VGND VPWR VPWR _6950_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_66_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5901_ _7037_/Q _5645_/X _5899_/X _5900_/X VGND VGND VPWR VPWR _5901_/X sky130_fd_sc_hd__a211o_1
X_6881_ _6881_/CLK hold99/X fanout523/X VGND VGND VPWR VPWR _6881_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_34_342 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_662 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5832_ _6645_/Q _5918_/A2 _5828_/X _5829_/X _5831_/X VGND VGND VPWR VPWR _5832_/X
+ sky130_fd_sc_hd__a2111o_1
XFILLER_22_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_148_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5763_ _5763_/A _5763_/B VGND VGND VPWR VPWR _5763_/X sky130_fd_sc_hd__or2_1
X_4714_ _4714_/A _4714_/B _4714_/C _5017_/B VGND VGND VPWR VPWR _4714_/X sky130_fd_sc_hd__or4b_1
XFILLER_147_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5694_ _7004_/Q _5912_/A2 _5618_/X _6876_/Q VGND VGND VPWR VPWR _5694_/X sky130_fd_sc_hd__a22o_1
XFILLER_187_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4645_ _5043_/B _4962_/C _4575_/X _4597_/Y VGND VGND VPWR VPWR _4645_/X sky130_fd_sc_hd__a31o_1
XFILLER_135_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_163_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold700 _5331_/X VGND VGND VPWR VPWR _6895_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_146_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4576_ _4692_/C _4748_/B VGND VGND VPWR VPWR _4576_/X sky130_fd_sc_hd__or2_1
Xhold711 _6957_/Q VGND VGND VPWR VPWR hold711/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold722 _5457_/X VGND VGND VPWR VPWR _7007_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_115_130 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold733 _7021_/Q VGND VGND VPWR VPWR hold733/X sky130_fd_sc_hd__dlygate4sd3_1
X_6315_ _3433_/X _6315_/A1 _6316_/S VGND VGND VPWR VPWR _7139_/D sky130_fd_sc_hd__mux2_1
Xhold744 _5259_/X VGND VGND VPWR VPWR _6831_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3527_ _3563_/A _3538_/B VGND VGND VPWR VPWR _4032_/A sky130_fd_sc_hd__nor2_8
Xhold755 _7013_/Q VGND VGND VPWR VPWR hold755/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_190_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmax_cap474 _3817_/C VGND VGND VPWR VPWR _3685_/S sky130_fd_sc_hd__buf_2
Xhold766 _5196_/X VGND VGND VPWR VPWR _6775_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold777 _6467_/Q VGND VGND VPWR VPWR hold777/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_103_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold788 _4270_/X VGND VGND VPWR VPWR _6672_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold799 _6677_/Q VGND VGND VPWR VPWR hold799/X sky130_fd_sc_hd__dlygate4sd3_1
X_6246_ _6462_/Q _5943_/Y _5948_/X _6547_/Q VGND VGND VPWR VPWR _6246_/X sky130_fd_sc_hd__a22o_1
XFILLER_89_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_196 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3458_ input40/X _4092_/S _5388_/A _6951_/Q VGND VGND VPWR VPWR _3458_/X sky130_fd_sc_hd__a22o_1
XFILLER_69_250 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6177_ _6177_/A _6177_/B _6177_/C _5975_/X VGND VGND VPWR VPWR _6177_/X sky130_fd_sc_hd__or4b_1
Xhold1400 _6598_/Q VGND VGND VPWR VPWR _4189_/A1 sky130_fd_sc_hd__dlygate4sd3_1
X_3389_ _3503_/A _3706_/A VGND VGND VPWR VPWR _5397_/A sky130_fd_sc_hd__nor2_8
Xhold1411 _6594_/Q VGND VGND VPWR VPWR _4185_/A1 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1422 _5183_/A VGND VGND VPWR VPWR _5180_/A1 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1433 _7137_/Q VGND VGND VPWR VPWR _6313_/A1 sky130_fd_sc_hd__dlygate4sd3_1
X_5128_ _5102_/X _5106_/Y _5113_/X _5127_/X VGND VGND VPWR VPWR _6725_/D sky130_fd_sc_hd__a211o_1
Xhold1444 _7150_/Q VGND VGND VPWR VPWR _6351_/A2 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_45_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1455 _6576_/Q VGND VGND VPWR VPWR _4164_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_55_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1466 hold25/A VGND VGND VPWR VPWR _3250_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_29_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1477 _7123_/Q VGND VGND VPWR VPWR _6129_/A1 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1488 _7113_/Q VGND VGND VPWR VPWR _5823_/A1 sky130_fd_sc_hd__dlygate4sd3_1
X_5059_ _6723_/Q _4222_/X _5119_/A _5058_/X _5039_/X VGND VGND VPWR VPWR _5059_/X
+ sky130_fd_sc_hd__a221o_1
XTAP_2905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1499 _3244_/X VGND VGND VPWR VPWR _7169_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_84_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_187_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_178_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_126_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_154_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_181_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_758 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_623 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold60 hold60/A VGND VGND VPWR VPWR hold60/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold71 hold71/A VGND VGND VPWR VPWR hold71/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold82 hold82/A VGND VGND VPWR VPWR hold82/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_48_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold93 hold93/A VGND VGND VPWR VPWR hold93/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_29_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_492 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_542 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_117_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4430_ _4901_/A _4894_/A _4430_/C VGND VGND VPWR VPWR _4557_/B sky130_fd_sc_hd__nor3_4
XANTENNA_2 _3975_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_144_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4361_ _4901_/A _4471_/A VGND VGND VPWR VPWR _4622_/A sky130_fd_sc_hd__or2_4
XFILLER_98_323 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6100_ _6838_/Q _5946_/X _6296_/B1 _6902_/Q _6099_/X VGND VGND VPWR VPWR _6100_/X
+ sky130_fd_sc_hd__a221o_1
X_3312_ hold60/X VGND VGND VPWR VPWR _3313_/B sky130_fd_sc_hd__inv_2
Xfanout509 fanout510/X VGND VGND VPWR VPWR fanout509/X sky130_fd_sc_hd__buf_8
X_7080_ _7080_/CLK _7080_/D fanout514/X VGND VGND VPWR VPWR _7080_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_98_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_656 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_291 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4292_ _4292_/A0 _5521_/A1 _4296_/S VGND VGND VPWR VPWR _4292_/X sky130_fd_sc_hd__mux2_1
XFILLER_98_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6031_ _6844_/Q _5939_/X _6284_/B1 _6860_/Q VGND VGND VPWR VPWR _6031_/X sky130_fd_sc_hd__a22o_1
X_3243_ _7169_/Q _3246_/A _3245_/B VGND VGND VPWR VPWR _3243_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_100_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3174_ _6507_/Q VGND VGND VPWR VPWR _3174_/Y sky130_fd_sc_hd__inv_6
XFILLER_27_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6933_ _7082_/CLK _6933_/D fanout519/X VGND VGND VPWR VPWR _6933_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6864_ _7058_/CLK _6864_/D fanout521/X VGND VGND VPWR VPWR _6864_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_50_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5815_ _6881_/Q _5618_/X _5915_/A2 _6961_/Q VGND VGND VPWR VPWR _5815_/X sky130_fd_sc_hd__a22o_1
XFILLER_50_654 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6795_ _7056_/CLK _6795_/D fanout504/X VGND VGND VPWR VPWR _6795_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_179_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_148_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5746_ _6958_/Q _5915_/A2 _5915_/B1 _6862_/Q _5745_/X VGND VGND VPWR VPWR _5754_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_41_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5677_ _6899_/Q _5918_/A2 _5918_/B1 _6851_/Q _5676_/X VGND VGND VPWR VPWR _5677_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_148_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_439 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4628_ _4985_/A _4649_/B VGND VGND VPWR VPWR _4793_/B sky130_fd_sc_hd__nor2_1
Xhold530 _4131_/X VGND VGND VPWR VPWR _6548_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold541 _6421_/Q VGND VGND VPWR VPWR hold541/X sky130_fd_sc_hd__dlygate4sd3_1
X_4559_ _4959_/C _4854_/A _4942_/B _4559_/D VGND VGND VPWR VPWR _4559_/X sky130_fd_sc_hd__and4bb_1
Xhold552 _4272_/X VGND VGND VPWR VPWR _6674_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_9_8 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold563 _6656_/Q VGND VGND VPWR VPWR hold563/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold574 _4031_/X VGND VGND VPWR VPWR _6474_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold585 _7051_/Q VGND VGND VPWR VPWR hold585/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold596 _6678_/Q VGND VGND VPWR VPWR hold596/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_106_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6229_ _7127_/Q _5612_/A _5612_/B VGND VGND VPWR VPWR _6229_/X sky130_fd_sc_hd__o21a_1
XFILLER_77_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1230 _4215_/X VGND VGND VPWR VPWR _6619_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1241 _6978_/Q VGND VGND VPWR VPWR _5425_/A0 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1252 _5218_/X VGND VGND VPWR VPWR _6794_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_66_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_702 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_415 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1263 _6565_/Q VGND VGND VPWR VPWR _4152_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_85_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1274 _5357_/X VGND VGND VPWR VPWR _6918_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1285 _6886_/Q VGND VGND VPWR VPWR _5321_/A0 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1296 _5465_/X VGND VGND VPWR VPWR _7014_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_154_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_139_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput150 wb_dat_i[26] VGND VGND VPWR VPWR _6330_/A2 sky130_fd_sc_hd__clkbuf_1
XFILLER_49_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput161 wb_dat_i[7] VGND VGND VPWR VPWR _6345_/B1 sky130_fd_sc_hd__clkbuf_1
XFILLER_48_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3930_ _6517_/Q user_clock _6766_/Q VGND VGND VPWR VPWR _3930_/X sky130_fd_sc_hd__mux2_1
XFILLER_16_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_177_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3861_ _3904_/B1 _3179_/Y _3825_/B _6405_/Q VGND VGND VPWR VPWR _3861_/X sky130_fd_sc_hd__a31o_1
XFILLER_31_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_189_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5600_ _5962_/B _5981_/B VGND VGND VPWR VPWR _5980_/B sky130_fd_sc_hd__nand2_8
XFILLER_32_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6580_ _6633_/CLK _6580_/D _6370_/A VGND VGND VPWR VPWR _6580_/Q sky130_fd_sc_hd__dfstp_1
X_3792_ _3792_/A _3792_/B _3792_/C _3792_/D VGND VGND VPWR VPWR _3815_/B sky130_fd_sc_hd__nor4_1
XFILLER_176_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5531_ hold891/X _5531_/A1 _5537_/S VGND VGND VPWR VPWR _5531_/X sky130_fd_sc_hd__mux2_1
XFILLER_117_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5462_ _5462_/A0 _5495_/A1 _5468_/S VGND VGND VPWR VPWR _5462_/X sky130_fd_sc_hd__mux2_1
XFILLER_172_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4413_ _4542_/A _5022_/A VGND VGND VPWR VPWR _4947_/A sky130_fd_sc_hd__nor2_1
XFILLER_145_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_160_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5393_ _5393_/A0 _5543_/A1 _5396_/S VGND VGND VPWR VPWR _5393_/X sky130_fd_sc_hd__mux2_1
X_7132_ _7150_/CLK _7132_/D _6308_/B VGND VGND VPWR VPWR _7132_/Q sky130_fd_sc_hd__dfrtp_4
X_4344_ _4541_/B _4345_/C _4544_/A VGND VGND VPWR VPWR _4346_/A sky130_fd_sc_hd__a21oi_1
XFILLER_99_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7063_ _7063_/CLK _7063_/D fanout495/X VGND VGND VPWR VPWR _7063_/Q sky130_fd_sc_hd__dfstp_1
X_4275_ hold877/X _5189_/A1 _4278_/S VGND VGND VPWR VPWR _4275_/X sky130_fd_sc_hd__mux2_1
XFILLER_98_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6014_ _7064_/Q _6283_/A2 _5980_/Y _7019_/Q VGND VGND VPWR VPWR _6014_/X sky130_fd_sc_hd__a22o_1
X_3226_ _4614_/A VGND VGND VPWR VPWR _4630_/A sky130_fd_sc_hd__clkinv_2
XFILLER_39_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_264 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6916_ _7073_/CLK _6916_/D fanout498/X VGND VGND VPWR VPWR _6916_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_52_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6847_ _7042_/CLK _6847_/D fanout524/X VGND VGND VPWR VPWR _6847_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_23_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6778_ _7069_/CLK _6778_/D fanout516/X VGND VGND VPWR VPWR _6778_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_139_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5729_ _6949_/Q _5924_/B2 _5912_/B1 _7029_/Q VGND VGND VPWR VPWR _5729_/X sky130_fd_sc_hd__a22o_1
XFILLER_109_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_136_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_190_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold360 _5515_/X VGND VGND VPWR VPWR _7058_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold371 _6916_/Q VGND VGND VPWR VPWR hold371/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold382 _5238_/X VGND VGND VPWR VPWR _6812_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold393 _6430_/Q VGND VGND VPWR VPWR hold393/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_117_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1060 _6435_/Q VGND VGND VPWR VPWR _3986_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_100_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1071 _5170_/X VGND VGND VPWR VPWR _5171_/B1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_85_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1082 _4078_/X VGND VGND VPWR VPWR _6505_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_200 _5974_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1093 _6768_/Q VGND VGND VPWR VPWR _5188_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_211 hold114/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_222 _5533_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_146_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_115_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_515 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4060_ _4111_/A0 hold27/X _4103_/B VGND VGND VPWR VPWR _4060_/X sky130_fd_sc_hd__mux2_1
XFILLER_96_679 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_584 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_278 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4962_ _4965_/A _4965_/B _4962_/C VGND VGND VPWR VPWR _4962_/X sky130_fd_sc_hd__and3_1
XFILLER_51_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6701_ _7034_/CLK _6701_/D fanout490/X VGND VGND VPWR VPWR _6701_/Q sky130_fd_sc_hd__dfrtp_1
X_3913_ _6522_/Q input89/X _3915_/S VGND VGND VPWR VPWR _3913_/X sky130_fd_sc_hd__mux2_2
XFILLER_32_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4893_ _4407_/X _5025_/B _4911_/B _4911_/C VGND VGND VPWR VPWR _4893_/Y sky130_fd_sc_hd__a211oi_1
XFILLER_149_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6632_ _6632_/CLK _6632_/D _3264_/A VGND VGND VPWR VPWR _6632_/Q sky130_fd_sc_hd__dfstp_2
X_3844_ _3856_/S _3847_/B VGND VGND VPWR VPWR _3844_/Y sky130_fd_sc_hd__nor2_1
XFILLER_149_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6563_ _6633_/CLK _6563_/D _6370_/A VGND VGND VPWR VPWR _6563_/Q sky130_fd_sc_hd__dfrtp_1
X_3775_ _6802_/Q _5226_/A _4297_/A _6695_/Q VGND VGND VPWR VPWR _3775_/X sky130_fd_sc_hd__a22o_1
XFILLER_164_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5514_ hold455/X _5541_/A1 _5519_/S VGND VGND VPWR VPWR _5514_/X sky130_fd_sc_hd__mux2_1
XFILLER_118_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6494_ _7041_/CLK _6494_/D fanout518/X VGND VGND VPWR VPWR _7185_/A sky130_fd_sc_hd__dfrtp_1
XFILLER_106_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5445_ hold377/X _5532_/A1 _5450_/S VGND VGND VPWR VPWR _5445_/X sky130_fd_sc_hd__mux2_1
XFILLER_105_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5376_ hold489/X _5526_/A1 hold42/X VGND VGND VPWR VPWR _5376_/X sky130_fd_sc_hd__mux2_1
XFILLER_154_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7115_ _7130_/CLK _7115_/D fanout485/X VGND VGND VPWR VPWR _7115_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_160_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4327_ _4554_/A _4596_/B VGND VGND VPWR VPWR _4575_/A sky130_fd_sc_hd__nand2_4
XFILLER_99_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7046_ _7046_/CLK _7046_/D fanout501/X VGND VGND VPWR VPWR _7046_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_47_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4258_ hold789/X _5505_/A1 _4260_/S VGND VGND VPWR VPWR _4258_/X sky130_fd_sc_hd__mux2_1
XFILLER_101_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3209_ _6885_/Q VGND VGND VPWR VPWR _3209_/Y sky130_fd_sc_hd__inv_2
X_4189_ _3396_/X _4189_/A1 _4189_/S VGND VGND VPWR VPWR _6598_/D sky130_fd_sc_hd__mux2_1
XFILLER_28_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_635 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_534 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_331 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_124_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold190 _5535_/X VGND VGND VPWR VPWR _7076_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_78_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_554 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_8_csclk _6684_/CLK VGND VGND VPWR VPWR _6683_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_46_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_186_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3560_ _5183_/A _3560_/B VGND VGND VPWR VPWR _4121_/A sky130_fd_sc_hd__nor2_8
XFILLER_127_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_161_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3491_ _6982_/Q _5424_/A _4225_/A _6629_/Q VGND VGND VPWR VPWR _3491_/X sky130_fd_sc_hd__a22o_1
XFILLER_115_537 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5230_ _5230_/A0 _5533_/A1 _5234_/S VGND VGND VPWR VPWR _5230_/X sky130_fd_sc_hd__mux2_1
XFILLER_154_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5161_ _5168_/A _5161_/B _5187_/B VGND VGND VPWR VPWR _5162_/S sky130_fd_sc_hd__or3b_1
XFILLER_170_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4112_ _6399_/B _4112_/B _5187_/B VGND VGND VPWR VPWR _4120_/S sky130_fd_sc_hd__and3b_4
XFILLER_111_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5092_ _4640_/B _4515_/B _5026_/B _4513_/A VGND VGND VPWR VPWR _5094_/A sky130_fd_sc_hd__o22a_1
XFILLER_68_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4043_ hold463/X _6357_/A1 _4043_/S VGND VGND VPWR VPWR _4043_/X sky130_fd_sc_hd__mux2_1
XFILLER_25_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5994_ _7047_/Q _5975_/C _5977_/X _6922_/Q VGND VGND VPWR VPWR _5994_/X sky130_fd_sc_hd__a22o_1
XFILLER_24_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4945_ _4679_/B _4629_/B _4944_/X VGND VGND VPWR VPWR _4958_/A sky130_fd_sc_hd__a21o_1
XFILLER_20_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4876_ _4748_/B _4597_/Y _4620_/B _4717_/B VGND VGND VPWR VPWR _4877_/D sky130_fd_sc_hd__o22a_1
X_6615_ _6686_/CLK _6615_/D fanout492/X VGND VGND VPWR VPWR _6615_/Q sky130_fd_sc_hd__dfrtp_2
X_3827_ _6485_/Q _3856_/S VGND VGND VPWR VPWR _3842_/B sky130_fd_sc_hd__nand2b_1
XFILLER_192_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6546_ _6746_/CLK _6546_/D fanout489/X VGND VGND VPWR VPWR _6546_/Q sky130_fd_sc_hd__dfrtp_4
X_3758_ input11/X _3355_/Y _3754_/X _3755_/X _3757_/X VGND VGND VPWR VPWR _3816_/A
+ sky130_fd_sc_hd__a2111o_1
XFILLER_145_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6477_ _6697_/CLK _6477_/D fanout486/X VGND VGND VPWR VPWR _6477_/Q sky130_fd_sc_hd__dfstp_1
X_3689_ _6931_/Q hold41/A _4267_/A _6671_/Q VGND VGND VPWR VPWR _3689_/X sky130_fd_sc_hd__a22o_1
XFILLER_173_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5428_ hold183/X hold46/X _5432_/S VGND VGND VPWR VPWR _5428_/X sky130_fd_sc_hd__mux2_1
Xoutput240 _3913_/X VGND VGND VPWR VPWR mgmt_gpio_out[36] sky130_fd_sc_hd__buf_12
Xoutput251 _3945_/X VGND VGND VPWR VPWR pad_flash_io0_do sky130_fd_sc_hd__buf_12
Xoutput262 _6737_/Q VGND VGND VPWR VPWR pll_div[0] sky130_fd_sc_hd__buf_12
XFILLER_160_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput273 _6429_/Q VGND VGND VPWR VPWR pll_trim[11] sky130_fd_sc_hd__buf_12
XFILLER_121_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput284 _6423_/Q VGND VGND VPWR VPWR pll_trim[21] sky130_fd_sc_hd__buf_12
X_5359_ hold610/X _5545_/A1 _5360_/S VGND VGND VPWR VPWR _5359_/X sky130_fd_sc_hd__mux2_1
XFILLER_160_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput295 _6426_/Q VGND VGND VPWR VPWR pll_trim[8] sky130_fd_sc_hd__buf_12
XFILLER_99_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_160_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7029_ _7029_/CLK _7029_/D fanout519/X VGND VGND VPWR VPWR _7029_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_43_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_168_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_183_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_172 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_323 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_376 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_20 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4730_ _4529_/X _4669_/Y _4729_/X _5040_/B _4730_/B2 VGND VGND VPWR VPWR _6720_/D
+ sky130_fd_sc_hd__o32a_1
XFILLER_14_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4661_ _4719_/B _4973_/A _4972_/A _4595_/Y VGND VGND VPWR VPWR _4662_/C sky130_fd_sc_hd__a31o_1
X_6400_ _6400_/A _6401_/B VGND VGND VPWR VPWR _6400_/X sky130_fd_sc_hd__and2_1
X_3612_ _6473_/Q _4026_/A _4285_/A _6688_/Q VGND VGND VPWR VPWR _3612_/X sky130_fd_sc_hd__a22o_2
XFILLER_175_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4592_ _4592_/A _4592_/B VGND VGND VPWR VPWR _4671_/B sky130_fd_sc_hd__nand2_4
XFILLER_190_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold904 _4204_/X VGND VGND VPWR VPWR _6610_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6331_ _6330_/X _6331_/A1 _6346_/S VGND VGND VPWR VPWR _7143_/D sky130_fd_sc_hd__mux2_1
X_3543_ _6926_/Q _5361_/A _5388_/A _6950_/Q _3542_/X VGND VGND VPWR VPWR _3548_/B
+ sky130_fd_sc_hd__a221o_1
Xhold915 _6905_/Q VGND VGND VPWR VPWR hold915/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold926 _4147_/X VGND VGND VPWR VPWR _6561_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold937 _6600_/Q VGND VGND VPWR VPWR hold937/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_115_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold948 _5336_/X VGND VGND VPWR VPWR _6899_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold959 _6671_/Q VGND VGND VPWR VPWR hold959/X sky130_fd_sc_hd__dlygate4sd3_1
X_6262_ _6683_/Q _5949_/X _5963_/X _6568_/Q _6261_/X VGND VGND VPWR VPWR _6268_/C
+ sky130_fd_sc_hd__a221o_1
X_3474_ _3533_/A _5161_/B VGND VGND VPWR VPWR _4166_/A sky130_fd_sc_hd__nor2_4
XFILLER_89_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_143_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_170_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5213_ hold225/X hold23/X _5216_/S VGND VGND VPWR VPWR _5213_/X sky130_fd_sc_hd__mux2_1
X_6193_ _6625_/Q _5973_/A _5971_/B _6609_/Q _6192_/X VGND VGND VPWR VPWR _6201_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_142_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5144_ hold941/X _6354_/A1 _5144_/S VGND VGND VPWR VPWR _5144_/X sky130_fd_sc_hd__mux2_1
XFILLER_96_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_318 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5075_ _4901_/A _4465_/B _4901_/B _5014_/D VGND VGND VPWR VPWR _5101_/B sky130_fd_sc_hd__o31a_1
XFILLER_56_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4026_ _4026_/A _5187_/B VGND VGND VPWR VPWR _4031_/S sky130_fd_sc_hd__and2_2
XFILLER_65_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5977_ _5977_/A _5981_/B _5981_/C VGND VGND VPWR VPWR _5977_/X sky130_fd_sc_hd__and3_4
X_4928_ _4479_/A _5026_/A _4962_/C _4676_/B _4813_/B VGND VGND VPWR VPWR _4932_/B
+ sky130_fd_sc_hd__o221a_1
XFILLER_60_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4859_ _4501_/B _4965_/C _5081_/A _4857_/X _4858_/X VGND VGND VPWR VPWR _4879_/B
+ sky130_fd_sc_hd__o2111a_1
XFILLER_166_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_176_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_176_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_621 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6529_ _7041_/CLK _6529_/D fanout518/X VGND VGND VPWR VPWR _6529_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_106_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_192_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_134_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_73_csclk clkbuf_3_2_0_csclk/X VGND VGND VPWR VPWR _6978_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_85_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_11_csclk _6684_/CLK VGND VGND VPWR VPWR _6633_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_8_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_157_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_137_481 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_26_csclk clkbuf_3_7_0_csclk/X VGND VGND VPWR VPWR _7022_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_166_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_98_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3190_ _7029_/Q VGND VGND VPWR VPWR _3190_/Y sky130_fd_sc_hd__inv_2
XFILLER_182_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5900_ _6668_/Q _5633_/X _5646_/X _6483_/Q VGND VGND VPWR VPWR _5900_/X sky130_fd_sc_hd__a22o_1
XFILLER_81_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6880_ _6881_/CLK _6880_/D fanout524/X VGND VGND VPWR VPWR _6880_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_62_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_179_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5831_ _6465_/Q _5629_/X _5630_/X _6705_/Q _5830_/X VGND VGND VPWR VPWR _5831_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_34_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_179_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5762_ _6959_/Q _5915_/A2 _5816_/B1 _6943_/Q VGND VGND VPWR VPWR _5763_/B sky130_fd_sc_hd__a22o_1
X_4713_ _4713_/A _4715_/B VGND VGND VPWR VPWR _4714_/C sky130_fd_sc_hd__nor2_1
XFILLER_147_201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5693_ _6916_/Q _5923_/B VGND VGND VPWR VPWR _5693_/X sky130_fd_sc_hd__and2b_1
XFILLER_148_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4644_ _4799_/A _4788_/A _4595_/Y _4631_/X _4984_/A VGND VGND VPWR VPWR _4644_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_135_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_621 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold701 _6839_/Q VGND VGND VPWR VPWR hold701/X sky130_fd_sc_hd__dlygate4sd3_1
X_4575_ _4575_/A _4575_/B VGND VGND VPWR VPWR _4575_/X sky130_fd_sc_hd__or2_2
Xmax_cap420 _5617_/X VGND VGND VPWR VPWR _5928_/A2 sky130_fd_sc_hd__buf_8
XFILLER_128_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold712 _5401_/X VGND VGND VPWR VPWR _6957_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold723 _6991_/Q VGND VGND VPWR VPWR hold723/X sky130_fd_sc_hd__dlygate4sd3_1
X_3526_ _6430_/Q _3975_/A _4214_/A _6623_/Q _3524_/X VGND VGND VPWR VPWR _3535_/B
+ sky130_fd_sc_hd__a221o_1
X_6314_ _3471_/X _6314_/A1 _6316_/S VGND VGND VPWR VPWR _7138_/D sky130_fd_sc_hd__mux2_1
Xhold734 _5473_/X VGND VGND VPWR VPWR _7021_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_142 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold745 _7029_/Q VGND VGND VPWR VPWR hold745/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold756 _5464_/X VGND VGND VPWR VPWR _7013_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold767 _6887_/Q VGND VGND VPWR VPWR hold767/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold778 _4023_/X VGND VGND VPWR VPWR _6467_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6245_ _6472_/Q _5941_/Y _6285_/A2 _6632_/Q _6244_/X VGND VGND VPWR VPWR _6251_/C
+ sky130_fd_sc_hd__a221o_1
Xhold789 _6662_/Q VGND VGND VPWR VPWR hold789/X sky130_fd_sc_hd__dlygate4sd3_1
X_3457_ _6847_/Q _5271_/A _5343_/A _6911_/Q _3456_/X VGND VGND VPWR VPWR _3460_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_103_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6176_ _6985_/Q _6176_/A2 _6173_/X _6175_/X VGND VGND VPWR VPWR _6177_/C sky130_fd_sc_hd__a211o_1
XFILLER_162_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3388_ _6865_/Q _5289_/A _5244_/A _6825_/Q _3385_/X VGND VGND VPWR VPWR _3395_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_69_262 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1401 _6596_/Q VGND VGND VPWR VPWR _4187_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_85_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1412 _7139_/Q VGND VGND VPWR VPWR _6315_/A1 sky130_fd_sc_hd__dlygate4sd3_1
X_5127_ _6725_/Q _4222_/X _5121_/X _5126_/X _5120_/Y VGND VGND VPWR VPWR _5127_/X
+ sky130_fd_sc_hd__a221o_1
Xhold1423 _5180_/X VGND VGND VPWR VPWR hold664/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_84_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_593 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1434 _7165_/Q VGND VGND VPWR VPWR hold112/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1445 _6727_/Q VGND VGND VPWR VPWR _3818_/A1 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1456 _6486_/Q VGND VGND VPWR VPWR _3904_/B1 sky130_fd_sc_hd__dlygate4sd3_1
X_5058_ _5058_/A _5058_/B _5055_/X VGND VGND VPWR VPWR _5058_/X sky130_fd_sc_hd__or3b_1
Xhold1467 _7147_/Q VGND VGND VPWR VPWR _6343_/A1 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1478 _6105_/X VGND VGND VPWR VPWR _7123_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_84_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1489 _5823_/X VGND VGND VPWR VPWR _7113_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4009_ _4009_/A0 _5488_/A1 _4013_/S VGND VGND VPWR VPWR _4009_/X sky130_fd_sc_hd__mux2_1
XTAP_2928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_696 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_470 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_161_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_161_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_156 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold50 hold50/A VGND VGND VPWR VPWR hold50/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_152_40 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold61 hold61/A VGND VGND VPWR VPWR hold61/X sky130_fd_sc_hd__buf_12
Xhold72 hold72/A VGND VGND VPWR VPWR hold72/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold83 hold83/A VGND VGND VPWR VPWR hold83/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_63_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold94 hold94/A VGND VGND VPWR VPWR hold94/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_35_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_151 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_346 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_188_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_598 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_3 _3975_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_184_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4360_ _4345_/C _4351_/Y _4886_/A _4888_/B VGND VGND VPWR VPWR _4471_/A sky130_fd_sc_hd__o211ai_4
XFILLER_6_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3311_ hold59/X hold31/X VGND VGND VPWR VPWR hold60/A sky130_fd_sc_hd__nand2b_1
XFILLER_98_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4291_ _4291_/A hold7/X VGND VGND VPWR VPWR _4296_/S sky130_fd_sc_hd__and2_2
XFILLER_112_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6030_ _6054_/A2 _6305_/A2 _6028_/X _6029_/X VGND VGND VPWR VPWR _7120_/D sky130_fd_sc_hd__o22a_1
XFILLER_113_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3242_ _3242_/A _3249_/S VGND VGND VPWR VPWR _3246_/A sky130_fd_sc_hd__nor2_1
XFILLER_79_571 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3173_ _6509_/Q VGND VGND VPWR VPWR _3876_/A sky130_fd_sc_hd__inv_2
XFILLER_66_276 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6932_ _6948_/CLK _6932_/D fanout514/X VGND VGND VPWR VPWR _6932_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_19_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6863_ _6999_/CLK _6863_/D fanout523/X VGND VGND VPWR VPWR _6863_/Q sky130_fd_sc_hd__dfrtp_1
X_5814_ _7017_/Q _5921_/A2 _5912_/B1 _7033_/Q _5813_/X VGND VGND VPWR VPWR _5817_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_167_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6794_ _7039_/CLK _6794_/D fanout498/X VGND VGND VPWR VPWR _6794_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_50_666 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5745_ _6846_/Q _5922_/B1 _5651_/X _6798_/Q VGND VGND VPWR VPWR _5745_/X sky130_fd_sc_hd__a22o_1
X_5676_ _6867_/Q _5928_/B1 _5913_/B1 _6883_/Q VGND VGND VPWR VPWR _5676_/X sky130_fd_sc_hd__a22o_1
XFILLER_163_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4627_ _4924_/B _4779_/A _4784_/A VGND VGND VPWR VPWR _4649_/B sky130_fd_sc_hd__or3b_1
XFILLER_135_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_190_343 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_259 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold520 _5203_/X VGND VGND VPWR VPWR _6781_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold531 _6564_/Q VGND VGND VPWR VPWR hold531/X sky130_fd_sc_hd__dlygate4sd3_1
X_4558_ _4447_/Y _4898_/B _4542_/A VGND VGND VPWR VPWR _4559_/D sky130_fd_sc_hd__a21o_1
XFILLER_190_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold542 _3966_/X VGND VGND VPWR VPWR _6421_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold553 _6628_/Q VGND VGND VPWR VPWR hold553/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold564 _4251_/X VGND VGND VPWR VPWR _6656_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_103_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3509_ _3525_/A _3560_/B VGND VGND VPWR VPWR _4249_/A sky130_fd_sc_hd__nor2_4
XFILLER_89_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold575 _6699_/Q VGND VGND VPWR VPWR hold575/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_143_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_173_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold586 _5507_/X VGND VGND VPWR VPWR _7051_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4489_ _4947_/A _4489_/B VGND VGND VPWR VPWR _5106_/A sky130_fd_sc_hd__nand2_2
Xhold597 _4277_/X VGND VGND VPWR VPWR _6678_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6228_ _6541_/Q _6004_/B _6218_/X _6227_/X _5610_/A VGND VGND VPWR VPWR _6228_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_103_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6159_ _6913_/Q _5972_/A _6283_/A2 _7070_/Q VGND VGND VPWR VPWR _6159_/X sky130_fd_sc_hd__a22o_1
Xhold1220 _4209_/X VGND VGND VPWR VPWR _6614_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1231 _6470_/Q VGND VGND VPWR VPWR _4027_/A0 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1242 _5425_/X VGND VGND VPWR VPWR _6978_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1253 _7010_/Q VGND VGND VPWR VPWR _5461_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_73_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1264 _4152_/X VGND VGND VPWR VPWR _6565_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1275 _6874_/Q VGND VGND VPWR VPWR _5308_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_122_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_427 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1286 _5321_/X VGND VGND VPWR VPWR _6886_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_45_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1297 _6878_/Q VGND VGND VPWR VPWR _5312_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_154_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput140 wb_dat_i[17] VGND VGND VPWR VPWR _6326_/A2 sky130_fd_sc_hd__clkbuf_1
Xinput151 wb_dat_i[27] VGND VGND VPWR VPWR _6332_/A2 sky130_fd_sc_hd__clkbuf_1
Xinput162 wb_dat_i[8] VGND VGND VPWR VPWR _6323_/B1 sky130_fd_sc_hd__clkbuf_1
XFILLER_36_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3860_ _3904_/A2 _6406_/Q _3860_/S VGND VGND VPWR VPWR _6406_/D sky130_fd_sc_hd__mux2_1
XFILLER_31_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3791_ _6599_/Q _4190_/A _4208_/A _6614_/Q _3790_/X VGND VGND VPWR VPWR _3792_/D
+ sky130_fd_sc_hd__a221o_1
XPHY_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5530_ _5530_/A0 _5530_/A1 _5537_/S VGND VGND VPWR VPWR _5530_/X sky130_fd_sc_hd__mux2_1
XFILLER_75_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_204 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5461_ _5461_/A0 _5530_/A1 _5468_/S VGND VGND VPWR VPWR _5461_/X sky130_fd_sc_hd__mux2_1
XFILLER_117_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4412_ _4679_/A _4554_/A _4691_/A VGND VGND VPWR VPWR _5022_/A sky130_fd_sc_hd__nand3_4
X_7200_ _7200_/A VGND VGND VPWR VPWR _7200_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_172_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5392_ hold859/X _5542_/A1 _5396_/S VGND VGND VPWR VPWR _5392_/X sky130_fd_sc_hd__mux2_1
X_7131_ _7131_/CLK _7131_/D fanout497/X VGND VGND VPWR VPWR _7131_/Q sky130_fd_sc_hd__dfrtp_1
X_4343_ _4617_/B _4888_/A _4356_/B _4592_/A VGND VGND VPWR VPWR _4345_/C sky130_fd_sc_hd__and4_2
XFILLER_125_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7062_ _7078_/CLK _7062_/D fanout507/X VGND VGND VPWR VPWR _7062_/Q sky130_fd_sc_hd__dfrtp_1
X_4274_ _4274_/A0 _6353_/A1 _4278_/S VGND VGND VPWR VPWR _4274_/X sky130_fd_sc_hd__mux2_1
X_6013_ _7011_/Q _5976_/Y _5979_/X _6971_/Q _6010_/X VGND VGND VPWR VPWR _6027_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_86_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3225_ _4596_/B VGND VGND VPWR VPWR _4691_/A sky130_fd_sc_hd__inv_6
XFILLER_100_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6915_ _7046_/CLK _6915_/D fanout497/X VGND VGND VPWR VPWR _6915_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_82_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6846_ _7041_/CLK _6846_/D fanout520/X VGND VGND VPWR VPWR _6846_/Q sky130_fd_sc_hd__dfrtp_2
X_6777_ _6881_/CLK _6777_/D fanout523/X VGND VGND VPWR VPWR _7196_/A sky130_fd_sc_hd__dfrtp_1
X_3989_ hold389/X _5534_/A1 _3992_/S VGND VGND VPWR VPWR _3989_/X sky130_fd_sc_hd__mux2_1
X_5728_ _6957_/Q _5915_/A2 _5816_/B1 _6941_/Q VGND VGND VPWR VPWR _5728_/X sky130_fd_sc_hd__a22o_1
XFILLER_6_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_148_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5659_ _6946_/Q _5626_/X _5648_/X _6962_/Q VGND VGND VPWR VPWR _5659_/X sky130_fd_sc_hd__a22o_1
XFILLER_136_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold350 _5320_/X VGND VGND VPWR VPWR _6885_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold361 _6924_/Q VGND VGND VPWR VPWR hold361/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold372 _5355_/X VGND VGND VPWR VPWR _6916_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold383 _6759_/Q VGND VGND VPWR VPWR hold383/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold394 _3980_/X VGND VGND VPWR VPWR _6430_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_132_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_117_98 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_295 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1050 _7027_/Q VGND VGND VPWR VPWR _5480_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_133_64 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1061 _3986_/X VGND VGND VPWR VPWR _6435_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1072 _5171_/X VGND VGND VPWR VPWR _6756_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_100_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1083 _7018_/Q VGND VGND VPWR VPWR _5470_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1094 _5188_/X VGND VGND VPWR VPWR _6768_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_93_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_201 _5928_/B1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_212 hold114/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_655 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_154_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_174_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_179 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_596 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_408 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4961_ _5022_/A _4556_/A _5043_/B _4789_/B _4668_/X VGND VGND VPWR VPWR _4961_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_17_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6700_ _7034_/CLK _6700_/D fanout490/X VGND VGND VPWR VPWR _6700_/Q sky130_fd_sc_hd__dfrtp_1
X_3912_ _6523_/Q input91/X _3915_/S VGND VGND VPWR VPWR _3912_/X sky130_fd_sc_hd__mux2_2
X_4892_ _4892_/A _4892_/B VGND VGND VPWR VPWR _4911_/C sky130_fd_sc_hd__nor2_1
X_6631_ _6632_/CLK _6631_/D _3264_/A VGND VGND VPWR VPWR _6631_/Q sky130_fd_sc_hd__dfrtp_4
X_3843_ _3843_/A _3843_/B VGND VGND VPWR VPWR _6412_/D sky130_fd_sc_hd__xor2_1
XFILLER_20_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3774_ _7018_/Q hold18/A hold62/A _6650_/Q _3773_/X VGND VGND VPWR VPWR _3777_/C
+ sky130_fd_sc_hd__a221o_1
X_6562_ _6689_/CLK _6562_/D _6370_/A VGND VGND VPWR VPWR _6562_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_118_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5513_ hold945/X _5531_/A1 _5519_/S VGND VGND VPWR VPWR _5513_/X sky130_fd_sc_hd__mux2_1
XFILLER_157_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6493_ _6527_/CLK _6493_/D fanout524/X VGND VGND VPWR VPWR _7184_/A sky130_fd_sc_hd__dfrtp_1
XFILLER_118_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_133_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5444_ hold982/X _5495_/A1 _5450_/S VGND VGND VPWR VPWR _5444_/X sky130_fd_sc_hd__mux2_1
XFILLER_105_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5375_ _5375_/A0 _5543_/A1 hold42/X VGND VGND VPWR VPWR _5375_/X sky130_fd_sc_hd__mux2_1
X_7114_ _7130_/CLK _7114_/D fanout485/X VGND VGND VPWR VPWR _7114_/Q sky130_fd_sc_hd__dfrtp_1
X_4326_ hold309/X _6357_/A1 _4326_/S VGND VGND VPWR VPWR _4326_/X sky130_fd_sc_hd__mux2_1
XFILLER_101_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4257_ hold791/X _4299_/A1 _4260_/S VGND VGND VPWR VPWR _4257_/X sky130_fd_sc_hd__mux2_1
X_7045_ _7072_/CLK _7045_/D fanout506/X VGND VGND VPWR VPWR _7045_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_101_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3208_ _6893_/Q VGND VGND VPWR VPWR _3208_/Y sky130_fd_sc_hd__inv_2
XFILLER_170_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4188_ _3433_/X _4188_/A1 _4189_/S VGND VGND VPWR VPWR _6597_/D sky130_fd_sc_hd__mux2_1
XFILLER_28_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6829_ _7078_/CLK _6829_/D fanout515/X VGND VGND VPWR VPWR _6829_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_11_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_647 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_149_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_183_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_546 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_343 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold180 _6535_/Q VGND VGND VPWR VPWR hold180/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold191 _6431_/Q VGND VGND VPWR VPWR hold191/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_77_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_63 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_160_40 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3490_ hold61/X _3538_/B VGND VGND VPWR VPWR _4225_/A sky130_fd_sc_hd__nor2_8
XFILLER_170_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5160_ _5160_/A0 _6354_/A1 _5160_/S VGND VGND VPWR VPWR _5160_/X sky130_fd_sc_hd__mux2_1
XFILLER_38_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4111_ _4111_/A0 hold27/X _4111_/S VGND VGND VPWR VPWR hold28/A sky130_fd_sc_hd__mux2_1
XFILLER_96_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5091_ _5091_/A VGND VGND VPWR VPWR _5121_/C sky130_fd_sc_hd__clkinv_2
XFILLER_96_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4042_ hold600/X _4289_/A1 _4043_/S VGND VGND VPWR VPWR _4042_/X sky130_fd_sc_hd__mux2_1
XFILLER_96_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_341 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5993_ _6442_/Q _6295_/A2 _6288_/A2 _6914_/Q _5982_/X VGND VGND VPWR VPWR _5996_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_40_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4944_ _4944_/A _4944_/B _4946_/C VGND VGND VPWR VPWR _4944_/X sky130_fd_sc_hd__and3_1
XFILLER_177_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4875_ _4901_/B _4973_/A _4972_/A _4748_/B VGND VGND VPWR VPWR _4877_/C sky130_fd_sc_hd__o22a_1
X_6614_ _6630_/CLK _6614_/D fanout492/X VGND VGND VPWR VPWR _6614_/Q sky130_fd_sc_hd__dfrtp_4
X_3826_ _3826_/A _3826_/B VGND VGND VPWR VPWR _6415_/D sky130_fd_sc_hd__nor2_1
XFILLER_165_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_192_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_146_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6545_ _6697_/CLK _6545_/D fanout489/X VGND VGND VPWR VPWR _6545_/Q sky130_fd_sc_hd__dfrtp_2
X_3757_ _6426_/Q _3975_/A _4279_/A _6680_/Q _3756_/X VGND VGND VPWR VPWR _3757_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_146_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_118_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6476_ _6769_/CLK _6476_/D _6399_/A VGND VGND VPWR VPWR _6476_/Q sky130_fd_sc_hd__dfrtp_2
X_3688_ _6651_/Q hold62/A _4038_/A _6481_/Q _3687_/X VGND VGND VPWR VPWR _3713_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_145_184 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5427_ hold453/X _5541_/A1 _5432_/S VGND VGND VPWR VPWR _5427_/X sky130_fd_sc_hd__mux2_1
Xoutput230 _7192_/X VGND VGND VPWR VPWR mgmt_gpio_out[27] sky130_fd_sc_hd__buf_12
Xoutput241 _3912_/X VGND VGND VPWR VPWR mgmt_gpio_out[37] sky130_fd_sc_hd__buf_12
Xoutput252 _3942_/A VGND VGND VPWR VPWR pad_flash_io0_ieb sky130_fd_sc_hd__buf_12
Xoutput263 _6738_/Q VGND VGND VPWR VPWR pll_div[1] sky130_fd_sc_hd__buf_12
XFILLER_161_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput274 _6430_/Q VGND VGND VPWR VPWR pll_trim[12] sky130_fd_sc_hd__buf_12
XFILLER_160_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5358_ hold159/X hold142/X _5360_/S VGND VGND VPWR VPWR _5358_/X sky130_fd_sc_hd__mux2_1
Xoutput285 _6424_/Q VGND VGND VPWR VPWR pll_trim[22] sky130_fd_sc_hd__buf_12
XFILLER_58_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_411 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput296 _6427_/Q VGND VGND VPWR VPWR pll_trim[9] sky130_fd_sc_hd__buf_12
XFILLER_59_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4309_ _4309_/A _6352_/B VGND VGND VPWR VPWR _4314_/S sky130_fd_sc_hd__and2_2
X_5289_ _5289_/A _5529_/B VGND VGND VPWR VPWR _5297_/S sky130_fd_sc_hd__and2_4
XFILLER_75_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7028_ _7083_/CLK _7028_/D fanout518/X VGND VGND VPWR VPWR _7028_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_28_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire346 _3489_/Y VGND VGND VPWR VPWR _3567_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_137_630 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_136_184 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_335 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout490 fanout526/X VGND VGND VPWR VPWR fanout490/X sky130_fd_sc_hd__buf_12
XFILLER_48_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_171_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_330 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_514 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_32 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_147_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_187_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4660_ _4789_/B _4649_/A _4594_/X _4721_/B _4659_/X VGND VGND VPWR VPWR _4662_/B
+ sky130_fd_sc_hd__o221a_1
XFILLER_30_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3611_ _6421_/Q _3958_/A _3984_/A _6437_/Q _3610_/X VGND VGND VPWR VPWR _3614_/C
+ sky130_fd_sc_hd__a221o_2
X_4591_ _4799_/A _4985_/A _6643_/Q VGND VGND VPWR VPWR _4915_/B sky130_fd_sc_hd__o21a_1
XFILLER_190_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6330_ _6644_/Q _6330_/A2 _6330_/B1 _6643_/Q _6329_/X VGND VGND VPWR VPWR _6330_/X
+ sky130_fd_sc_hd__a221o_1
Xhold905 _7012_/Q VGND VGND VPWR VPWR hold905/X sky130_fd_sc_hd__dlygate4sd3_1
X_3542_ _7014_/Q _5460_/A _6352_/A _7155_/Q VGND VGND VPWR VPWR _3542_/X sky130_fd_sc_hd__a22o_1
Xhold916 _5342_/X VGND VGND VPWR VPWR _6905_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold927 _7003_/Q VGND VGND VPWR VPWR hold927/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold938 _4192_/X VGND VGND VPWR VPWR _6600_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_127_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold949 _6701_/Q VGND VGND VPWR VPWR hold949/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3473_ _3472_/X _3473_/A1 _3749_/S VGND VGND VPWR VPWR _3473_/X sky130_fd_sc_hd__mux2_1
X_6261_ _6602_/Q _5939_/X _5943_/Y _6463_/Q VGND VGND VPWR VPWR _6261_/X sky130_fd_sc_hd__a22o_1
X_5212_ hold239/X _5533_/A1 _5216_/S VGND VGND VPWR VPWR _5212_/X sky130_fd_sc_hd__mux2_1
XFILLER_170_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6192_ _6578_/Q _5946_/X _5959_/Y _6614_/Q VGND VGND VPWR VPWR _6192_/X sky130_fd_sc_hd__a22o_1
XFILLER_69_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5143_ _5143_/A0 _6353_/A1 _5144_/S VGND VGND VPWR VPWR _5143_/X sky130_fd_sc_hd__mux2_1
XFILLER_97_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5074_ _5074_/A _5074_/B _5074_/C VGND VGND VPWR VPWR _5102_/B sky130_fd_sc_hd__and3_1
XFILLER_111_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4025_ hold449/X _5534_/A1 _4025_/S VGND VGND VPWR VPWR _4025_/X sky130_fd_sc_hd__mux2_1
XFILLER_25_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_344 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5976_ _5976_/A _5980_/B VGND VGND VPWR VPWR _5976_/Y sky130_fd_sc_hd__nor2_8
XFILLER_52_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4927_ _4984_/C _5064_/B _5108_/B VGND VGND VPWR VPWR _4927_/X sky130_fd_sc_hd__and3_1
XFILLER_33_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_178_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4858_ _4861_/B _4620_/B _4684_/Y VGND VGND VPWR VPWR _4858_/X sky130_fd_sc_hd__o21ba_1
XFILLER_166_736 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3809_ _6922_/Q _5361_/A _6352_/A _7151_/Q VGND VGND VPWR VPWR _3809_/X sky130_fd_sc_hd__a22o_1
X_4789_ _4789_/A _4789_/B VGND VGND VPWR VPWR _5081_/B sky130_fd_sc_hd__or2_1
XFILLER_180_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6528_ _7041_/CLK _6528_/D fanout518/X VGND VGND VPWR VPWR _6528_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_118_173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_7_csclk clkbuf_3_1_0_csclk/X VGND VGND VPWR VPWR _6565_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_106_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6459_ _6565_/CLK _6459_/D fanout495/X VGND VGND VPWR VPWR _6459_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_133_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_121_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_198 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_163 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_169_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_129_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_169_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_98_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_263 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5830_ _6475_/Q _5620_/X _5639_/X _6550_/Q VGND VGND VPWR VPWR _5830_/X sky130_fd_sc_hd__a22o_1
XFILLER_62_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5761_ _7007_/Q _5912_/A2 _5618_/X _6879_/Q VGND VGND VPWR VPWR _5763_/A sky130_fd_sc_hd__a22o_1
X_4712_ _4603_/Y _4673_/Y _4767_/B _4711_/X VGND VGND VPWR VPWR _4714_/B sky130_fd_sc_hd__a211o_1
XFILLER_147_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5692_ _6964_/Q _5925_/B1 _5650_/X _6892_/Q VGND VGND VPWR VPWR _5692_/X sky130_fd_sc_hd__a22o_1
XFILLER_187_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4643_ _4799_/A _4788_/A VGND VGND VPWR VPWR _5067_/A sky130_fd_sc_hd__nor2_1
XFILLER_175_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmax_cap410 _5630_/X VGND VGND VPWR VPWR _5915_/A2 sky130_fd_sc_hd__buf_12
X_4574_ _4574_/A _4574_/B VGND VGND VPWR VPWR _4574_/Y sky130_fd_sc_hd__nor2_1
Xhold702 _5268_/X VGND VGND VPWR VPWR _6839_/D sky130_fd_sc_hd__dlygate4sd3_1
Xmax_cap421 _5614_/X VGND VGND VPWR VPWR _5912_/A2 sky130_fd_sc_hd__buf_12
XFILLER_116_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold713 _7082_/Q VGND VGND VPWR VPWR hold713/X sky130_fd_sc_hd__dlygate4sd3_1
X_6313_ _6313_/A0 _6313_/A1 _6316_/S VGND VGND VPWR VPWR _7137_/D sky130_fd_sc_hd__mux2_1
XFILLER_115_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold724 _5439_/X VGND VGND VPWR VPWR _6991_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3525_ _3525_/A hold53/A VGND VGND VPWR VPWR _4214_/A sky130_fd_sc_hd__nor2_4
Xhold735 _6917_/Q VGND VGND VPWR VPWR hold735/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold746 _5482_/X VGND VGND VPWR VPWR _7029_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_154 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold757 _6879_/Q VGND VGND VPWR VPWR hold757/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_103_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold768 _5322_/X VGND VGND VPWR VPWR _6887_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold779 _7036_/Q VGND VGND VPWR VPWR hold779/X sky130_fd_sc_hd__dlygate4sd3_1
X_6244_ _6552_/Q _5973_/B _5963_/X _6567_/Q VGND VGND VPWR VPWR _6244_/X sky130_fd_sc_hd__a22o_1
X_3456_ _6887_/Q hold83/A _5334_/A _6903_/Q VGND VGND VPWR VPWR _3456_/X sky130_fd_sc_hd__a22o_1
X_6175_ _6801_/Q _6299_/A2 _6294_/A2 _7086_/Q _6174_/X VGND VGND VPWR VPWR _6175_/X
+ sky130_fd_sc_hd__a221o_1
X_3387_ hold82/A _3523_/A VGND VGND VPWR VPWR _5244_/A sky130_fd_sc_hd__nor2_8
XFILLER_97_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1402 _6589_/Q VGND VGND VPWR VPWR _4179_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_69_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1413 _7135_/Q VGND VGND VPWR VPWR _6311_/A1 sky130_fd_sc_hd__dlygate4sd3_1
X_5126_ _5126_/A _5134_/B VGND VGND VPWR VPWR _5126_/X sky130_fd_sc_hd__or2_1
Xhold1424 _6574_/Q VGND VGND VPWR VPWR _4162_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_57_436 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1435 _3971_/X VGND VGND VPWR VPWR hold113/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1446 _6734_/Q VGND VGND VPWR VPWR _3399_/A1 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1457 _3861_/X VGND VGND VPWR VPWR _6405_/D sky130_fd_sc_hd__dlygate4sd3_1
X_5057_ _5057_/A _5058_/B VGND VGND VPWR VPWR _5116_/B sky130_fd_sc_hd__nor2_1
Xhold1468 hold67/A VGND VGND VPWR VPWR _6337_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_55_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1479 _6414_/Q VGND VGND VPWR VPWR _3835_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_44_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4008_ _4008_/A _6352_/B VGND VGND VPWR VPWR _4013_/S sky130_fd_sc_hd__and2_2
XTAP_2918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5959_ _5959_/A _5965_/B VGND VGND VPWR VPWR _5959_/Y sky130_fd_sc_hd__nor2_8
XFILLER_40_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_482 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_162_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold40 hold40/A VGND VGND VPWR VPWR hold40/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_29_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold51 hold51/A VGND VGND VPWR VPWR hold51/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold62 hold62/A VGND VGND VPWR VPWR hold62/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_152_52 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold73 hold73/A VGND VGND VPWR VPWR hold73/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold84 hold84/A VGND VGND VPWR VPWR hold84/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_152_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold95 hold95/A VGND VGND VPWR VPWR hold95/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_63_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_358 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_176_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_543 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_144_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_4 _5208_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3310_ hold58/X hold16/X VGND VGND VPWR VPWR hold59/A sky130_fd_sc_hd__or2_1
X_4290_ hold535/X _6357_/A1 _4290_/S VGND VGND VPWR VPWR _4290_/X sky130_fd_sc_hd__mux2_1
XFILLER_113_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_140_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3241_ _3867_/A _3828_/B _3256_/S _3235_/Y VGND VGND VPWR VPWR _3249_/S sky130_fd_sc_hd__o31a_1
XFILLER_79_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3172_ _3172_/A VGND VGND VPWR VPWR _5570_/A sky130_fd_sc_hd__inv_2
XFILLER_79_583 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_436 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_288 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6931_ _7074_/CLK _6931_/D fanout505/X VGND VGND VPWR VPWR _6931_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_81_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_236 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6862_ _7083_/CLK _6862_/D fanout518/X VGND VGND VPWR VPWR _6862_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_179_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5813_ _6953_/Q _5924_/B2 _5926_/A2 _6809_/Q VGND VGND VPWR VPWR _5813_/X sky130_fd_sc_hd__a22o_1
XFILLER_50_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6793_ _7072_/CLK _6793_/D fanout507/X VGND VGND VPWR VPWR _6793_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_167_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_509 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_678 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5744_ _6894_/Q _5650_/X _5740_/X _5741_/X _5743_/X VGND VGND VPWR VPWR _5744_/X
+ sky130_fd_sc_hd__a2111o_1
XFILLER_188_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5675_ _6979_/Q _5642_/X _5644_/X _6971_/Q _5670_/Y VGND VGND VPWR VPWR _5675_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_136_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_190_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_148_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4626_ _4799_/A _4778_/C _4778_/B VGND VGND VPWR VPWR _4924_/B sky130_fd_sc_hd__a21bo_1
Xhold510 _5365_/X VGND VGND VPWR VPWR _6925_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_190_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold521 _6451_/Q VGND VGND VPWR VPWR hold521/X sky130_fd_sc_hd__dlygate4sd3_1
X_4557_ _5025_/A _4557_/B VGND VGND VPWR VPWR _4898_/B sky130_fd_sc_hd__nand2_1
Xhold532 _4150_/X VGND VGND VPWR VPWR _6564_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold543 _6582_/Q VGND VGND VPWR VPWR hold543/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_190_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold554 _4229_/X VGND VGND VPWR VPWR _6628_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold565 _6456_/Q VGND VGND VPWR VPWR hold565/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3508_ _6830_/Q _5253_/A _4273_/A _6679_/Q VGND VGND VPWR VPWR _3508_/X sky130_fd_sc_hd__a22o_1
XFILLER_131_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold576 _4302_/X VGND VGND VPWR VPWR _6699_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4488_ _5025_/B _4489_/B VGND VGND VPWR VPWR _4523_/A sky130_fd_sc_hd__nand2_1
Xhold587 _7141_/Q VGND VGND VPWR VPWR hold587/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold598 _6688_/Q VGND VGND VPWR VPWR hold598/X sky130_fd_sc_hd__dlygate4sd3_1
X_6227_ _6227_/A _6227_/B _6227_/C _6004_/B VGND VGND VPWR VPWR _6227_/X sky130_fd_sc_hd__or4b_1
XFILLER_104_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3439_ _7118_/Q _6760_/Q _6762_/Q VGND VGND VPWR VPWR _3439_/X sky130_fd_sc_hd__mux2_2
XFILLER_58_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_211 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6158_ _7001_/Q _6282_/A2 _6300_/B1 _6881_/Q _6157_/X VGND VGND VPWR VPWR _6168_/A
+ sky130_fd_sc_hd__a221o_1
XTAP_881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1210 _4310_/X VGND VGND VPWR VPWR _6705_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1221 _6685_/Q VGND VGND VPWR VPWR _4286_/A0 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_10_csclk _6684_/CLK VGND VGND VPWR VPWR _6689_/CLK sky130_fd_sc_hd__clkbuf_16
Xhold1232 _4027_/X VGND VGND VPWR VPWR _6470_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1243 _7055_/Q VGND VGND VPWR VPWR _5512_/A0 sky130_fd_sc_hd__dlygate4sd3_1
X_5109_ _4988_/A _4788_/A _4786_/Y _4631_/X _4725_/B VGND VGND VPWR VPWR _5110_/C
+ sky130_fd_sc_hd__o32a_1
Xhold1254 _5461_/X VGND VGND VPWR VPWR _7010_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6089_ _7067_/Q _6283_/A2 _5981_/X _6934_/Q _6088_/X VGND VGND VPWR VPWR _6092_/A
+ sky130_fd_sc_hd__a221o_1
Xhold1265 _6906_/Q VGND VGND VPWR VPWR _5344_/A0 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1276 _5308_/X VGND VGND VPWR VPWR _6874_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_72_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1287 _6798_/Q VGND VGND VPWR VPWR _5222_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1298 _5312_/X VGND VGND VPWR VPWR _6878_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_122_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_25_csclk clkbuf_3_7_0_csclk/X VGND VGND VPWR VPWR _7084_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_53_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_186_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_154_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_107_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_606 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput130 wb_adr_i[9] VGND VGND VPWR VPWR _4336_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_163_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput141 wb_dat_i[18] VGND VGND VPWR VPWR _6329_/A2 sky130_fd_sc_hd__clkbuf_1
Xinput152 wb_dat_i[28] VGND VGND VPWR VPWR _6336_/A2 sky130_fd_sc_hd__clkbuf_1
Xinput163 wb_dat_i[9] VGND VGND VPWR VPWR _6326_/B1 sky130_fd_sc_hd__clkbuf_1
XFILLER_36_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_612 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_177_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_155 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3790_ _6906_/Q _5343_/A _3789_/Y _6750_/Q VGND VGND VPWR VPWR _3790_/X sky130_fd_sc_hd__a22o_1
XFILLER_176_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_191_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5460_ _5460_/A _5511_/B VGND VGND VPWR VPWR _5468_/S sky130_fd_sc_hd__and2_4
XFILLER_117_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4411_ _4679_/A _4554_/A _4691_/A VGND VGND VPWR VPWR _5025_/A sky130_fd_sc_hd__and3_4
X_5391_ hold411/X _5541_/A1 _5396_/S VGND VGND VPWR VPWR _5391_/X sky130_fd_sc_hd__mux2_1
X_7130_ _7130_/CLK _7130_/D fanout488/X VGND VGND VPWR VPWR _7130_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_113_411 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4342_ _4617_/B _4356_/B _4592_/A VGND VGND VPWR VPWR _4352_/B sky130_fd_sc_hd__and3_1
X_7061_ _7069_/CLK _7061_/D fanout516/X VGND VGND VPWR VPWR _7061_/Q sky130_fd_sc_hd__dfrtp_1
X_4273_ _4273_/A _5187_/B VGND VGND VPWR VPWR _4278_/S sky130_fd_sc_hd__and2_2
XFILLER_101_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_140_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6012_ _6851_/Q wire390/X _6270_/B1 _6931_/Q _6011_/X VGND VGND VPWR VPWR _6012_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_98_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_140_274 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3224_ _6921_/Q VGND VGND VPWR VPWR _3224_/Y sky130_fd_sc_hd__inv_2
.ends

