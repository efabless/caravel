magic
tech sky130A
magscale 1 2
timestamp 1665668947
<< viali >>
rect 1409 13481 1443 13515
rect 4721 13481 4755 13515
rect 9505 13481 9539 13515
rect 10241 13481 10275 13515
rect 6377 13413 6411 13447
rect 6745 13413 6779 13447
rect 8125 13413 8159 13447
rect 10609 13413 10643 13447
rect 2329 13345 2363 13379
rect 2973 13345 3007 13379
rect 4169 13345 4203 13379
rect 5089 13345 5123 13379
rect 5641 13345 5675 13379
rect 5825 13345 5859 13379
rect 12725 13345 12759 13379
rect 1593 13277 1627 13311
rect 2421 13277 2455 13311
rect 3065 13277 3099 13311
rect 3985 13277 4019 13311
rect 6561 13277 6595 13311
rect 6877 13277 6911 13311
rect 7021 13277 7055 13311
rect 7297 13277 7331 13311
rect 7389 13277 7423 13311
rect 8304 13277 8338 13311
rect 8677 13277 8711 13311
rect 9137 13277 9171 13311
rect 10885 13277 10919 13311
rect 11069 13277 11103 13311
rect 11161 13277 11195 13311
rect 12081 13277 12115 13311
rect 12173 13277 12207 13311
rect 13093 13277 13127 13311
rect 13461 13277 13495 13311
rect 2053 13209 2087 13243
rect 2145 13209 2179 13243
rect 2881 13209 2915 13243
rect 3525 13209 3559 13243
rect 3617 13209 3651 13243
rect 4077 13209 4111 13243
rect 4997 13209 5031 13243
rect 5549 13209 5583 13243
rect 6009 13209 6043 13243
rect 7113 13209 7147 13243
rect 7849 13209 7883 13243
rect 7941 13209 7975 13243
rect 8401 13209 8435 13243
rect 8493 13209 8527 13243
rect 9321 13209 9355 13243
rect 9505 13209 9539 13243
rect 10701 13209 10735 13243
rect 11529 13209 11563 13243
rect 11621 13209 11655 13243
rect 12633 13209 12667 13243
rect 13369 13209 13403 13243
rect 3801 13141 3835 13175
rect 4445 13141 4479 13175
rect 4905 13141 4939 13175
rect 6101 13141 6135 13175
rect 8953 13141 8987 13175
rect 9689 13141 9723 13175
rect 9873 13141 9907 13175
rect 9965 13141 9999 13175
rect 10425 13141 10459 13175
rect 11345 13141 11379 13175
rect 12909 13141 12943 13175
rect 13185 13141 13219 13175
rect 6377 12937 6411 12971
rect 1593 12869 1627 12903
rect 4261 12869 4295 12903
rect 4353 12869 4387 12903
rect 6837 12869 6871 12903
rect 7297 12869 7331 12903
rect 7665 12869 7699 12903
rect 8585 12869 8619 12903
rect 10701 12869 10735 12903
rect 13093 12869 13127 12903
rect 13369 12869 13403 12903
rect 1685 12801 1719 12835
rect 1869 12801 1903 12835
rect 2053 12801 2087 12835
rect 2237 12801 2271 12835
rect 3617 12801 3651 12835
rect 4117 12801 4151 12835
rect 4537 12801 4571 12835
rect 4629 12801 4663 12835
rect 5733 12801 5767 12835
rect 6561 12801 6595 12835
rect 6745 12801 6779 12835
rect 6934 12801 6968 12835
rect 7481 12801 7515 12835
rect 7849 12801 7883 12835
rect 8769 12801 8803 12835
rect 8861 12801 8895 12835
rect 9045 12801 9079 12835
rect 9965 12801 9999 12835
rect 10793 12801 10827 12835
rect 10977 12801 11011 12835
rect 11529 12801 11563 12835
rect 12449 12801 12483 12835
rect 10609 12733 10643 12767
rect 3525 12665 3559 12699
rect 3985 12665 4019 12699
rect 5917 12665 5951 12699
rect 13185 12665 13219 12699
rect 1409 12597 1443 12631
rect 7113 12597 7147 12631
rect 11161 12597 11195 12631
rect 2421 12393 2455 12427
rect 3985 12393 4019 12427
rect 7665 12393 7699 12427
rect 8033 12393 8067 12427
rect 9045 12393 9079 12427
rect 6009 12325 6043 12359
rect 7297 12325 7331 12359
rect 5917 12257 5951 12291
rect 6469 12257 6503 12291
rect 8476 12257 8510 12291
rect 9413 12257 9447 12291
rect 9965 12257 9999 12291
rect 10592 12257 10626 12291
rect 10793 12257 10827 12291
rect 1409 12189 1443 12223
rect 2053 12189 2087 12223
rect 2605 12189 2639 12223
rect 2697 12189 2731 12223
rect 3433 12189 3467 12223
rect 3617 12189 3651 12223
rect 4353 12189 4387 12223
rect 4813 12189 4847 12223
rect 4905 12189 4939 12223
rect 5549 12189 5583 12223
rect 5825 12189 5859 12223
rect 6745 12189 6779 12223
rect 6929 12189 6963 12223
rect 7118 12189 7152 12223
rect 7941 12189 7975 12223
rect 8769 12189 8803 12223
rect 9321 12189 9355 12223
rect 9873 12189 9907 12223
rect 10333 12189 10367 12223
rect 10885 12189 10919 12223
rect 10977 12189 11011 12223
rect 11621 12189 11655 12223
rect 11897 12189 11931 12223
rect 11989 12189 12023 12223
rect 13001 12189 13035 12223
rect 2329 12121 2363 12155
rect 3893 12121 3927 12155
rect 4537 12121 4571 12155
rect 7021 12121 7055 12155
rect 7481 12121 7515 12155
rect 8217 12121 8251 12155
rect 9137 12121 9171 12155
rect 10149 12121 10183 12155
rect 13553 12121 13587 12155
rect 6561 12053 6595 12087
rect 7665 12053 7699 12087
rect 8585 12053 8619 12087
rect 8677 12053 8711 12087
rect 10701 12053 10735 12087
rect 1777 11849 1811 11883
rect 3433 11849 3467 11883
rect 6469 11849 6503 11883
rect 6837 11849 6871 11883
rect 8401 11849 8435 11883
rect 8953 11849 8987 11883
rect 9229 11849 9263 11883
rect 10517 11849 10551 11883
rect 12081 11849 12115 11883
rect 13461 11849 13495 11883
rect 1501 11781 1535 11815
rect 2605 11781 2639 11815
rect 3801 11781 3835 11815
rect 5549 11781 5583 11815
rect 7481 11781 7515 11815
rect 8033 11781 8067 11815
rect 8585 11781 8619 11815
rect 8769 11781 8803 11815
rect 10333 11781 10367 11815
rect 10885 11781 10919 11815
rect 12725 11781 12759 11815
rect 13369 11781 13403 11815
rect 2513 11713 2547 11747
rect 2789 11713 2823 11747
rect 5181 11713 5215 11747
rect 5791 11713 5825 11747
rect 5917 11713 5951 11747
rect 6009 11713 6043 11747
rect 6193 11713 6227 11747
rect 7021 11713 7055 11747
rect 7113 11713 7147 11747
rect 7389 11713 7423 11747
rect 7665 11713 7699 11747
rect 7849 11713 7883 11747
rect 8217 11713 8251 11747
rect 8493 11713 8527 11747
rect 9505 11713 9539 11747
rect 9688 11713 9722 11747
rect 9873 11713 9907 11747
rect 10057 11713 10091 11747
rect 11069 11713 11103 11747
rect 11253 11713 11287 11747
rect 11529 11713 11563 11747
rect 11713 11713 11747 11747
rect 12633 11713 12667 11747
rect 13277 11713 13311 11747
rect 1685 11645 1719 11679
rect 1869 11645 1903 11679
rect 2421 11645 2455 11679
rect 2973 11645 3007 11679
rect 4261 11645 4295 11679
rect 4813 11645 4847 11679
rect 5365 11645 5399 11679
rect 9781 11645 9815 11679
rect 10241 11645 10275 11679
rect 12173 11645 12207 11679
rect 12817 11645 12851 11679
rect 1961 11577 1995 11611
rect 4077 11577 4111 11611
rect 4353 11577 4387 11611
rect 6653 11577 6687 11611
rect 3157 11509 3191 11543
rect 3525 11509 3559 11543
rect 3893 11509 3927 11543
rect 4905 11509 4939 11543
rect 7297 11509 7331 11543
rect 8769 11509 8803 11543
rect 9413 11509 9447 11543
rect 10517 11509 10551 11543
rect 10701 11509 10735 11543
rect 11805 11509 11839 11543
rect 8677 11305 8711 11339
rect 8953 11305 8987 11339
rect 9137 11305 9171 11339
rect 9413 11305 9447 11339
rect 10149 11305 10183 11339
rect 10885 11305 10919 11339
rect 11989 11305 12023 11339
rect 2881 11237 2915 11271
rect 5089 11237 5123 11271
rect 5641 11237 5675 11271
rect 7665 11237 7699 11271
rect 8217 11237 8251 11271
rect 9873 11237 9907 11271
rect 5897 11169 5931 11203
rect 6193 11169 6227 11203
rect 8125 11169 8159 11203
rect 9321 11169 9355 11203
rect 11069 11169 11103 11203
rect 11161 11169 11195 11203
rect 13553 11169 13587 11203
rect 1409 11101 1443 11135
rect 2421 11101 2455 11135
rect 3065 11101 3099 11135
rect 3801 11101 3835 11135
rect 4721 11101 4755 11135
rect 5641 11101 5675 11135
rect 6560 11079 6594 11113
rect 6652 11079 6686 11113
rect 6763 11101 6797 11135
rect 6929 11101 6963 11135
rect 7021 11101 7055 11135
rect 7205 11101 7239 11135
rect 7298 11079 7332 11113
rect 7423 11101 7457 11135
rect 8401 11101 8435 11135
rect 8493 11101 8527 11135
rect 9597 11101 9631 11135
rect 9689 11101 9723 11135
rect 10333 11101 10367 11135
rect 10609 11101 10643 11135
rect 10706 11101 10740 11135
rect 11391 11101 11425 11135
rect 11805 11101 11839 11135
rect 12081 11101 12115 11135
rect 13001 11101 13035 11135
rect 13277 11101 13311 11135
rect 3525 11033 3559 11067
rect 3617 11033 3651 11067
rect 6101 11033 6135 11067
rect 6285 11033 6319 11067
rect 10517 11033 10551 11067
rect 11621 11033 11655 11067
rect 12817 11033 12851 11067
rect 6009 10965 6043 10999
rect 7849 10965 7883 10999
rect 11253 10965 11287 10999
rect 13185 10965 13219 10999
rect 2421 10761 2455 10795
rect 3709 10761 3743 10795
rect 5365 10761 5399 10795
rect 5825 10761 5859 10795
rect 6009 10761 6043 10795
rect 8677 10761 8711 10795
rect 9413 10761 9447 10795
rect 10425 10761 10459 10795
rect 11604 10761 11638 10795
rect 2881 10693 2915 10727
rect 3341 10693 3375 10727
rect 3801 10693 3835 10727
rect 3985 10693 4019 10727
rect 4353 10693 4387 10727
rect 6193 10693 6227 10727
rect 7021 10693 7055 10727
rect 7389 10693 7423 10727
rect 7941 10693 7975 10727
rect 8033 10693 8067 10727
rect 9965 10693 9999 10727
rect 10793 10693 10827 10727
rect 11253 10693 11287 10727
rect 13461 10693 13495 10727
rect 1633 10625 1667 10659
rect 1777 10625 1811 10659
rect 1869 10625 1903 10659
rect 2053 10625 2087 10659
rect 2513 10625 2547 10659
rect 2973 10625 3007 10659
rect 3157 10625 3191 10659
rect 4077 10625 4111 10659
rect 4997 10625 5031 10659
rect 5273 10625 5307 10659
rect 5549 10625 5583 10659
rect 6929 10625 6963 10659
rect 7205 10625 7239 10659
rect 7844 10625 7878 10659
rect 8217 10625 8251 10659
rect 8309 10625 8343 10659
rect 8401 10625 8435 10659
rect 9137 10625 9171 10659
rect 9321 10625 9355 10659
rect 9597 10625 9631 10659
rect 9781 10625 9815 10659
rect 10057 10625 10091 10659
rect 10609 10625 10643 10659
rect 11345 10625 11379 10659
rect 11800 10625 11834 10659
rect 11897 10625 11931 10659
rect 11989 10625 12023 10659
rect 12173 10625 12207 10659
rect 12725 10625 12759 10659
rect 8953 10557 8987 10591
rect 10149 10557 10183 10591
rect 12265 10557 12299 10591
rect 12817 10557 12851 10591
rect 12909 10557 12943 10591
rect 6653 10489 6687 10523
rect 13369 10489 13403 10523
rect 1501 10421 1535 10455
rect 2145 10421 2179 10455
rect 2789 10421 2823 10455
rect 5181 10421 5215 10455
rect 6009 10421 6043 10455
rect 6469 10421 6503 10455
rect 7665 10421 7699 10455
rect 8493 10421 8527 10455
rect 10057 10421 10091 10455
rect 10885 10421 10919 10455
rect 1409 10217 1443 10251
rect 1685 10217 1719 10251
rect 7113 10217 7147 10251
rect 8677 10217 8711 10251
rect 9413 10217 9447 10251
rect 8217 10149 8251 10183
rect 9873 10149 9907 10183
rect 13369 10149 13403 10183
rect 1777 10081 1811 10115
rect 3893 10081 3927 10115
rect 4629 10081 4663 10115
rect 4813 10081 4847 10115
rect 6745 10081 6779 10115
rect 10221 10081 10255 10115
rect 10517 10081 10551 10115
rect 10977 10081 11011 10115
rect 2329 10013 2363 10047
rect 2421 10013 2455 10047
rect 2881 10013 2915 10047
rect 3341 10013 3375 10047
rect 3525 10013 3559 10047
rect 4077 10013 4111 10047
rect 5365 10013 5399 10047
rect 5549 10013 5583 10047
rect 5733 10013 5767 10047
rect 5825 10013 5859 10047
rect 6245 10013 6279 10047
rect 6653 10013 6687 10047
rect 6837 10013 6871 10047
rect 6929 10013 6963 10047
rect 7389 10013 7423 10047
rect 7573 10013 7607 10047
rect 7757 10013 7791 10047
rect 7850 9991 7884 10025
rect 7975 10013 8009 10047
rect 8585 10013 8619 10047
rect 8769 10013 8803 10047
rect 9229 10013 9263 10047
rect 9413 10013 9447 10047
rect 9505 10013 9539 10047
rect 10609 10013 10643 10047
rect 10793 10013 10827 10047
rect 11069 10013 11103 10047
rect 11345 10013 11379 10047
rect 11713 10013 11747 10047
rect 11897 10013 11931 10047
rect 12817 10013 12851 10047
rect 2237 9945 2271 9979
rect 2973 9945 3007 9979
rect 3069 9945 3103 9979
rect 3801 9945 3835 9979
rect 4537 9945 4571 9979
rect 4997 9945 5031 9979
rect 5181 9945 5215 9979
rect 6009 9945 6043 9979
rect 6101 9945 6135 9979
rect 9965 9945 9999 9979
rect 10309 9945 10343 9979
rect 10425 9945 10459 9979
rect 11437 9945 11471 9979
rect 3157 9877 3191 9911
rect 6394 9877 6428 9911
rect 9045 9877 9079 9911
rect 9597 9877 9631 9911
rect 11621 9877 11655 9911
rect 7205 9673 7239 9707
rect 8217 9673 8251 9707
rect 8861 9673 8895 9707
rect 9137 9673 9171 9707
rect 10793 9673 10827 9707
rect 1409 9605 1443 9639
rect 3525 9605 3559 9639
rect 5457 9605 5491 9639
rect 7941 9605 7975 9639
rect 10701 9605 10735 9639
rect 11621 9605 11655 9639
rect 12817 9605 12851 9639
rect 13277 9605 13311 9639
rect 1593 9537 1627 9571
rect 3065 9537 3099 9571
rect 3341 9537 3375 9571
rect 3709 9537 3743 9571
rect 5181 9537 5215 9571
rect 6193 9537 6227 9571
rect 6648 9537 6682 9571
rect 6748 9537 6782 9571
rect 6883 9537 6917 9571
rect 7021 9537 7055 9571
rect 7573 9537 7607 9571
rect 8392 9549 8426 9583
rect 8492 9537 8526 9571
rect 8677 9537 8711 9571
rect 8764 9537 8798 9571
rect 9505 9537 9539 9571
rect 9781 9537 9815 9571
rect 10057 9537 10091 9571
rect 10333 9537 10367 9571
rect 10517 9537 10551 9571
rect 11161 9537 11195 9571
rect 11345 9537 11379 9571
rect 11529 9537 11563 9571
rect 11897 9537 11931 9571
rect 12173 9537 12207 9571
rect 13093 9537 13127 9571
rect 5365 9469 5399 9503
rect 5917 9469 5951 9503
rect 7757 9469 7791 9503
rect 9413 9469 9447 9503
rect 10149 9469 10183 9503
rect 11713 9469 11747 9503
rect 2881 9401 2915 9435
rect 4997 9401 5031 9435
rect 6009 9401 6043 9435
rect 7573 9401 7607 9435
rect 11253 9401 11287 9435
rect 13461 9401 13495 9435
rect 6469 9333 6503 9367
rect 9413 9333 9447 9367
rect 9689 9333 9723 9367
rect 1501 9129 1535 9163
rect 3341 9129 3375 9163
rect 6653 9129 6687 9163
rect 7297 9129 7331 9163
rect 8217 9129 8251 9163
rect 9137 9129 9171 9163
rect 9689 9129 9723 9163
rect 10885 9129 10919 9163
rect 11161 9129 11195 9163
rect 12081 9129 12115 9163
rect 11805 9061 11839 9095
rect 8033 8993 8067 9027
rect 9045 8993 9079 9027
rect 10333 8993 10367 9027
rect 12633 8993 12667 9027
rect 1961 8925 1995 8959
rect 2329 8925 2363 8959
rect 2973 8925 3007 8959
rect 3249 8925 3283 8959
rect 3525 8925 3559 8959
rect 3893 8925 3927 8959
rect 4077 8925 4111 8959
rect 4537 8925 4571 8959
rect 4997 8925 5031 8959
rect 5641 8925 5675 8959
rect 6101 8925 6135 8959
rect 6285 8925 6319 8959
rect 6561 8925 6595 8959
rect 6653 8925 6687 8959
rect 6929 8925 6963 8959
rect 7113 8925 7147 8959
rect 7849 8925 7883 8959
rect 8125 8925 8159 8959
rect 9229 8925 9263 8959
rect 9781 8925 9815 8959
rect 9965 8925 9999 8959
rect 10149 8925 10183 8959
rect 10701 8925 10735 8959
rect 10977 8925 11011 8959
rect 11253 8925 11287 8959
rect 11626 8925 11660 8959
rect 12265 8925 12299 8959
rect 13461 8925 13495 8959
rect 3801 8857 3835 8891
rect 4261 8857 4295 8891
rect 4721 8857 4755 8891
rect 6837 8857 6871 8891
rect 7665 8857 7699 8891
rect 8953 8857 8987 8891
rect 9873 8857 9907 8891
rect 10517 8857 10551 8891
rect 11437 8857 11471 8891
rect 11529 8857 11563 8891
rect 12449 8857 12483 8891
rect 12541 8857 12575 8891
rect 13093 8857 13127 8891
rect 13185 8857 13219 8891
rect 1777 8789 1811 8823
rect 2145 8789 2179 8823
rect 4629 8789 4663 8823
rect 5733 8789 5767 8823
rect 6193 8789 6227 8823
rect 9413 8789 9447 8823
rect 13277 8789 13311 8823
rect 9505 8585 9539 8619
rect 11253 8585 11287 8619
rect 12265 8585 12299 8619
rect 5181 8517 5215 8551
rect 5457 8517 5491 8551
rect 6377 8517 6411 8551
rect 11529 8517 11563 8551
rect 11897 8517 11931 8551
rect 13093 8517 13127 8551
rect 13369 8517 13403 8551
rect 1501 8449 1535 8483
rect 3617 8449 3651 8483
rect 5089 8449 5123 8483
rect 5273 8449 5307 8483
rect 6193 8449 6227 8483
rect 6561 8449 6595 8483
rect 6745 8449 6779 8483
rect 7021 8449 7055 8483
rect 7389 8449 7423 8483
rect 8217 8449 8251 8483
rect 9137 8449 9171 8483
rect 9393 8449 9427 8483
rect 10149 8449 10183 8483
rect 11713 8449 11747 8483
rect 12081 8449 12115 8483
rect 12357 8449 12391 8483
rect 13277 8449 13311 8483
rect 6929 8381 6963 8415
rect 8033 8381 8067 8415
rect 8861 8381 8895 8415
rect 9597 8381 9631 8415
rect 9689 8381 9723 8415
rect 10241 8381 10275 8415
rect 10885 8381 10919 8415
rect 11161 8381 11195 8415
rect 2973 8313 3007 8347
rect 13461 8313 13495 8347
rect 3433 8245 3467 8279
rect 7297 8245 7331 8279
rect 8953 8245 8987 8279
rect 1501 8041 1535 8075
rect 5917 8041 5951 8075
rect 7849 8041 7883 8075
rect 13461 8041 13495 8075
rect 5181 7973 5215 8007
rect 10241 7973 10275 8007
rect 4169 7905 4203 7939
rect 4721 7905 4755 7939
rect 5641 7905 5675 7939
rect 7021 7905 7055 7939
rect 7941 7905 7975 7939
rect 8217 7905 8251 7939
rect 8769 7905 8803 7939
rect 9597 7905 9631 7939
rect 1777 7837 1811 7871
rect 2881 7837 2915 7871
rect 3065 7837 3099 7871
rect 3893 7837 3927 7871
rect 3985 7837 4019 7871
rect 4813 7837 4847 7871
rect 6745 7837 6779 7871
rect 7573 7837 7607 7871
rect 7665 7837 7699 7871
rect 8125 7837 8159 7871
rect 8584 7837 8618 7871
rect 9505 7837 9539 7871
rect 10483 7837 10517 7871
rect 10609 7837 10643 7871
rect 10701 7837 10735 7871
rect 10885 7837 10919 7871
rect 11345 7837 11379 7871
rect 11713 7837 11747 7871
rect 11805 7837 11839 7871
rect 13277 7837 13311 7871
rect 3157 7769 3191 7803
rect 3341 7769 3375 7803
rect 3525 7769 3559 7803
rect 4629 7769 4663 7803
rect 5089 7769 5123 7803
rect 5825 7769 5859 7803
rect 11529 7769 11563 7803
rect 13369 7769 13403 7803
rect 2789 7701 2823 7735
rect 4997 7701 5031 7735
rect 6101 7701 6135 7735
rect 7389 7701 7423 7735
rect 10149 7701 10183 7735
rect 2421 7497 2455 7531
rect 6469 7497 6503 7531
rect 7481 7497 7515 7531
rect 9689 7497 9723 7531
rect 12817 7497 12851 7531
rect 2329 7429 2363 7463
rect 6929 7429 6963 7463
rect 12357 7429 12391 7463
rect 1685 7361 1719 7395
rect 1777 7361 1811 7395
rect 4721 7361 4755 7395
rect 4905 7361 4939 7395
rect 5457 7361 5491 7395
rect 5641 7361 5675 7395
rect 5825 7361 5859 7395
rect 6009 7361 6043 7395
rect 6653 7361 6687 7395
rect 6837 7361 6871 7395
rect 7113 7361 7147 7395
rect 7369 7361 7403 7395
rect 7665 7361 7699 7395
rect 9229 7361 9263 7395
rect 9413 7361 9447 7395
rect 9965 7361 9999 7395
rect 10241 7361 10275 7395
rect 11805 7361 11839 7395
rect 12265 7361 12299 7395
rect 2605 7293 2639 7327
rect 2789 7293 2823 7327
rect 3065 7293 3099 7327
rect 7573 7293 7607 7327
rect 8033 7293 8067 7327
rect 8861 7293 8895 7327
rect 9781 7293 9815 7327
rect 9873 7293 9907 7327
rect 12449 7293 12483 7327
rect 12817 7293 12851 7327
rect 12909 7293 12943 7327
rect 4813 7225 4847 7259
rect 5641 7225 5675 7259
rect 1501 7157 1535 7191
rect 1961 7157 1995 7191
rect 4537 7157 4571 7191
rect 5273 7157 5307 7191
rect 1764 6953 1798 6987
rect 3249 6953 3283 6987
rect 4261 6953 4295 6987
rect 5904 6953 5938 6987
rect 13277 6885 13311 6919
rect 1501 6817 1535 6851
rect 4537 6817 4571 6851
rect 5641 6817 5675 6851
rect 7389 6817 7423 6851
rect 7757 6817 7791 6851
rect 8769 6817 8803 6851
rect 9321 6817 9355 6851
rect 11805 6817 11839 6851
rect 3433 6749 3467 6783
rect 3893 6749 3927 6783
rect 4169 6749 4203 6783
rect 5273 6749 5307 6783
rect 7941 6749 7975 6783
rect 8125 6749 8159 6783
rect 8217 6749 8251 6783
rect 8401 6749 8435 6783
rect 9505 6749 9539 6783
rect 9597 6749 9631 6783
rect 10057 6749 10091 6783
rect 11989 6749 12023 6783
rect 13461 6749 13495 6783
rect 8677 6681 8711 6715
rect 10333 6681 10367 6715
rect 4077 6613 4111 6647
rect 9965 6613 9999 6647
rect 3525 6409 3559 6443
rect 3893 6409 3927 6443
rect 6101 6409 6135 6443
rect 6561 6409 6595 6443
rect 10149 6409 10183 6443
rect 6929 6341 6963 6375
rect 7113 6341 7147 6375
rect 11161 6341 11195 6375
rect 11989 6341 12023 6375
rect 13185 6341 13219 6375
rect 1777 6273 1811 6307
rect 1943 6273 1977 6307
rect 2054 6295 2088 6329
rect 2146 6263 2180 6297
rect 2513 6273 2547 6307
rect 2697 6273 2731 6307
rect 3249 6273 3283 6307
rect 3433 6273 3467 6307
rect 4353 6273 4387 6307
rect 6515 6273 6549 6307
rect 6653 6273 6687 6307
rect 7941 6273 7975 6307
rect 8677 6273 8711 6307
rect 8861 6273 8895 6307
rect 10701 6273 10735 6307
rect 10793 6273 10827 6307
rect 10977 6273 11011 6307
rect 11713 6273 11747 6307
rect 11805 6273 11839 6307
rect 12081 6273 12115 6307
rect 12265 6273 12299 6307
rect 12725 6273 12759 6307
rect 3985 6205 4019 6239
rect 4077 6205 4111 6239
rect 4629 6205 4663 6239
rect 7757 6205 7791 6239
rect 9689 6205 9723 6239
rect 10241 6205 10275 6239
rect 10333 6205 10367 6239
rect 10881 6205 10915 6239
rect 13277 6205 13311 6239
rect 2421 6137 2455 6171
rect 3157 6137 3191 6171
rect 11621 6137 11655 6171
rect 1409 6069 1443 6103
rect 1593 6069 1627 6103
rect 2881 6069 2915 6103
rect 9781 6069 9815 6103
rect 12449 6069 12483 6103
rect 13369 6069 13403 6103
rect 5365 5865 5399 5899
rect 8033 5865 8067 5899
rect 10149 5865 10183 5899
rect 13277 5865 13311 5899
rect 2329 5797 2363 5831
rect 3801 5797 3835 5831
rect 8493 5797 8527 5831
rect 2145 5729 2179 5763
rect 5549 5729 5583 5763
rect 5733 5729 5767 5763
rect 6009 5729 6043 5763
rect 10333 5729 10367 5763
rect 10609 5729 10643 5763
rect 1501 5661 1535 5695
rect 1593 5661 1627 5695
rect 1777 5661 1811 5695
rect 2421 5661 2455 5695
rect 2605 5661 2639 5695
rect 2973 5661 3007 5695
rect 3433 5661 3467 5695
rect 3525 5661 3559 5695
rect 4721 5661 4755 5695
rect 4905 5661 4939 5695
rect 5825 5661 5859 5695
rect 6193 5661 6227 5695
rect 6285 5661 6319 5695
rect 8585 5661 8619 5695
rect 8769 5661 8803 5695
rect 8953 5661 8987 5695
rect 9045 5661 9079 5695
rect 9321 5661 9355 5695
rect 9719 5661 9753 5695
rect 10241 5661 10275 5695
rect 12357 5661 12391 5695
rect 12541 5661 12575 5695
rect 2789 5593 2823 5627
rect 3249 5593 3283 5627
rect 3985 5593 4019 5627
rect 4353 5593 4387 5627
rect 4537 5593 4571 5627
rect 8125 5593 8159 5627
rect 8309 5593 8343 5627
rect 12265 5593 12299 5627
rect 1961 5525 1995 5559
rect 3157 5525 3191 5559
rect 4077 5525 4111 5559
rect 4169 5525 4203 5559
rect 9597 5525 9631 5559
rect 9781 5525 9815 5559
rect 12081 5525 12115 5559
rect 12725 5525 12759 5559
rect 13185 5525 13219 5559
rect 8401 5321 8435 5355
rect 12182 5321 12216 5355
rect 1409 5253 1443 5287
rect 3525 5253 3559 5287
rect 3617 5253 3651 5287
rect 4445 5253 4479 5287
rect 4629 5253 4663 5287
rect 4997 5253 5031 5287
rect 5181 5253 5215 5287
rect 8861 5253 8895 5287
rect 11713 5253 11747 5287
rect 13277 5253 13311 5287
rect 1501 5185 1535 5219
rect 1685 5185 1719 5219
rect 2145 5185 2179 5219
rect 2329 5185 2363 5219
rect 2421 5185 2455 5219
rect 2789 5185 2823 5219
rect 3341 5185 3375 5219
rect 3709 5185 3743 5219
rect 4077 5185 4111 5219
rect 4353 5185 4387 5219
rect 5365 5185 5399 5219
rect 5641 5185 5675 5219
rect 6009 5185 6043 5219
rect 6377 5185 6411 5219
rect 6561 5185 6595 5219
rect 7113 5185 7147 5219
rect 7573 5185 7607 5219
rect 8953 5185 8987 5219
rect 9137 5185 9171 5219
rect 11805 5185 11839 5219
rect 12633 5185 12667 5219
rect 13553 5185 13587 5219
rect 2973 5117 3007 5151
rect 4813 5117 4847 5151
rect 6745 5117 6779 5151
rect 7941 5117 7975 5151
rect 8493 5117 8527 5151
rect 8585 5117 8619 5151
rect 9505 5117 9539 5151
rect 9781 5117 9815 5151
rect 2513 5049 2547 5083
rect 11253 5049 11287 5083
rect 1961 4981 1995 5015
rect 2329 4981 2363 5015
rect 3157 4981 3191 5015
rect 3801 4981 3835 5015
rect 6009 4981 6043 5015
rect 8033 4981 8067 5015
rect 12173 4981 12207 5015
rect 12357 4981 12391 5015
rect 1409 4777 1443 4811
rect 8677 4777 8711 4811
rect 9505 4777 9539 4811
rect 11989 4777 12023 4811
rect 13185 4709 13219 4743
rect 2329 4641 2363 4675
rect 3433 4641 3467 4675
rect 5641 4641 5675 4675
rect 6929 4641 6963 4675
rect 7205 4641 7239 4675
rect 10241 4641 10275 4675
rect 10517 4641 10551 4675
rect 1593 4573 1627 4607
rect 1777 4573 1811 4607
rect 2145 4573 2179 4607
rect 2421 4573 2455 4607
rect 3137 4573 3171 4607
rect 3341 4573 3375 4607
rect 5733 4573 5767 4607
rect 5917 4573 5951 4607
rect 6009 4573 6043 4607
rect 6135 4573 6169 4607
rect 6561 4573 6595 4607
rect 6745 4573 6779 4607
rect 9045 4573 9079 4607
rect 9137 4573 9171 4607
rect 9505 4573 9539 4607
rect 12725 4573 12759 4607
rect 13553 4573 13587 4607
rect 2697 4505 2731 4539
rect 2881 4505 2915 4539
rect 5365 4505 5399 4539
rect 6377 4505 6411 4539
rect 13277 4505 13311 4539
rect 2237 4437 2271 4471
rect 3249 4437 3283 4471
rect 3525 4437 3559 4471
rect 3893 4437 3927 4471
rect 6745 4437 6779 4471
rect 9689 4437 9723 4471
rect 13369 4437 13403 4471
rect 3341 4233 3375 4267
rect 4629 4233 4663 4267
rect 5089 4233 5123 4267
rect 5549 4233 5583 4267
rect 6469 4233 6503 4267
rect 9689 4233 9723 4267
rect 11161 4233 11195 4267
rect 11253 4233 11287 4267
rect 11621 4233 11655 4267
rect 6193 4165 6227 4199
rect 12541 4165 12575 4199
rect 1869 4097 1903 4131
rect 2053 4097 2087 4131
rect 2237 4097 2271 4131
rect 2329 4097 2363 4131
rect 2697 4097 2731 4131
rect 2881 4097 2915 4131
rect 3341 4097 3375 4131
rect 3525 4097 3559 4131
rect 3985 4097 4019 4131
rect 4077 4097 4111 4131
rect 4261 4097 4295 4131
rect 4537 4097 4571 4131
rect 4721 4097 4755 4131
rect 5181 4097 5215 4131
rect 5825 4097 5859 4131
rect 6101 4097 6135 4131
rect 8217 4097 8251 4131
rect 8769 4097 8803 4131
rect 9045 4097 9079 4131
rect 9505 4097 9539 4131
rect 9597 4097 9631 4131
rect 9965 4097 9999 4131
rect 10057 4097 10091 4131
rect 10793 4097 10827 4131
rect 10885 4097 10919 4131
rect 11621 4097 11655 4131
rect 11805 4097 11839 4131
rect 12081 4097 12115 4131
rect 12265 4097 12299 4131
rect 12725 4097 12759 4131
rect 12909 4097 12943 4131
rect 13001 4097 13035 4131
rect 1777 4029 1811 4063
rect 4905 4029 4939 4063
rect 7941 4029 7975 4063
rect 10241 4029 10275 4063
rect 10609 4029 10643 4063
rect 11989 4029 12023 4063
rect 13093 4029 13127 4063
rect 1501 3961 1535 3995
rect 2145 3961 2179 3995
rect 3065 3961 3099 3995
rect 3801 3961 3835 3995
rect 5733 3961 5767 3995
rect 8585 3961 8619 3995
rect 9321 3961 9355 3995
rect 9873 3961 9907 3995
rect 1869 3893 1903 3927
rect 2513 3893 2547 3927
rect 8953 3893 8987 3927
rect 10425 3893 10459 3927
rect 13369 3893 13403 3927
rect 1501 3689 1535 3723
rect 2237 3689 2271 3723
rect 6469 3689 6503 3723
rect 6653 3689 6687 3723
rect 9597 3689 9631 3723
rect 9781 3689 9815 3723
rect 11805 3689 11839 3723
rect 6009 3621 6043 3655
rect 1869 3553 1903 3587
rect 2605 3553 2639 3587
rect 3433 3553 3467 3587
rect 3801 3553 3835 3587
rect 4169 3553 4203 3587
rect 5549 3553 5583 3587
rect 6377 3553 6411 3587
rect 8769 3553 8803 3587
rect 10057 3553 10091 3587
rect 10333 3553 10367 3587
rect 12909 3553 12943 3587
rect 13093 3553 13127 3587
rect 1501 3485 1535 3519
rect 1593 3485 1627 3519
rect 2237 3485 2271 3519
rect 3341 3485 3375 3519
rect 4353 3485 4387 3519
rect 4445 3485 4479 3519
rect 4629 3485 4663 3519
rect 4721 3485 4755 3519
rect 5181 3485 5215 3519
rect 5365 3485 5399 3519
rect 5733 3485 5767 3519
rect 5917 3485 5951 3519
rect 9045 3485 9079 3519
rect 9229 3485 9263 3519
rect 12081 3485 12115 3519
rect 12265 3485 12299 3519
rect 12449 3485 12483 3519
rect 12633 3485 12667 3519
rect 4997 3417 5031 3451
rect 8493 3417 8527 3451
rect 9965 3417 9999 3451
rect 11989 3417 12023 3451
rect 12817 3417 12851 3451
rect 2053 3349 2087 3383
rect 4813 3349 4847 3383
rect 7021 3349 7055 3383
rect 9045 3349 9079 3383
rect 9781 3349 9815 3383
rect 1593 3145 1627 3179
rect 2329 3145 2363 3179
rect 5181 3145 5215 3179
rect 7481 3145 7515 3179
rect 10793 3145 10827 3179
rect 11345 3145 11379 3179
rect 2789 3077 2823 3111
rect 3341 3077 3375 3111
rect 3709 3077 3743 3111
rect 5733 3077 5767 3111
rect 5917 3077 5951 3111
rect 8033 3077 8067 3111
rect 1777 3009 1811 3043
rect 1869 3009 1903 3043
rect 2513 3009 2547 3043
rect 2881 3009 2915 3043
rect 3157 3009 3191 3043
rect 3525 3009 3559 3043
rect 3801 3009 3835 3043
rect 4721 3009 4755 3043
rect 5365 3009 5399 3043
rect 5549 3009 5583 3043
rect 6561 3009 6595 3043
rect 7021 3009 7055 3043
rect 7205 3009 7239 3043
rect 7665 3009 7699 3043
rect 7849 3009 7883 3043
rect 8309 3009 8343 3043
rect 10701 3009 10735 3043
rect 11529 3009 11563 3043
rect 11805 3009 11839 3043
rect 12909 3009 12943 3043
rect 13093 3009 13127 3043
rect 2145 2941 2179 2975
rect 2697 2941 2731 2975
rect 3893 2941 3927 2975
rect 4629 2941 4663 2975
rect 6377 2941 6411 2975
rect 6929 2941 6963 2975
rect 7573 2941 7607 2975
rect 8585 2941 8619 2975
rect 10057 2941 10091 2975
rect 10977 2941 11011 2975
rect 12081 2941 12115 2975
rect 2053 2873 2087 2907
rect 6837 2873 6871 2907
rect 11805 2873 11839 2907
rect 5917 2805 5951 2839
rect 6101 2805 6135 2839
rect 10333 2805 10367 2839
rect 2697 2601 2731 2635
rect 4169 2601 4203 2635
rect 8953 2601 8987 2635
rect 12081 2601 12115 2635
rect 9873 2533 9907 2567
rect 1961 2465 1995 2499
rect 3525 2465 3559 2499
rect 4537 2465 4571 2499
rect 5641 2465 5675 2499
rect 9597 2465 9631 2499
rect 12265 2465 12299 2499
rect 1593 2397 1627 2431
rect 1685 2397 1719 2431
rect 2145 2397 2179 2431
rect 2329 2397 2363 2431
rect 2605 2397 2639 2431
rect 2789 2397 2823 2431
rect 3341 2397 3375 2431
rect 3893 2397 3927 2431
rect 3985 2397 4019 2431
rect 5457 2397 5491 2431
rect 7573 2397 7607 2431
rect 7757 2397 7791 2431
rect 8125 2397 8159 2431
rect 9321 2397 9355 2431
rect 9965 2397 9999 2431
rect 10057 2397 10091 2431
rect 10333 2397 10367 2431
rect 13277 2397 13311 2431
rect 1869 2329 1903 2363
rect 5917 2329 5951 2363
rect 9413 2329 9447 2363
rect 10609 2329 10643 2363
rect 2881 2261 2915 2295
rect 3249 2261 3283 2295
rect 7389 2261 7423 2295
rect 8033 2261 8067 2295
rect 8309 2261 8343 2295
rect 8677 2261 8711 2295
rect 1593 2057 1627 2091
rect 1777 2057 1811 2091
rect 3617 2057 3651 2091
rect 5549 2057 5583 2091
rect 6101 2057 6135 2091
rect 6469 2057 6503 2091
rect 10333 2057 10367 2091
rect 13277 2057 13311 2091
rect 3249 1989 3283 2023
rect 8217 1989 8251 2023
rect 10517 1989 10551 2023
rect 3525 1921 3559 1955
rect 3801 1921 3835 1955
rect 5917 1921 5951 1955
rect 6101 1921 6135 1955
rect 10701 1921 10735 1955
rect 10793 1921 10827 1955
rect 11161 1921 11195 1955
rect 11253 1921 11287 1955
rect 4077 1853 4111 1887
rect 8493 1853 8527 1887
rect 8585 1853 8619 1887
rect 8861 1853 8895 1887
rect 11529 1853 11563 1887
rect 11805 1853 11839 1887
rect 11069 1785 11103 1819
rect 6745 1717 6779 1751
rect 13461 1717 13495 1751
rect 4077 1513 4111 1547
rect 8493 1513 8527 1547
rect 8677 1513 8711 1547
rect 9768 1513 9802 1547
rect 13277 1513 13311 1547
rect 8953 1445 8987 1479
rect 1409 1377 1443 1411
rect 5273 1377 5307 1411
rect 5917 1377 5951 1411
rect 7297 1377 7331 1411
rect 7757 1377 7791 1411
rect 7941 1377 7975 1411
rect 9505 1377 9539 1411
rect 11529 1377 11563 1411
rect 3157 1309 3191 1343
rect 3617 1309 3651 1343
rect 3893 1309 3927 1343
rect 4077 1309 4111 1343
rect 4261 1309 4295 1343
rect 4445 1309 4479 1343
rect 4629 1309 4663 1343
rect 5181 1309 5215 1343
rect 5549 1309 5583 1343
rect 5733 1309 5767 1343
rect 6193 1309 6227 1343
rect 6561 1309 6595 1343
rect 7021 1309 7055 1343
rect 8033 1309 8067 1343
rect 8309 1309 8343 1343
rect 9137 1309 9171 1343
rect 13461 1309 13495 1343
rect 3249 1241 3283 1275
rect 3433 1241 3467 1275
rect 9321 1241 9355 1275
rect 11805 1241 11839 1275
rect 4721 1173 4755 1207
rect 5089 1173 5123 1207
rect 6377 1173 6411 1207
rect 11253 1173 11287 1207
<< metal1 >>
rect 6638 13920 6644 13932
rect 2746 13892 6644 13920
rect 2314 13744 2320 13796
rect 2372 13784 2378 13796
rect 2746 13784 2774 13892
rect 6638 13880 6644 13892
rect 6696 13880 6702 13932
rect 11238 13852 11244 13864
rect 2372 13756 2774 13784
rect 4908 13824 11244 13852
rect 2372 13744 2378 13756
rect 1578 13676 1584 13728
rect 1636 13716 1642 13728
rect 4908 13716 4936 13824
rect 11238 13812 11244 13824
rect 11296 13812 11302 13864
rect 1636 13688 4936 13716
rect 1636 13676 1642 13688
rect 5074 13676 5080 13728
rect 5132 13716 5138 13728
rect 8110 13716 8116 13728
rect 5132 13688 8116 13716
rect 5132 13676 5138 13688
rect 8110 13676 8116 13688
rect 8168 13676 8174 13728
rect 1104 13626 13892 13648
rect 1104 13574 4214 13626
rect 4266 13574 4278 13626
rect 4330 13574 4342 13626
rect 4394 13574 4406 13626
rect 4458 13574 4470 13626
rect 4522 13574 12214 13626
rect 12266 13574 12278 13626
rect 12330 13574 12342 13626
rect 12394 13574 12406 13626
rect 12458 13574 12470 13626
rect 12522 13574 13892 13626
rect 1104 13552 13892 13574
rect 1394 13512 1400 13524
rect 1355 13484 1400 13512
rect 1394 13472 1400 13484
rect 1452 13512 1458 13524
rect 4062 13512 4068 13524
rect 1452 13484 4068 13512
rect 1452 13472 1458 13484
rect 4062 13472 4068 13484
rect 4120 13472 4126 13524
rect 4709 13515 4767 13521
rect 4709 13481 4721 13515
rect 4755 13512 4767 13515
rect 6914 13512 6920 13524
rect 4755 13484 6920 13512
rect 4755 13481 4767 13484
rect 4709 13475 4767 13481
rect 1670 13404 1676 13456
rect 1728 13444 1734 13456
rect 4724 13444 4752 13475
rect 6914 13472 6920 13484
rect 6972 13472 6978 13524
rect 8036 13484 8616 13512
rect 6365 13447 6423 13453
rect 6365 13444 6377 13447
rect 1728 13416 4752 13444
rect 5644 13416 6377 13444
rect 1728 13404 1734 13416
rect 842 13336 848 13388
rect 900 13376 906 13388
rect 2314 13376 2320 13388
rect 900 13348 2320 13376
rect 900 13336 906 13348
rect 2314 13336 2320 13348
rect 2372 13336 2378 13388
rect 2961 13379 3019 13385
rect 2961 13345 2973 13379
rect 3007 13376 3019 13379
rect 4157 13379 4215 13385
rect 4157 13376 4169 13379
rect 3007 13348 4169 13376
rect 3007 13345 3019 13348
rect 2961 13339 3019 13345
rect 4157 13345 4169 13348
rect 4203 13345 4215 13379
rect 5074 13376 5080 13388
rect 5035 13348 5080 13376
rect 4157 13339 4215 13345
rect 5074 13336 5080 13348
rect 5132 13336 5138 13388
rect 5644 13385 5672 13416
rect 6365 13413 6377 13416
rect 6411 13413 6423 13447
rect 6365 13407 6423 13413
rect 6733 13447 6791 13453
rect 6733 13413 6745 13447
rect 6779 13444 6791 13447
rect 8036 13444 8064 13484
rect 6779 13416 8064 13444
rect 6779 13413 6791 13416
rect 6733 13407 6791 13413
rect 8110 13404 8116 13456
rect 8168 13444 8174 13456
rect 8588 13444 8616 13484
rect 8662 13472 8668 13524
rect 8720 13512 8726 13524
rect 9493 13515 9551 13521
rect 9493 13512 9505 13515
rect 8720 13484 9505 13512
rect 8720 13472 8726 13484
rect 9493 13481 9505 13484
rect 9539 13481 9551 13515
rect 9493 13475 9551 13481
rect 10229 13515 10287 13521
rect 10229 13481 10241 13515
rect 10275 13512 10287 13515
rect 14366 13512 14372 13524
rect 10275 13484 14372 13512
rect 10275 13481 10287 13484
rect 10229 13475 10287 13481
rect 9030 13444 9036 13456
rect 8168 13416 8213 13444
rect 8588 13416 9036 13444
rect 8168 13404 8174 13416
rect 9030 13404 9036 13416
rect 9088 13404 9094 13456
rect 5629 13379 5687 13385
rect 5629 13345 5641 13379
rect 5675 13345 5687 13379
rect 5629 13339 5687 13345
rect 5813 13379 5871 13385
rect 5813 13345 5825 13379
rect 5859 13376 5871 13379
rect 5859 13348 7052 13376
rect 5859 13345 5871 13348
rect 5813 13339 5871 13345
rect 7024 13320 7052 13348
rect 7098 13336 7104 13388
rect 7156 13376 7162 13388
rect 8202 13376 8208 13388
rect 7156 13348 8208 13376
rect 7156 13336 7162 13348
rect 8202 13336 8208 13348
rect 8260 13336 8266 13388
rect 10244 13376 10272 13475
rect 14366 13472 14372 13484
rect 14424 13472 14430 13524
rect 10597 13447 10655 13453
rect 10597 13413 10609 13447
rect 10643 13444 10655 13447
rect 10643 13416 12434 13444
rect 10643 13413 10655 13416
rect 10597 13407 10655 13413
rect 11882 13376 11888 13388
rect 8312 13348 10272 13376
rect 11164 13348 11888 13376
rect 1578 13308 1584 13320
rect 1539 13280 1584 13308
rect 1578 13268 1584 13280
rect 1636 13268 1642 13320
rect 2222 13268 2228 13320
rect 2280 13308 2286 13320
rect 2409 13311 2467 13317
rect 2409 13308 2421 13311
rect 2280 13280 2421 13308
rect 2280 13268 2286 13280
rect 2409 13277 2421 13280
rect 2455 13277 2467 13311
rect 2409 13271 2467 13277
rect 2682 13268 2688 13320
rect 2740 13308 2746 13320
rect 3053 13311 3111 13317
rect 3053 13308 3065 13311
rect 2740 13280 3065 13308
rect 2740 13268 2746 13280
rect 3053 13277 3065 13280
rect 3099 13277 3111 13311
rect 3053 13271 3111 13277
rect 3528 13280 3740 13308
rect 2038 13240 2044 13252
rect 1999 13212 2044 13240
rect 2038 13200 2044 13212
rect 2096 13200 2102 13252
rect 2130 13200 2136 13252
rect 2188 13240 2194 13252
rect 2866 13240 2872 13252
rect 2188 13212 2233 13240
rect 2827 13212 2872 13240
rect 2188 13200 2194 13212
rect 2866 13200 2872 13212
rect 2924 13200 2930 13252
rect 3418 13200 3424 13252
rect 3476 13240 3482 13252
rect 3528 13249 3556 13280
rect 3513 13243 3571 13249
rect 3513 13240 3525 13243
rect 3476 13212 3525 13240
rect 3476 13200 3482 13212
rect 3513 13209 3525 13212
rect 3559 13209 3571 13243
rect 3513 13203 3571 13209
rect 3605 13243 3663 13249
rect 3605 13209 3617 13243
rect 3651 13209 3663 13243
rect 3712 13240 3740 13280
rect 3878 13268 3884 13320
rect 3936 13308 3942 13320
rect 3973 13311 4031 13317
rect 3973 13308 3985 13311
rect 3936 13280 3985 13308
rect 3936 13268 3942 13280
rect 3973 13277 3985 13280
rect 4019 13277 4031 13311
rect 3973 13271 4031 13277
rect 5718 13268 5724 13320
rect 5776 13308 5782 13320
rect 6086 13308 6092 13320
rect 5776 13280 6092 13308
rect 5776 13268 5782 13280
rect 6086 13268 6092 13280
rect 6144 13308 6150 13320
rect 6549 13311 6607 13317
rect 6549 13308 6561 13311
rect 6144 13280 6561 13308
rect 6144 13268 6150 13280
rect 6549 13277 6561 13280
rect 6595 13277 6607 13311
rect 6549 13271 6607 13277
rect 6638 13268 6644 13320
rect 6696 13308 6702 13320
rect 6865 13311 6923 13317
rect 6865 13308 6877 13311
rect 6696 13280 6877 13308
rect 6696 13268 6702 13280
rect 6865 13277 6877 13280
rect 6911 13277 6923 13311
rect 6865 13271 6923 13277
rect 7006 13268 7012 13320
rect 7064 13308 7070 13320
rect 7282 13308 7288 13320
rect 7064 13280 7109 13308
rect 7243 13280 7288 13308
rect 7064 13268 7070 13280
rect 7282 13268 7288 13280
rect 7340 13268 7346 13320
rect 7377 13311 7435 13317
rect 7377 13277 7389 13311
rect 7423 13308 7435 13311
rect 7742 13308 7748 13320
rect 7423 13280 7748 13308
rect 7423 13277 7435 13280
rect 7377 13271 7435 13277
rect 7742 13268 7748 13280
rect 7800 13268 7806 13320
rect 8312 13317 8340 13348
rect 8292 13311 8350 13317
rect 8292 13277 8304 13311
rect 8338 13277 8350 13311
rect 8662 13308 8668 13320
rect 8623 13280 8668 13308
rect 8292 13271 8350 13277
rect 8662 13268 8668 13280
rect 8720 13268 8726 13320
rect 8754 13268 8760 13320
rect 8812 13308 8818 13320
rect 9125 13311 9183 13317
rect 9125 13308 9137 13311
rect 8812 13280 9137 13308
rect 8812 13268 8818 13280
rect 9125 13277 9137 13280
rect 9171 13277 9183 13311
rect 9125 13271 9183 13277
rect 10594 13268 10600 13320
rect 10652 13308 10658 13320
rect 11164 13317 11192 13348
rect 11882 13336 11888 13348
rect 11940 13336 11946 13388
rect 12406 13376 12434 13416
rect 12713 13379 12771 13385
rect 12713 13376 12725 13379
rect 12406 13348 12725 13376
rect 12713 13345 12725 13348
rect 12759 13345 12771 13379
rect 12713 13339 12771 13345
rect 10873 13311 10931 13317
rect 10873 13308 10885 13311
rect 10652 13280 10885 13308
rect 10652 13268 10658 13280
rect 10873 13277 10885 13280
rect 10919 13277 10931 13311
rect 10873 13271 10931 13277
rect 11057 13311 11115 13317
rect 11057 13277 11069 13311
rect 11103 13308 11115 13311
rect 11149 13311 11207 13317
rect 11149 13308 11161 13311
rect 11103 13280 11161 13308
rect 11103 13277 11115 13280
rect 11057 13271 11115 13277
rect 11149 13277 11161 13280
rect 11195 13277 11207 13311
rect 12066 13308 12072 13320
rect 11149 13271 11207 13277
rect 11348 13280 11652 13308
rect 12027 13280 12072 13308
rect 4065 13243 4123 13249
rect 4065 13240 4077 13243
rect 3712 13212 4077 13240
rect 3605 13203 3663 13209
rect 4065 13209 4077 13212
rect 4111 13209 4123 13243
rect 4065 13203 4123 13209
rect 4985 13243 5043 13249
rect 4985 13209 4997 13243
rect 5031 13240 5043 13243
rect 5534 13240 5540 13252
rect 5031 13212 5540 13240
rect 5031 13209 5043 13212
rect 4985 13203 5043 13209
rect 3620 13172 3648 13203
rect 5534 13200 5540 13212
rect 5592 13200 5598 13252
rect 5994 13240 6000 13252
rect 5955 13212 6000 13240
rect 5994 13200 6000 13212
rect 6052 13200 6058 13252
rect 6178 13200 6184 13252
rect 6236 13240 6242 13252
rect 7098 13240 7104 13252
rect 6236 13212 7104 13240
rect 6236 13200 6242 13212
rect 7098 13200 7104 13212
rect 7156 13200 7162 13252
rect 7834 13240 7840 13252
rect 7795 13212 7840 13240
rect 7834 13200 7840 13212
rect 7892 13200 7898 13252
rect 7929 13243 7987 13249
rect 7929 13209 7941 13243
rect 7975 13209 7987 13243
rect 7929 13203 7987 13209
rect 3789 13175 3847 13181
rect 3789 13172 3801 13175
rect 3620 13144 3801 13172
rect 3789 13141 3801 13144
rect 3835 13141 3847 13175
rect 3789 13135 3847 13141
rect 4246 13132 4252 13184
rect 4304 13172 4310 13184
rect 4433 13175 4491 13181
rect 4433 13172 4445 13175
rect 4304 13144 4445 13172
rect 4304 13132 4310 13144
rect 4433 13141 4445 13144
rect 4479 13141 4491 13175
rect 4433 13135 4491 13141
rect 4893 13175 4951 13181
rect 4893 13141 4905 13175
rect 4939 13172 4951 13175
rect 5626 13172 5632 13184
rect 4939 13144 5632 13172
rect 4939 13141 4951 13144
rect 4893 13135 4951 13141
rect 5626 13132 5632 13144
rect 5684 13132 5690 13184
rect 6089 13175 6147 13181
rect 6089 13141 6101 13175
rect 6135 13172 6147 13175
rect 7650 13172 7656 13184
rect 6135 13144 7656 13172
rect 6135 13141 6147 13144
rect 6089 13135 6147 13141
rect 7650 13132 7656 13144
rect 7708 13132 7714 13184
rect 7944 13172 7972 13203
rect 8110 13200 8116 13252
rect 8168 13240 8174 13252
rect 8389 13243 8447 13249
rect 8389 13240 8401 13243
rect 8168 13212 8401 13240
rect 8168 13200 8174 13212
rect 8389 13209 8401 13212
rect 8435 13209 8447 13243
rect 8389 13203 8447 13209
rect 8478 13200 8484 13252
rect 8536 13240 8542 13252
rect 9309 13243 9367 13249
rect 9309 13240 9321 13243
rect 8536 13212 9321 13240
rect 8536 13200 8542 13212
rect 9309 13209 9321 13212
rect 9355 13209 9367 13243
rect 9309 13203 9367 13209
rect 9493 13243 9551 13249
rect 9493 13209 9505 13243
rect 9539 13240 9551 13243
rect 10042 13240 10048 13252
rect 9539 13212 10048 13240
rect 9539 13209 9551 13212
rect 9493 13203 9551 13209
rect 10042 13200 10048 13212
rect 10100 13200 10106 13252
rect 10689 13243 10747 13249
rect 10689 13209 10701 13243
rect 10735 13240 10747 13243
rect 11348 13240 11376 13280
rect 11624 13252 11652 13280
rect 12066 13268 12072 13280
rect 12124 13268 12130 13320
rect 12158 13268 12164 13320
rect 12216 13308 12222 13320
rect 12216 13280 12261 13308
rect 12216 13268 12222 13280
rect 12986 13268 12992 13320
rect 13044 13308 13050 13320
rect 13081 13311 13139 13317
rect 13081 13308 13093 13311
rect 13044 13280 13093 13308
rect 13044 13268 13050 13280
rect 13081 13277 13093 13280
rect 13127 13277 13139 13311
rect 13081 13271 13139 13277
rect 13170 13268 13176 13320
rect 13228 13308 13234 13320
rect 13449 13311 13507 13317
rect 13449 13308 13461 13311
rect 13228 13280 13461 13308
rect 13228 13268 13234 13280
rect 13449 13277 13461 13280
rect 13495 13277 13507 13311
rect 13449 13271 13507 13277
rect 10735 13212 11376 13240
rect 11517 13243 11575 13249
rect 10735 13209 10747 13212
rect 10689 13203 10747 13209
rect 11517 13209 11529 13243
rect 11563 13209 11575 13243
rect 11517 13203 11575 13209
rect 8941 13175 8999 13181
rect 8941 13172 8953 13175
rect 7944 13144 8953 13172
rect 8941 13141 8953 13144
rect 8987 13141 8999 13175
rect 9674 13172 9680 13184
rect 9635 13144 9680 13172
rect 8941 13135 8999 13141
rect 9674 13132 9680 13144
rect 9732 13132 9738 13184
rect 9858 13172 9864 13184
rect 9819 13144 9864 13172
rect 9858 13132 9864 13144
rect 9916 13132 9922 13184
rect 9950 13132 9956 13184
rect 10008 13172 10014 13184
rect 10410 13172 10416 13184
rect 10008 13144 10053 13172
rect 10371 13144 10416 13172
rect 10008 13132 10014 13144
rect 10410 13132 10416 13144
rect 10468 13132 10474 13184
rect 11333 13175 11391 13181
rect 11333 13141 11345 13175
rect 11379 13172 11391 13175
rect 11532 13172 11560 13203
rect 11606 13200 11612 13252
rect 11664 13240 11670 13252
rect 12618 13240 12624 13252
rect 11664 13212 11709 13240
rect 12579 13212 12624 13240
rect 11664 13200 11670 13212
rect 12618 13200 12624 13212
rect 12676 13200 12682 13252
rect 13354 13240 13360 13252
rect 13315 13212 13360 13240
rect 13354 13200 13360 13212
rect 13412 13200 13418 13252
rect 12894 13172 12900 13184
rect 11379 13144 11560 13172
rect 12855 13144 12900 13172
rect 11379 13141 11391 13144
rect 11333 13135 11391 13141
rect 12894 13132 12900 13144
rect 12952 13132 12958 13184
rect 13078 13132 13084 13184
rect 13136 13172 13142 13184
rect 13173 13175 13231 13181
rect 13173 13172 13185 13175
rect 13136 13144 13185 13172
rect 13136 13132 13142 13144
rect 13173 13141 13185 13144
rect 13219 13141 13231 13175
rect 13173 13135 13231 13141
rect 1104 13082 13892 13104
rect 1104 13030 8214 13082
rect 8266 13030 8278 13082
rect 8330 13030 8342 13082
rect 8394 13030 8406 13082
rect 8458 13030 8470 13082
rect 8522 13030 13892 13082
rect 1104 13008 13892 13030
rect 3142 12928 3148 12980
rect 3200 12968 3206 12980
rect 6365 12971 6423 12977
rect 6365 12968 6377 12971
rect 3200 12940 6377 12968
rect 3200 12928 3206 12940
rect 6365 12937 6377 12940
rect 6411 12968 6423 12971
rect 7098 12968 7104 12980
rect 6411 12940 7104 12968
rect 6411 12937 6423 12940
rect 6365 12931 6423 12937
rect 7098 12928 7104 12940
rect 7156 12928 7162 12980
rect 7834 12928 7840 12980
rect 7892 12968 7898 12980
rect 7892 12940 8616 12968
rect 7892 12928 7898 12940
rect 1486 12860 1492 12912
rect 1544 12900 1550 12912
rect 1581 12903 1639 12909
rect 1581 12900 1593 12903
rect 1544 12872 1593 12900
rect 1544 12860 1550 12872
rect 1581 12869 1593 12872
rect 1627 12900 1639 12903
rect 3234 12900 3240 12912
rect 1627 12872 3240 12900
rect 1627 12869 1639 12872
rect 1581 12863 1639 12869
rect 3234 12860 3240 12872
rect 3292 12860 3298 12912
rect 3694 12860 3700 12912
rect 3752 12900 3758 12912
rect 4246 12900 4252 12912
rect 3752 12872 4252 12900
rect 3752 12860 3758 12872
rect 4246 12860 4252 12872
rect 4304 12860 4310 12912
rect 4341 12903 4399 12909
rect 4341 12869 4353 12903
rect 4387 12900 4399 12903
rect 6638 12900 6644 12912
rect 4387 12872 6644 12900
rect 4387 12869 4399 12872
rect 4341 12863 4399 12869
rect 6638 12860 6644 12872
rect 6696 12860 6702 12912
rect 6825 12903 6883 12909
rect 6825 12869 6837 12903
rect 6871 12900 6883 12903
rect 7006 12900 7012 12912
rect 6871 12872 7012 12900
rect 6871 12869 6883 12872
rect 6825 12863 6883 12869
rect 7006 12860 7012 12872
rect 7064 12860 7070 12912
rect 7282 12900 7288 12912
rect 7243 12872 7288 12900
rect 7282 12860 7288 12872
rect 7340 12860 7346 12912
rect 7653 12903 7711 12909
rect 7653 12869 7665 12903
rect 7699 12900 7711 12903
rect 8478 12900 8484 12912
rect 7699 12872 8484 12900
rect 7699 12869 7711 12872
rect 7653 12863 7711 12869
rect 8478 12860 8484 12872
rect 8536 12860 8542 12912
rect 8588 12909 8616 12940
rect 9674 12928 9680 12980
rect 9732 12968 9738 12980
rect 10502 12968 10508 12980
rect 9732 12940 10508 12968
rect 9732 12928 9738 12940
rect 10502 12928 10508 12940
rect 10560 12968 10566 12980
rect 10560 12940 11008 12968
rect 10560 12928 10566 12940
rect 8573 12903 8631 12909
rect 8573 12869 8585 12903
rect 8619 12900 8631 12903
rect 9858 12900 9864 12912
rect 8619 12872 9864 12900
rect 8619 12869 8631 12872
rect 8573 12863 8631 12869
rect 9858 12860 9864 12872
rect 9916 12860 9922 12912
rect 10226 12860 10232 12912
rect 10284 12900 10290 12912
rect 10689 12903 10747 12909
rect 10689 12900 10701 12903
rect 10284 12872 10701 12900
rect 10284 12860 10290 12872
rect 10689 12869 10701 12872
rect 10735 12900 10747 12903
rect 10870 12900 10876 12912
rect 10735 12872 10876 12900
rect 10735 12869 10747 12872
rect 10689 12863 10747 12869
rect 10870 12860 10876 12872
rect 10928 12860 10934 12912
rect 1394 12792 1400 12844
rect 1452 12832 1458 12844
rect 1673 12835 1731 12841
rect 1673 12832 1685 12835
rect 1452 12804 1685 12832
rect 1452 12792 1458 12804
rect 1673 12801 1685 12804
rect 1719 12801 1731 12835
rect 1854 12832 1860 12844
rect 1815 12804 1860 12832
rect 1673 12795 1731 12801
rect 1854 12792 1860 12804
rect 1912 12792 1918 12844
rect 2041 12835 2099 12841
rect 2041 12801 2053 12835
rect 2087 12832 2099 12835
rect 2222 12832 2228 12844
rect 2087 12804 2228 12832
rect 2087 12801 2099 12804
rect 2041 12795 2099 12801
rect 2222 12792 2228 12804
rect 2280 12792 2286 12844
rect 3605 12835 3663 12841
rect 3605 12801 3617 12835
rect 3651 12832 3663 12835
rect 3878 12832 3884 12844
rect 3651 12804 3884 12832
rect 3651 12801 3663 12804
rect 3605 12795 3663 12801
rect 3878 12792 3884 12804
rect 3936 12792 3942 12844
rect 4062 12792 4068 12844
rect 4120 12841 4126 12844
rect 4120 12835 4163 12841
rect 4151 12801 4163 12835
rect 4120 12795 4163 12801
rect 4120 12792 4126 12795
rect 4430 12792 4436 12844
rect 4488 12832 4494 12844
rect 4525 12835 4583 12841
rect 4525 12832 4537 12835
rect 4488 12804 4537 12832
rect 4488 12792 4494 12804
rect 4525 12801 4537 12804
rect 4571 12801 4583 12835
rect 4525 12795 4583 12801
rect 4617 12835 4675 12841
rect 4617 12801 4629 12835
rect 4663 12832 4675 12835
rect 5718 12832 5724 12844
rect 4663 12804 5028 12832
rect 5679 12804 5724 12832
rect 4663 12801 4675 12804
rect 4617 12795 4675 12801
rect 2866 12656 2872 12708
rect 2924 12696 2930 12708
rect 3513 12699 3571 12705
rect 3513 12696 3525 12699
rect 2924 12668 3525 12696
rect 2924 12656 2930 12668
rect 3513 12665 3525 12668
rect 3559 12696 3571 12699
rect 3786 12696 3792 12708
rect 3559 12668 3792 12696
rect 3559 12665 3571 12668
rect 3513 12659 3571 12665
rect 3786 12656 3792 12668
rect 3844 12656 3850 12708
rect 3973 12699 4031 12705
rect 3973 12665 3985 12699
rect 4019 12696 4031 12699
rect 4632 12696 4660 12795
rect 5000 12764 5028 12804
rect 5718 12792 5724 12804
rect 5776 12792 5782 12844
rect 6549 12835 6607 12841
rect 6549 12801 6561 12835
rect 6595 12801 6607 12835
rect 6730 12832 6736 12844
rect 6691 12804 6736 12832
rect 6549 12795 6607 12801
rect 6454 12764 6460 12776
rect 5000 12736 6460 12764
rect 6454 12724 6460 12736
rect 6512 12724 6518 12776
rect 6564 12764 6592 12795
rect 6730 12792 6736 12804
rect 6788 12792 6794 12844
rect 6914 12832 6920 12844
rect 6972 12841 6978 12844
rect 6880 12804 6920 12832
rect 6914 12792 6920 12804
rect 6972 12795 6980 12841
rect 6972 12792 6978 12795
rect 7374 12792 7380 12844
rect 7432 12832 7438 12844
rect 7469 12835 7527 12841
rect 7469 12832 7481 12835
rect 7432 12804 7481 12832
rect 7432 12792 7438 12804
rect 7469 12801 7481 12804
rect 7515 12801 7527 12835
rect 7469 12795 7527 12801
rect 7742 12792 7748 12844
rect 7800 12832 7806 12844
rect 7837 12835 7895 12841
rect 7837 12832 7849 12835
rect 7800 12804 7849 12832
rect 7800 12792 7806 12804
rect 7837 12801 7849 12804
rect 7883 12801 7895 12835
rect 8754 12832 8760 12844
rect 8667 12804 8760 12832
rect 7837 12795 7895 12801
rect 8754 12792 8760 12804
rect 8812 12792 8818 12844
rect 8846 12792 8852 12844
rect 8904 12832 8910 12844
rect 9030 12832 9036 12844
rect 8904 12804 8949 12832
rect 8991 12804 9036 12832
rect 8904 12792 8910 12804
rect 9030 12792 9036 12804
rect 9088 12792 9094 12844
rect 9953 12835 10011 12841
rect 9953 12801 9965 12835
rect 9999 12801 10011 12835
rect 9953 12795 10011 12801
rect 7282 12764 7288 12776
rect 6564 12736 7288 12764
rect 7282 12724 7288 12736
rect 7340 12724 7346 12776
rect 7650 12724 7656 12776
rect 7708 12764 7714 12776
rect 8772 12764 8800 12792
rect 9968 12764 9996 12795
rect 10410 12792 10416 12844
rect 10468 12832 10474 12844
rect 10980 12841 11008 12940
rect 11882 12860 11888 12912
rect 11940 12900 11946 12912
rect 11940 12872 12480 12900
rect 11940 12860 11946 12872
rect 10781 12835 10839 12841
rect 10781 12832 10793 12835
rect 10468 12804 10793 12832
rect 10468 12792 10474 12804
rect 10781 12801 10793 12804
rect 10827 12801 10839 12835
rect 10781 12795 10839 12801
rect 10965 12835 11023 12841
rect 10965 12801 10977 12835
rect 11011 12801 11023 12835
rect 10965 12795 11023 12801
rect 11517 12835 11575 12841
rect 11517 12801 11529 12835
rect 11563 12832 11575 12835
rect 12158 12832 12164 12844
rect 11563 12804 12164 12832
rect 11563 12801 11575 12804
rect 11517 12795 11575 12801
rect 10594 12764 10600 12776
rect 7708 12736 9996 12764
rect 10555 12736 10600 12764
rect 7708 12724 7714 12736
rect 10594 12724 10600 12736
rect 10652 12724 10658 12776
rect 10796 12764 10824 12795
rect 11790 12764 11796 12776
rect 10796 12736 11796 12764
rect 11790 12724 11796 12736
rect 11848 12724 11854 12776
rect 4019 12668 4660 12696
rect 5905 12699 5963 12705
rect 4019 12665 4031 12668
rect 3973 12659 4031 12665
rect 5905 12665 5917 12699
rect 5951 12696 5963 12699
rect 5994 12696 6000 12708
rect 5951 12668 6000 12696
rect 5951 12665 5963 12668
rect 5905 12659 5963 12665
rect 5994 12656 6000 12668
rect 6052 12656 6058 12708
rect 8478 12696 8484 12708
rect 7024 12668 8484 12696
rect 1394 12628 1400 12640
rect 1355 12600 1400 12628
rect 1394 12588 1400 12600
rect 1452 12588 1458 12640
rect 4430 12588 4436 12640
rect 4488 12628 4494 12640
rect 7024 12628 7052 12668
rect 8478 12656 8484 12668
rect 8536 12696 8542 12708
rect 8938 12696 8944 12708
rect 8536 12668 8944 12696
rect 8536 12656 8542 12668
rect 8938 12656 8944 12668
rect 8996 12656 9002 12708
rect 9858 12656 9864 12708
rect 9916 12696 9922 12708
rect 10612 12696 10640 12724
rect 11900 12696 11928 12804
rect 12158 12792 12164 12804
rect 12216 12792 12222 12844
rect 12452 12841 12480 12872
rect 12618 12860 12624 12912
rect 12676 12900 12682 12912
rect 13081 12903 13139 12909
rect 13081 12900 13093 12903
rect 12676 12872 13093 12900
rect 12676 12860 12682 12872
rect 13081 12869 13093 12872
rect 13127 12900 13139 12903
rect 13357 12903 13415 12909
rect 13357 12900 13369 12903
rect 13127 12872 13369 12900
rect 13127 12869 13139 12872
rect 13081 12863 13139 12869
rect 13357 12869 13369 12872
rect 13403 12869 13415 12903
rect 13357 12863 13415 12869
rect 12437 12835 12495 12841
rect 12437 12801 12449 12835
rect 12483 12801 12495 12835
rect 12437 12795 12495 12801
rect 9916 12668 10640 12696
rect 11072 12668 11928 12696
rect 9916 12656 9922 12668
rect 4488 12600 7052 12628
rect 7101 12631 7159 12637
rect 4488 12588 4494 12600
rect 7101 12597 7113 12631
rect 7147 12628 7159 12631
rect 11072 12628 11100 12668
rect 12986 12656 12992 12708
rect 13044 12696 13050 12708
rect 13173 12699 13231 12705
rect 13173 12696 13185 12699
rect 13044 12668 13185 12696
rect 13044 12656 13050 12668
rect 13173 12665 13185 12668
rect 13219 12665 13231 12699
rect 13173 12659 13231 12665
rect 7147 12600 11100 12628
rect 11149 12631 11207 12637
rect 7147 12597 7159 12600
rect 7101 12591 7159 12597
rect 11149 12597 11161 12631
rect 11195 12628 11207 12631
rect 11238 12628 11244 12640
rect 11195 12600 11244 12628
rect 11195 12597 11207 12600
rect 11149 12591 11207 12597
rect 11238 12588 11244 12600
rect 11296 12588 11302 12640
rect 1104 12538 13892 12560
rect 1104 12486 4214 12538
rect 4266 12486 4278 12538
rect 4330 12486 4342 12538
rect 4394 12486 4406 12538
rect 4458 12486 4470 12538
rect 4522 12486 12214 12538
rect 12266 12486 12278 12538
rect 12330 12486 12342 12538
rect 12394 12486 12406 12538
rect 12458 12486 12470 12538
rect 12522 12486 13892 12538
rect 1104 12464 13892 12486
rect 2130 12384 2136 12436
rect 2188 12424 2194 12436
rect 2409 12427 2467 12433
rect 2409 12424 2421 12427
rect 2188 12396 2421 12424
rect 2188 12384 2194 12396
rect 2409 12393 2421 12396
rect 2455 12393 2467 12427
rect 2409 12387 2467 12393
rect 3878 12384 3884 12436
rect 3936 12424 3942 12436
rect 3973 12427 4031 12433
rect 3973 12424 3985 12427
rect 3936 12396 3985 12424
rect 3936 12384 3942 12396
rect 3973 12393 3985 12396
rect 4019 12393 4031 12427
rect 7650 12424 7656 12436
rect 7611 12396 7656 12424
rect 3973 12387 4031 12393
rect 7650 12384 7656 12396
rect 7708 12384 7714 12436
rect 7742 12384 7748 12436
rect 7800 12424 7806 12436
rect 8021 12427 8079 12433
rect 8021 12424 8033 12427
rect 7800 12396 8033 12424
rect 7800 12384 7806 12396
rect 8021 12393 8033 12396
rect 8067 12393 8079 12427
rect 8021 12387 8079 12393
rect 8662 12384 8668 12436
rect 8720 12424 8726 12436
rect 9033 12427 9091 12433
rect 9033 12424 9045 12427
rect 8720 12396 9045 12424
rect 8720 12384 8726 12396
rect 9033 12393 9045 12396
rect 9079 12424 9091 12427
rect 9490 12424 9496 12436
rect 9079 12396 9496 12424
rect 9079 12393 9091 12396
rect 9033 12387 9091 12393
rect 9490 12384 9496 12396
rect 9548 12384 9554 12436
rect 10686 12384 10692 12436
rect 10744 12424 10750 12436
rect 11974 12424 11980 12436
rect 10744 12396 11980 12424
rect 10744 12384 10750 12396
rect 11974 12384 11980 12396
rect 12032 12384 12038 12436
rect 1397 12223 1455 12229
rect 1397 12189 1409 12223
rect 1443 12220 1455 12223
rect 1578 12220 1584 12232
rect 1443 12192 1584 12220
rect 1443 12189 1455 12192
rect 1397 12183 1455 12189
rect 1578 12180 1584 12192
rect 1636 12180 1642 12232
rect 2038 12220 2044 12232
rect 1999 12192 2044 12220
rect 2038 12180 2044 12192
rect 2096 12180 2102 12232
rect 2593 12223 2651 12229
rect 2593 12220 2605 12223
rect 2424 12192 2605 12220
rect 2424 12164 2452 12192
rect 2593 12189 2605 12192
rect 2639 12189 2651 12223
rect 2593 12183 2651 12189
rect 2682 12180 2688 12232
rect 2740 12220 2746 12232
rect 3418 12220 3424 12232
rect 2740 12192 2785 12220
rect 3379 12192 3424 12220
rect 2740 12180 2746 12192
rect 3418 12180 3424 12192
rect 3476 12180 3482 12232
rect 3605 12223 3663 12229
rect 3605 12189 3617 12223
rect 3651 12220 3663 12223
rect 3896 12220 3924 12384
rect 5994 12356 6000 12368
rect 5955 12328 6000 12356
rect 5994 12316 6000 12328
rect 6052 12316 6058 12368
rect 6638 12316 6644 12368
rect 6696 12356 6702 12368
rect 6914 12356 6920 12368
rect 6696 12328 6920 12356
rect 6696 12316 6702 12328
rect 6914 12316 6920 12328
rect 6972 12356 6978 12368
rect 7285 12359 7343 12365
rect 6972 12328 7236 12356
rect 6972 12316 6978 12328
rect 5626 12248 5632 12300
rect 5684 12288 5690 12300
rect 5905 12291 5963 12297
rect 5905 12288 5917 12291
rect 5684 12260 5917 12288
rect 5684 12248 5690 12260
rect 5905 12257 5917 12260
rect 5951 12257 5963 12291
rect 6454 12288 6460 12300
rect 6415 12260 6460 12288
rect 5905 12251 5963 12257
rect 6454 12248 6460 12260
rect 6512 12248 6518 12300
rect 6656 12260 6960 12288
rect 3651 12192 3924 12220
rect 3651 12189 3663 12192
rect 3605 12183 3663 12189
rect 4062 12180 4068 12232
rect 4120 12220 4126 12232
rect 4341 12223 4399 12229
rect 4341 12220 4353 12223
rect 4120 12192 4353 12220
rect 4120 12180 4126 12192
rect 4341 12189 4353 12192
rect 4387 12189 4399 12223
rect 4798 12220 4804 12232
rect 4759 12192 4804 12220
rect 4341 12183 4399 12189
rect 4798 12180 4804 12192
rect 4856 12180 4862 12232
rect 4893 12223 4951 12229
rect 4893 12189 4905 12223
rect 4939 12220 4951 12223
rect 5074 12220 5080 12232
rect 4939 12192 5080 12220
rect 4939 12189 4951 12192
rect 4893 12183 4951 12189
rect 5074 12180 5080 12192
rect 5132 12180 5138 12232
rect 5534 12220 5540 12232
rect 5495 12192 5540 12220
rect 5534 12180 5540 12192
rect 5592 12180 5598 12232
rect 5810 12220 5816 12232
rect 5723 12192 5816 12220
rect 5810 12180 5816 12192
rect 5868 12220 5874 12232
rect 6086 12220 6092 12232
rect 5868 12192 6092 12220
rect 5868 12180 5874 12192
rect 6086 12180 6092 12192
rect 6144 12180 6150 12232
rect 6270 12180 6276 12232
rect 6328 12220 6334 12232
rect 6656 12220 6684 12260
rect 6328 12192 6684 12220
rect 6733 12223 6791 12229
rect 6328 12180 6334 12192
rect 6733 12189 6745 12223
rect 6779 12220 6791 12223
rect 6822 12220 6828 12232
rect 6779 12192 6828 12220
rect 6779 12189 6791 12192
rect 6733 12183 6791 12189
rect 6822 12180 6828 12192
rect 6880 12180 6886 12232
rect 6932 12229 6960 12260
rect 6917 12223 6975 12229
rect 6917 12189 6929 12223
rect 6963 12189 6975 12223
rect 7098 12220 7104 12232
rect 7156 12229 7162 12232
rect 7064 12192 7104 12220
rect 6917 12183 6975 12189
rect 7098 12180 7104 12192
rect 7156 12183 7164 12229
rect 7156 12180 7162 12183
rect 2317 12155 2375 12161
rect 2317 12121 2329 12155
rect 2363 12152 2375 12155
rect 2406 12152 2412 12164
rect 2363 12124 2412 12152
rect 2363 12121 2375 12124
rect 2317 12115 2375 12121
rect 2406 12112 2412 12124
rect 2464 12112 2470 12164
rect 2866 12112 2872 12164
rect 2924 12152 2930 12164
rect 3881 12155 3939 12161
rect 3881 12152 3893 12155
rect 2924 12124 3893 12152
rect 2924 12112 2930 12124
rect 3881 12121 3893 12124
rect 3927 12121 3939 12155
rect 3881 12115 3939 12121
rect 4525 12155 4583 12161
rect 4525 12121 4537 12155
rect 4571 12152 4583 12155
rect 6638 12152 6644 12164
rect 4571 12124 6644 12152
rect 4571 12121 4583 12124
rect 4525 12115 4583 12121
rect 6638 12112 6644 12124
rect 6696 12112 6702 12164
rect 7006 12152 7012 12164
rect 6919 12124 7012 12152
rect 7006 12112 7012 12124
rect 7064 12112 7070 12164
rect 7208 12152 7236 12328
rect 7285 12325 7297 12359
rect 7331 12356 7343 12359
rect 7331 12328 12020 12356
rect 7331 12325 7343 12328
rect 7285 12319 7343 12325
rect 8464 12291 8522 12297
rect 8464 12257 8476 12291
rect 8510 12288 8522 12291
rect 8846 12288 8852 12300
rect 8510 12260 8852 12288
rect 8510 12257 8522 12260
rect 8464 12251 8522 12257
rect 8846 12248 8852 12260
rect 8904 12248 8910 12300
rect 9030 12248 9036 12300
rect 9088 12288 9094 12300
rect 9401 12291 9459 12297
rect 9401 12288 9413 12291
rect 9088 12260 9413 12288
rect 9088 12248 9094 12260
rect 9401 12257 9413 12260
rect 9447 12257 9459 12291
rect 9950 12288 9956 12300
rect 9911 12260 9956 12288
rect 9401 12251 9459 12257
rect 9950 12248 9956 12260
rect 10008 12248 10014 12300
rect 10580 12291 10638 12297
rect 10580 12257 10592 12291
rect 10626 12288 10638 12291
rect 10686 12288 10692 12300
rect 10626 12260 10692 12288
rect 10626 12257 10638 12260
rect 10580 12251 10638 12257
rect 10686 12248 10692 12260
rect 10744 12248 10750 12300
rect 10781 12291 10839 12297
rect 10781 12257 10793 12291
rect 10827 12288 10839 12291
rect 11330 12288 11336 12300
rect 10827 12260 11336 12288
rect 10827 12257 10839 12260
rect 10781 12251 10839 12257
rect 11330 12248 11336 12260
rect 11388 12248 11394 12300
rect 7929 12223 7987 12229
rect 7929 12189 7941 12223
rect 7975 12220 7987 12223
rect 8662 12220 8668 12232
rect 7975 12192 8668 12220
rect 7975 12189 7987 12192
rect 7929 12183 7987 12189
rect 8662 12180 8668 12192
rect 8720 12180 8726 12232
rect 8757 12223 8815 12229
rect 8757 12189 8769 12223
rect 8803 12220 8815 12223
rect 9306 12220 9312 12232
rect 8803 12192 8984 12220
rect 9267 12192 9312 12220
rect 8803 12189 8815 12192
rect 8757 12183 8815 12189
rect 7469 12155 7527 12161
rect 7469 12152 7481 12155
rect 7208 12124 7481 12152
rect 7469 12121 7481 12124
rect 7515 12121 7527 12155
rect 8110 12152 8116 12164
rect 7469 12115 7527 12121
rect 7576 12124 8116 12152
rect 1854 12044 1860 12096
rect 1912 12084 1918 12096
rect 5442 12084 5448 12096
rect 1912 12056 5448 12084
rect 1912 12044 1918 12056
rect 5442 12044 5448 12056
rect 5500 12044 5506 12096
rect 6546 12084 6552 12096
rect 6507 12056 6552 12084
rect 6546 12044 6552 12056
rect 6604 12084 6610 12096
rect 7024 12084 7052 12112
rect 7576 12084 7604 12124
rect 8110 12112 8116 12124
rect 8168 12152 8174 12164
rect 8205 12155 8263 12161
rect 8205 12152 8217 12155
rect 8168 12124 8217 12152
rect 8168 12112 8174 12124
rect 8205 12121 8217 12124
rect 8251 12121 8263 12155
rect 8205 12115 8263 12121
rect 6604 12056 7604 12084
rect 7653 12087 7711 12093
rect 6604 12044 6610 12056
rect 7653 12053 7665 12087
rect 7699 12084 7711 12087
rect 7742 12084 7748 12096
rect 7699 12056 7748 12084
rect 7699 12053 7711 12056
rect 7653 12047 7711 12053
rect 7742 12044 7748 12056
rect 7800 12044 7806 12096
rect 8478 12044 8484 12096
rect 8536 12084 8542 12096
rect 8573 12087 8631 12093
rect 8573 12084 8585 12087
rect 8536 12056 8585 12084
rect 8536 12044 8542 12056
rect 8573 12053 8585 12056
rect 8619 12053 8631 12087
rect 8573 12047 8631 12053
rect 8662 12044 8668 12096
rect 8720 12084 8726 12096
rect 8956 12084 8984 12192
rect 9306 12180 9312 12192
rect 9364 12180 9370 12232
rect 9858 12220 9864 12232
rect 9819 12192 9864 12220
rect 9858 12180 9864 12192
rect 9916 12180 9922 12232
rect 10321 12223 10379 12229
rect 10321 12189 10333 12223
rect 10367 12220 10379 12223
rect 10410 12220 10416 12232
rect 10367 12192 10416 12220
rect 10367 12189 10379 12192
rect 10321 12183 10379 12189
rect 10410 12180 10416 12192
rect 10468 12180 10474 12232
rect 10870 12220 10876 12232
rect 10831 12192 10876 12220
rect 10870 12180 10876 12192
rect 10928 12180 10934 12232
rect 10965 12223 11023 12229
rect 10965 12189 10977 12223
rect 11011 12220 11023 12223
rect 11238 12220 11244 12232
rect 11011 12192 11244 12220
rect 11011 12189 11023 12192
rect 10965 12183 11023 12189
rect 11238 12180 11244 12192
rect 11296 12220 11302 12232
rect 11606 12220 11612 12232
rect 11296 12192 11376 12220
rect 11567 12192 11612 12220
rect 11296 12180 11302 12192
rect 9122 12152 9128 12164
rect 9083 12124 9128 12152
rect 9122 12112 9128 12124
rect 9180 12112 9186 12164
rect 9214 12112 9220 12164
rect 9272 12152 9278 12164
rect 10137 12155 10195 12161
rect 10137 12152 10149 12155
rect 9272 12124 10149 12152
rect 9272 12112 9278 12124
rect 10137 12121 10149 12124
rect 10183 12121 10195 12155
rect 11348 12152 11376 12192
rect 11606 12180 11612 12192
rect 11664 12180 11670 12232
rect 11882 12220 11888 12232
rect 11843 12192 11888 12220
rect 11882 12180 11888 12192
rect 11940 12180 11946 12232
rect 11992 12229 12020 12328
rect 11977 12223 12035 12229
rect 11977 12189 11989 12223
rect 12023 12220 12035 12223
rect 12802 12220 12808 12232
rect 12023 12192 12808 12220
rect 12023 12189 12035 12192
rect 11977 12183 12035 12189
rect 12802 12180 12808 12192
rect 12860 12180 12866 12232
rect 12986 12220 12992 12232
rect 12947 12192 12992 12220
rect 12986 12180 12992 12192
rect 13044 12180 13050 12232
rect 12066 12152 12072 12164
rect 10137 12115 10195 12121
rect 10520 12124 11100 12152
rect 11348 12124 12072 12152
rect 10520 12084 10548 12124
rect 10686 12084 10692 12096
rect 8720 12056 8765 12084
rect 8956 12056 10548 12084
rect 10647 12056 10692 12084
rect 8720 12044 8726 12056
rect 10686 12044 10692 12056
rect 10744 12044 10750 12096
rect 11072 12084 11100 12124
rect 12066 12112 12072 12124
rect 12124 12112 12130 12164
rect 13262 12112 13268 12164
rect 13320 12152 13326 12164
rect 13541 12155 13599 12161
rect 13541 12152 13553 12155
rect 13320 12124 13553 12152
rect 13320 12112 13326 12124
rect 13541 12121 13553 12124
rect 13587 12121 13599 12155
rect 13541 12115 13599 12121
rect 11422 12084 11428 12096
rect 11072 12056 11428 12084
rect 11422 12044 11428 12056
rect 11480 12044 11486 12096
rect 1104 11994 13892 12016
rect 1104 11942 8214 11994
rect 8266 11942 8278 11994
rect 8330 11942 8342 11994
rect 8394 11942 8406 11994
rect 8458 11942 8470 11994
rect 8522 11942 13892 11994
rect 1104 11920 13892 11942
rect 1765 11883 1823 11889
rect 1765 11849 1777 11883
rect 1811 11880 1823 11883
rect 2038 11880 2044 11892
rect 1811 11852 2044 11880
rect 1811 11849 1823 11852
rect 1765 11843 1823 11849
rect 2038 11840 2044 11852
rect 2096 11840 2102 11892
rect 3421 11883 3479 11889
rect 3421 11849 3433 11883
rect 3467 11880 3479 11883
rect 4062 11880 4068 11892
rect 3467 11852 4068 11880
rect 3467 11849 3479 11852
rect 3421 11843 3479 11849
rect 4062 11840 4068 11852
rect 4120 11840 4126 11892
rect 6457 11883 6515 11889
rect 6457 11849 6469 11883
rect 6503 11880 6515 11883
rect 6546 11880 6552 11892
rect 6503 11852 6552 11880
rect 6503 11849 6515 11852
rect 6457 11843 6515 11849
rect 6546 11840 6552 11852
rect 6604 11840 6610 11892
rect 6822 11880 6828 11892
rect 6783 11852 6828 11880
rect 6822 11840 6828 11852
rect 6880 11840 6886 11892
rect 7834 11880 7840 11892
rect 7024 11852 7840 11880
rect 1394 11772 1400 11824
rect 1452 11812 1458 11824
rect 1489 11815 1547 11821
rect 1489 11812 1501 11815
rect 1452 11784 1501 11812
rect 1452 11772 1458 11784
rect 1489 11781 1501 11784
rect 1535 11812 1547 11815
rect 2593 11815 2651 11821
rect 2593 11812 2605 11815
rect 1535 11784 2605 11812
rect 1535 11781 1547 11784
rect 1489 11775 1547 11781
rect 2593 11781 2605 11784
rect 2639 11812 2651 11815
rect 3142 11812 3148 11824
rect 2639 11784 3148 11812
rect 2639 11781 2651 11784
rect 2593 11775 2651 11781
rect 3142 11772 3148 11784
rect 3200 11772 3206 11824
rect 3786 11812 3792 11824
rect 3747 11784 3792 11812
rect 3786 11772 3792 11784
rect 3844 11772 3850 11824
rect 5442 11772 5448 11824
rect 5500 11812 5506 11824
rect 5537 11815 5595 11821
rect 5537 11812 5549 11815
rect 5500 11784 5549 11812
rect 5500 11772 5506 11784
rect 5537 11781 5549 11784
rect 5583 11781 5595 11815
rect 7024 11812 7052 11852
rect 7834 11840 7840 11852
rect 7892 11880 7898 11892
rect 8386 11880 8392 11892
rect 7892 11852 8294 11880
rect 8347 11852 8392 11880
rect 7892 11840 7898 11852
rect 5537 11775 5595 11781
rect 6012 11784 7052 11812
rect 6012 11756 6040 11784
rect 2498 11744 2504 11756
rect 2459 11716 2504 11744
rect 2498 11704 2504 11716
rect 2556 11704 2562 11756
rect 2682 11704 2688 11756
rect 2740 11744 2746 11756
rect 2777 11747 2835 11753
rect 2777 11744 2789 11747
rect 2740 11716 2789 11744
rect 2740 11704 2746 11716
rect 2777 11713 2789 11716
rect 2823 11713 2835 11747
rect 2777 11707 2835 11713
rect 5074 11704 5080 11756
rect 5132 11744 5138 11756
rect 5169 11747 5227 11753
rect 5169 11744 5181 11747
rect 5132 11716 5181 11744
rect 5132 11704 5138 11716
rect 5169 11713 5181 11716
rect 5215 11713 5227 11747
rect 5169 11707 5227 11713
rect 5779 11747 5837 11753
rect 5779 11713 5791 11747
rect 5825 11744 5837 11747
rect 5905 11747 5963 11753
rect 5825 11713 5855 11744
rect 5779 11707 5855 11713
rect 5905 11713 5917 11747
rect 5951 11713 5963 11747
rect 5905 11707 5963 11713
rect 1673 11679 1731 11685
rect 1673 11645 1685 11679
rect 1719 11676 1731 11679
rect 1857 11679 1915 11685
rect 1857 11676 1869 11679
rect 1719 11648 1869 11676
rect 1719 11645 1731 11648
rect 1673 11639 1731 11645
rect 1857 11645 1869 11648
rect 1903 11645 1915 11679
rect 1857 11639 1915 11645
rect 2222 11636 2228 11688
rect 2280 11676 2286 11688
rect 2409 11679 2467 11685
rect 2409 11676 2421 11679
rect 2280 11648 2421 11676
rect 2280 11636 2286 11648
rect 2409 11645 2421 11648
rect 2455 11676 2467 11679
rect 2961 11679 3019 11685
rect 2961 11676 2973 11679
rect 2455 11648 2973 11676
rect 2455 11645 2467 11648
rect 2409 11639 2467 11645
rect 2961 11645 2973 11648
rect 3007 11645 3019 11679
rect 2961 11639 3019 11645
rect 4249 11679 4307 11685
rect 4249 11645 4261 11679
rect 4295 11676 4307 11679
rect 4706 11676 4712 11688
rect 4295 11648 4712 11676
rect 4295 11645 4307 11648
rect 4249 11639 4307 11645
rect 4706 11636 4712 11648
rect 4764 11636 4770 11688
rect 4801 11679 4859 11685
rect 4801 11645 4813 11679
rect 4847 11676 4859 11679
rect 4982 11676 4988 11688
rect 4847 11648 4988 11676
rect 4847 11645 4859 11648
rect 4801 11639 4859 11645
rect 4982 11636 4988 11648
rect 5040 11636 5046 11688
rect 5353 11679 5411 11685
rect 5353 11645 5365 11679
rect 5399 11676 5411 11679
rect 5626 11676 5632 11688
rect 5399 11648 5632 11676
rect 5399 11645 5411 11648
rect 5353 11639 5411 11645
rect 5626 11636 5632 11648
rect 5684 11636 5690 11688
rect 1949 11611 2007 11617
rect 1949 11577 1961 11611
rect 1995 11608 2007 11611
rect 2866 11608 2872 11620
rect 1995 11580 2872 11608
rect 1995 11577 2007 11580
rect 1949 11571 2007 11577
rect 2866 11568 2872 11580
rect 2924 11568 2930 11620
rect 3694 11608 3700 11620
rect 3528 11580 3700 11608
rect 3142 11540 3148 11552
rect 3103 11512 3148 11540
rect 3142 11500 3148 11512
rect 3200 11540 3206 11552
rect 3528 11549 3556 11580
rect 3694 11568 3700 11580
rect 3752 11608 3758 11620
rect 4065 11611 4123 11617
rect 4065 11608 4077 11611
rect 3752 11580 4077 11608
rect 3752 11568 3758 11580
rect 4065 11577 4077 11580
rect 4111 11577 4123 11611
rect 4065 11571 4123 11577
rect 4341 11611 4399 11617
rect 4341 11577 4353 11611
rect 4387 11608 4399 11611
rect 4614 11608 4620 11620
rect 4387 11580 4620 11608
rect 4387 11577 4399 11580
rect 4341 11571 4399 11577
rect 3513 11543 3571 11549
rect 3513 11540 3525 11543
rect 3200 11512 3525 11540
rect 3200 11500 3206 11512
rect 3513 11509 3525 11512
rect 3559 11509 3571 11543
rect 3878 11540 3884 11552
rect 3839 11512 3884 11540
rect 3513 11503 3571 11509
rect 3878 11500 3884 11512
rect 3936 11500 3942 11552
rect 4080 11540 4108 11571
rect 4614 11568 4620 11580
rect 4672 11568 4678 11620
rect 5534 11568 5540 11620
rect 5592 11608 5598 11620
rect 5827 11608 5855 11707
rect 5920 11676 5948 11707
rect 5994 11704 6000 11756
rect 6052 11744 6058 11756
rect 6052 11716 6097 11744
rect 6052 11704 6058 11716
rect 6178 11704 6184 11756
rect 6236 11744 6242 11756
rect 6730 11744 6736 11756
rect 6236 11716 6736 11744
rect 6236 11704 6242 11716
rect 6730 11704 6736 11716
rect 6788 11704 6794 11756
rect 7024 11753 7052 11784
rect 7282 11772 7288 11824
rect 7340 11812 7346 11824
rect 7469 11815 7527 11821
rect 7469 11812 7481 11815
rect 7340 11784 7481 11812
rect 7340 11772 7346 11784
rect 7469 11781 7481 11784
rect 7515 11781 7527 11815
rect 7469 11775 7527 11781
rect 7742 11772 7748 11824
rect 7800 11812 7806 11824
rect 8021 11815 8079 11821
rect 8021 11812 8033 11815
rect 7800 11784 8033 11812
rect 7800 11772 7806 11784
rect 8021 11781 8033 11784
rect 8067 11781 8079 11815
rect 8266 11812 8294 11852
rect 8386 11840 8392 11852
rect 8444 11840 8450 11892
rect 8662 11840 8668 11892
rect 8720 11880 8726 11892
rect 8941 11883 8999 11889
rect 8941 11880 8953 11883
rect 8720 11852 8953 11880
rect 8720 11840 8726 11852
rect 8941 11849 8953 11852
rect 8987 11849 8999 11883
rect 8941 11843 8999 11849
rect 9217 11883 9275 11889
rect 9217 11849 9229 11883
rect 9263 11880 9275 11883
rect 10505 11883 10563 11889
rect 9263 11852 10456 11880
rect 9263 11849 9275 11852
rect 9217 11843 9275 11849
rect 8573 11815 8631 11821
rect 8266 11784 8524 11812
rect 8021 11775 8079 11781
rect 7009 11747 7067 11753
rect 7009 11713 7021 11747
rect 7055 11713 7067 11747
rect 7009 11707 7067 11713
rect 7101 11747 7159 11753
rect 7101 11713 7113 11747
rect 7147 11713 7159 11747
rect 7374 11744 7380 11756
rect 7335 11716 7380 11744
rect 7101 11707 7159 11713
rect 6454 11676 6460 11688
rect 5920 11648 6460 11676
rect 6454 11636 6460 11648
rect 6512 11636 6518 11688
rect 5592 11580 5855 11608
rect 5592 11568 5598 11580
rect 6546 11568 6552 11620
rect 6604 11608 6610 11620
rect 6641 11611 6699 11617
rect 6641 11608 6653 11611
rect 6604 11580 6653 11608
rect 6604 11568 6610 11580
rect 6641 11577 6653 11580
rect 6687 11608 6699 11611
rect 6730 11608 6736 11620
rect 6687 11580 6736 11608
rect 6687 11577 6699 11580
rect 6641 11571 6699 11577
rect 6730 11568 6736 11580
rect 6788 11568 6794 11620
rect 7116 11608 7144 11707
rect 7374 11704 7380 11716
rect 7432 11744 7438 11756
rect 7650 11744 7656 11756
rect 7432 11716 7656 11744
rect 7432 11704 7438 11716
rect 7650 11704 7656 11716
rect 7708 11704 7714 11756
rect 7834 11744 7840 11756
rect 7795 11716 7840 11744
rect 7834 11704 7840 11716
rect 7892 11704 7898 11756
rect 8202 11744 8208 11756
rect 8163 11716 8208 11744
rect 8202 11704 8208 11716
rect 8260 11704 8266 11756
rect 8496 11753 8524 11784
rect 8573 11781 8585 11815
rect 8619 11781 8631 11815
rect 8754 11812 8760 11824
rect 8715 11784 8760 11812
rect 8573 11775 8631 11781
rect 8481 11747 8539 11753
rect 8481 11713 8493 11747
rect 8527 11713 8539 11747
rect 8481 11707 8539 11713
rect 7742 11636 7748 11688
rect 7800 11676 7806 11688
rect 8588 11676 8616 11775
rect 8754 11772 8760 11784
rect 8812 11772 8818 11824
rect 9582 11772 9588 11824
rect 9640 11812 9646 11824
rect 10321 11815 10379 11821
rect 10321 11812 10333 11815
rect 9640 11784 10333 11812
rect 9640 11772 9646 11784
rect 10321 11781 10333 11784
rect 10367 11781 10379 11815
rect 10428 11812 10456 11852
rect 10505 11849 10517 11883
rect 10551 11880 10563 11883
rect 10778 11880 10784 11892
rect 10551 11852 10784 11880
rect 10551 11849 10563 11852
rect 10505 11843 10563 11849
rect 10778 11840 10784 11852
rect 10836 11840 10842 11892
rect 11974 11840 11980 11892
rect 12032 11880 12038 11892
rect 12069 11883 12127 11889
rect 12069 11880 12081 11883
rect 12032 11852 12081 11880
rect 12032 11840 12038 11852
rect 12069 11849 12081 11852
rect 12115 11880 12127 11883
rect 13170 11880 13176 11892
rect 12115 11852 13176 11880
rect 12115 11849 12127 11852
rect 12069 11843 12127 11849
rect 13170 11840 13176 11852
rect 13228 11840 13234 11892
rect 13446 11880 13452 11892
rect 13407 11852 13452 11880
rect 13446 11840 13452 11852
rect 13504 11840 13510 11892
rect 10594 11812 10600 11824
rect 10428 11784 10600 11812
rect 10321 11775 10379 11781
rect 10594 11772 10600 11784
rect 10652 11772 10658 11824
rect 10686 11772 10692 11824
rect 10744 11812 10750 11824
rect 10873 11815 10931 11821
rect 10873 11812 10885 11815
rect 10744 11784 10885 11812
rect 10744 11772 10750 11784
rect 10873 11781 10885 11784
rect 10919 11781 10931 11815
rect 10873 11775 10931 11781
rect 12713 11815 12771 11821
rect 12713 11781 12725 11815
rect 12759 11812 12771 11815
rect 12894 11812 12900 11824
rect 12759 11784 12900 11812
rect 12759 11781 12771 11784
rect 12713 11775 12771 11781
rect 12894 11772 12900 11784
rect 12952 11772 12958 11824
rect 13354 11812 13360 11824
rect 13315 11784 13360 11812
rect 13354 11772 13360 11784
rect 13412 11772 13418 11824
rect 9490 11744 9496 11756
rect 9451 11716 9496 11744
rect 9490 11704 9496 11716
rect 9548 11704 9554 11756
rect 9674 11704 9680 11756
rect 9732 11744 9738 11756
rect 9858 11744 9864 11756
rect 9732 11716 9776 11744
rect 9819 11716 9864 11744
rect 9732 11704 9738 11716
rect 9858 11704 9864 11716
rect 9916 11704 9922 11756
rect 9950 11704 9956 11756
rect 10008 11744 10014 11756
rect 10045 11747 10103 11753
rect 10045 11744 10057 11747
rect 10008 11716 10057 11744
rect 10008 11704 10014 11716
rect 10045 11713 10057 11716
rect 10091 11713 10103 11747
rect 11057 11747 11115 11753
rect 11057 11744 11069 11747
rect 10045 11707 10103 11713
rect 10152 11716 11069 11744
rect 7800 11648 8616 11676
rect 7800 11636 7806 11648
rect 9398 11636 9404 11688
rect 9456 11676 9462 11688
rect 9769 11679 9827 11685
rect 9769 11676 9781 11679
rect 9456 11648 9781 11676
rect 9456 11636 9462 11648
rect 9769 11645 9781 11648
rect 9815 11645 9827 11679
rect 10152 11676 10180 11716
rect 11057 11713 11069 11716
rect 11103 11713 11115 11747
rect 11057 11707 11115 11713
rect 11146 11704 11152 11756
rect 11204 11744 11210 11756
rect 11241 11747 11299 11753
rect 11241 11744 11253 11747
rect 11204 11716 11253 11744
rect 11204 11704 11210 11716
rect 11241 11713 11253 11716
rect 11287 11744 11299 11747
rect 11517 11747 11575 11753
rect 11517 11744 11529 11747
rect 11287 11716 11529 11744
rect 11287 11713 11299 11716
rect 11241 11707 11299 11713
rect 11517 11713 11529 11716
rect 11563 11713 11575 11747
rect 11698 11744 11704 11756
rect 11659 11716 11704 11744
rect 11517 11707 11575 11713
rect 11698 11704 11704 11716
rect 11756 11704 11762 11756
rect 12621 11747 12679 11753
rect 12621 11713 12633 11747
rect 12667 11744 12679 11747
rect 13078 11744 13084 11756
rect 12667 11716 13084 11744
rect 12667 11713 12679 11716
rect 12621 11707 12679 11713
rect 13078 11704 13084 11716
rect 13136 11704 13142 11756
rect 13262 11744 13268 11756
rect 13223 11716 13268 11744
rect 13262 11704 13268 11716
rect 13320 11704 13326 11756
rect 9769 11639 9827 11645
rect 9968 11648 10180 11676
rect 10229 11679 10287 11685
rect 8202 11608 8208 11620
rect 7116 11580 8208 11608
rect 8202 11568 8208 11580
rect 8260 11568 8266 11620
rect 9214 11568 9220 11620
rect 9272 11608 9278 11620
rect 9968 11608 9996 11648
rect 10229 11645 10241 11679
rect 10275 11676 10287 11679
rect 11330 11676 11336 11688
rect 10275 11648 11336 11676
rect 10275 11645 10287 11648
rect 10229 11639 10287 11645
rect 11330 11636 11336 11648
rect 11388 11636 11394 11688
rect 12066 11636 12072 11688
rect 12124 11676 12130 11688
rect 12161 11679 12219 11685
rect 12161 11676 12173 11679
rect 12124 11648 12173 11676
rect 12124 11636 12130 11648
rect 12161 11645 12173 11648
rect 12207 11645 12219 11679
rect 12802 11676 12808 11688
rect 12763 11648 12808 11676
rect 12161 11639 12219 11645
rect 12802 11636 12808 11648
rect 12860 11636 12866 11688
rect 9272 11580 9996 11608
rect 9272 11568 9278 11580
rect 10042 11568 10048 11620
rect 10100 11608 10106 11620
rect 10100 11580 10548 11608
rect 10100 11568 10106 11580
rect 4798 11540 4804 11552
rect 4080 11512 4804 11540
rect 4798 11500 4804 11512
rect 4856 11540 4862 11552
rect 4893 11543 4951 11549
rect 4893 11540 4905 11543
rect 4856 11512 4905 11540
rect 4856 11500 4862 11512
rect 4893 11509 4905 11512
rect 4939 11509 4951 11543
rect 4893 11503 4951 11509
rect 6454 11500 6460 11552
rect 6512 11540 6518 11552
rect 7285 11543 7343 11549
rect 7285 11540 7297 11543
rect 6512 11512 7297 11540
rect 6512 11500 6518 11512
rect 7285 11509 7297 11512
rect 7331 11540 7343 11543
rect 7374 11540 7380 11552
rect 7331 11512 7380 11540
rect 7331 11509 7343 11512
rect 7285 11503 7343 11509
rect 7374 11500 7380 11512
rect 7432 11540 7438 11552
rect 8386 11540 8392 11552
rect 7432 11512 8392 11540
rect 7432 11500 7438 11512
rect 8386 11500 8392 11512
rect 8444 11500 8450 11552
rect 8662 11500 8668 11552
rect 8720 11540 8726 11552
rect 8757 11543 8815 11549
rect 8757 11540 8769 11543
rect 8720 11512 8769 11540
rect 8720 11500 8726 11512
rect 8757 11509 8769 11512
rect 8803 11509 8815 11543
rect 8757 11503 8815 11509
rect 9030 11500 9036 11552
rect 9088 11540 9094 11552
rect 9401 11543 9459 11549
rect 9401 11540 9413 11543
rect 9088 11512 9413 11540
rect 9088 11500 9094 11512
rect 9401 11509 9413 11512
rect 9447 11540 9459 11543
rect 9490 11540 9496 11552
rect 9447 11512 9496 11540
rect 9447 11509 9459 11512
rect 9401 11503 9459 11509
rect 9490 11500 9496 11512
rect 9548 11500 9554 11552
rect 10520 11549 10548 11580
rect 10505 11543 10563 11549
rect 10505 11509 10517 11543
rect 10551 11509 10563 11543
rect 10686 11540 10692 11552
rect 10647 11512 10692 11540
rect 10505 11503 10563 11509
rect 10686 11500 10692 11512
rect 10744 11540 10750 11552
rect 10870 11540 10876 11552
rect 10744 11512 10876 11540
rect 10744 11500 10750 11512
rect 10870 11500 10876 11512
rect 10928 11500 10934 11552
rect 11054 11500 11060 11552
rect 11112 11540 11118 11552
rect 11793 11543 11851 11549
rect 11793 11540 11805 11543
rect 11112 11512 11805 11540
rect 11112 11500 11118 11512
rect 11793 11509 11805 11512
rect 11839 11509 11851 11543
rect 11793 11503 11851 11509
rect 1104 11450 13892 11472
rect 1104 11398 4214 11450
rect 4266 11398 4278 11450
rect 4330 11398 4342 11450
rect 4394 11398 4406 11450
rect 4458 11398 4470 11450
rect 4522 11398 12214 11450
rect 12266 11398 12278 11450
rect 12330 11398 12342 11450
rect 12394 11398 12406 11450
rect 12458 11398 12470 11450
rect 12522 11398 13892 11450
rect 1104 11376 13892 11398
rect 8662 11336 8668 11348
rect 8623 11308 8668 11336
rect 8662 11296 8668 11308
rect 8720 11296 8726 11348
rect 8846 11296 8852 11348
rect 8904 11336 8910 11348
rect 8941 11339 8999 11345
rect 8941 11336 8953 11339
rect 8904 11308 8953 11336
rect 8904 11296 8910 11308
rect 8941 11305 8953 11308
rect 8987 11305 8999 11339
rect 9122 11336 9128 11348
rect 9083 11308 9128 11336
rect 8941 11299 8999 11305
rect 9122 11296 9128 11308
rect 9180 11296 9186 11348
rect 9306 11336 9312 11348
rect 9232 11308 9312 11336
rect 2866 11268 2872 11280
rect 2827 11240 2872 11268
rect 2866 11228 2872 11240
rect 2924 11228 2930 11280
rect 3510 11228 3516 11280
rect 3568 11268 3574 11280
rect 5074 11268 5080 11280
rect 3568 11240 5080 11268
rect 3568 11228 3574 11240
rect 5074 11228 5080 11240
rect 5132 11228 5138 11280
rect 5629 11271 5687 11277
rect 5629 11237 5641 11271
rect 5675 11268 5687 11271
rect 6086 11268 6092 11280
rect 5675 11240 6092 11268
rect 5675 11237 5687 11240
rect 5629 11231 5687 11237
rect 6086 11228 6092 11240
rect 6144 11228 6150 11280
rect 7653 11271 7711 11277
rect 6196 11240 7144 11268
rect 4522 11160 4528 11212
rect 4580 11200 4586 11212
rect 5166 11200 5172 11212
rect 4580 11172 5172 11200
rect 4580 11160 4586 11172
rect 5166 11160 5172 11172
rect 5224 11200 5230 11212
rect 6196 11209 6224 11240
rect 5885 11203 5943 11209
rect 5885 11200 5897 11203
rect 5224 11172 5897 11200
rect 5224 11160 5230 11172
rect 5885 11169 5897 11172
rect 5931 11169 5943 11203
rect 5885 11163 5943 11169
rect 6181 11203 6239 11209
rect 6181 11169 6193 11203
rect 6227 11169 6239 11203
rect 6181 11163 6239 11169
rect 6380 11172 6868 11200
rect 1397 11135 1455 11141
rect 1397 11101 1409 11135
rect 1443 11132 1455 11135
rect 2222 11132 2228 11144
rect 1443 11104 2228 11132
rect 1443 11101 1455 11104
rect 1397 11095 1455 11101
rect 2222 11092 2228 11104
rect 2280 11092 2286 11144
rect 2406 11132 2412 11144
rect 2367 11104 2412 11132
rect 2406 11092 2412 11104
rect 2464 11092 2470 11144
rect 3053 11135 3111 11141
rect 3053 11101 3065 11135
rect 3099 11132 3111 11135
rect 3326 11132 3332 11144
rect 3099 11104 3332 11132
rect 3099 11101 3111 11104
rect 3053 11095 3111 11101
rect 3326 11092 3332 11104
rect 3384 11132 3390 11144
rect 3789 11135 3847 11141
rect 3789 11132 3801 11135
rect 3384 11104 3801 11132
rect 3384 11092 3390 11104
rect 3789 11101 3801 11104
rect 3835 11101 3847 11135
rect 3789 11095 3847 11101
rect 3878 11092 3884 11144
rect 3936 11132 3942 11144
rect 4709 11135 4767 11141
rect 4709 11132 4721 11135
rect 3936 11104 4721 11132
rect 3936 11092 3942 11104
rect 4709 11101 4721 11104
rect 4755 11101 4767 11135
rect 4709 11095 4767 11101
rect 4798 11092 4804 11144
rect 4856 11132 4862 11144
rect 5629 11135 5687 11141
rect 5629 11132 5641 11135
rect 4856 11104 5641 11132
rect 4856 11092 4862 11104
rect 5629 11101 5641 11104
rect 5675 11101 5687 11135
rect 6380 11132 6408 11172
rect 5629 11095 5687 11101
rect 6104 11104 6408 11132
rect 6104 11076 6132 11104
rect 6546 11092 6552 11144
rect 6604 11092 6610 11144
rect 6751 11135 6809 11141
rect 6640 11113 6698 11119
rect 6548 11079 6560 11092
rect 6594 11079 6606 11092
rect 3510 11064 3516 11076
rect 3471 11036 3516 11064
rect 3510 11024 3516 11036
rect 3568 11024 3574 11076
rect 3602 11024 3608 11076
rect 3660 11064 3666 11076
rect 5902 11064 5908 11076
rect 3660 11036 3705 11064
rect 5815 11036 5908 11064
rect 3660 11024 3666 11036
rect 2682 10956 2688 11008
rect 2740 10996 2746 11008
rect 5828 10996 5856 11036
rect 5902 11024 5908 11036
rect 5960 11064 5966 11076
rect 6086 11064 6092 11076
rect 5960 11036 6092 11064
rect 5960 11024 5966 11036
rect 6086 11024 6092 11036
rect 6144 11024 6150 11076
rect 6270 11064 6276 11076
rect 6231 11036 6276 11064
rect 6270 11024 6276 11036
rect 6328 11024 6334 11076
rect 6548 11073 6606 11079
rect 6640 11079 6652 11113
rect 6686 11079 6698 11113
rect 6751 11101 6763 11135
rect 6797 11132 6809 11135
rect 6840 11132 6868 11172
rect 6797 11104 6868 11132
rect 6917 11135 6975 11141
rect 6797 11101 6809 11104
rect 6751 11095 6809 11101
rect 6917 11101 6929 11135
rect 6963 11101 6975 11135
rect 6917 11095 6975 11101
rect 6640 11073 6698 11079
rect 5994 10996 6000 11008
rect 2740 10968 5856 10996
rect 5955 10968 6000 10996
rect 2740 10956 2746 10968
rect 5994 10956 6000 10968
rect 6052 10996 6058 11008
rect 6655 10996 6683 11073
rect 6932 11064 6960 11095
rect 7006 11092 7012 11144
rect 7064 11132 7070 11144
rect 7116 11132 7144 11240
rect 7653 11237 7665 11271
rect 7699 11268 7711 11271
rect 7742 11268 7748 11280
rect 7699 11240 7748 11268
rect 7699 11237 7711 11240
rect 7653 11231 7711 11237
rect 7742 11228 7748 11240
rect 7800 11228 7806 11280
rect 7834 11228 7840 11280
rect 7892 11268 7898 11280
rect 8205 11271 8263 11277
rect 8205 11268 8217 11271
rect 7892 11240 8217 11268
rect 7892 11228 7898 11240
rect 8205 11237 8217 11240
rect 8251 11268 8263 11271
rect 8570 11268 8576 11280
rect 8251 11240 8576 11268
rect 8251 11237 8263 11240
rect 8205 11231 8263 11237
rect 8570 11228 8576 11240
rect 8628 11228 8634 11280
rect 7282 11200 7288 11212
rect 7208 11172 7288 11200
rect 7208 11141 7236 11172
rect 7282 11160 7288 11172
rect 7340 11160 7346 11212
rect 7558 11160 7564 11212
rect 7616 11200 7622 11212
rect 8113 11203 8171 11209
rect 8113 11200 8125 11203
rect 7616 11172 8125 11200
rect 7616 11160 7622 11172
rect 8113 11169 8125 11172
rect 8159 11169 8171 11203
rect 8113 11163 8171 11169
rect 8294 11160 8300 11212
rect 8352 11200 8358 11212
rect 8662 11200 8668 11212
rect 8352 11172 8668 11200
rect 8352 11160 8358 11172
rect 7193 11135 7251 11141
rect 7064 11104 7157 11132
rect 7064 11092 7070 11104
rect 7193 11101 7205 11135
rect 7239 11101 7251 11135
rect 7411 11135 7469 11141
rect 7193 11095 7251 11101
rect 7286 11113 7344 11119
rect 7208 11064 7236 11095
rect 7286 11079 7298 11113
rect 7332 11079 7344 11113
rect 7411 11101 7423 11135
rect 7457 11132 7469 11135
rect 8018 11132 8024 11144
rect 7457 11104 8024 11132
rect 7457 11101 7469 11104
rect 7411 11095 7469 11101
rect 8018 11092 8024 11104
rect 8076 11132 8082 11144
rect 8404 11141 8432 11172
rect 8662 11160 8668 11172
rect 8720 11200 8726 11212
rect 9122 11200 9128 11212
rect 8720 11172 9128 11200
rect 8720 11160 8726 11172
rect 9122 11160 9128 11172
rect 9180 11160 9186 11212
rect 8389 11135 8447 11141
rect 8076 11104 8340 11132
rect 8076 11092 8082 11104
rect 7286 11076 7344 11079
rect 6932 11036 7236 11064
rect 7282 11024 7288 11076
rect 7340 11024 7346 11076
rect 7558 11024 7564 11076
rect 7616 11064 7622 11076
rect 8312 11064 8340 11104
rect 8389 11101 8401 11135
rect 8435 11101 8447 11135
rect 8389 11095 8447 11101
rect 8481 11135 8539 11141
rect 8481 11101 8493 11135
rect 8527 11132 8539 11135
rect 9030 11132 9036 11144
rect 8527 11104 9036 11132
rect 8527 11101 8539 11104
rect 8481 11095 8539 11101
rect 9030 11092 9036 11104
rect 9088 11132 9094 11144
rect 9232 11132 9260 11308
rect 9306 11296 9312 11308
rect 9364 11336 9370 11348
rect 9401 11339 9459 11345
rect 9401 11336 9413 11339
rect 9364 11308 9413 11336
rect 9364 11296 9370 11308
rect 9401 11305 9413 11308
rect 9447 11305 9459 11339
rect 9401 11299 9459 11305
rect 9766 11296 9772 11348
rect 9824 11336 9830 11348
rect 10137 11339 10195 11345
rect 10137 11336 10149 11339
rect 9824 11308 10149 11336
rect 9824 11296 9830 11308
rect 10137 11305 10149 11308
rect 10183 11305 10195 11339
rect 10137 11299 10195 11305
rect 10873 11339 10931 11345
rect 10873 11305 10885 11339
rect 10919 11336 10931 11339
rect 11238 11336 11244 11348
rect 10919 11308 11244 11336
rect 10919 11305 10931 11308
rect 10873 11299 10931 11305
rect 11238 11296 11244 11308
rect 11296 11296 11302 11348
rect 11974 11336 11980 11348
rect 11935 11308 11980 11336
rect 11974 11296 11980 11308
rect 12032 11296 12038 11348
rect 9861 11271 9919 11277
rect 9861 11237 9873 11271
rect 9907 11268 9919 11271
rect 10042 11268 10048 11280
rect 9907 11240 10048 11268
rect 9907 11237 9919 11240
rect 9861 11231 9919 11237
rect 10042 11228 10048 11240
rect 10100 11228 10106 11280
rect 10686 11228 10692 11280
rect 10744 11268 10750 11280
rect 10744 11240 11192 11268
rect 10744 11228 10750 11240
rect 9306 11160 9312 11212
rect 9364 11200 9370 11212
rect 11054 11200 11060 11212
rect 9364 11172 9409 11200
rect 9600 11172 10088 11200
rect 11015 11172 11060 11200
rect 9364 11160 9370 11172
rect 9600 11144 9628 11172
rect 10060 11144 10088 11172
rect 11054 11160 11060 11172
rect 11112 11160 11118 11212
rect 11164 11209 11192 11240
rect 11790 11228 11796 11280
rect 11848 11268 11854 11280
rect 13446 11268 13452 11280
rect 11848 11240 13452 11268
rect 11848 11228 11854 11240
rect 13446 11228 13452 11240
rect 13504 11228 13510 11280
rect 11149 11203 11207 11209
rect 11149 11169 11161 11203
rect 11195 11169 11207 11203
rect 13538 11200 13544 11212
rect 11149 11163 11207 11169
rect 11256 11172 13544 11200
rect 9582 11132 9588 11144
rect 9088 11104 9260 11132
rect 9543 11104 9588 11132
rect 9088 11092 9094 11104
rect 9582 11092 9588 11104
rect 9640 11092 9646 11144
rect 9674 11092 9680 11144
rect 9732 11132 9738 11144
rect 9732 11104 9777 11132
rect 9732 11092 9738 11104
rect 10042 11092 10048 11144
rect 10100 11092 10106 11144
rect 10318 11132 10324 11144
rect 10279 11104 10324 11132
rect 10318 11092 10324 11104
rect 10376 11092 10382 11144
rect 10594 11132 10600 11144
rect 10555 11104 10600 11132
rect 10594 11092 10600 11104
rect 10652 11092 10658 11144
rect 10694 11135 10752 11141
rect 10694 11101 10706 11135
rect 10740 11126 10752 11135
rect 11256 11132 11284 11172
rect 13538 11160 13544 11172
rect 13596 11160 13602 11212
rect 10888 11126 11284 11132
rect 10740 11104 11284 11126
rect 11379 11135 11437 11141
rect 10740 11101 10916 11104
rect 10694 11098 10916 11101
rect 11379 11101 11391 11135
rect 11425 11132 11437 11135
rect 11793 11135 11851 11141
rect 11425 11104 11560 11132
rect 11425 11101 11437 11104
rect 10694 11095 10752 11098
rect 11379 11095 11437 11101
rect 9950 11064 9956 11076
rect 7616 11036 8064 11064
rect 8312 11036 9956 11064
rect 7616 11024 7622 11036
rect 6052 10968 6683 10996
rect 6052 10956 6058 10968
rect 6730 10956 6736 11008
rect 6788 10996 6794 11008
rect 7837 10999 7895 11005
rect 7837 10996 7849 10999
rect 6788 10968 7849 10996
rect 6788 10956 6794 10968
rect 7837 10965 7849 10968
rect 7883 10996 7895 10999
rect 7926 10996 7932 11008
rect 7883 10968 7932 10996
rect 7883 10965 7895 10968
rect 7837 10959 7895 10965
rect 7926 10956 7932 10968
rect 7984 10956 7990 11008
rect 8036 10996 8064 11036
rect 9950 11024 9956 11036
rect 10008 11024 10014 11076
rect 10502 11064 10508 11076
rect 10463 11036 10508 11064
rect 10502 11024 10508 11036
rect 10560 11024 10566 11076
rect 10962 11024 10968 11076
rect 11020 11064 11026 11076
rect 11532 11064 11560 11104
rect 11793 11101 11805 11135
rect 11839 11132 11851 11135
rect 12066 11132 12072 11144
rect 11839 11104 12072 11132
rect 11839 11101 11851 11104
rect 11793 11095 11851 11101
rect 12066 11092 12072 11104
rect 12124 11092 12130 11144
rect 12986 11132 12992 11144
rect 12947 11104 12992 11132
rect 12986 11092 12992 11104
rect 13044 11092 13050 11144
rect 13262 11132 13268 11144
rect 13223 11104 13268 11132
rect 13262 11092 13268 11104
rect 13320 11092 13326 11144
rect 11020 11036 11560 11064
rect 11020 11024 11026 11036
rect 9030 10996 9036 11008
rect 8036 10968 9036 10996
rect 9030 10956 9036 10968
rect 9088 10996 9094 11008
rect 10686 10996 10692 11008
rect 9088 10968 10692 10996
rect 9088 10956 9094 10968
rect 10686 10956 10692 10968
rect 10744 10956 10750 11008
rect 11241 10999 11299 11005
rect 11241 10965 11253 10999
rect 11287 10996 11299 10999
rect 11330 10996 11336 11008
rect 11287 10968 11336 10996
rect 11287 10965 11299 10968
rect 11241 10959 11299 10965
rect 11330 10956 11336 10968
rect 11388 10956 11394 11008
rect 11532 10996 11560 11036
rect 11609 11067 11667 11073
rect 11609 11033 11621 11067
rect 11655 11064 11667 11067
rect 11974 11064 11980 11076
rect 11655 11036 11980 11064
rect 11655 11033 11667 11036
rect 11609 11027 11667 11033
rect 11974 11024 11980 11036
rect 12032 11064 12038 11076
rect 12250 11064 12256 11076
rect 12032 11036 12256 11064
rect 12032 11024 12038 11036
rect 12250 11024 12256 11036
rect 12308 11024 12314 11076
rect 12805 11067 12863 11073
rect 12805 11033 12817 11067
rect 12851 11064 12863 11067
rect 13078 11064 13084 11076
rect 12851 11036 13084 11064
rect 12851 11033 12863 11036
rect 12805 11027 12863 11033
rect 13078 11024 13084 11036
rect 13136 11024 13142 11076
rect 12526 10996 12532 11008
rect 11532 10968 12532 10996
rect 12526 10956 12532 10968
rect 12584 10956 12590 11008
rect 12710 10956 12716 11008
rect 12768 10996 12774 11008
rect 13173 10999 13231 11005
rect 13173 10996 13185 10999
rect 12768 10968 13185 10996
rect 12768 10956 12774 10968
rect 13173 10965 13185 10968
rect 13219 10965 13231 10999
rect 13173 10959 13231 10965
rect 1104 10906 13892 10928
rect 1104 10854 8214 10906
rect 8266 10854 8278 10906
rect 8330 10854 8342 10906
rect 8394 10854 8406 10906
rect 8458 10854 8470 10906
rect 8522 10854 13892 10906
rect 1104 10832 13892 10854
rect 2406 10792 2412 10804
rect 2367 10764 2412 10792
rect 2406 10752 2412 10764
rect 2464 10752 2470 10804
rect 2774 10752 2780 10804
rect 2832 10792 2838 10804
rect 3697 10795 3755 10801
rect 2832 10764 2912 10792
rect 2832 10752 2838 10764
rect 2682 10724 2688 10736
rect 2056 10696 2688 10724
rect 1578 10616 1584 10668
rect 1636 10665 1642 10668
rect 2056 10665 2084 10696
rect 2682 10684 2688 10696
rect 2740 10684 2746 10736
rect 2884 10733 2912 10764
rect 3697 10761 3709 10795
rect 3743 10792 3755 10795
rect 4522 10792 4528 10804
rect 3743 10764 4528 10792
rect 3743 10761 3755 10764
rect 3697 10755 3755 10761
rect 4522 10752 4528 10764
rect 4580 10752 4586 10804
rect 4706 10752 4712 10804
rect 4764 10792 4770 10804
rect 5353 10795 5411 10801
rect 5353 10792 5365 10795
rect 4764 10764 5365 10792
rect 4764 10752 4770 10764
rect 5353 10761 5365 10764
rect 5399 10761 5411 10795
rect 5810 10792 5816 10804
rect 5771 10764 5816 10792
rect 5353 10755 5411 10761
rect 5810 10752 5816 10764
rect 5868 10752 5874 10804
rect 5902 10752 5908 10804
rect 5960 10792 5966 10804
rect 5997 10795 6055 10801
rect 5997 10792 6009 10795
rect 5960 10764 6009 10792
rect 5960 10752 5966 10764
rect 5997 10761 6009 10764
rect 6043 10761 6055 10795
rect 5997 10755 6055 10761
rect 6270 10752 6276 10804
rect 6328 10792 6334 10804
rect 6328 10764 8064 10792
rect 6328 10752 6334 10764
rect 2869 10727 2927 10733
rect 2869 10693 2881 10727
rect 2915 10693 2927 10727
rect 3326 10724 3332 10736
rect 3287 10696 3332 10724
rect 2869 10687 2927 10693
rect 3326 10684 3332 10696
rect 3384 10684 3390 10736
rect 3602 10684 3608 10736
rect 3660 10724 3666 10736
rect 3789 10727 3847 10733
rect 3789 10724 3801 10727
rect 3660 10696 3801 10724
rect 3660 10684 3666 10696
rect 3789 10693 3801 10696
rect 3835 10693 3847 10727
rect 3789 10687 3847 10693
rect 3973 10727 4031 10733
rect 3973 10693 3985 10727
rect 4019 10724 4031 10727
rect 4341 10727 4399 10733
rect 4341 10724 4353 10727
rect 4019 10696 4353 10724
rect 4019 10693 4031 10696
rect 3973 10687 4031 10693
rect 4341 10693 4353 10696
rect 4387 10724 4399 10727
rect 4614 10724 4620 10736
rect 4387 10696 4620 10724
rect 4387 10693 4399 10696
rect 4341 10687 4399 10693
rect 4614 10684 4620 10696
rect 4672 10684 4678 10736
rect 6181 10727 6239 10733
rect 6181 10693 6193 10727
rect 6227 10724 6239 10727
rect 6454 10724 6460 10736
rect 6227 10696 6460 10724
rect 6227 10693 6239 10696
rect 6181 10687 6239 10693
rect 6454 10684 6460 10696
rect 6512 10684 6518 10736
rect 7006 10724 7012 10736
rect 6967 10696 7012 10724
rect 7006 10684 7012 10696
rect 7064 10684 7070 10736
rect 7374 10724 7380 10736
rect 7335 10696 7380 10724
rect 7374 10684 7380 10696
rect 7432 10684 7438 10736
rect 7926 10724 7932 10736
rect 7887 10696 7932 10724
rect 7926 10684 7932 10696
rect 7984 10684 7990 10736
rect 8036 10733 8064 10764
rect 8386 10752 8392 10804
rect 8444 10752 8450 10804
rect 8665 10795 8723 10801
rect 8665 10761 8677 10795
rect 8711 10792 8723 10795
rect 8938 10792 8944 10804
rect 8711 10764 8944 10792
rect 8711 10761 8723 10764
rect 8665 10755 8723 10761
rect 8938 10752 8944 10764
rect 8996 10752 9002 10804
rect 9401 10795 9459 10801
rect 9401 10792 9413 10795
rect 9048 10764 9413 10792
rect 8021 10727 8079 10733
rect 8021 10693 8033 10727
rect 8067 10693 8079 10727
rect 8021 10687 8079 10693
rect 1636 10659 1679 10665
rect 1667 10625 1679 10659
rect 1636 10619 1679 10625
rect 1765 10659 1823 10665
rect 1765 10625 1777 10659
rect 1811 10625 1823 10659
rect 1765 10619 1823 10625
rect 1857 10659 1915 10665
rect 1857 10625 1869 10659
rect 1903 10625 1915 10659
rect 1857 10619 1915 10625
rect 2041 10659 2099 10665
rect 2041 10625 2053 10659
rect 2087 10625 2099 10659
rect 2041 10619 2099 10625
rect 2501 10659 2559 10665
rect 2501 10625 2513 10659
rect 2547 10656 2559 10659
rect 2774 10656 2780 10668
rect 2547 10628 2780 10656
rect 2547 10625 2559 10628
rect 2501 10619 2559 10625
rect 1636 10616 1642 10619
rect 1394 10480 1400 10532
rect 1452 10520 1458 10532
rect 1780 10520 1808 10619
rect 1872 10588 1900 10619
rect 2774 10616 2780 10628
rect 2832 10616 2838 10668
rect 2961 10659 3019 10665
rect 2961 10625 2973 10659
rect 3007 10625 3019 10659
rect 2961 10619 3019 10625
rect 3145 10659 3203 10665
rect 3145 10625 3157 10659
rect 3191 10625 3203 10659
rect 3145 10619 3203 10625
rect 2682 10588 2688 10600
rect 1872 10560 2688 10588
rect 2682 10548 2688 10560
rect 2740 10548 2746 10600
rect 2976 10520 3004 10619
rect 1452 10492 3004 10520
rect 3160 10520 3188 10619
rect 3878 10616 3884 10668
rect 3936 10656 3942 10668
rect 4065 10659 4123 10665
rect 4065 10656 4077 10659
rect 3936 10628 4077 10656
rect 3936 10616 3942 10628
rect 4065 10625 4077 10628
rect 4111 10625 4123 10659
rect 4982 10656 4988 10668
rect 4943 10628 4988 10656
rect 4065 10619 4123 10625
rect 4080 10588 4108 10619
rect 4982 10616 4988 10628
rect 5040 10616 5046 10668
rect 5258 10656 5264 10668
rect 5219 10628 5264 10656
rect 5258 10616 5264 10628
rect 5316 10616 5322 10668
rect 5537 10659 5595 10665
rect 5537 10625 5549 10659
rect 5583 10625 5595 10659
rect 5537 10619 5595 10625
rect 5552 10588 5580 10619
rect 6730 10616 6736 10668
rect 6788 10656 6794 10668
rect 6917 10659 6975 10665
rect 6917 10656 6929 10659
rect 6788 10628 6929 10656
rect 6788 10616 6794 10628
rect 6917 10625 6929 10628
rect 6963 10625 6975 10659
rect 6917 10619 6975 10625
rect 7193 10659 7251 10665
rect 7193 10625 7205 10659
rect 7239 10656 7251 10659
rect 7650 10656 7656 10668
rect 7239 10628 7656 10656
rect 7239 10625 7251 10628
rect 7193 10619 7251 10625
rect 7650 10616 7656 10628
rect 7708 10616 7714 10668
rect 7834 10665 7840 10668
rect 7832 10656 7840 10665
rect 7795 10628 7840 10656
rect 7832 10619 7840 10628
rect 7834 10616 7840 10619
rect 7892 10616 7898 10668
rect 8202 10656 8208 10668
rect 8163 10628 8208 10656
rect 8202 10616 8208 10628
rect 8260 10616 8266 10668
rect 8404 10665 8432 10752
rect 8754 10684 8760 10736
rect 8812 10724 8818 10736
rect 9048 10724 9076 10764
rect 9401 10761 9413 10764
rect 9447 10761 9459 10795
rect 9401 10755 9459 10761
rect 9508 10764 10088 10792
rect 8812 10696 9076 10724
rect 8812 10684 8818 10696
rect 9214 10684 9220 10736
rect 9272 10724 9278 10736
rect 9508 10724 9536 10764
rect 9272 10696 9536 10724
rect 9272 10684 9278 10696
rect 9674 10684 9680 10736
rect 9732 10724 9738 10736
rect 9953 10727 10011 10733
rect 9953 10724 9965 10727
rect 9732 10696 9965 10724
rect 9732 10684 9738 10696
rect 9953 10693 9965 10696
rect 9999 10693 10011 10727
rect 10060 10724 10088 10764
rect 10318 10752 10324 10804
rect 10376 10792 10382 10804
rect 10413 10795 10471 10801
rect 10413 10792 10425 10795
rect 10376 10764 10425 10792
rect 10376 10752 10382 10764
rect 10413 10761 10425 10764
rect 10459 10761 10471 10795
rect 11592 10795 11650 10801
rect 11592 10792 11604 10795
rect 10413 10755 10471 10761
rect 10520 10764 11604 10792
rect 10520 10724 10548 10764
rect 11592 10761 11604 10764
rect 11638 10761 11650 10795
rect 11592 10755 11650 10761
rect 11716 10764 13492 10792
rect 10060 10696 10548 10724
rect 9953 10687 10011 10693
rect 8297 10659 8355 10665
rect 8297 10625 8309 10659
rect 8343 10625 8355 10659
rect 8297 10619 8355 10625
rect 8389 10659 8447 10665
rect 8389 10625 8401 10659
rect 8435 10625 8447 10659
rect 9122 10656 9128 10668
rect 9083 10628 9128 10656
rect 8389 10619 8447 10625
rect 4080 10560 5580 10588
rect 5902 10548 5908 10600
rect 5960 10588 5966 10600
rect 6822 10588 6828 10600
rect 5960 10560 6592 10588
rect 5960 10548 5966 10560
rect 6270 10520 6276 10532
rect 3160 10492 6276 10520
rect 1452 10480 1458 10492
rect 1486 10452 1492 10464
rect 1447 10424 1492 10452
rect 1486 10412 1492 10424
rect 1544 10412 1550 10464
rect 2130 10452 2136 10464
rect 2091 10424 2136 10452
rect 2130 10412 2136 10424
rect 2188 10412 2194 10464
rect 2777 10455 2835 10461
rect 2777 10421 2789 10455
rect 2823 10452 2835 10455
rect 2976 10452 3004 10492
rect 6270 10480 6276 10492
rect 6328 10480 6334 10532
rect 3142 10452 3148 10464
rect 2823 10424 3148 10452
rect 2823 10421 2835 10424
rect 2777 10415 2835 10421
rect 3142 10412 3148 10424
rect 3200 10412 3206 10464
rect 4614 10412 4620 10464
rect 4672 10452 4678 10464
rect 5169 10455 5227 10461
rect 5169 10452 5181 10455
rect 4672 10424 5181 10452
rect 4672 10412 4678 10424
rect 5169 10421 5181 10424
rect 5215 10421 5227 10455
rect 5169 10415 5227 10421
rect 5350 10412 5356 10464
rect 5408 10452 5414 10464
rect 5994 10452 6000 10464
rect 5408 10424 6000 10452
rect 5408 10412 5414 10424
rect 5994 10412 6000 10424
rect 6052 10412 6058 10464
rect 6178 10412 6184 10464
rect 6236 10452 6242 10464
rect 6457 10455 6515 10461
rect 6457 10452 6469 10455
rect 6236 10424 6469 10452
rect 6236 10412 6242 10424
rect 6457 10421 6469 10424
rect 6503 10421 6515 10455
rect 6564 10452 6592 10560
rect 6656 10560 6828 10588
rect 6656 10529 6684 10560
rect 6822 10548 6828 10560
rect 6880 10588 6886 10600
rect 7098 10588 7104 10600
rect 6880 10560 7104 10588
rect 6880 10548 6886 10560
rect 7098 10548 7104 10560
rect 7156 10588 7162 10600
rect 7282 10588 7288 10600
rect 7156 10560 7288 10588
rect 7156 10548 7162 10560
rect 7282 10548 7288 10560
rect 7340 10588 7346 10600
rect 8307 10588 8335 10619
rect 9122 10616 9128 10628
rect 9180 10616 9186 10668
rect 9309 10659 9367 10665
rect 9309 10625 9321 10659
rect 9355 10656 9367 10659
rect 9398 10656 9404 10668
rect 9355 10628 9404 10656
rect 9355 10625 9367 10628
rect 9309 10619 9367 10625
rect 9398 10616 9404 10628
rect 9456 10616 9462 10668
rect 9582 10656 9588 10668
rect 9543 10628 9588 10656
rect 9582 10616 9588 10628
rect 9640 10616 9646 10668
rect 9769 10659 9827 10665
rect 9769 10625 9781 10659
rect 9815 10625 9827 10659
rect 9968 10656 9996 10687
rect 10686 10684 10692 10736
rect 10744 10724 10750 10736
rect 10781 10727 10839 10733
rect 10781 10724 10793 10727
rect 10744 10696 10793 10724
rect 10744 10684 10750 10696
rect 10781 10693 10793 10696
rect 10827 10693 10839 10727
rect 10781 10687 10839 10693
rect 11241 10727 11299 10733
rect 11241 10693 11253 10727
rect 11287 10724 11299 10727
rect 11716 10724 11744 10764
rect 12250 10724 12256 10736
rect 11287 10696 11744 10724
rect 11900 10696 12256 10724
rect 11287 10693 11299 10696
rect 11241 10687 11299 10693
rect 10045 10659 10103 10665
rect 10045 10656 10057 10659
rect 9968 10628 10057 10656
rect 9769 10619 9827 10625
rect 10045 10625 10057 10628
rect 10091 10656 10103 10659
rect 10597 10659 10655 10665
rect 10597 10656 10609 10659
rect 10091 10628 10609 10656
rect 10091 10625 10103 10628
rect 10045 10619 10103 10625
rect 10597 10625 10609 10628
rect 10643 10625 10655 10659
rect 11330 10656 11336 10668
rect 11291 10628 11336 10656
rect 10597 10619 10655 10625
rect 8938 10588 8944 10600
rect 7340 10560 8335 10588
rect 8899 10560 8944 10588
rect 7340 10548 7346 10560
rect 8938 10548 8944 10560
rect 8996 10548 9002 10600
rect 6641 10523 6699 10529
rect 6641 10489 6653 10523
rect 6687 10489 6699 10523
rect 6641 10483 6699 10489
rect 7374 10480 7380 10532
rect 7432 10520 7438 10532
rect 8386 10520 8392 10532
rect 7432 10492 8392 10520
rect 7432 10480 7438 10492
rect 8386 10480 8392 10492
rect 8444 10480 8450 10532
rect 8570 10480 8576 10532
rect 8628 10520 8634 10532
rect 9784 10520 9812 10619
rect 11330 10616 11336 10628
rect 11388 10616 11394 10668
rect 11790 10665 11796 10668
rect 11788 10656 11796 10665
rect 11751 10628 11796 10656
rect 11788 10619 11796 10628
rect 11790 10616 11796 10619
rect 11848 10616 11854 10668
rect 11900 10665 11928 10696
rect 12250 10684 12256 10696
rect 12308 10684 12314 10736
rect 13464 10733 13492 10764
rect 13449 10727 13507 10733
rect 13449 10693 13461 10727
rect 13495 10693 13507 10727
rect 13449 10687 13507 10693
rect 11885 10659 11943 10665
rect 11885 10625 11897 10659
rect 11931 10625 11943 10659
rect 11885 10619 11943 10625
rect 11977 10659 12035 10665
rect 11977 10625 11989 10659
rect 12023 10625 12035 10659
rect 12158 10656 12164 10668
rect 12119 10628 12164 10656
rect 11977 10619 12035 10625
rect 9858 10548 9864 10600
rect 9916 10588 9922 10600
rect 10137 10591 10195 10597
rect 10137 10588 10149 10591
rect 9916 10560 10149 10588
rect 9916 10548 9922 10560
rect 10137 10557 10149 10560
rect 10183 10588 10195 10591
rect 11238 10588 11244 10600
rect 10183 10560 11244 10588
rect 10183 10557 10195 10560
rect 10137 10551 10195 10557
rect 11238 10548 11244 10560
rect 11296 10548 11302 10600
rect 11992 10520 12020 10619
rect 12158 10616 12164 10628
rect 12216 10616 12222 10668
rect 12618 10616 12624 10668
rect 12676 10656 12682 10668
rect 12713 10659 12771 10665
rect 12713 10656 12725 10659
rect 12676 10628 12725 10656
rect 12676 10616 12682 10628
rect 12713 10625 12725 10628
rect 12759 10625 12771 10659
rect 12713 10619 12771 10625
rect 12066 10548 12072 10600
rect 12124 10588 12130 10600
rect 12253 10591 12311 10597
rect 12253 10588 12265 10591
rect 12124 10560 12265 10588
rect 12124 10548 12130 10560
rect 12253 10557 12265 10560
rect 12299 10557 12311 10591
rect 12253 10551 12311 10557
rect 12342 10548 12348 10600
rect 12400 10588 12406 10600
rect 12805 10591 12863 10597
rect 12805 10588 12817 10591
rect 12400 10560 12817 10588
rect 12400 10548 12406 10560
rect 12805 10557 12817 10560
rect 12851 10557 12863 10591
rect 12805 10551 12863 10557
rect 12894 10548 12900 10600
rect 12952 10588 12958 10600
rect 12952 10560 12997 10588
rect 12952 10548 12958 10560
rect 13354 10520 13360 10532
rect 8628 10492 10640 10520
rect 8628 10480 8634 10492
rect 10612 10464 10640 10492
rect 11716 10492 12020 10520
rect 13315 10492 13360 10520
rect 11716 10464 11744 10492
rect 13354 10480 13360 10492
rect 13412 10480 13418 10532
rect 7653 10455 7711 10461
rect 7653 10452 7665 10455
rect 6564 10424 7665 10452
rect 6457 10415 6515 10421
rect 7653 10421 7665 10424
rect 7699 10421 7711 10455
rect 7653 10415 7711 10421
rect 8481 10455 8539 10461
rect 8481 10421 8493 10455
rect 8527 10452 8539 10455
rect 9950 10452 9956 10464
rect 8527 10424 9956 10452
rect 8527 10421 8539 10424
rect 8481 10415 8539 10421
rect 9950 10412 9956 10424
rect 10008 10452 10014 10464
rect 10045 10455 10103 10461
rect 10045 10452 10057 10455
rect 10008 10424 10057 10452
rect 10008 10412 10014 10424
rect 10045 10421 10057 10424
rect 10091 10421 10103 10455
rect 10045 10415 10103 10421
rect 10594 10412 10600 10464
rect 10652 10412 10658 10464
rect 10870 10452 10876 10464
rect 10831 10424 10876 10452
rect 10870 10412 10876 10424
rect 10928 10412 10934 10464
rect 11698 10412 11704 10464
rect 11756 10412 11762 10464
rect 11974 10412 11980 10464
rect 12032 10452 12038 10464
rect 12250 10452 12256 10464
rect 12032 10424 12256 10452
rect 12032 10412 12038 10424
rect 12250 10412 12256 10424
rect 12308 10412 12314 10464
rect 1104 10362 13892 10384
rect 1104 10310 4214 10362
rect 4266 10310 4278 10362
rect 4330 10310 4342 10362
rect 4394 10310 4406 10362
rect 4458 10310 4470 10362
rect 4522 10310 12214 10362
rect 12266 10310 12278 10362
rect 12330 10310 12342 10362
rect 12394 10310 12406 10362
rect 12458 10310 12470 10362
rect 12522 10310 13892 10362
rect 1104 10288 13892 10310
rect 1394 10248 1400 10260
rect 1355 10220 1400 10248
rect 1394 10208 1400 10220
rect 1452 10208 1458 10260
rect 1673 10251 1731 10257
rect 1673 10217 1685 10251
rect 1719 10248 1731 10251
rect 2866 10248 2872 10260
rect 1719 10220 2872 10248
rect 1719 10217 1731 10220
rect 1673 10211 1731 10217
rect 2866 10208 2872 10220
rect 2924 10208 2930 10260
rect 3326 10208 3332 10260
rect 3384 10248 3390 10260
rect 5810 10248 5816 10260
rect 3384 10220 5816 10248
rect 3384 10208 3390 10220
rect 5810 10208 5816 10220
rect 5868 10208 5874 10260
rect 7101 10251 7159 10257
rect 7101 10217 7113 10251
rect 7147 10248 7159 10251
rect 7190 10248 7196 10260
rect 7147 10220 7196 10248
rect 7147 10217 7159 10220
rect 7101 10211 7159 10217
rect 7190 10208 7196 10220
rect 7248 10208 7254 10260
rect 8478 10208 8484 10260
rect 8536 10248 8542 10260
rect 8665 10251 8723 10257
rect 8665 10248 8677 10251
rect 8536 10220 8677 10248
rect 8536 10208 8542 10220
rect 8665 10217 8677 10220
rect 8711 10217 8723 10251
rect 8665 10211 8723 10217
rect 9401 10251 9459 10257
rect 9401 10217 9413 10251
rect 9447 10248 9459 10251
rect 9490 10248 9496 10260
rect 9447 10220 9496 10248
rect 9447 10217 9459 10220
rect 9401 10211 9459 10217
rect 9490 10208 9496 10220
rect 9548 10208 9554 10260
rect 10962 10248 10968 10260
rect 9691 10220 10968 10248
rect 2148 10152 2636 10180
rect 1486 10072 1492 10124
rect 1544 10112 1550 10124
rect 1765 10115 1823 10121
rect 1765 10112 1777 10115
rect 1544 10084 1777 10112
rect 1544 10072 1550 10084
rect 1765 10081 1777 10084
rect 1811 10081 1823 10115
rect 1765 10075 1823 10081
rect 2148 10044 2176 10152
rect 2608 10112 2636 10152
rect 2682 10140 2688 10192
rect 2740 10180 2746 10192
rect 8202 10180 8208 10192
rect 2740 10152 4752 10180
rect 2740 10140 2746 10152
rect 3881 10115 3939 10121
rect 3881 10112 3893 10115
rect 2608 10084 3893 10112
rect 3881 10081 3893 10084
rect 3927 10081 3939 10115
rect 4614 10112 4620 10124
rect 4575 10084 4620 10112
rect 3881 10075 3939 10081
rect 4614 10072 4620 10084
rect 4672 10072 4678 10124
rect 2317 10047 2375 10053
rect 2317 10044 2329 10047
rect 2148 10016 2329 10044
rect 2317 10013 2329 10016
rect 2363 10013 2375 10047
rect 2317 10007 2375 10013
rect 2406 10004 2412 10056
rect 2464 10044 2470 10056
rect 2866 10044 2872 10056
rect 2464 10016 2509 10044
rect 2779 10016 2872 10044
rect 2464 10004 2470 10016
rect 2866 10004 2872 10016
rect 2924 10044 2930 10056
rect 2924 10016 3280 10044
rect 2924 10004 2930 10016
rect 2225 9979 2283 9985
rect 2225 9945 2237 9979
rect 2271 9976 2283 9979
rect 2774 9976 2780 9988
rect 2271 9948 2780 9976
rect 2271 9945 2283 9948
rect 2225 9939 2283 9945
rect 2774 9936 2780 9948
rect 2832 9936 2838 9988
rect 2958 9976 2964 9988
rect 2919 9948 2964 9976
rect 2958 9936 2964 9948
rect 3016 9936 3022 9988
rect 3057 9979 3115 9985
rect 3057 9945 3069 9979
rect 3103 9945 3115 9979
rect 3252 9976 3280 10016
rect 3326 10004 3332 10056
rect 3384 10044 3390 10056
rect 3513 10047 3571 10053
rect 3384 10016 3429 10044
rect 3384 10004 3390 10016
rect 3513 10013 3525 10047
rect 3559 10044 3571 10047
rect 3694 10044 3700 10056
rect 3559 10016 3700 10044
rect 3559 10013 3571 10016
rect 3513 10007 3571 10013
rect 3694 10004 3700 10016
rect 3752 10044 3758 10056
rect 4065 10047 4123 10053
rect 4065 10044 4077 10047
rect 3752 10016 4077 10044
rect 3752 10004 3758 10016
rect 4065 10013 4077 10016
rect 4111 10013 4123 10047
rect 4724 10044 4752 10152
rect 7668 10152 8064 10180
rect 8163 10152 8208 10180
rect 7668 10124 7696 10152
rect 4801 10115 4859 10121
rect 4801 10081 4813 10115
rect 4847 10112 4859 10115
rect 6733 10115 6791 10121
rect 4847 10084 5948 10112
rect 4847 10081 4859 10084
rect 4801 10075 4859 10081
rect 5350 10044 5356 10056
rect 4724 10016 5356 10044
rect 4065 10007 4123 10013
rect 5350 10004 5356 10016
rect 5408 10004 5414 10056
rect 5534 10044 5540 10056
rect 5495 10016 5540 10044
rect 5534 10004 5540 10016
rect 5592 10004 5598 10056
rect 5721 10047 5779 10053
rect 5721 10013 5733 10047
rect 5767 10044 5779 10047
rect 5813 10047 5871 10053
rect 5813 10044 5825 10047
rect 5767 10016 5825 10044
rect 5767 10013 5779 10016
rect 5721 10007 5779 10013
rect 5813 10013 5825 10016
rect 5859 10013 5871 10047
rect 5920 10044 5948 10084
rect 6733 10081 6745 10115
rect 6779 10112 6791 10115
rect 7650 10112 7656 10124
rect 6779 10084 7656 10112
rect 6779 10081 6791 10084
rect 6733 10075 6791 10081
rect 7650 10072 7656 10084
rect 7708 10072 7714 10124
rect 7834 10072 7840 10124
rect 7892 10072 7898 10124
rect 8036 10112 8064 10152
rect 8202 10140 8208 10152
rect 8260 10140 8266 10192
rect 8478 10112 8484 10124
rect 8036 10084 8484 10112
rect 8478 10072 8484 10084
rect 8536 10072 8542 10124
rect 8938 10112 8944 10124
rect 8772 10084 8944 10112
rect 6233 10047 6291 10053
rect 6233 10044 6245 10047
rect 5920 10016 6245 10044
rect 5813 10007 5871 10013
rect 6233 10013 6245 10016
rect 6279 10044 6291 10047
rect 6362 10044 6368 10056
rect 6279 10016 6368 10044
rect 6279 10013 6291 10016
rect 6233 10007 6291 10013
rect 6362 10004 6368 10016
rect 6420 10004 6426 10056
rect 6638 10044 6644 10056
rect 6599 10016 6644 10044
rect 6638 10004 6644 10016
rect 6696 10004 6702 10056
rect 6822 10044 6828 10056
rect 6783 10016 6828 10044
rect 6822 10004 6828 10016
rect 6880 10004 6886 10056
rect 6917 10047 6975 10053
rect 6917 10013 6929 10047
rect 6963 10044 6975 10047
rect 7098 10044 7104 10056
rect 6963 10016 7104 10044
rect 6963 10013 6975 10016
rect 6917 10007 6975 10013
rect 3789 9979 3847 9985
rect 3789 9976 3801 9979
rect 3252 9948 3801 9976
rect 3057 9939 3115 9945
rect 3789 9945 3801 9948
rect 3835 9945 3847 9979
rect 4522 9976 4528 9988
rect 4483 9948 4528 9976
rect 3789 9939 3847 9945
rect 2130 9868 2136 9920
rect 2188 9908 2194 9920
rect 3068 9908 3096 9939
rect 4522 9936 4528 9948
rect 4580 9936 4586 9988
rect 4982 9976 4988 9988
rect 4943 9948 4988 9976
rect 4982 9936 4988 9948
rect 5040 9936 5046 9988
rect 5166 9976 5172 9988
rect 5127 9948 5172 9976
rect 5166 9936 5172 9948
rect 5224 9936 5230 9988
rect 5997 9979 6055 9985
rect 5997 9945 6009 9979
rect 6043 9945 6055 9979
rect 5997 9939 6055 9945
rect 6089 9979 6147 9985
rect 6089 9945 6101 9979
rect 6135 9976 6147 9979
rect 6730 9976 6736 9988
rect 6135 9948 6736 9976
rect 6135 9945 6147 9948
rect 6089 9939 6147 9945
rect 2188 9880 3096 9908
rect 2188 9868 2194 9880
rect 3142 9868 3148 9920
rect 3200 9908 3206 9920
rect 3970 9908 3976 9920
rect 3200 9880 3976 9908
rect 3200 9868 3206 9880
rect 3970 9868 3976 9880
rect 4028 9868 4034 9920
rect 6012 9908 6040 9939
rect 6730 9936 6736 9948
rect 6788 9976 6794 9988
rect 6932 9976 6960 10007
rect 7098 10004 7104 10016
rect 7156 10044 7162 10056
rect 7377 10047 7435 10053
rect 7377 10044 7389 10047
rect 7156 10016 7389 10044
rect 7156 10004 7162 10016
rect 7377 10013 7389 10016
rect 7423 10013 7435 10047
rect 7558 10044 7564 10056
rect 7519 10016 7564 10044
rect 7377 10007 7435 10013
rect 7558 10004 7564 10016
rect 7616 10004 7622 10056
rect 7742 10044 7748 10056
rect 7703 10016 7748 10044
rect 7742 10004 7748 10016
rect 7800 10004 7806 10056
rect 7853 10031 7881 10072
rect 7963 10047 8021 10053
rect 7838 10025 7896 10031
rect 7838 9991 7850 10025
rect 7884 9991 7896 10025
rect 7963 10013 7975 10047
rect 8009 10013 8021 10047
rect 8570 10044 8576 10056
rect 8531 10016 8576 10044
rect 7963 10007 8021 10013
rect 7838 9985 7896 9991
rect 6788 9948 6960 9976
rect 7978 9976 8006 10007
rect 8570 10004 8576 10016
rect 8628 10004 8634 10056
rect 8772 10053 8800 10084
rect 8938 10072 8944 10084
rect 8996 10112 9002 10124
rect 9691 10112 9719 10220
rect 10962 10208 10968 10220
rect 11020 10208 11026 10260
rect 9858 10180 9864 10192
rect 9819 10152 9864 10180
rect 9858 10140 9864 10152
rect 9916 10140 9922 10192
rect 11054 10140 11060 10192
rect 11112 10180 11118 10192
rect 12894 10180 12900 10192
rect 11112 10152 12900 10180
rect 11112 10140 11118 10152
rect 8996 10084 9719 10112
rect 8996 10072 9002 10084
rect 9766 10072 9772 10124
rect 9824 10112 9830 10124
rect 10209 10115 10267 10121
rect 10209 10112 10221 10115
rect 9824 10084 10221 10112
rect 9824 10072 9830 10084
rect 10209 10081 10221 10084
rect 10255 10081 10267 10115
rect 10209 10075 10267 10081
rect 10410 10072 10416 10124
rect 10468 10072 10474 10124
rect 10505 10115 10563 10121
rect 10505 10081 10517 10115
rect 10551 10112 10563 10115
rect 10686 10112 10692 10124
rect 10551 10084 10692 10112
rect 10551 10081 10563 10084
rect 10505 10075 10563 10081
rect 10686 10072 10692 10084
rect 10744 10072 10750 10124
rect 10965 10115 11023 10121
rect 10965 10112 10977 10115
rect 10888 10084 10977 10112
rect 8757 10047 8815 10053
rect 8757 10013 8769 10047
rect 8803 10013 8815 10047
rect 8757 10007 8815 10013
rect 9217 10047 9275 10053
rect 9217 10013 9229 10047
rect 9263 10013 9275 10047
rect 9217 10007 9275 10013
rect 9401 10047 9459 10053
rect 9401 10013 9413 10047
rect 9447 10013 9459 10047
rect 9401 10007 9459 10013
rect 9493 10047 9551 10053
rect 9493 10013 9505 10047
rect 9539 10044 9551 10047
rect 9582 10044 9588 10056
rect 9539 10016 9588 10044
rect 9539 10013 9551 10016
rect 9493 10007 9551 10013
rect 9232 9976 9260 10007
rect 9416 9976 9444 10007
rect 9582 10004 9588 10016
rect 9640 10044 9646 10056
rect 10428 10044 10456 10072
rect 10594 10044 10600 10056
rect 9640 10016 10456 10044
rect 10555 10016 10600 10044
rect 9640 10004 9646 10016
rect 10594 10004 10600 10016
rect 10652 10004 10658 10056
rect 10778 10044 10784 10056
rect 10739 10016 10784 10044
rect 10778 10004 10784 10016
rect 10836 10004 10842 10056
rect 9766 9976 9772 9988
rect 7978 9948 9352 9976
rect 9416 9948 9772 9976
rect 6788 9936 6794 9948
rect 6178 9908 6184 9920
rect 6012 9880 6184 9908
rect 6178 9868 6184 9880
rect 6236 9868 6242 9920
rect 6382 9911 6440 9917
rect 6382 9877 6394 9911
rect 6428 9908 6440 9911
rect 7190 9908 7196 9920
rect 6428 9880 7196 9908
rect 6428 9877 6440 9880
rect 6382 9871 6440 9877
rect 7190 9868 7196 9880
rect 7248 9868 7254 9920
rect 7834 9868 7840 9920
rect 7892 9908 7898 9920
rect 7978 9908 8006 9948
rect 9324 9920 9352 9948
rect 9766 9936 9772 9948
rect 9824 9936 9830 9988
rect 9953 9979 10011 9985
rect 9953 9945 9965 9979
rect 9999 9976 10011 9979
rect 10134 9976 10140 9988
rect 9999 9948 10140 9976
rect 9999 9945 10011 9948
rect 9953 9939 10011 9945
rect 10134 9936 10140 9948
rect 10192 9936 10198 9988
rect 10318 9985 10324 9988
rect 10297 9979 10324 9985
rect 10297 9945 10309 9979
rect 10297 9939 10324 9945
rect 10318 9936 10324 9939
rect 10376 9936 10382 9988
rect 10413 9979 10471 9985
rect 10413 9945 10425 9979
rect 10459 9976 10471 9979
rect 10888 9976 10916 10084
rect 10965 10081 10977 10084
rect 11011 10112 11023 10115
rect 11790 10112 11796 10124
rect 11011 10084 11796 10112
rect 11011 10081 11023 10084
rect 10965 10075 11023 10081
rect 11790 10072 11796 10084
rect 11848 10072 11854 10124
rect 11054 10044 11060 10056
rect 11015 10016 11060 10044
rect 11054 10004 11060 10016
rect 11112 10004 11118 10056
rect 11146 10004 11152 10056
rect 11204 10044 11210 10056
rect 11900 10053 11928 10152
rect 12894 10140 12900 10152
rect 12952 10140 12958 10192
rect 13354 10180 13360 10192
rect 13315 10152 13360 10180
rect 13354 10140 13360 10152
rect 13412 10140 13418 10192
rect 11333 10047 11391 10053
rect 11333 10044 11345 10047
rect 11204 10016 11345 10044
rect 11204 10004 11210 10016
rect 11333 10013 11345 10016
rect 11379 10044 11391 10047
rect 11701 10047 11759 10053
rect 11701 10044 11713 10047
rect 11379 10016 11713 10044
rect 11379 10013 11391 10016
rect 11333 10007 11391 10013
rect 11701 10013 11713 10016
rect 11747 10044 11759 10047
rect 11885 10047 11943 10053
rect 11747 10016 11836 10044
rect 11747 10013 11759 10016
rect 11701 10007 11759 10013
rect 11808 9988 11836 10016
rect 11885 10013 11897 10047
rect 11931 10013 11943 10047
rect 11885 10007 11943 10013
rect 12710 10004 12716 10056
rect 12768 10044 12774 10056
rect 12805 10047 12863 10053
rect 12805 10044 12817 10047
rect 12768 10016 12817 10044
rect 12768 10004 12774 10016
rect 12805 10013 12817 10016
rect 12851 10013 12863 10047
rect 12805 10007 12863 10013
rect 10459 9948 10916 9976
rect 10459 9945 10471 9948
rect 10413 9939 10471 9945
rect 11238 9936 11244 9988
rect 11296 9976 11302 9988
rect 11425 9979 11483 9985
rect 11425 9976 11437 9979
rect 11296 9948 11437 9976
rect 11296 9936 11302 9948
rect 11425 9945 11437 9948
rect 11471 9945 11483 9979
rect 11425 9939 11483 9945
rect 11790 9936 11796 9988
rect 11848 9936 11854 9988
rect 7892 9880 8006 9908
rect 7892 9868 7898 9880
rect 8386 9868 8392 9920
rect 8444 9908 8450 9920
rect 9033 9911 9091 9917
rect 9033 9908 9045 9911
rect 8444 9880 9045 9908
rect 8444 9868 8450 9880
rect 9033 9877 9045 9880
rect 9079 9877 9091 9911
rect 9033 9871 9091 9877
rect 9306 9868 9312 9920
rect 9364 9868 9370 9920
rect 9490 9868 9496 9920
rect 9548 9908 9554 9920
rect 9585 9911 9643 9917
rect 9585 9908 9597 9911
rect 9548 9880 9597 9908
rect 9548 9868 9554 9880
rect 9585 9877 9597 9880
rect 9631 9877 9643 9911
rect 9585 9871 9643 9877
rect 10594 9868 10600 9920
rect 10652 9908 10658 9920
rect 11609 9911 11667 9917
rect 11609 9908 11621 9911
rect 10652 9880 11621 9908
rect 10652 9868 10658 9880
rect 11609 9877 11621 9880
rect 11655 9877 11667 9911
rect 11609 9871 11667 9877
rect 1104 9818 13892 9840
rect 1104 9766 8214 9818
rect 8266 9766 8278 9818
rect 8330 9766 8342 9818
rect 8394 9766 8406 9818
rect 8458 9766 8470 9818
rect 8522 9766 13892 9818
rect 1104 9744 13892 9766
rect 6454 9664 6460 9716
rect 6512 9704 6518 9716
rect 7006 9704 7012 9716
rect 6512 9676 7012 9704
rect 6512 9664 6518 9676
rect 7006 9664 7012 9676
rect 7064 9664 7070 9716
rect 7193 9707 7251 9713
rect 7193 9673 7205 9707
rect 7239 9704 7251 9707
rect 7466 9704 7472 9716
rect 7239 9676 7472 9704
rect 7239 9673 7251 9676
rect 7193 9667 7251 9673
rect 7466 9664 7472 9676
rect 7524 9664 7530 9716
rect 7742 9664 7748 9716
rect 7800 9704 7806 9716
rect 8205 9707 8263 9713
rect 8205 9704 8217 9707
rect 7800 9676 8217 9704
rect 7800 9664 7806 9676
rect 8205 9673 8217 9676
rect 8251 9673 8263 9707
rect 8386 9704 8392 9716
rect 8205 9667 8263 9673
rect 8312 9676 8392 9704
rect 1397 9639 1455 9645
rect 1397 9605 1409 9639
rect 1443 9636 1455 9639
rect 1762 9636 1768 9648
rect 1443 9608 1768 9636
rect 1443 9605 1455 9608
rect 1397 9599 1455 9605
rect 1762 9596 1768 9608
rect 1820 9596 1826 9648
rect 3513 9639 3571 9645
rect 3513 9605 3525 9639
rect 3559 9636 3571 9639
rect 4522 9636 4528 9648
rect 3559 9608 4528 9636
rect 3559 9605 3571 9608
rect 3513 9599 3571 9605
rect 4522 9596 4528 9608
rect 4580 9596 4586 9648
rect 5258 9596 5264 9648
rect 5316 9636 5322 9648
rect 5445 9639 5503 9645
rect 5445 9636 5457 9639
rect 5316 9608 5457 9636
rect 5316 9596 5322 9608
rect 5445 9605 5457 9608
rect 5491 9605 5503 9639
rect 5445 9599 5503 9605
rect 7929 9639 7987 9645
rect 7929 9605 7941 9639
rect 7975 9636 7987 9639
rect 8312 9636 8340 9676
rect 8386 9664 8392 9676
rect 8444 9664 8450 9716
rect 8846 9704 8852 9716
rect 8807 9676 8852 9704
rect 8846 9664 8852 9676
rect 8904 9664 8910 9716
rect 9125 9707 9183 9713
rect 9125 9673 9137 9707
rect 9171 9674 9183 9707
rect 9214 9674 9220 9716
rect 9171 9673 9220 9674
rect 9125 9667 9220 9673
rect 9140 9664 9220 9667
rect 9272 9664 9278 9716
rect 9766 9704 9772 9716
rect 9428 9676 9772 9704
rect 9140 9646 9260 9664
rect 7975 9608 8340 9636
rect 8680 9608 8984 9636
rect 7975 9605 7987 9608
rect 7929 9599 7987 9605
rect 8380 9583 8438 9589
rect 8380 9580 8392 9583
rect 1486 9528 1492 9580
rect 1544 9568 1550 9580
rect 1581 9571 1639 9577
rect 1581 9568 1593 9571
rect 1544 9540 1593 9568
rect 1544 9528 1550 9540
rect 1581 9537 1593 9540
rect 1627 9537 1639 9571
rect 1581 9531 1639 9537
rect 3053 9571 3111 9577
rect 3053 9537 3065 9571
rect 3099 9568 3111 9571
rect 3234 9568 3240 9580
rect 3099 9540 3240 9568
rect 3099 9537 3111 9540
rect 3053 9531 3111 9537
rect 3234 9528 3240 9540
rect 3292 9568 3298 9580
rect 3329 9571 3387 9577
rect 3329 9568 3341 9571
rect 3292 9540 3341 9568
rect 3292 9528 3298 9540
rect 3329 9537 3341 9540
rect 3375 9537 3387 9571
rect 3694 9568 3700 9580
rect 3655 9540 3700 9568
rect 3329 9531 3387 9537
rect 3694 9528 3700 9540
rect 3752 9528 3758 9580
rect 5166 9568 5172 9580
rect 5079 9540 5172 9568
rect 5166 9528 5172 9540
rect 5224 9568 5230 9580
rect 6638 9577 6644 9580
rect 6181 9571 6239 9577
rect 6181 9568 6193 9571
rect 5224 9540 6193 9568
rect 5224 9528 5230 9540
rect 6181 9537 6193 9540
rect 6227 9537 6239 9571
rect 6636 9568 6644 9577
rect 6599 9540 6644 9568
rect 6181 9531 6239 9537
rect 6636 9531 6644 9540
rect 6638 9528 6644 9531
rect 6696 9528 6702 9580
rect 6730 9528 6736 9580
rect 6788 9568 6794 9580
rect 6871 9571 6929 9577
rect 6788 9540 6833 9568
rect 6788 9528 6794 9540
rect 6871 9537 6883 9571
rect 6917 9537 6929 9571
rect 6871 9531 6929 9537
rect 7009 9571 7067 9577
rect 7009 9537 7021 9571
rect 7055 9537 7067 9571
rect 7009 9531 7067 9537
rect 7561 9571 7619 9577
rect 7561 9537 7573 9571
rect 7607 9568 7619 9571
rect 7650 9568 7656 9580
rect 7607 9540 7656 9568
rect 7607 9537 7619 9540
rect 7561 9531 7619 9537
rect 5353 9503 5411 9509
rect 5353 9469 5365 9503
rect 5399 9500 5411 9503
rect 5902 9500 5908 9512
rect 5399 9472 5672 9500
rect 5863 9472 5908 9500
rect 5399 9469 5411 9472
rect 5353 9463 5411 9469
rect 2774 9392 2780 9444
rect 2832 9432 2838 9444
rect 2869 9435 2927 9441
rect 2869 9432 2881 9435
rect 2832 9404 2881 9432
rect 2832 9392 2838 9404
rect 2869 9401 2881 9404
rect 2915 9401 2927 9435
rect 2869 9395 2927 9401
rect 4522 9392 4528 9444
rect 4580 9432 4586 9444
rect 4985 9435 5043 9441
rect 4985 9432 4997 9435
rect 4580 9404 4997 9432
rect 4580 9392 4586 9404
rect 4985 9401 4997 9404
rect 5031 9401 5043 9435
rect 5644 9432 5672 9472
rect 5902 9460 5908 9472
rect 5960 9460 5966 9512
rect 5997 9435 6055 9441
rect 5997 9432 6009 9435
rect 5644 9404 6009 9432
rect 4985 9395 5043 9401
rect 5997 9401 6009 9404
rect 6043 9401 6055 9435
rect 5997 9395 6055 9401
rect 6822 9392 6828 9444
rect 6880 9404 6908 9531
rect 7024 9500 7052 9531
rect 7650 9528 7656 9540
rect 7708 9528 7714 9580
rect 8110 9528 8116 9580
rect 8168 9568 8174 9580
rect 8307 9568 8392 9580
rect 8168 9552 8392 9568
rect 8168 9540 8335 9552
rect 8380 9549 8392 9552
rect 8426 9549 8438 9583
rect 8380 9543 8438 9549
rect 8168 9528 8174 9540
rect 8478 9528 8484 9580
rect 8536 9568 8542 9580
rect 8680 9577 8708 9608
rect 8754 9577 8760 9580
rect 8665 9571 8723 9577
rect 8536 9540 8580 9568
rect 8536 9528 8542 9540
rect 8665 9537 8677 9571
rect 8711 9537 8723 9571
rect 8665 9531 8723 9537
rect 8752 9531 8760 9577
rect 8812 9568 8818 9580
rect 8956 9568 8984 9608
rect 9428 9568 9456 9676
rect 9766 9664 9772 9676
rect 9824 9664 9830 9716
rect 10134 9664 10140 9716
rect 10192 9704 10198 9716
rect 10778 9704 10784 9716
rect 10192 9676 10784 9704
rect 10192 9664 10198 9676
rect 10778 9664 10784 9676
rect 10836 9704 10842 9716
rect 11238 9704 11244 9716
rect 10836 9676 11244 9704
rect 10836 9664 10842 9676
rect 11238 9664 11244 9676
rect 11296 9664 11302 9716
rect 9858 9636 9864 9648
rect 9779 9608 9864 9636
rect 9779 9577 9807 9608
rect 9858 9596 9864 9608
rect 9916 9596 9922 9648
rect 10686 9636 10692 9648
rect 10647 9608 10692 9636
rect 10686 9596 10692 9608
rect 10744 9596 10750 9648
rect 11609 9639 11667 9645
rect 11609 9636 11621 9639
rect 11348 9608 11621 9636
rect 8812 9540 8852 9568
rect 8956 9540 9456 9568
rect 9493 9571 9551 9577
rect 8754 9528 8760 9531
rect 8812 9528 8818 9540
rect 9493 9537 9505 9571
rect 9539 9537 9551 9571
rect 9493 9531 9551 9537
rect 9769 9571 9827 9577
rect 9769 9537 9781 9571
rect 9815 9537 9827 9571
rect 9769 9531 9827 9537
rect 10045 9571 10103 9577
rect 10045 9537 10057 9571
rect 10091 9537 10103 9571
rect 10045 9531 10103 9537
rect 10321 9571 10379 9577
rect 10321 9537 10333 9571
rect 10367 9537 10379 9571
rect 10321 9531 10379 9537
rect 9508 9530 9544 9531
rect 7190 9500 7196 9512
rect 7024 9472 7196 9500
rect 7190 9460 7196 9472
rect 7248 9460 7254 9512
rect 7745 9503 7803 9509
rect 7745 9469 7757 9503
rect 7791 9500 7803 9503
rect 7834 9500 7840 9512
rect 7791 9472 7840 9500
rect 7791 9469 7803 9472
rect 7745 9463 7803 9469
rect 7834 9460 7840 9472
rect 7892 9460 7898 9512
rect 8128 9500 8156 9528
rect 7944 9472 8156 9500
rect 7558 9432 7564 9444
rect 7519 9404 7564 9432
rect 6880 9392 6886 9404
rect 7558 9392 7564 9404
rect 7616 9392 7622 9444
rect 7944 9432 7972 9472
rect 9306 9460 9312 9512
rect 9364 9500 9370 9512
rect 9401 9503 9459 9509
rect 9401 9500 9413 9503
rect 9364 9472 9413 9500
rect 9364 9460 9370 9472
rect 9401 9469 9413 9472
rect 9447 9469 9459 9503
rect 9516 9500 9544 9530
rect 9674 9500 9680 9512
rect 9516 9472 9680 9500
rect 9401 9463 9459 9469
rect 9674 9460 9680 9472
rect 9732 9460 9738 9512
rect 9950 9460 9956 9512
rect 10008 9500 10014 9512
rect 10060 9500 10088 9531
rect 10008 9472 10088 9500
rect 10137 9503 10195 9509
rect 10008 9460 10014 9472
rect 10137 9469 10149 9503
rect 10183 9500 10195 9503
rect 10226 9500 10232 9512
rect 10183 9472 10232 9500
rect 10183 9469 10195 9472
rect 10137 9463 10195 9469
rect 10226 9460 10232 9472
rect 10284 9460 10290 9512
rect 7668 9404 7972 9432
rect 6178 9324 6184 9376
rect 6236 9364 6242 9376
rect 6457 9367 6515 9373
rect 6457 9364 6469 9367
rect 6236 9336 6469 9364
rect 6236 9324 6242 9336
rect 6457 9333 6469 9336
rect 6503 9333 6515 9367
rect 6457 9327 6515 9333
rect 6638 9324 6644 9376
rect 6696 9364 6702 9376
rect 7668 9364 7696 9404
rect 8018 9392 8024 9444
rect 8076 9432 8082 9444
rect 9858 9432 9864 9444
rect 8076 9404 9864 9432
rect 8076 9392 8082 9404
rect 9858 9392 9864 9404
rect 9916 9392 9922 9444
rect 10042 9392 10048 9444
rect 10100 9432 10106 9444
rect 10336 9432 10364 9531
rect 10410 9528 10416 9580
rect 10468 9568 10474 9580
rect 10505 9571 10563 9577
rect 10505 9568 10517 9571
rect 10468 9540 10517 9568
rect 10468 9528 10474 9540
rect 10505 9537 10517 9540
rect 10551 9537 10563 9571
rect 11146 9568 11152 9580
rect 11107 9540 11152 9568
rect 10505 9531 10563 9537
rect 10520 9500 10548 9531
rect 11146 9528 11152 9540
rect 11204 9528 11210 9580
rect 11348 9577 11376 9608
rect 11609 9605 11621 9608
rect 11655 9605 11667 9639
rect 12802 9636 12808 9648
rect 12763 9608 12808 9636
rect 11609 9599 11667 9605
rect 12802 9596 12808 9608
rect 12860 9596 12866 9648
rect 13265 9639 13323 9645
rect 13265 9605 13277 9639
rect 13311 9636 13323 9639
rect 13354 9636 13360 9648
rect 13311 9608 13360 9636
rect 13311 9605 13323 9608
rect 13265 9599 13323 9605
rect 13354 9596 13360 9608
rect 13412 9596 13418 9648
rect 11333 9571 11391 9577
rect 11333 9537 11345 9571
rect 11379 9537 11391 9571
rect 11333 9531 11391 9537
rect 11517 9571 11575 9577
rect 11517 9537 11529 9571
rect 11563 9537 11575 9571
rect 11517 9531 11575 9537
rect 11885 9571 11943 9577
rect 11885 9537 11897 9571
rect 11931 9537 11943 9571
rect 11885 9531 11943 9537
rect 11532 9500 11560 9531
rect 10520 9472 11560 9500
rect 11606 9460 11612 9512
rect 11664 9500 11670 9512
rect 11701 9503 11759 9509
rect 11701 9500 11713 9503
rect 11664 9472 11713 9500
rect 11664 9460 11670 9472
rect 11701 9469 11713 9472
rect 11747 9469 11759 9503
rect 11701 9463 11759 9469
rect 10100 9404 10364 9432
rect 11241 9435 11299 9441
rect 10100 9392 10106 9404
rect 11241 9401 11253 9435
rect 11287 9432 11299 9435
rect 11422 9432 11428 9444
rect 11287 9404 11428 9432
rect 11287 9401 11299 9404
rect 11241 9395 11299 9401
rect 11422 9392 11428 9404
rect 11480 9392 11486 9444
rect 6696 9336 7696 9364
rect 6696 9324 6702 9336
rect 7926 9324 7932 9376
rect 7984 9364 7990 9376
rect 8846 9364 8852 9376
rect 7984 9336 8852 9364
rect 7984 9324 7990 9336
rect 8846 9324 8852 9336
rect 8904 9324 8910 9376
rect 9398 9364 9404 9376
rect 9359 9336 9404 9364
rect 9398 9324 9404 9336
rect 9456 9324 9462 9376
rect 9677 9367 9735 9373
rect 9677 9333 9689 9367
rect 9723 9364 9735 9367
rect 10134 9364 10140 9376
rect 9723 9336 10140 9364
rect 9723 9333 9735 9336
rect 9677 9327 9735 9333
rect 10134 9324 10140 9336
rect 10192 9324 10198 9376
rect 11330 9324 11336 9376
rect 11388 9364 11394 9376
rect 11900 9364 11928 9531
rect 12066 9528 12072 9580
rect 12124 9568 12130 9580
rect 12161 9571 12219 9577
rect 12161 9568 12173 9571
rect 12124 9540 12173 9568
rect 12124 9528 12130 9540
rect 12161 9537 12173 9540
rect 12207 9537 12219 9571
rect 12161 9531 12219 9537
rect 12710 9528 12716 9580
rect 12768 9568 12774 9580
rect 13081 9571 13139 9577
rect 13081 9568 13093 9571
rect 12768 9540 13093 9568
rect 12768 9528 12774 9540
rect 13081 9537 13093 9540
rect 13127 9537 13139 9571
rect 13081 9531 13139 9537
rect 13446 9432 13452 9444
rect 13407 9404 13452 9432
rect 13446 9392 13452 9404
rect 13504 9392 13510 9444
rect 11388 9336 11928 9364
rect 11388 9324 11394 9336
rect 1104 9274 13892 9296
rect 1104 9222 4214 9274
rect 4266 9222 4278 9274
rect 4330 9222 4342 9274
rect 4394 9222 4406 9274
rect 4458 9222 4470 9274
rect 4522 9222 12214 9274
rect 12266 9222 12278 9274
rect 12330 9222 12342 9274
rect 12394 9222 12406 9274
rect 12458 9222 12470 9274
rect 12522 9222 13892 9274
rect 1104 9200 13892 9222
rect 1489 9163 1547 9169
rect 1489 9129 1501 9163
rect 1535 9160 1547 9163
rect 1578 9160 1584 9172
rect 1535 9132 1584 9160
rect 1535 9129 1547 9132
rect 1489 9123 1547 9129
rect 1578 9120 1584 9132
rect 1636 9120 1642 9172
rect 2958 9120 2964 9172
rect 3016 9160 3022 9172
rect 3329 9163 3387 9169
rect 3329 9160 3341 9163
rect 3016 9132 3341 9160
rect 3016 9120 3022 9132
rect 3329 9129 3341 9132
rect 3375 9129 3387 9163
rect 3329 9123 3387 9129
rect 6546 9120 6552 9172
rect 6604 9160 6610 9172
rect 6641 9163 6699 9169
rect 6641 9160 6653 9163
rect 6604 9132 6653 9160
rect 6604 9120 6610 9132
rect 6641 9129 6653 9132
rect 6687 9129 6699 9163
rect 7098 9160 7104 9172
rect 6641 9123 6699 9129
rect 6840 9132 7104 9160
rect 3510 9092 3516 9104
rect 1964 9064 3516 9092
rect 1964 8965 1992 9064
rect 3510 9052 3516 9064
rect 3568 9052 3574 9104
rect 5718 9052 5724 9104
rect 5776 9092 5782 9104
rect 6840 9092 6868 9132
rect 7098 9120 7104 9132
rect 7156 9160 7162 9172
rect 7285 9163 7343 9169
rect 7285 9160 7297 9163
rect 7156 9132 7297 9160
rect 7156 9120 7162 9132
rect 7285 9129 7297 9132
rect 7331 9129 7343 9163
rect 7285 9123 7343 9129
rect 8018 9120 8024 9172
rect 8076 9160 8082 9172
rect 8205 9163 8263 9169
rect 8205 9160 8217 9163
rect 8076 9132 8217 9160
rect 8076 9120 8082 9132
rect 8205 9129 8217 9132
rect 8251 9129 8263 9163
rect 8205 9123 8263 9129
rect 8386 9120 8392 9172
rect 8444 9160 8450 9172
rect 8938 9160 8944 9172
rect 8444 9132 8944 9160
rect 8444 9120 8450 9132
rect 8938 9120 8944 9132
rect 8996 9120 9002 9172
rect 9122 9160 9128 9172
rect 9083 9132 9128 9160
rect 9122 9120 9128 9132
rect 9180 9160 9186 9172
rect 9674 9160 9680 9172
rect 9180 9132 9680 9160
rect 9180 9120 9186 9132
rect 9674 9120 9680 9132
rect 9732 9120 9738 9172
rect 9950 9120 9956 9172
rect 10008 9160 10014 9172
rect 10873 9163 10931 9169
rect 10873 9160 10885 9163
rect 10008 9132 10885 9160
rect 10008 9120 10014 9132
rect 10873 9129 10885 9132
rect 10919 9129 10931 9163
rect 10873 9123 10931 9129
rect 11149 9163 11207 9169
rect 11149 9129 11161 9163
rect 11195 9160 11207 9163
rect 11238 9160 11244 9172
rect 11195 9132 11244 9160
rect 11195 9129 11207 9132
rect 11149 9123 11207 9129
rect 11238 9120 11244 9132
rect 11296 9160 11302 9172
rect 12066 9160 12072 9172
rect 11296 9132 11744 9160
rect 12027 9132 12072 9160
rect 11296 9120 11302 9132
rect 8662 9092 8668 9104
rect 5776 9064 6868 9092
rect 6932 9064 8668 9092
rect 5776 9052 5782 9064
rect 6454 9024 6460 9036
rect 2746 8996 3924 9024
rect 1949 8959 2007 8965
rect 1949 8925 1961 8959
rect 1995 8925 2007 8959
rect 1949 8919 2007 8925
rect 2317 8959 2375 8965
rect 2317 8925 2329 8959
rect 2363 8956 2375 8959
rect 2590 8956 2596 8968
rect 2363 8928 2596 8956
rect 2363 8925 2375 8928
rect 2317 8919 2375 8925
rect 2590 8916 2596 8928
rect 2648 8916 2654 8968
rect 1762 8820 1768 8832
rect 1723 8792 1768 8820
rect 1762 8780 1768 8792
rect 1820 8780 1826 8832
rect 2130 8820 2136 8832
rect 2091 8792 2136 8820
rect 2130 8780 2136 8792
rect 2188 8820 2194 8832
rect 2746 8820 2774 8996
rect 2866 8916 2872 8968
rect 2924 8956 2930 8968
rect 2961 8959 3019 8965
rect 2961 8956 2973 8959
rect 2924 8928 2973 8956
rect 2924 8916 2930 8928
rect 2961 8925 2973 8928
rect 3007 8925 3019 8959
rect 3234 8956 3240 8968
rect 3195 8928 3240 8956
rect 2961 8919 3019 8925
rect 3234 8916 3240 8928
rect 3292 8956 3298 8968
rect 3896 8965 3924 8996
rect 4080 8996 5396 9024
rect 4080 8965 4108 8996
rect 3513 8959 3571 8965
rect 3513 8956 3525 8959
rect 3292 8928 3525 8956
rect 3292 8916 3298 8928
rect 3513 8925 3525 8928
rect 3559 8925 3571 8959
rect 3513 8919 3571 8925
rect 3881 8959 3939 8965
rect 3881 8925 3893 8959
rect 3927 8925 3939 8959
rect 3881 8919 3939 8925
rect 4065 8959 4123 8965
rect 4065 8925 4077 8959
rect 4111 8925 4123 8959
rect 4065 8919 4123 8925
rect 4525 8959 4583 8965
rect 4525 8925 4537 8959
rect 4571 8956 4583 8959
rect 4614 8956 4620 8968
rect 4571 8928 4620 8956
rect 4571 8925 4583 8928
rect 4525 8919 4583 8925
rect 4614 8916 4620 8928
rect 4672 8916 4678 8968
rect 4985 8959 5043 8965
rect 4985 8925 4997 8959
rect 5031 8956 5043 8959
rect 5258 8956 5264 8968
rect 5031 8928 5264 8956
rect 5031 8925 5043 8928
rect 4985 8919 5043 8925
rect 5258 8916 5264 8928
rect 5316 8916 5322 8968
rect 3789 8891 3847 8897
rect 3789 8857 3801 8891
rect 3835 8888 3847 8891
rect 3970 8888 3976 8900
rect 3835 8860 3976 8888
rect 3835 8857 3847 8860
rect 3789 8851 3847 8857
rect 3970 8848 3976 8860
rect 4028 8848 4034 8900
rect 4246 8888 4252 8900
rect 4207 8860 4252 8888
rect 4246 8848 4252 8860
rect 4304 8848 4310 8900
rect 4709 8891 4767 8897
rect 4709 8857 4721 8891
rect 4755 8888 4767 8891
rect 5166 8888 5172 8900
rect 4755 8860 5172 8888
rect 4755 8857 4767 8860
rect 4709 8851 4767 8857
rect 5166 8848 5172 8860
rect 5224 8848 5230 8900
rect 5368 8888 5396 8996
rect 6104 8996 6460 9024
rect 5629 8959 5687 8965
rect 5629 8925 5641 8959
rect 5675 8956 5687 8959
rect 5902 8956 5908 8968
rect 5675 8928 5908 8956
rect 5675 8925 5687 8928
rect 5629 8919 5687 8925
rect 5902 8916 5908 8928
rect 5960 8916 5966 8968
rect 6104 8965 6132 8996
rect 6454 8984 6460 8996
rect 6512 8984 6518 9036
rect 6932 9024 6960 9064
rect 6656 8996 6960 9024
rect 6089 8959 6147 8965
rect 6089 8925 6101 8959
rect 6135 8925 6147 8959
rect 6089 8919 6147 8925
rect 6273 8959 6331 8965
rect 6273 8925 6285 8959
rect 6319 8956 6331 8959
rect 6546 8956 6552 8968
rect 6319 8928 6552 8956
rect 6319 8925 6331 8928
rect 6273 8919 6331 8925
rect 6546 8916 6552 8928
rect 6604 8916 6610 8968
rect 6656 8965 6684 8996
rect 7006 8984 7012 9036
rect 7064 9024 7070 9036
rect 8021 9027 8079 9033
rect 8021 9024 8033 9027
rect 7064 8996 8033 9024
rect 7064 8984 7070 8996
rect 8021 8993 8033 8996
rect 8067 8993 8079 9027
rect 8021 8987 8079 8993
rect 6641 8959 6699 8965
rect 6641 8925 6653 8959
rect 6687 8925 6699 8959
rect 6641 8919 6699 8925
rect 6917 8959 6975 8965
rect 6917 8925 6929 8959
rect 6963 8925 6975 8959
rect 7098 8956 7104 8968
rect 7059 8928 7104 8956
rect 6917 8919 6975 8925
rect 6822 8888 6828 8900
rect 5368 8860 6828 8888
rect 6822 8848 6828 8860
rect 6880 8848 6886 8900
rect 6937 8888 6965 8919
rect 7098 8916 7104 8928
rect 7156 8916 7162 8968
rect 7834 8956 7840 8968
rect 7795 8928 7840 8956
rect 7834 8916 7840 8928
rect 7892 8916 7898 8968
rect 8113 8959 8171 8965
rect 8113 8925 8125 8959
rect 8159 8956 8171 8959
rect 8202 8956 8208 8968
rect 8159 8928 8208 8956
rect 8159 8925 8171 8928
rect 8113 8919 8171 8925
rect 8202 8916 8208 8928
rect 8260 8916 8266 8968
rect 6937 8860 7144 8888
rect 2188 8792 2774 8820
rect 4617 8823 4675 8829
rect 2188 8780 2194 8792
rect 4617 8789 4629 8823
rect 4663 8820 4675 8823
rect 5442 8820 5448 8832
rect 4663 8792 5448 8820
rect 4663 8789 4675 8792
rect 4617 8783 4675 8789
rect 5442 8780 5448 8792
rect 5500 8780 5506 8832
rect 5718 8820 5724 8832
rect 5679 8792 5724 8820
rect 5718 8780 5724 8792
rect 5776 8780 5782 8832
rect 6181 8823 6239 8829
rect 6181 8789 6193 8823
rect 6227 8820 6239 8823
rect 7116 8820 7144 8860
rect 7558 8848 7564 8900
rect 7616 8888 7622 8900
rect 7653 8891 7711 8897
rect 7653 8888 7665 8891
rect 7616 8860 7665 8888
rect 7616 8848 7622 8860
rect 7653 8857 7665 8860
rect 7699 8857 7711 8891
rect 8496 8888 8524 9064
rect 8662 9052 8668 9064
rect 8720 9052 8726 9104
rect 8846 9052 8852 9104
rect 8904 9092 8910 9104
rect 9398 9092 9404 9104
rect 8904 9064 9404 9092
rect 8904 9052 8910 9064
rect 9398 9052 9404 9064
rect 9456 9052 9462 9104
rect 9766 9092 9772 9104
rect 9679 9064 9772 9092
rect 9766 9052 9772 9064
rect 9824 9092 9830 9104
rect 11606 9092 11612 9104
rect 9824 9064 11612 9092
rect 9824 9052 9830 9064
rect 11606 9052 11612 9064
rect 11664 9052 11670 9104
rect 9030 9024 9036 9036
rect 8991 8996 9036 9024
rect 9030 8984 9036 8996
rect 9088 8984 9094 9036
rect 9306 8984 9312 9036
rect 9364 9024 9370 9036
rect 9582 9024 9588 9036
rect 9364 8996 9588 9024
rect 9364 8984 9370 8996
rect 9582 8984 9588 8996
rect 9640 8984 9646 9036
rect 8570 8916 8576 8968
rect 8628 8956 8634 8968
rect 8754 8956 8760 8968
rect 8628 8928 8760 8956
rect 8628 8916 8634 8928
rect 8754 8916 8760 8928
rect 8812 8956 8818 8968
rect 9784 8965 9812 9052
rect 10042 8984 10048 9036
rect 10100 9024 10106 9036
rect 10321 9027 10379 9033
rect 10321 9024 10333 9027
rect 10100 8996 10333 9024
rect 10100 8984 10106 8996
rect 10321 8993 10333 8996
rect 10367 8993 10379 9027
rect 10321 8987 10379 8993
rect 10870 8984 10876 9036
rect 10928 9024 10934 9036
rect 10928 8996 11284 9024
rect 10928 8984 10934 8996
rect 9217 8959 9275 8965
rect 9217 8956 9229 8959
rect 8812 8928 9229 8956
rect 8812 8916 8818 8928
rect 9217 8925 9229 8928
rect 9263 8925 9275 8959
rect 9217 8919 9275 8925
rect 9769 8959 9827 8965
rect 9769 8925 9781 8959
rect 9815 8925 9827 8959
rect 9769 8919 9827 8925
rect 9953 8959 10011 8965
rect 9953 8925 9965 8959
rect 9999 8925 10011 8959
rect 10134 8956 10140 8968
rect 10095 8928 10140 8956
rect 9953 8919 10011 8925
rect 8941 8891 8999 8897
rect 8941 8888 8953 8891
rect 8496 8860 8953 8888
rect 7653 8851 7711 8857
rect 8941 8857 8953 8860
rect 8987 8888 8999 8891
rect 9861 8891 9919 8897
rect 9861 8888 9873 8891
rect 8987 8860 9873 8888
rect 8987 8857 8999 8860
rect 8941 8851 8999 8857
rect 9861 8857 9873 8860
rect 9907 8857 9919 8891
rect 9968 8888 9996 8919
rect 10134 8916 10140 8928
rect 10192 8956 10198 8968
rect 11256 8965 11284 8996
rect 10689 8959 10747 8965
rect 10689 8956 10701 8959
rect 10192 8928 10701 8956
rect 10192 8916 10198 8928
rect 10689 8925 10701 8928
rect 10735 8956 10747 8959
rect 10965 8959 11023 8965
rect 10965 8956 10977 8959
rect 10735 8928 10977 8956
rect 10735 8925 10747 8928
rect 10689 8919 10747 8925
rect 10965 8925 10977 8928
rect 11011 8925 11023 8959
rect 10965 8919 11023 8925
rect 11241 8959 11299 8965
rect 11241 8925 11253 8959
rect 11287 8925 11299 8959
rect 11241 8919 11299 8925
rect 11330 8916 11336 8968
rect 11388 8956 11394 8968
rect 11614 8959 11672 8965
rect 11614 8956 11626 8959
rect 11388 8928 11626 8956
rect 11388 8916 11394 8928
rect 11614 8925 11626 8928
rect 11660 8925 11672 8959
rect 11614 8919 11672 8925
rect 10226 8888 10232 8900
rect 9968 8860 10232 8888
rect 9861 8851 9919 8857
rect 10226 8848 10232 8860
rect 10284 8888 10290 8900
rect 10505 8891 10563 8897
rect 10505 8888 10517 8891
rect 10284 8860 10517 8888
rect 10284 8848 10290 8860
rect 10505 8857 10517 8860
rect 10551 8888 10563 8891
rect 10551 8860 10824 8888
rect 10551 8857 10563 8860
rect 10505 8851 10563 8857
rect 9122 8820 9128 8832
rect 6227 8792 9128 8820
rect 6227 8789 6239 8792
rect 6181 8783 6239 8789
rect 9122 8780 9128 8792
rect 9180 8780 9186 8832
rect 9401 8823 9459 8829
rect 9401 8789 9413 8823
rect 9447 8820 9459 8823
rect 10686 8820 10692 8832
rect 9447 8792 10692 8820
rect 9447 8789 9459 8792
rect 9401 8783 9459 8789
rect 10686 8780 10692 8792
rect 10744 8780 10750 8832
rect 10796 8820 10824 8860
rect 10870 8848 10876 8900
rect 10928 8888 10934 8900
rect 11425 8891 11483 8897
rect 11425 8888 11437 8891
rect 10928 8860 11437 8888
rect 10928 8848 10934 8860
rect 11425 8857 11437 8860
rect 11471 8857 11483 8891
rect 11425 8851 11483 8857
rect 11517 8891 11575 8897
rect 11517 8857 11529 8891
rect 11563 8888 11575 8891
rect 11716 8888 11744 9132
rect 12066 9120 12072 9132
rect 12124 9120 12130 9172
rect 11793 9095 11851 9101
rect 11793 9061 11805 9095
rect 11839 9092 11851 9095
rect 12342 9092 12348 9104
rect 11839 9064 12348 9092
rect 11839 9061 11851 9064
rect 11793 9055 11851 9061
rect 12342 9052 12348 9064
rect 12400 9092 12406 9104
rect 12400 9064 12664 9092
rect 12400 9052 12406 9064
rect 12636 9033 12664 9064
rect 12621 9027 12679 9033
rect 12621 8993 12633 9027
rect 12667 8993 12679 9027
rect 12621 8987 12679 8993
rect 11882 8916 11888 8968
rect 11940 8956 11946 8968
rect 12253 8959 12311 8965
rect 12253 8956 12265 8959
rect 11940 8928 12265 8956
rect 11940 8916 11946 8928
rect 12253 8925 12265 8928
rect 12299 8925 12311 8959
rect 12253 8919 12311 8925
rect 13262 8916 13268 8968
rect 13320 8956 13326 8968
rect 13449 8959 13507 8965
rect 13449 8956 13461 8959
rect 13320 8928 13461 8956
rect 13320 8916 13326 8928
rect 13449 8925 13461 8928
rect 13495 8925 13507 8959
rect 13449 8919 13507 8925
rect 12437 8891 12495 8897
rect 12437 8888 12449 8891
rect 11563 8860 12449 8888
rect 11563 8857 11575 8860
rect 11517 8851 11575 8857
rect 12437 8857 12449 8860
rect 12483 8857 12495 8891
rect 12437 8851 12495 8857
rect 12529 8891 12587 8897
rect 12529 8857 12541 8891
rect 12575 8888 12587 8891
rect 12894 8888 12900 8900
rect 12575 8860 12900 8888
rect 12575 8857 12587 8860
rect 12529 8851 12587 8857
rect 12894 8848 12900 8860
rect 12952 8848 12958 8900
rect 13078 8888 13084 8900
rect 13039 8860 13084 8888
rect 13078 8848 13084 8860
rect 13136 8848 13142 8900
rect 13173 8891 13231 8897
rect 13173 8857 13185 8891
rect 13219 8857 13231 8891
rect 13173 8851 13231 8857
rect 11330 8820 11336 8832
rect 10796 8792 11336 8820
rect 11330 8780 11336 8792
rect 11388 8780 11394 8832
rect 13188 8820 13216 8851
rect 13265 8823 13323 8829
rect 13265 8820 13277 8823
rect 13188 8792 13277 8820
rect 13265 8789 13277 8792
rect 13311 8789 13323 8823
rect 13265 8783 13323 8789
rect 1104 8730 13892 8752
rect 1104 8678 8214 8730
rect 8266 8678 8278 8730
rect 8330 8678 8342 8730
rect 8394 8678 8406 8730
rect 8458 8678 8470 8730
rect 8522 8678 13892 8730
rect 1104 8656 13892 8678
rect 5534 8576 5540 8628
rect 5592 8616 5598 8628
rect 6546 8616 6552 8628
rect 5592 8588 6552 8616
rect 5592 8576 5598 8588
rect 6546 8576 6552 8588
rect 6604 8616 6610 8628
rect 6604 8588 7052 8616
rect 6604 8576 6610 8588
rect 4982 8508 4988 8560
rect 5040 8548 5046 8560
rect 5169 8551 5227 8557
rect 5169 8548 5181 8551
rect 5040 8520 5181 8548
rect 5040 8508 5046 8520
rect 5169 8517 5181 8520
rect 5215 8517 5227 8551
rect 5442 8548 5448 8560
rect 5403 8520 5448 8548
rect 5169 8511 5227 8517
rect 5442 8508 5448 8520
rect 5500 8508 5506 8560
rect 6365 8551 6423 8557
rect 6365 8517 6377 8551
rect 6411 8548 6423 8551
rect 6822 8548 6828 8560
rect 6411 8520 6828 8548
rect 6411 8517 6423 8520
rect 6365 8511 6423 8517
rect 6822 8508 6828 8520
rect 6880 8508 6886 8560
rect 7024 8548 7052 8588
rect 7558 8576 7564 8628
rect 7616 8616 7622 8628
rect 9306 8616 9312 8628
rect 7616 8588 9312 8616
rect 7616 8576 7622 8588
rect 9306 8576 9312 8588
rect 9364 8576 9370 8628
rect 9490 8616 9496 8628
rect 9451 8588 9496 8616
rect 9490 8576 9496 8588
rect 9548 8576 9554 8628
rect 9582 8576 9588 8628
rect 9640 8616 9646 8628
rect 9640 8588 11100 8616
rect 9640 8576 9646 8588
rect 8110 8548 8116 8560
rect 7024 8520 8116 8548
rect 8110 8508 8116 8520
rect 8168 8508 8174 8560
rect 9950 8548 9956 8560
rect 8220 8520 9956 8548
rect 1486 8480 1492 8492
rect 1447 8452 1492 8480
rect 1486 8440 1492 8452
rect 1544 8440 1550 8492
rect 3605 8483 3663 8489
rect 3605 8449 3617 8483
rect 3651 8480 3663 8483
rect 4246 8480 4252 8492
rect 3651 8452 4252 8480
rect 3651 8449 3663 8452
rect 3605 8443 3663 8449
rect 4246 8440 4252 8452
rect 4304 8440 4310 8492
rect 5077 8483 5135 8489
rect 5077 8449 5089 8483
rect 5123 8480 5135 8483
rect 5258 8480 5264 8492
rect 5123 8452 5264 8480
rect 5123 8449 5135 8452
rect 5077 8443 5135 8449
rect 5258 8440 5264 8452
rect 5316 8440 5322 8492
rect 6178 8480 6184 8492
rect 6139 8452 6184 8480
rect 6178 8440 6184 8452
rect 6236 8440 6242 8492
rect 6546 8480 6552 8492
rect 6507 8452 6552 8480
rect 6546 8440 6552 8452
rect 6604 8440 6610 8492
rect 6733 8483 6791 8489
rect 6733 8449 6745 8483
rect 6779 8449 6791 8483
rect 7006 8480 7012 8492
rect 6967 8452 7012 8480
rect 6733 8443 6791 8449
rect 2958 8344 2964 8356
rect 2919 8316 2964 8344
rect 2958 8304 2964 8316
rect 3016 8304 3022 8356
rect 6748 8344 6776 8443
rect 7006 8440 7012 8452
rect 7064 8440 7070 8492
rect 7377 8483 7435 8489
rect 7377 8449 7389 8483
rect 7423 8480 7435 8483
rect 7834 8480 7840 8492
rect 7423 8452 7840 8480
rect 7423 8449 7435 8452
rect 7377 8443 7435 8449
rect 7834 8440 7840 8452
rect 7892 8440 7898 8492
rect 8220 8489 8248 8520
rect 9950 8508 9956 8520
rect 10008 8508 10014 8560
rect 11072 8548 11100 8588
rect 11146 8576 11152 8628
rect 11204 8616 11210 8628
rect 11241 8619 11299 8625
rect 11241 8616 11253 8619
rect 11204 8588 11253 8616
rect 11204 8576 11210 8588
rect 11241 8585 11253 8588
rect 11287 8585 11299 8619
rect 11698 8616 11704 8628
rect 11241 8579 11299 8585
rect 11440 8588 11704 8616
rect 11440 8548 11468 8588
rect 11698 8576 11704 8588
rect 11756 8616 11762 8628
rect 11756 8588 11928 8616
rect 11756 8576 11762 8588
rect 11072 8520 11468 8548
rect 11517 8551 11575 8557
rect 11517 8517 11529 8551
rect 11563 8548 11575 8551
rect 11606 8548 11612 8560
rect 11563 8520 11612 8548
rect 11563 8517 11575 8520
rect 11517 8511 11575 8517
rect 11606 8508 11612 8520
rect 11664 8508 11670 8560
rect 11900 8557 11928 8588
rect 11974 8576 11980 8628
rect 12032 8616 12038 8628
rect 12253 8619 12311 8625
rect 12253 8616 12265 8619
rect 12032 8588 12265 8616
rect 12032 8576 12038 8588
rect 12253 8585 12265 8588
rect 12299 8585 12311 8619
rect 12253 8579 12311 8585
rect 11885 8551 11943 8557
rect 11885 8517 11897 8551
rect 11931 8517 11943 8551
rect 12710 8548 12716 8560
rect 11885 8511 11943 8517
rect 12084 8520 12716 8548
rect 8205 8483 8263 8489
rect 8205 8449 8217 8483
rect 8251 8449 8263 8483
rect 9125 8483 9183 8489
rect 9125 8480 9137 8483
rect 8205 8443 8263 8449
rect 8312 8452 9137 8480
rect 6914 8412 6920 8424
rect 6875 8384 6920 8412
rect 6914 8372 6920 8384
rect 6972 8372 6978 8424
rect 8018 8412 8024 8424
rect 7979 8384 8024 8412
rect 8018 8372 8024 8384
rect 8076 8412 8082 8424
rect 8312 8412 8340 8452
rect 9125 8449 9137 8452
rect 9171 8449 9183 8483
rect 9125 8443 9183 8449
rect 9381 8483 9439 8489
rect 9381 8449 9393 8483
rect 9427 8480 9439 8483
rect 9427 8452 9807 8480
rect 9427 8449 9439 8452
rect 9381 8443 9439 8449
rect 8076 8384 8340 8412
rect 8849 8415 8907 8421
rect 8076 8372 8082 8384
rect 8849 8381 8861 8415
rect 8895 8412 8907 8415
rect 9490 8412 9496 8424
rect 8895 8384 9496 8412
rect 8895 8381 8907 8384
rect 8849 8375 8907 8381
rect 9490 8372 9496 8384
rect 9548 8412 9554 8424
rect 9585 8415 9643 8421
rect 9585 8412 9597 8415
rect 9548 8384 9597 8412
rect 9548 8372 9554 8384
rect 9585 8381 9597 8384
rect 9631 8381 9643 8415
rect 9585 8375 9643 8381
rect 9677 8415 9735 8421
rect 9677 8381 9689 8415
rect 9723 8381 9735 8415
rect 9779 8412 9807 8452
rect 9858 8440 9864 8492
rect 9916 8480 9922 8492
rect 10137 8483 10195 8489
rect 10137 8480 10149 8483
rect 9916 8452 10149 8480
rect 9916 8440 9922 8452
rect 10137 8449 10149 8452
rect 10183 8449 10195 8483
rect 10137 8443 10195 8449
rect 10410 8440 10416 8492
rect 10468 8480 10474 8492
rect 12084 8489 12112 8520
rect 12710 8508 12716 8520
rect 12768 8508 12774 8560
rect 13078 8548 13084 8560
rect 13039 8520 13084 8548
rect 13078 8508 13084 8520
rect 13136 8548 13142 8560
rect 13357 8551 13415 8557
rect 13357 8548 13369 8551
rect 13136 8520 13369 8548
rect 13136 8508 13142 8520
rect 13357 8517 13369 8520
rect 13403 8517 13415 8551
rect 13357 8511 13415 8517
rect 11701 8483 11759 8489
rect 11701 8480 11713 8483
rect 10468 8452 11713 8480
rect 10468 8440 10474 8452
rect 11701 8449 11713 8452
rect 11747 8449 11759 8483
rect 11701 8443 11759 8449
rect 12069 8483 12127 8489
rect 12069 8449 12081 8483
rect 12115 8449 12127 8483
rect 12342 8480 12348 8492
rect 12303 8452 12348 8480
rect 12069 8443 12127 8449
rect 12342 8440 12348 8452
rect 12400 8440 12406 8492
rect 13262 8480 13268 8492
rect 13223 8452 13268 8480
rect 13262 8440 13268 8452
rect 13320 8440 13326 8492
rect 10042 8412 10048 8424
rect 9779 8384 10048 8412
rect 9677 8375 9735 8381
rect 9214 8344 9220 8356
rect 6748 8316 9220 8344
rect 9214 8304 9220 8316
rect 9272 8304 9278 8356
rect 9692 8288 9720 8375
rect 10042 8372 10048 8384
rect 10100 8372 10106 8424
rect 10226 8412 10232 8424
rect 10187 8384 10232 8412
rect 10226 8372 10232 8384
rect 10284 8372 10290 8424
rect 10594 8372 10600 8424
rect 10652 8412 10658 8424
rect 10873 8415 10931 8421
rect 10873 8412 10885 8415
rect 10652 8384 10885 8412
rect 10652 8372 10658 8384
rect 10873 8381 10885 8384
rect 10919 8381 10931 8415
rect 10873 8375 10931 8381
rect 11149 8415 11207 8421
rect 11149 8381 11161 8415
rect 11195 8412 11207 8415
rect 11238 8412 11244 8424
rect 11195 8384 11244 8412
rect 11195 8381 11207 8384
rect 11149 8375 11207 8381
rect 11238 8372 11244 8384
rect 11296 8372 11302 8424
rect 12066 8304 12072 8356
rect 12124 8344 12130 8356
rect 13449 8347 13507 8353
rect 13449 8344 13461 8347
rect 12124 8316 13461 8344
rect 12124 8304 12130 8316
rect 13449 8313 13461 8316
rect 13495 8313 13507 8347
rect 13449 8307 13507 8313
rect 3050 8236 3056 8288
rect 3108 8276 3114 8288
rect 3421 8279 3479 8285
rect 3421 8276 3433 8279
rect 3108 8248 3433 8276
rect 3108 8236 3114 8248
rect 3421 8245 3433 8248
rect 3467 8245 3479 8279
rect 3421 8239 3479 8245
rect 7285 8279 7343 8285
rect 7285 8245 7297 8279
rect 7331 8276 7343 8279
rect 7650 8276 7656 8288
rect 7331 8248 7656 8276
rect 7331 8245 7343 8248
rect 7285 8239 7343 8245
rect 7650 8236 7656 8248
rect 7708 8236 7714 8288
rect 8938 8276 8944 8288
rect 8899 8248 8944 8276
rect 8938 8236 8944 8248
rect 8996 8236 9002 8288
rect 9674 8236 9680 8288
rect 9732 8236 9738 8288
rect 1104 8186 13892 8208
rect 1104 8134 4214 8186
rect 4266 8134 4278 8186
rect 4330 8134 4342 8186
rect 4394 8134 4406 8186
rect 4458 8134 4470 8186
rect 4522 8134 12214 8186
rect 12266 8134 12278 8186
rect 12330 8134 12342 8186
rect 12394 8134 12406 8186
rect 12458 8134 12470 8186
rect 12522 8134 13892 8186
rect 1104 8112 13892 8134
rect 1486 8072 1492 8084
rect 1447 8044 1492 8072
rect 1486 8032 1492 8044
rect 1544 8032 1550 8084
rect 5258 8072 5264 8084
rect 4816 8044 5264 8072
rect 3786 7936 3792 7948
rect 2884 7908 3792 7936
rect 1762 7868 1768 7880
rect 1723 7840 1768 7868
rect 1762 7828 1768 7840
rect 1820 7828 1826 7880
rect 2884 7877 2912 7908
rect 3786 7896 3792 7908
rect 3844 7896 3850 7948
rect 4062 7896 4068 7948
rect 4120 7936 4126 7948
rect 4157 7939 4215 7945
rect 4157 7936 4169 7939
rect 4120 7908 4169 7936
rect 4120 7896 4126 7908
rect 4157 7905 4169 7908
rect 4203 7905 4215 7939
rect 4157 7899 4215 7905
rect 4614 7896 4620 7948
rect 4672 7936 4678 7948
rect 4709 7939 4767 7945
rect 4709 7936 4721 7939
rect 4672 7908 4721 7936
rect 4672 7896 4678 7908
rect 4709 7905 4721 7908
rect 4755 7905 4767 7939
rect 4709 7899 4767 7905
rect 2869 7871 2927 7877
rect 2869 7837 2881 7871
rect 2915 7837 2927 7871
rect 3050 7868 3056 7880
rect 3011 7840 3056 7868
rect 2869 7831 2927 7837
rect 3050 7828 3056 7840
rect 3108 7868 3114 7880
rect 3881 7871 3939 7877
rect 3881 7868 3893 7871
rect 3108 7840 3893 7868
rect 3108 7828 3114 7840
rect 3881 7837 3893 7840
rect 3927 7868 3939 7871
rect 3970 7868 3976 7880
rect 3927 7840 3976 7868
rect 3927 7837 3939 7840
rect 3881 7831 3939 7837
rect 3970 7828 3976 7840
rect 4028 7828 4034 7880
rect 4816 7877 4844 8044
rect 5258 8032 5264 8044
rect 5316 8072 5322 8084
rect 5905 8075 5963 8081
rect 5905 8072 5917 8075
rect 5316 8044 5917 8072
rect 5316 8032 5322 8044
rect 5905 8041 5917 8044
rect 5951 8041 5963 8075
rect 7834 8072 7840 8084
rect 7795 8044 7840 8072
rect 5905 8035 5963 8041
rect 7834 8032 7840 8044
rect 7892 8032 7898 8084
rect 12894 8032 12900 8084
rect 12952 8072 12958 8084
rect 13449 8075 13507 8081
rect 13449 8072 13461 8075
rect 12952 8044 13461 8072
rect 12952 8032 12958 8044
rect 13449 8041 13461 8044
rect 13495 8072 13507 8075
rect 13538 8072 13544 8084
rect 13495 8044 13544 8072
rect 13495 8041 13507 8044
rect 13449 8035 13507 8041
rect 13538 8032 13544 8044
rect 13596 8032 13602 8084
rect 5169 8007 5227 8013
rect 5169 7973 5181 8007
rect 5215 8004 5227 8007
rect 5442 8004 5448 8016
rect 5215 7976 5448 8004
rect 5215 7973 5227 7976
rect 5169 7967 5227 7973
rect 5442 7964 5448 7976
rect 5500 7964 5506 8016
rect 10226 8004 10232 8016
rect 6748 7976 7788 8004
rect 10187 7976 10232 8004
rect 5629 7939 5687 7945
rect 5629 7905 5641 7939
rect 5675 7936 5687 7939
rect 6086 7936 6092 7948
rect 5675 7908 6092 7936
rect 5675 7905 5687 7908
rect 5629 7899 5687 7905
rect 6086 7896 6092 7908
rect 6144 7896 6150 7948
rect 4801 7871 4859 7877
rect 4801 7837 4813 7871
rect 4847 7837 4859 7871
rect 4801 7831 4859 7837
rect 4982 7828 4988 7880
rect 5040 7828 5046 7880
rect 6748 7877 6776 7976
rect 7760 7948 7788 7976
rect 10226 7964 10232 7976
rect 10284 7964 10290 8016
rect 7009 7939 7067 7945
rect 7009 7905 7021 7939
rect 7055 7936 7067 7939
rect 7190 7936 7196 7948
rect 7055 7908 7196 7936
rect 7055 7905 7067 7908
rect 7009 7899 7067 7905
rect 7190 7896 7196 7908
rect 7248 7896 7254 7948
rect 7742 7896 7748 7948
rect 7800 7936 7806 7948
rect 7929 7939 7987 7945
rect 7929 7936 7941 7939
rect 7800 7908 7941 7936
rect 7800 7896 7806 7908
rect 7929 7905 7941 7908
rect 7975 7905 7987 7939
rect 7929 7899 7987 7905
rect 8018 7896 8024 7948
rect 8076 7936 8082 7948
rect 8205 7939 8263 7945
rect 8205 7936 8217 7939
rect 8076 7908 8217 7936
rect 8076 7896 8082 7908
rect 8205 7905 8217 7908
rect 8251 7905 8263 7939
rect 8205 7899 8263 7905
rect 8757 7939 8815 7945
rect 8757 7905 8769 7939
rect 8803 7936 8815 7939
rect 9585 7939 9643 7945
rect 9585 7936 9597 7939
rect 8803 7908 9597 7936
rect 8803 7905 8815 7908
rect 8757 7899 8815 7905
rect 9585 7905 9597 7908
rect 9631 7936 9643 7939
rect 9674 7936 9680 7948
rect 9631 7908 9680 7936
rect 9631 7905 9643 7908
rect 9585 7899 9643 7905
rect 9674 7896 9680 7908
rect 9732 7936 9738 7948
rect 9732 7908 10640 7936
rect 9732 7896 9738 7908
rect 6733 7871 6791 7877
rect 6733 7837 6745 7871
rect 6779 7837 6791 7871
rect 6733 7831 6791 7837
rect 6822 7828 6828 7880
rect 6880 7868 6886 7880
rect 7561 7871 7619 7877
rect 7561 7868 7573 7871
rect 6880 7840 7573 7868
rect 6880 7828 6886 7840
rect 7561 7837 7573 7840
rect 7607 7837 7619 7871
rect 7561 7831 7619 7837
rect 7650 7828 7656 7880
rect 7708 7868 7714 7880
rect 8110 7868 8116 7880
rect 7708 7840 7753 7868
rect 8071 7840 8116 7868
rect 7708 7828 7714 7840
rect 8110 7828 8116 7840
rect 8168 7828 8174 7880
rect 8572 7871 8630 7877
rect 8572 7837 8584 7871
rect 8618 7868 8630 7871
rect 9030 7868 9036 7880
rect 8618 7840 9036 7868
rect 8618 7837 8630 7840
rect 8572 7831 8630 7837
rect 9030 7828 9036 7840
rect 9088 7828 9094 7880
rect 9490 7868 9496 7880
rect 9451 7840 9496 7868
rect 9490 7828 9496 7840
rect 9548 7828 9554 7880
rect 9950 7828 9956 7880
rect 10008 7868 10014 7880
rect 10612 7877 10640 7908
rect 10471 7871 10529 7877
rect 10471 7868 10483 7871
rect 10008 7840 10483 7868
rect 10008 7828 10014 7840
rect 10471 7837 10483 7840
rect 10517 7837 10529 7871
rect 10471 7831 10529 7837
rect 10597 7871 10655 7877
rect 10597 7837 10609 7871
rect 10643 7837 10655 7871
rect 10597 7831 10655 7837
rect 10686 7828 10692 7880
rect 10744 7868 10750 7880
rect 10744 7840 10789 7868
rect 10744 7828 10750 7840
rect 10870 7828 10876 7880
rect 10928 7868 10934 7880
rect 10928 7840 10973 7868
rect 10928 7828 10934 7840
rect 11054 7828 11060 7880
rect 11112 7868 11118 7880
rect 11333 7871 11391 7877
rect 11333 7868 11345 7871
rect 11112 7840 11345 7868
rect 11112 7828 11118 7840
rect 11333 7837 11345 7840
rect 11379 7837 11391 7871
rect 11333 7831 11391 7837
rect 11701 7871 11759 7877
rect 11701 7837 11713 7871
rect 11747 7868 11759 7871
rect 11793 7871 11851 7877
rect 11793 7868 11805 7871
rect 11747 7840 11805 7868
rect 11747 7837 11759 7840
rect 11701 7831 11759 7837
rect 11793 7837 11805 7840
rect 11839 7837 11851 7871
rect 13262 7868 13268 7880
rect 13223 7840 13268 7868
rect 11793 7831 11851 7837
rect 13262 7828 13268 7840
rect 13320 7828 13326 7880
rect 1670 7760 1676 7812
rect 1728 7800 1734 7812
rect 3145 7803 3203 7809
rect 3145 7800 3157 7803
rect 1728 7772 3157 7800
rect 1728 7760 1734 7772
rect 3145 7769 3157 7772
rect 3191 7769 3203 7803
rect 3145 7763 3203 7769
rect 3329 7803 3387 7809
rect 3329 7769 3341 7803
rect 3375 7769 3387 7803
rect 3510 7800 3516 7812
rect 3471 7772 3516 7800
rect 3329 7763 3387 7769
rect 2777 7735 2835 7741
rect 2777 7701 2789 7735
rect 2823 7732 2835 7735
rect 2866 7732 2872 7744
rect 2823 7704 2872 7732
rect 2823 7701 2835 7704
rect 2777 7695 2835 7701
rect 2866 7692 2872 7704
rect 2924 7692 2930 7744
rect 3050 7692 3056 7744
rect 3108 7732 3114 7744
rect 3344 7732 3372 7763
rect 3510 7760 3516 7772
rect 3568 7760 3574 7812
rect 4617 7803 4675 7809
rect 4617 7769 4629 7803
rect 4663 7800 4675 7803
rect 5000 7800 5028 7828
rect 4663 7772 5028 7800
rect 5077 7803 5135 7809
rect 4663 7769 4675 7772
rect 4617 7763 4675 7769
rect 5077 7769 5089 7803
rect 5123 7769 5135 7803
rect 5077 7763 5135 7769
rect 3694 7732 3700 7744
rect 3108 7704 3700 7732
rect 3108 7692 3114 7704
rect 3694 7692 3700 7704
rect 3752 7692 3758 7744
rect 4985 7735 5043 7741
rect 4985 7701 4997 7735
rect 5031 7732 5043 7735
rect 5092 7732 5120 7763
rect 5442 7760 5448 7812
rect 5500 7800 5506 7812
rect 5813 7803 5871 7809
rect 5813 7800 5825 7803
rect 5500 7772 5825 7800
rect 5500 7760 5506 7772
rect 5813 7769 5825 7772
rect 5859 7800 5871 7803
rect 11517 7803 11575 7809
rect 5859 7772 11468 7800
rect 5859 7769 5871 7772
rect 5813 7763 5871 7769
rect 5031 7704 5120 7732
rect 6089 7735 6147 7741
rect 5031 7701 5043 7704
rect 4985 7695 5043 7701
rect 6089 7701 6101 7735
rect 6135 7732 6147 7735
rect 6270 7732 6276 7744
rect 6135 7704 6276 7732
rect 6135 7701 6147 7704
rect 6089 7695 6147 7701
rect 6270 7692 6276 7704
rect 6328 7692 6334 7744
rect 7374 7732 7380 7744
rect 7335 7704 7380 7732
rect 7374 7692 7380 7704
rect 7432 7692 7438 7744
rect 10134 7732 10140 7744
rect 10095 7704 10140 7732
rect 10134 7692 10140 7704
rect 10192 7692 10198 7744
rect 11440 7732 11468 7772
rect 11517 7769 11529 7803
rect 11563 7800 11575 7803
rect 11974 7800 11980 7812
rect 11563 7772 11980 7800
rect 11563 7769 11575 7772
rect 11517 7763 11575 7769
rect 11974 7760 11980 7772
rect 12032 7760 12038 7812
rect 13357 7803 13415 7809
rect 13357 7800 13369 7803
rect 12406 7772 13369 7800
rect 12250 7732 12256 7744
rect 11440 7704 12256 7732
rect 12250 7692 12256 7704
rect 12308 7732 12314 7744
rect 12406 7732 12434 7772
rect 13357 7769 13369 7772
rect 13403 7769 13415 7803
rect 13357 7763 13415 7769
rect 12308 7704 12434 7732
rect 12308 7692 12314 7704
rect 1104 7642 13892 7664
rect 1104 7590 8214 7642
rect 8266 7590 8278 7642
rect 8330 7590 8342 7642
rect 8394 7590 8406 7642
rect 8458 7590 8470 7642
rect 8522 7590 13892 7642
rect 1104 7568 13892 7590
rect 2409 7531 2467 7537
rect 2409 7497 2421 7531
rect 2455 7528 2467 7531
rect 3418 7528 3424 7540
rect 2455 7500 3424 7528
rect 2455 7497 2467 7500
rect 2409 7491 2467 7497
rect 3418 7488 3424 7500
rect 3476 7488 3482 7540
rect 3694 7488 3700 7540
rect 3752 7528 3758 7540
rect 6457 7531 6515 7537
rect 3752 7500 4844 7528
rect 3752 7488 3758 7500
rect 2317 7463 2375 7469
rect 2317 7429 2329 7463
rect 2363 7460 2375 7463
rect 3050 7460 3056 7472
rect 2363 7432 3056 7460
rect 2363 7429 2375 7432
rect 2317 7423 2375 7429
rect 3050 7420 3056 7432
rect 3108 7420 3114 7472
rect 1670 7392 1676 7404
rect 1631 7364 1676 7392
rect 1670 7352 1676 7364
rect 1728 7352 1734 7404
rect 1762 7352 1768 7404
rect 1820 7392 1826 7404
rect 1820 7364 1865 7392
rect 1820 7352 1826 7364
rect 4154 7352 4160 7404
rect 4212 7352 4218 7404
rect 4709 7395 4767 7401
rect 4709 7361 4721 7395
rect 4755 7361 4767 7395
rect 4816 7392 4844 7500
rect 6457 7497 6469 7531
rect 6503 7528 6515 7531
rect 6822 7528 6828 7540
rect 6503 7500 6828 7528
rect 6503 7497 6515 7500
rect 6457 7491 6515 7497
rect 6822 7488 6828 7500
rect 6880 7488 6886 7540
rect 7466 7528 7472 7540
rect 7427 7500 7472 7528
rect 7466 7488 7472 7500
rect 7524 7488 7530 7540
rect 8110 7488 8116 7540
rect 8168 7528 8174 7540
rect 9677 7531 9735 7537
rect 8168 7500 9260 7528
rect 8168 7488 8174 7500
rect 6730 7460 6736 7472
rect 5644 7432 6736 7460
rect 4893 7395 4951 7401
rect 4893 7392 4905 7395
rect 4816 7364 4905 7392
rect 4709 7355 4767 7361
rect 4893 7361 4905 7364
rect 4939 7361 4951 7395
rect 5442 7392 5448 7404
rect 5403 7364 5448 7392
rect 4893 7355 4951 7361
rect 2590 7324 2596 7336
rect 2551 7296 2596 7324
rect 2590 7284 2596 7296
rect 2648 7284 2654 7336
rect 2774 7284 2780 7336
rect 2832 7324 2838 7336
rect 3050 7324 3056 7336
rect 2832 7296 2877 7324
rect 3011 7296 3056 7324
rect 2832 7284 2838 7296
rect 3050 7284 3056 7296
rect 3108 7284 3114 7336
rect 3510 7284 3516 7336
rect 3568 7324 3574 7336
rect 4724 7324 4752 7355
rect 3568 7296 4752 7324
rect 4908 7324 4936 7355
rect 5442 7352 5448 7364
rect 5500 7352 5506 7404
rect 5534 7352 5540 7404
rect 5592 7392 5598 7404
rect 5644 7401 5672 7432
rect 6730 7420 6736 7432
rect 6788 7420 6794 7472
rect 6914 7460 6920 7472
rect 6840 7432 6920 7460
rect 5629 7395 5687 7401
rect 5629 7392 5641 7395
rect 5592 7364 5641 7392
rect 5592 7352 5598 7364
rect 5629 7361 5641 7364
rect 5675 7361 5687 7395
rect 5629 7355 5687 7361
rect 5718 7352 5724 7404
rect 5776 7392 5782 7404
rect 5813 7395 5871 7401
rect 5813 7392 5825 7395
rect 5776 7364 5825 7392
rect 5776 7352 5782 7364
rect 5813 7361 5825 7364
rect 5859 7392 5871 7395
rect 5997 7395 6055 7401
rect 5997 7392 6009 7395
rect 5859 7364 6009 7392
rect 5859 7361 5871 7364
rect 5813 7355 5871 7361
rect 5997 7361 6009 7364
rect 6043 7361 6055 7395
rect 5997 7355 6055 7361
rect 6270 7352 6276 7404
rect 6328 7392 6334 7404
rect 6840 7401 6868 7432
rect 6914 7420 6920 7432
rect 6972 7420 6978 7472
rect 7558 7420 7564 7472
rect 7616 7420 7622 7472
rect 7668 7432 8524 7460
rect 6641 7395 6699 7401
rect 6641 7392 6653 7395
rect 6328 7364 6653 7392
rect 6328 7352 6334 7364
rect 6641 7361 6653 7364
rect 6687 7361 6699 7395
rect 6641 7355 6699 7361
rect 6825 7395 6883 7401
rect 6825 7361 6837 7395
rect 6871 7361 6883 7395
rect 6825 7355 6883 7361
rect 7101 7395 7159 7401
rect 7101 7361 7113 7395
rect 7147 7392 7159 7395
rect 7190 7392 7196 7404
rect 7147 7364 7196 7392
rect 7147 7361 7159 7364
rect 7101 7355 7159 7361
rect 6086 7324 6092 7336
rect 4908 7296 6092 7324
rect 3568 7284 3574 7296
rect 6086 7284 6092 7296
rect 6144 7284 6150 7336
rect 6656 7324 6684 7355
rect 7190 7352 7196 7364
rect 7248 7352 7254 7404
rect 7357 7395 7415 7401
rect 7357 7361 7369 7395
rect 7403 7392 7415 7395
rect 7576 7392 7604 7420
rect 7668 7401 7696 7432
rect 7403 7364 7604 7392
rect 7653 7395 7711 7401
rect 7403 7361 7415 7364
rect 7357 7355 7415 7361
rect 7653 7361 7665 7395
rect 7699 7361 7711 7395
rect 7653 7355 7711 7361
rect 8496 7392 8524 7432
rect 8938 7392 8944 7404
rect 8496 7364 8944 7392
rect 7006 7324 7012 7336
rect 6656 7296 7012 7324
rect 7006 7284 7012 7296
rect 7064 7284 7070 7336
rect 7561 7327 7619 7333
rect 7561 7293 7573 7327
rect 7607 7293 7619 7327
rect 7561 7287 7619 7293
rect 8021 7327 8079 7333
rect 8021 7293 8033 7327
rect 8067 7324 8079 7327
rect 8386 7324 8392 7336
rect 8067 7296 8392 7324
rect 8067 7293 8079 7296
rect 8021 7287 8079 7293
rect 1762 7216 1768 7268
rect 1820 7256 1826 7268
rect 4801 7259 4859 7265
rect 4801 7256 4813 7259
rect 1820 7228 2176 7256
rect 1820 7216 1826 7228
rect 1486 7188 1492 7200
rect 1447 7160 1492 7188
rect 1486 7148 1492 7160
rect 1544 7148 1550 7200
rect 1946 7188 1952 7200
rect 1907 7160 1952 7188
rect 1946 7148 1952 7160
rect 2004 7148 2010 7200
rect 2148 7188 2176 7228
rect 4080 7228 4813 7256
rect 4080 7188 4108 7228
rect 4801 7225 4813 7228
rect 4847 7225 4859 7259
rect 4801 7219 4859 7225
rect 5629 7259 5687 7265
rect 5629 7225 5641 7259
rect 5675 7256 5687 7259
rect 5718 7256 5724 7268
rect 5675 7228 5724 7256
rect 5675 7225 5687 7228
rect 5629 7219 5687 7225
rect 5718 7216 5724 7228
rect 5776 7216 5782 7268
rect 7576 7256 7604 7287
rect 8036 7256 8064 7287
rect 8386 7284 8392 7296
rect 8444 7284 8450 7336
rect 7576 7228 8064 7256
rect 8294 7216 8300 7268
rect 8352 7256 8358 7268
rect 8496 7256 8524 7364
rect 8938 7352 8944 7364
rect 8996 7352 9002 7404
rect 9232 7401 9260 7500
rect 9677 7497 9689 7531
rect 9723 7528 9735 7531
rect 10686 7528 10692 7540
rect 9723 7500 10692 7528
rect 9723 7497 9735 7500
rect 9677 7491 9735 7497
rect 10686 7488 10692 7500
rect 10744 7488 10750 7540
rect 12250 7488 12256 7540
rect 12308 7528 12314 7540
rect 12805 7531 12863 7537
rect 12805 7528 12817 7531
rect 12308 7500 12817 7528
rect 12308 7488 12314 7500
rect 12805 7497 12817 7500
rect 12851 7497 12863 7531
rect 12805 7491 12863 7497
rect 12066 7420 12072 7472
rect 12124 7460 12130 7472
rect 12345 7463 12403 7469
rect 12345 7460 12357 7463
rect 12124 7432 12357 7460
rect 12124 7420 12130 7432
rect 12345 7429 12357 7432
rect 12391 7429 12403 7463
rect 12345 7423 12403 7429
rect 9217 7395 9275 7401
rect 9217 7361 9229 7395
rect 9263 7361 9275 7395
rect 9217 7355 9275 7361
rect 9401 7395 9459 7401
rect 9401 7361 9413 7395
rect 9447 7392 9459 7395
rect 9953 7395 10011 7401
rect 9953 7392 9965 7395
rect 9447 7364 9965 7392
rect 9447 7361 9459 7364
rect 9401 7355 9459 7361
rect 9953 7361 9965 7364
rect 9999 7361 10011 7395
rect 10226 7392 10232 7404
rect 10187 7364 10232 7392
rect 9953 7355 10011 7361
rect 8846 7324 8852 7336
rect 8807 7296 8852 7324
rect 8846 7284 8852 7296
rect 8904 7284 8910 7336
rect 8352 7228 8524 7256
rect 8352 7216 8358 7228
rect 2148 7160 4108 7188
rect 4525 7191 4583 7197
rect 4525 7157 4537 7191
rect 4571 7188 4583 7191
rect 4614 7188 4620 7200
rect 4571 7160 4620 7188
rect 4571 7157 4583 7160
rect 4525 7151 4583 7157
rect 4614 7148 4620 7160
rect 4672 7148 4678 7200
rect 5258 7188 5264 7200
rect 5219 7160 5264 7188
rect 5258 7148 5264 7160
rect 5316 7148 5322 7200
rect 8018 7148 8024 7200
rect 8076 7188 8082 7200
rect 9416 7188 9444 7355
rect 9769 7327 9827 7333
rect 9769 7293 9781 7327
rect 9815 7324 9827 7327
rect 9861 7327 9919 7333
rect 9861 7324 9873 7327
rect 9815 7296 9873 7324
rect 9815 7293 9827 7296
rect 9769 7287 9827 7293
rect 9861 7293 9873 7296
rect 9907 7293 9919 7327
rect 9968 7324 9996 7355
rect 10226 7352 10232 7364
rect 10284 7352 10290 7404
rect 11054 7352 11060 7404
rect 11112 7392 11118 7404
rect 11793 7395 11851 7401
rect 11793 7392 11805 7395
rect 11112 7364 11805 7392
rect 11112 7352 11118 7364
rect 11793 7361 11805 7364
rect 11839 7361 11851 7395
rect 12250 7392 12256 7404
rect 12211 7364 12256 7392
rect 11793 7355 11851 7361
rect 12250 7352 12256 7364
rect 12308 7352 12314 7404
rect 10502 7324 10508 7336
rect 9968 7296 10508 7324
rect 9861 7287 9919 7293
rect 10502 7284 10508 7296
rect 10560 7284 10566 7336
rect 12066 7284 12072 7336
rect 12124 7324 12130 7336
rect 12437 7327 12495 7333
rect 12437 7324 12449 7327
rect 12124 7296 12449 7324
rect 12124 7284 12130 7296
rect 12437 7293 12449 7296
rect 12483 7293 12495 7327
rect 12437 7287 12495 7293
rect 12805 7327 12863 7333
rect 12805 7293 12817 7327
rect 12851 7324 12863 7327
rect 12897 7327 12955 7333
rect 12897 7324 12909 7327
rect 12851 7296 12909 7324
rect 12851 7293 12863 7296
rect 12805 7287 12863 7293
rect 12897 7293 12909 7296
rect 12943 7293 12955 7327
rect 12897 7287 12955 7293
rect 8076 7160 9444 7188
rect 8076 7148 8082 7160
rect 1104 7098 13892 7120
rect 1104 7046 4214 7098
rect 4266 7046 4278 7098
rect 4330 7046 4342 7098
rect 4394 7046 4406 7098
rect 4458 7046 4470 7098
rect 4522 7046 12214 7098
rect 12266 7046 12278 7098
rect 12330 7046 12342 7098
rect 12394 7046 12406 7098
rect 12458 7046 12470 7098
rect 12522 7046 13892 7098
rect 1104 7024 13892 7046
rect 1752 6987 1810 6993
rect 1752 6953 1764 6987
rect 1798 6984 1810 6987
rect 1946 6984 1952 6996
rect 1798 6956 1952 6984
rect 1798 6953 1810 6956
rect 1752 6947 1810 6953
rect 1946 6944 1952 6956
rect 2004 6944 2010 6996
rect 3237 6987 3295 6993
rect 3237 6953 3249 6987
rect 3283 6984 3295 6987
rect 3510 6984 3516 6996
rect 3283 6956 3516 6984
rect 3283 6953 3295 6956
rect 3237 6947 3295 6953
rect 3510 6944 3516 6956
rect 3568 6944 3574 6996
rect 3970 6944 3976 6996
rect 4028 6984 4034 6996
rect 4154 6984 4160 6996
rect 4028 6956 4160 6984
rect 4028 6944 4034 6956
rect 4154 6944 4160 6956
rect 4212 6984 4218 6996
rect 4249 6987 4307 6993
rect 4249 6984 4261 6987
rect 4212 6956 4261 6984
rect 4212 6944 4218 6956
rect 4249 6953 4261 6956
rect 4295 6984 4307 6987
rect 5626 6984 5632 6996
rect 4295 6956 5632 6984
rect 4295 6953 4307 6956
rect 4249 6947 4307 6953
rect 5626 6944 5632 6956
rect 5684 6944 5690 6996
rect 5892 6987 5950 6993
rect 5892 6953 5904 6987
rect 5938 6984 5950 6987
rect 7374 6984 7380 6996
rect 5938 6956 7380 6984
rect 5938 6953 5950 6956
rect 5892 6947 5950 6953
rect 7374 6944 7380 6956
rect 7432 6944 7438 6996
rect 5644 6916 5672 6944
rect 2792 6888 4200 6916
rect 5644 6888 5764 6916
rect 2792 6860 2820 6888
rect 3988 6860 4016 6888
rect 1489 6851 1547 6857
rect 1489 6817 1501 6851
rect 1535 6848 1547 6851
rect 2774 6848 2780 6860
rect 1535 6820 2780 6848
rect 1535 6817 1547 6820
rect 1489 6811 1547 6817
rect 2774 6808 2780 6820
rect 2832 6808 2838 6860
rect 3970 6808 3976 6860
rect 4028 6808 4034 6860
rect 4172 6848 4200 6888
rect 4525 6851 4583 6857
rect 4525 6848 4537 6851
rect 4172 6820 4537 6848
rect 4525 6817 4537 6820
rect 4571 6848 4583 6851
rect 5626 6848 5632 6860
rect 4571 6820 5632 6848
rect 4571 6817 4583 6820
rect 4525 6811 4583 6817
rect 5626 6808 5632 6820
rect 5684 6808 5690 6860
rect 5736 6848 5764 6888
rect 7834 6876 7840 6928
rect 7892 6916 7898 6928
rect 9674 6916 9680 6928
rect 7892 6888 9680 6916
rect 7892 6876 7898 6888
rect 6454 6848 6460 6860
rect 5736 6820 6460 6848
rect 6454 6808 6460 6820
rect 6512 6848 6518 6860
rect 6914 6848 6920 6860
rect 6512 6820 6920 6848
rect 6512 6808 6518 6820
rect 6914 6808 6920 6820
rect 6972 6808 6978 6860
rect 7377 6851 7435 6857
rect 7377 6817 7389 6851
rect 7423 6848 7435 6851
rect 7650 6848 7656 6860
rect 7423 6820 7656 6848
rect 7423 6817 7435 6820
rect 7377 6811 7435 6817
rect 7650 6808 7656 6820
rect 7708 6808 7714 6860
rect 7745 6851 7803 6857
rect 7745 6817 7757 6851
rect 7791 6848 7803 6851
rect 8570 6848 8576 6860
rect 7791 6820 8576 6848
rect 7791 6817 7803 6820
rect 7745 6811 7803 6817
rect 8570 6808 8576 6820
rect 8628 6848 8634 6860
rect 9324 6857 9352 6888
rect 9674 6876 9680 6888
rect 9732 6876 9738 6928
rect 13262 6916 13268 6928
rect 13223 6888 13268 6916
rect 13262 6876 13268 6888
rect 13320 6876 13326 6928
rect 8757 6851 8815 6857
rect 8757 6848 8769 6851
rect 8628 6820 8769 6848
rect 8628 6808 8634 6820
rect 8757 6817 8769 6820
rect 8803 6817 8815 6851
rect 8757 6811 8815 6817
rect 9309 6851 9367 6857
rect 9309 6817 9321 6851
rect 9355 6817 9367 6851
rect 11606 6848 11612 6860
rect 9309 6811 9367 6817
rect 9600 6820 11612 6848
rect 2866 6740 2872 6792
rect 2924 6740 2930 6792
rect 3326 6740 3332 6792
rect 3384 6780 3390 6792
rect 3421 6783 3479 6789
rect 3421 6780 3433 6783
rect 3384 6752 3433 6780
rect 3384 6740 3390 6752
rect 3421 6749 3433 6752
rect 3467 6749 3479 6783
rect 3421 6743 3479 6749
rect 3786 6740 3792 6792
rect 3844 6780 3850 6792
rect 3881 6783 3939 6789
rect 3881 6780 3893 6783
rect 3844 6752 3893 6780
rect 3844 6740 3850 6752
rect 3881 6749 3893 6752
rect 3927 6749 3939 6783
rect 4154 6780 4160 6792
rect 4115 6752 4160 6780
rect 3881 6743 3939 6749
rect 4154 6740 4160 6752
rect 4212 6740 4218 6792
rect 5258 6780 5264 6792
rect 5219 6752 5264 6780
rect 5258 6740 5264 6752
rect 5316 6740 5322 6792
rect 7190 6740 7196 6792
rect 7248 6780 7254 6792
rect 7929 6783 7987 6789
rect 7929 6780 7941 6783
rect 7248 6752 7941 6780
rect 7248 6740 7254 6752
rect 7760 6724 7788 6752
rect 7929 6749 7941 6752
rect 7975 6780 7987 6783
rect 8018 6780 8024 6792
rect 7975 6752 8024 6780
rect 7975 6749 7987 6752
rect 7929 6743 7987 6749
rect 8018 6740 8024 6752
rect 8076 6740 8082 6792
rect 8113 6783 8171 6789
rect 8113 6749 8125 6783
rect 8159 6749 8171 6783
rect 8113 6743 8171 6749
rect 8205 6783 8263 6789
rect 8205 6749 8217 6783
rect 8251 6780 8263 6783
rect 8294 6780 8300 6792
rect 8251 6752 8300 6780
rect 8251 6749 8263 6752
rect 8205 6743 8263 6749
rect 6546 6672 6552 6724
rect 6604 6672 6610 6724
rect 7742 6672 7748 6724
rect 7800 6672 7806 6724
rect 8128 6712 8156 6743
rect 8294 6740 8300 6752
rect 8352 6740 8358 6792
rect 8386 6740 8392 6792
rect 8444 6780 8450 6792
rect 8444 6752 8800 6780
rect 8444 6740 8450 6752
rect 8772 6724 8800 6752
rect 8846 6740 8852 6792
rect 8904 6780 8910 6792
rect 9600 6789 9628 6820
rect 11606 6808 11612 6820
rect 11664 6848 11670 6860
rect 11793 6851 11851 6857
rect 11793 6848 11805 6851
rect 11664 6820 11805 6848
rect 11664 6808 11670 6820
rect 11793 6817 11805 6820
rect 11839 6817 11851 6851
rect 11793 6811 11851 6817
rect 9493 6783 9551 6789
rect 9493 6780 9505 6783
rect 8904 6752 9505 6780
rect 8904 6740 8910 6752
rect 9493 6749 9505 6752
rect 9539 6749 9551 6783
rect 9493 6743 9551 6749
rect 9585 6783 9643 6789
rect 9585 6749 9597 6783
rect 9631 6749 9643 6783
rect 10042 6780 10048 6792
rect 10003 6752 10048 6780
rect 9585 6743 9643 6749
rect 8662 6712 8668 6724
rect 8128 6684 8524 6712
rect 8623 6684 8668 6712
rect 1486 6604 1492 6656
rect 1544 6644 1550 6656
rect 2498 6644 2504 6656
rect 1544 6616 2504 6644
rect 1544 6604 1550 6616
rect 2498 6604 2504 6616
rect 2556 6604 2562 6656
rect 4062 6644 4068 6656
rect 4023 6616 4068 6644
rect 4062 6604 4068 6616
rect 4120 6604 4126 6656
rect 8496 6644 8524 6684
rect 8662 6672 8668 6684
rect 8720 6672 8726 6724
rect 8754 6672 8760 6724
rect 8812 6672 8818 6724
rect 9306 6644 9312 6656
rect 8496 6616 9312 6644
rect 9306 6604 9312 6616
rect 9364 6644 9370 6656
rect 9600 6644 9628 6743
rect 10042 6740 10048 6752
rect 10100 6740 10106 6792
rect 11698 6740 11704 6792
rect 11756 6780 11762 6792
rect 11977 6783 12035 6789
rect 11977 6780 11989 6783
rect 11756 6752 11989 6780
rect 11756 6740 11762 6752
rect 11977 6749 11989 6752
rect 12023 6780 12035 6783
rect 12342 6780 12348 6792
rect 12023 6752 12348 6780
rect 12023 6749 12035 6752
rect 11977 6743 12035 6749
rect 12342 6740 12348 6752
rect 12400 6740 12406 6792
rect 13446 6780 13452 6792
rect 13407 6752 13452 6780
rect 13446 6740 13452 6752
rect 13504 6740 13510 6792
rect 10321 6715 10379 6721
rect 10321 6681 10333 6715
rect 10367 6681 10379 6715
rect 11882 6712 11888 6724
rect 11546 6684 11888 6712
rect 10321 6675 10379 6681
rect 9364 6616 9628 6644
rect 9953 6647 10011 6653
rect 9364 6604 9370 6616
rect 9953 6613 9965 6647
rect 9999 6644 10011 6647
rect 10336 6644 10364 6675
rect 11882 6672 11888 6684
rect 11940 6672 11946 6724
rect 9999 6616 10364 6644
rect 9999 6613 10011 6616
rect 9953 6607 10011 6613
rect 1104 6554 13892 6576
rect 1104 6502 8214 6554
rect 8266 6502 8278 6554
rect 8330 6502 8342 6554
rect 8394 6502 8406 6554
rect 8458 6502 8470 6554
rect 8522 6502 13892 6554
rect 1104 6480 13892 6502
rect 2038 6400 2044 6452
rect 2096 6400 2102 6452
rect 3050 6400 3056 6452
rect 3108 6440 3114 6452
rect 3513 6443 3571 6449
rect 3513 6440 3525 6443
rect 3108 6412 3525 6440
rect 3108 6400 3114 6412
rect 3513 6409 3525 6412
rect 3559 6409 3571 6443
rect 3513 6403 3571 6409
rect 3881 6443 3939 6449
rect 3881 6409 3893 6443
rect 3927 6440 3939 6443
rect 5534 6440 5540 6452
rect 3927 6412 5540 6440
rect 3927 6409 3939 6412
rect 3881 6403 3939 6409
rect 2057 6335 2085 6400
rect 2042 6329 2100 6335
rect 1762 6304 1768 6316
rect 1723 6276 1768 6304
rect 1762 6264 1768 6276
rect 1820 6264 1826 6316
rect 1946 6313 1952 6316
rect 1931 6307 1952 6313
rect 1931 6273 1943 6307
rect 1931 6267 1952 6273
rect 1946 6264 1952 6267
rect 2004 6264 2010 6316
rect 2042 6295 2054 6329
rect 2088 6295 2100 6329
rect 2498 6304 2504 6316
rect 2042 6289 2100 6295
rect 2134 6297 2192 6303
rect 2134 6263 2146 6297
rect 2180 6263 2192 6297
rect 2459 6276 2504 6304
rect 2498 6264 2504 6276
rect 2556 6264 2562 6316
rect 2682 6304 2688 6316
rect 2643 6276 2688 6304
rect 2682 6264 2688 6276
rect 2740 6264 2746 6316
rect 3237 6307 3295 6313
rect 3237 6273 3249 6307
rect 3283 6273 3295 6307
rect 3237 6267 3295 6273
rect 3421 6307 3479 6313
rect 3421 6273 3433 6307
rect 3467 6304 3479 6307
rect 3896 6304 3924 6403
rect 5534 6400 5540 6412
rect 5592 6400 5598 6452
rect 6086 6440 6092 6452
rect 6047 6412 6092 6440
rect 6086 6400 6092 6412
rect 6144 6400 6150 6452
rect 6546 6440 6552 6452
rect 6507 6412 6552 6440
rect 6546 6400 6552 6412
rect 6604 6400 6610 6452
rect 10137 6443 10195 6449
rect 10137 6409 10149 6443
rect 10183 6440 10195 6443
rect 10410 6440 10416 6452
rect 10183 6412 10416 6440
rect 10183 6409 10195 6412
rect 10137 6403 10195 6409
rect 10410 6400 10416 6412
rect 10468 6400 10474 6452
rect 10870 6400 10876 6452
rect 10928 6400 10934 6452
rect 12066 6440 12072 6452
rect 11808 6412 12072 6440
rect 3970 6332 3976 6384
rect 4028 6332 4034 6384
rect 6914 6372 6920 6384
rect 6875 6344 6920 6372
rect 6914 6332 6920 6344
rect 6972 6332 6978 6384
rect 7101 6375 7159 6381
rect 7101 6341 7113 6375
rect 7147 6372 7159 6375
rect 7466 6372 7472 6384
rect 7147 6344 7472 6372
rect 7147 6341 7159 6344
rect 7101 6335 7159 6341
rect 7466 6332 7472 6344
rect 7524 6372 7530 6384
rect 7524 6344 8892 6372
rect 7524 6332 7530 6344
rect 3467 6276 3924 6304
rect 3988 6304 4016 6332
rect 4341 6307 4399 6313
rect 4341 6304 4353 6307
rect 3988 6276 4353 6304
rect 3467 6273 3479 6276
rect 3421 6267 3479 6273
rect 4341 6273 4353 6276
rect 4387 6273 4399 6307
rect 4341 6267 4399 6273
rect 2134 6257 2192 6263
rect 1394 6100 1400 6112
rect 1355 6072 1400 6100
rect 1394 6060 1400 6072
rect 1452 6100 1458 6112
rect 1581 6103 1639 6109
rect 1581 6100 1593 6103
rect 1452 6072 1593 6100
rect 1452 6060 1458 6072
rect 1581 6069 1593 6072
rect 1627 6100 1639 6103
rect 2148 6100 2176 6257
rect 3252 6236 3280 6267
rect 5718 6264 5724 6316
rect 5776 6264 5782 6316
rect 6454 6264 6460 6316
rect 6512 6313 6518 6316
rect 6512 6307 6561 6313
rect 6512 6273 6515 6307
rect 6549 6273 6561 6307
rect 6512 6267 6561 6273
rect 6641 6307 6699 6313
rect 6641 6273 6653 6307
rect 6687 6273 6699 6307
rect 7926 6304 7932 6316
rect 7839 6276 7932 6304
rect 6641 6267 6699 6273
rect 6512 6264 6518 6267
rect 3973 6239 4031 6245
rect 3973 6236 3985 6239
rect 3252 6208 3985 6236
rect 3973 6205 3985 6208
rect 4019 6205 4031 6239
rect 3973 6199 4031 6205
rect 2222 6128 2228 6180
rect 2280 6168 2286 6180
rect 2409 6171 2467 6177
rect 2409 6168 2421 6171
rect 2280 6140 2421 6168
rect 2280 6128 2286 6140
rect 2409 6137 2421 6140
rect 2455 6137 2467 6171
rect 3142 6168 3148 6180
rect 3103 6140 3148 6168
rect 2409 6131 2467 6137
rect 3142 6128 3148 6140
rect 3200 6128 3206 6180
rect 1627 6072 2176 6100
rect 1627 6069 1639 6072
rect 1581 6063 1639 6069
rect 2314 6060 2320 6112
rect 2372 6100 2378 6112
rect 2869 6103 2927 6109
rect 2869 6100 2881 6103
rect 2372 6072 2881 6100
rect 2372 6060 2378 6072
rect 2869 6069 2881 6072
rect 2915 6069 2927 6103
rect 3988 6100 4016 6199
rect 4062 6196 4068 6248
rect 4120 6236 4126 6248
rect 4617 6239 4675 6245
rect 4120 6208 4165 6236
rect 4120 6196 4126 6208
rect 4617 6205 4629 6239
rect 4663 6236 4675 6239
rect 5350 6236 5356 6248
rect 4663 6208 5356 6236
rect 4663 6205 4675 6208
rect 4617 6199 4675 6205
rect 5350 6196 5356 6208
rect 5408 6196 5414 6248
rect 6656 6236 6684 6267
rect 7926 6264 7932 6276
rect 7984 6264 7990 6316
rect 8662 6304 8668 6316
rect 8623 6276 8668 6304
rect 8662 6264 8668 6276
rect 8720 6264 8726 6316
rect 8864 6313 8892 6344
rect 9674 6332 9680 6384
rect 9732 6372 9738 6384
rect 10888 6372 10916 6400
rect 11149 6375 11207 6381
rect 11149 6372 11161 6375
rect 9732 6344 11161 6372
rect 9732 6332 9738 6344
rect 8849 6307 8907 6313
rect 8849 6273 8861 6307
rect 8895 6273 8907 6307
rect 10244 6304 10272 6344
rect 11149 6341 11161 6344
rect 11195 6341 11207 6375
rect 11808 6372 11836 6412
rect 12066 6400 12072 6412
rect 12124 6400 12130 6452
rect 11149 6335 11207 6341
rect 11716 6344 11836 6372
rect 10686 6304 10692 6316
rect 10244 6276 10364 6304
rect 10647 6276 10692 6304
rect 8849 6267 8907 6273
rect 6730 6236 6736 6248
rect 6656 6208 6736 6236
rect 6730 6196 6736 6208
rect 6788 6196 6794 6248
rect 7742 6236 7748 6248
rect 7703 6208 7748 6236
rect 7742 6196 7748 6208
rect 7800 6196 7806 6248
rect 7944 6168 7972 6264
rect 10336 6245 10364 6276
rect 10686 6264 10692 6276
rect 10744 6264 10750 6316
rect 10778 6264 10784 6316
rect 10836 6304 10842 6316
rect 11716 6313 11744 6344
rect 11882 6332 11888 6384
rect 11940 6372 11946 6384
rect 11977 6375 12035 6381
rect 11977 6372 11989 6375
rect 11940 6344 11989 6372
rect 11940 6332 11946 6344
rect 11977 6341 11989 6344
rect 12023 6341 12035 6375
rect 11977 6335 12035 6341
rect 13173 6375 13231 6381
rect 13173 6341 13185 6375
rect 13219 6372 13231 6375
rect 13262 6372 13268 6384
rect 13219 6344 13268 6372
rect 13219 6341 13231 6344
rect 13173 6335 13231 6341
rect 13262 6332 13268 6344
rect 13320 6332 13326 6384
rect 10965 6307 11023 6313
rect 10836 6276 10881 6304
rect 10836 6264 10842 6276
rect 10965 6273 10977 6307
rect 11011 6273 11023 6307
rect 10965 6267 11023 6273
rect 11701 6307 11759 6313
rect 11701 6273 11713 6307
rect 11747 6273 11759 6307
rect 11701 6267 11759 6273
rect 11793 6307 11851 6313
rect 11793 6273 11805 6307
rect 11839 6273 11851 6307
rect 12066 6304 12072 6316
rect 12027 6276 12072 6304
rect 11793 6267 11851 6273
rect 9677 6239 9735 6245
rect 9677 6205 9689 6239
rect 9723 6236 9735 6239
rect 10229 6239 10287 6245
rect 10229 6236 10241 6239
rect 9723 6208 10241 6236
rect 9723 6205 9735 6208
rect 9677 6199 9735 6205
rect 10229 6205 10241 6208
rect 10275 6205 10287 6239
rect 10229 6199 10287 6205
rect 10321 6239 10379 6245
rect 10321 6205 10333 6239
rect 10367 6205 10379 6239
rect 10321 6199 10379 6205
rect 10502 6196 10508 6248
rect 10560 6236 10566 6248
rect 10869 6239 10927 6245
rect 10869 6236 10881 6239
rect 10560 6208 10881 6236
rect 10560 6196 10566 6208
rect 10869 6205 10881 6208
rect 10915 6205 10927 6239
rect 10869 6199 10927 6205
rect 10980 6168 11008 6267
rect 11146 6196 11152 6248
rect 11204 6236 11210 6248
rect 11808 6236 11836 6267
rect 12066 6264 12072 6276
rect 12124 6264 12130 6316
rect 12253 6307 12311 6313
rect 12253 6273 12265 6307
rect 12299 6273 12311 6307
rect 12253 6267 12311 6273
rect 12268 6236 12296 6267
rect 12342 6264 12348 6316
rect 12400 6304 12406 6316
rect 12713 6307 12771 6313
rect 12713 6304 12725 6307
rect 12400 6276 12725 6304
rect 12400 6264 12406 6276
rect 12713 6273 12725 6276
rect 12759 6273 12771 6307
rect 12713 6267 12771 6273
rect 13262 6236 13268 6248
rect 11204 6208 12296 6236
rect 13223 6208 13268 6236
rect 11204 6196 11210 6208
rect 11606 6168 11612 6180
rect 7944 6140 11008 6168
rect 11567 6140 11612 6168
rect 11606 6128 11612 6140
rect 11664 6128 11670 6180
rect 4614 6100 4620 6112
rect 3988 6072 4620 6100
rect 2869 6063 2927 6069
rect 4614 6060 4620 6072
rect 4672 6060 4678 6112
rect 9766 6100 9772 6112
rect 9727 6072 9772 6100
rect 9766 6060 9772 6072
rect 9824 6060 9830 6112
rect 12066 6060 12072 6112
rect 12124 6100 12130 6112
rect 12268 6100 12296 6208
rect 13262 6196 13268 6208
rect 13320 6196 13326 6248
rect 12437 6103 12495 6109
rect 12437 6100 12449 6103
rect 12124 6072 12449 6100
rect 12124 6060 12130 6072
rect 12437 6069 12449 6072
rect 12483 6100 12495 6103
rect 13357 6103 13415 6109
rect 13357 6100 13369 6103
rect 12483 6072 13369 6100
rect 12483 6069 12495 6072
rect 12437 6063 12495 6069
rect 13357 6069 13369 6072
rect 13403 6069 13415 6103
rect 13357 6063 13415 6069
rect 1104 6010 13892 6032
rect 1104 5958 4214 6010
rect 4266 5958 4278 6010
rect 4330 5958 4342 6010
rect 4394 5958 4406 6010
rect 4458 5958 4470 6010
rect 4522 5958 12214 6010
rect 12266 5958 12278 6010
rect 12330 5958 12342 6010
rect 12394 5958 12406 6010
rect 12458 5958 12470 6010
rect 12522 5958 13892 6010
rect 1104 5936 13892 5958
rect 1578 5856 1584 5908
rect 1636 5896 1642 5908
rect 2682 5896 2688 5908
rect 1636 5868 2688 5896
rect 1636 5856 1642 5868
rect 2682 5856 2688 5868
rect 2740 5896 2746 5908
rect 5350 5896 5356 5908
rect 2740 5868 3832 5896
rect 5311 5868 5356 5896
rect 2740 5856 2746 5868
rect 2314 5828 2320 5840
rect 2275 5800 2320 5828
rect 2314 5788 2320 5800
rect 2372 5788 2378 5840
rect 3804 5837 3832 5868
rect 5350 5856 5356 5868
rect 5408 5856 5414 5908
rect 5718 5896 5724 5908
rect 5552 5868 5724 5896
rect 3789 5831 3847 5837
rect 3789 5797 3801 5831
rect 3835 5797 3847 5831
rect 3789 5791 3847 5797
rect 4062 5788 4068 5840
rect 4120 5828 4126 5840
rect 5552 5828 5580 5868
rect 5718 5856 5724 5868
rect 5776 5856 5782 5908
rect 8021 5899 8079 5905
rect 8021 5865 8033 5899
rect 8067 5896 8079 5899
rect 8110 5896 8116 5908
rect 8067 5868 8116 5896
rect 8067 5865 8079 5868
rect 8021 5859 8079 5865
rect 8110 5856 8116 5868
rect 8168 5856 8174 5908
rect 10137 5899 10195 5905
rect 10137 5865 10149 5899
rect 10183 5896 10195 5899
rect 10318 5896 10324 5908
rect 10183 5868 10324 5896
rect 10183 5865 10195 5868
rect 10137 5859 10195 5865
rect 10318 5856 10324 5868
rect 10376 5896 10382 5908
rect 10686 5896 10692 5908
rect 10376 5868 10692 5896
rect 10376 5856 10382 5868
rect 10686 5856 10692 5868
rect 10744 5856 10750 5908
rect 13262 5896 13268 5908
rect 13223 5868 13268 5896
rect 13262 5856 13268 5868
rect 13320 5856 13326 5908
rect 4120 5800 5580 5828
rect 4120 5788 4126 5800
rect 1394 5720 1400 5772
rect 1452 5760 1458 5772
rect 2133 5763 2191 5769
rect 2133 5760 2145 5763
rect 1452 5732 2145 5760
rect 1452 5720 1458 5732
rect 2133 5729 2145 5732
rect 2179 5729 2191 5763
rect 2774 5760 2780 5772
rect 2133 5723 2191 5729
rect 2746 5720 2780 5760
rect 2832 5720 2838 5772
rect 3142 5720 3148 5772
rect 3200 5760 3206 5772
rect 4614 5760 4620 5772
rect 3200 5732 4620 5760
rect 3200 5720 3206 5732
rect 1486 5692 1492 5704
rect 1447 5664 1492 5692
rect 1486 5652 1492 5664
rect 1544 5652 1550 5704
rect 1578 5652 1584 5704
rect 1636 5692 1642 5704
rect 1765 5695 1823 5701
rect 1636 5664 1681 5692
rect 1636 5652 1642 5664
rect 1765 5661 1777 5695
rect 1811 5692 1823 5695
rect 2038 5692 2044 5704
rect 1811 5664 2044 5692
rect 1811 5661 1823 5664
rect 1765 5655 1823 5661
rect 2038 5652 2044 5664
rect 2096 5692 2102 5704
rect 2409 5695 2467 5701
rect 2409 5692 2421 5695
rect 2096 5664 2421 5692
rect 2096 5652 2102 5664
rect 2409 5661 2421 5664
rect 2455 5661 2467 5695
rect 2409 5655 2467 5661
rect 2593 5695 2651 5701
rect 2593 5661 2605 5695
rect 2639 5692 2651 5695
rect 2746 5692 2774 5720
rect 3436 5701 3464 5732
rect 4614 5720 4620 5732
rect 4672 5720 4678 5772
rect 5552 5769 5580 5800
rect 8481 5831 8539 5837
rect 8481 5797 8493 5831
rect 8527 5828 8539 5831
rect 8754 5828 8760 5840
rect 8527 5800 8760 5828
rect 8527 5797 8539 5800
rect 8481 5791 8539 5797
rect 8754 5788 8760 5800
rect 8812 5788 8818 5840
rect 5537 5763 5595 5769
rect 5537 5729 5549 5763
rect 5583 5729 5595 5763
rect 5537 5723 5595 5729
rect 5721 5763 5779 5769
rect 5721 5729 5733 5763
rect 5767 5760 5779 5763
rect 5994 5760 6000 5772
rect 5767 5732 6000 5760
rect 5767 5729 5779 5732
rect 5721 5723 5779 5729
rect 5994 5720 6000 5732
rect 6052 5720 6058 5772
rect 7742 5720 7748 5772
rect 7800 5760 7806 5772
rect 7800 5732 9076 5760
rect 7800 5720 7806 5732
rect 2961 5695 3019 5701
rect 2961 5692 2973 5695
rect 2639 5664 2973 5692
rect 2639 5661 2651 5664
rect 2593 5655 2651 5661
rect 2961 5661 2973 5664
rect 3007 5661 3019 5695
rect 2961 5655 3019 5661
rect 3421 5695 3479 5701
rect 3421 5661 3433 5695
rect 3467 5661 3479 5695
rect 3421 5655 3479 5661
rect 3513 5695 3571 5701
rect 3513 5661 3525 5695
rect 3559 5692 3571 5695
rect 4706 5692 4712 5704
rect 3559 5664 4200 5692
rect 4667 5664 4712 5692
rect 3559 5661 3571 5664
rect 3513 5655 3571 5661
rect 2777 5627 2835 5633
rect 2777 5593 2789 5627
rect 2823 5624 2835 5627
rect 2866 5624 2872 5636
rect 2823 5596 2872 5624
rect 2823 5593 2835 5596
rect 2777 5587 2835 5593
rect 2866 5584 2872 5596
rect 2924 5584 2930 5636
rect 3237 5627 3295 5633
rect 3237 5593 3249 5627
rect 3283 5624 3295 5627
rect 3283 5596 3464 5624
rect 3283 5593 3295 5596
rect 3237 5587 3295 5593
rect 3436 5568 3464 5596
rect 3602 5584 3608 5636
rect 3660 5624 3666 5636
rect 3970 5624 3976 5636
rect 3660 5596 3976 5624
rect 3660 5584 3666 5596
rect 3970 5584 3976 5596
rect 4028 5584 4034 5636
rect 1949 5559 2007 5565
rect 1949 5525 1961 5559
rect 1995 5556 2007 5559
rect 2222 5556 2228 5568
rect 1995 5528 2228 5556
rect 1995 5525 2007 5528
rect 1949 5519 2007 5525
rect 2222 5516 2228 5528
rect 2280 5516 2286 5568
rect 3145 5559 3203 5565
rect 3145 5525 3157 5559
rect 3191 5556 3203 5559
rect 3326 5556 3332 5568
rect 3191 5528 3332 5556
rect 3191 5525 3203 5528
rect 3145 5519 3203 5525
rect 3326 5516 3332 5528
rect 3384 5516 3390 5568
rect 3418 5516 3424 5568
rect 3476 5516 3482 5568
rect 4062 5556 4068 5568
rect 4023 5528 4068 5556
rect 4062 5516 4068 5528
rect 4120 5516 4126 5568
rect 4172 5565 4200 5664
rect 4706 5652 4712 5664
rect 4764 5652 4770 5704
rect 4893 5695 4951 5701
rect 4893 5661 4905 5695
rect 4939 5661 4951 5695
rect 4893 5655 4951 5661
rect 5813 5695 5871 5701
rect 5813 5661 5825 5695
rect 5859 5692 5871 5695
rect 5902 5692 5908 5704
rect 5859 5664 5908 5692
rect 5859 5661 5871 5664
rect 5813 5655 5871 5661
rect 4341 5627 4399 5633
rect 4341 5593 4353 5627
rect 4387 5624 4399 5627
rect 4430 5624 4436 5636
rect 4387 5596 4436 5624
rect 4387 5593 4399 5596
rect 4341 5587 4399 5593
rect 4430 5584 4436 5596
rect 4488 5624 4494 5636
rect 4525 5627 4583 5633
rect 4525 5624 4537 5627
rect 4488 5596 4537 5624
rect 4488 5584 4494 5596
rect 4525 5593 4537 5596
rect 4571 5593 4583 5627
rect 4908 5624 4936 5655
rect 5902 5652 5908 5664
rect 5960 5652 5966 5704
rect 6178 5692 6184 5704
rect 6139 5664 6184 5692
rect 6178 5652 6184 5664
rect 6236 5652 6242 5704
rect 6273 5695 6331 5701
rect 6273 5661 6285 5695
rect 6319 5661 6331 5695
rect 8570 5692 8576 5704
rect 8531 5664 8576 5692
rect 6273 5655 6331 5661
rect 6086 5624 6092 5636
rect 4908 5596 6092 5624
rect 4525 5587 4583 5593
rect 5552 5568 5580 5596
rect 6086 5584 6092 5596
rect 6144 5624 6150 5636
rect 6288 5624 6316 5655
rect 8570 5652 8576 5664
rect 8628 5652 8634 5704
rect 9048 5701 9076 5732
rect 10042 5720 10048 5772
rect 10100 5760 10106 5772
rect 10321 5763 10379 5769
rect 10321 5760 10333 5763
rect 10100 5732 10333 5760
rect 10100 5720 10106 5732
rect 10321 5729 10333 5732
rect 10367 5729 10379 5763
rect 10594 5760 10600 5772
rect 10555 5732 10600 5760
rect 10321 5723 10379 5729
rect 10594 5720 10600 5732
rect 10652 5720 10658 5772
rect 8757 5695 8815 5701
rect 8757 5661 8769 5695
rect 8803 5692 8815 5695
rect 8941 5695 8999 5701
rect 8941 5692 8953 5695
rect 8803 5664 8953 5692
rect 8803 5661 8815 5664
rect 8757 5655 8815 5661
rect 8941 5661 8953 5664
rect 8987 5661 8999 5695
rect 8941 5655 8999 5661
rect 9033 5695 9091 5701
rect 9033 5661 9045 5695
rect 9079 5661 9091 5695
rect 9306 5692 9312 5704
rect 9267 5664 9312 5692
rect 9033 5655 9091 5661
rect 9306 5652 9312 5664
rect 9364 5652 9370 5704
rect 9674 5652 9680 5704
rect 9732 5701 9738 5704
rect 9732 5695 9765 5701
rect 9753 5692 9765 5695
rect 9858 5692 9864 5704
rect 9753 5664 9864 5692
rect 9753 5661 9765 5664
rect 9732 5655 9765 5661
rect 9732 5652 9738 5655
rect 9858 5652 9864 5664
rect 9916 5652 9922 5704
rect 10226 5692 10232 5704
rect 10187 5664 10232 5692
rect 10226 5652 10232 5664
rect 10284 5652 10290 5704
rect 11974 5652 11980 5704
rect 12032 5692 12038 5704
rect 12345 5695 12403 5701
rect 12345 5692 12357 5695
rect 12032 5664 12357 5692
rect 12032 5652 12038 5664
rect 12345 5661 12357 5664
rect 12391 5661 12403 5695
rect 12345 5655 12403 5661
rect 12529 5695 12587 5701
rect 12529 5661 12541 5695
rect 12575 5661 12587 5695
rect 12529 5655 12587 5661
rect 6144 5596 6316 5624
rect 8113 5627 8171 5633
rect 6144 5584 6150 5596
rect 8113 5593 8125 5627
rect 8159 5593 8171 5627
rect 8113 5587 8171 5593
rect 8297 5627 8355 5633
rect 8297 5593 8309 5627
rect 8343 5624 8355 5627
rect 9398 5624 9404 5636
rect 8343 5596 9404 5624
rect 8343 5593 8355 5596
rect 8297 5587 8355 5593
rect 4157 5559 4215 5565
rect 4157 5525 4169 5559
rect 4203 5525 4215 5559
rect 4157 5519 4215 5525
rect 5534 5516 5540 5568
rect 5592 5516 5598 5568
rect 8128 5556 8156 5587
rect 9398 5584 9404 5596
rect 9456 5584 9462 5636
rect 11606 5584 11612 5636
rect 11664 5584 11670 5636
rect 11882 5584 11888 5636
rect 11940 5624 11946 5636
rect 12253 5627 12311 5633
rect 12253 5624 12265 5627
rect 11940 5596 12265 5624
rect 11940 5584 11946 5596
rect 12253 5593 12265 5596
rect 12299 5593 12311 5627
rect 12253 5587 12311 5593
rect 8570 5556 8576 5568
rect 8128 5528 8576 5556
rect 8570 5516 8576 5528
rect 8628 5516 8634 5568
rect 9585 5559 9643 5565
rect 9585 5525 9597 5559
rect 9631 5556 9643 5559
rect 9674 5556 9680 5568
rect 9631 5528 9680 5556
rect 9631 5525 9643 5528
rect 9585 5519 9643 5525
rect 9674 5516 9680 5528
rect 9732 5516 9738 5568
rect 9769 5559 9827 5565
rect 9769 5525 9781 5559
rect 9815 5556 9827 5559
rect 10134 5556 10140 5568
rect 9815 5528 10140 5556
rect 9815 5525 9827 5528
rect 9769 5519 9827 5525
rect 10134 5516 10140 5528
rect 10192 5516 10198 5568
rect 11422 5516 11428 5568
rect 11480 5556 11486 5568
rect 12069 5559 12127 5565
rect 12069 5556 12081 5559
rect 11480 5528 12081 5556
rect 11480 5516 11486 5528
rect 12069 5525 12081 5528
rect 12115 5525 12127 5559
rect 12069 5519 12127 5525
rect 12158 5516 12164 5568
rect 12216 5556 12222 5568
rect 12544 5556 12572 5655
rect 12713 5559 12771 5565
rect 12713 5556 12725 5559
rect 12216 5528 12725 5556
rect 12216 5516 12222 5528
rect 12713 5525 12725 5528
rect 12759 5525 12771 5559
rect 13170 5556 13176 5568
rect 13131 5528 13176 5556
rect 12713 5519 12771 5525
rect 13170 5516 13176 5528
rect 13228 5516 13234 5568
rect 1104 5466 13892 5488
rect 1104 5414 8214 5466
rect 8266 5414 8278 5466
rect 8330 5414 8342 5466
rect 8394 5414 8406 5466
rect 8458 5414 8470 5466
rect 8522 5414 13892 5466
rect 1104 5392 13892 5414
rect 2774 5352 2780 5364
rect 2746 5312 2780 5352
rect 2832 5312 2838 5364
rect 4062 5312 4068 5364
rect 4120 5352 4126 5364
rect 8389 5355 8447 5361
rect 4120 5324 5028 5352
rect 4120 5312 4126 5324
rect 1397 5287 1455 5293
rect 1397 5253 1409 5287
rect 1443 5284 1455 5287
rect 1946 5284 1952 5296
rect 1443 5256 1952 5284
rect 1443 5253 1455 5256
rect 1397 5247 1455 5253
rect 1946 5244 1952 5256
rect 2004 5244 2010 5296
rect 2746 5284 2774 5312
rect 2424 5256 2774 5284
rect 3513 5287 3571 5293
rect 1486 5216 1492 5228
rect 1447 5188 1492 5216
rect 1486 5176 1492 5188
rect 1544 5176 1550 5228
rect 1578 5176 1584 5228
rect 1636 5216 1642 5228
rect 1673 5219 1731 5225
rect 1673 5216 1685 5219
rect 1636 5188 1685 5216
rect 1636 5176 1642 5188
rect 1673 5185 1685 5188
rect 1719 5185 1731 5219
rect 2130 5216 2136 5228
rect 2091 5188 2136 5216
rect 1673 5179 1731 5185
rect 2130 5176 2136 5188
rect 2188 5176 2194 5228
rect 2314 5216 2320 5228
rect 2275 5188 2320 5216
rect 2314 5176 2320 5188
rect 2372 5176 2378 5228
rect 2424 5225 2452 5256
rect 3513 5253 3525 5287
rect 3559 5253 3571 5287
rect 3513 5247 3571 5253
rect 2409 5219 2467 5225
rect 2409 5185 2421 5219
rect 2455 5185 2467 5219
rect 2409 5179 2467 5185
rect 2777 5219 2835 5225
rect 2777 5185 2789 5219
rect 2823 5216 2835 5219
rect 3234 5216 3240 5228
rect 2823 5188 3240 5216
rect 2823 5185 2835 5188
rect 2777 5179 2835 5185
rect 3234 5176 3240 5188
rect 3292 5176 3298 5228
rect 3329 5219 3387 5225
rect 3329 5185 3341 5219
rect 3375 5185 3387 5219
rect 3329 5179 3387 5185
rect 3528 5206 3556 5247
rect 3602 5244 3608 5296
rect 3660 5284 3666 5296
rect 4080 5284 4108 5312
rect 4430 5284 4436 5296
rect 3660 5256 3705 5284
rect 3804 5256 4108 5284
rect 4391 5256 4436 5284
rect 3660 5244 3666 5256
rect 3697 5222 3755 5225
rect 3804 5222 3832 5256
rect 4430 5244 4436 5256
rect 4488 5244 4494 5296
rect 4614 5284 4620 5296
rect 4575 5256 4620 5284
rect 4614 5244 4620 5256
rect 4672 5244 4678 5296
rect 5000 5293 5028 5324
rect 8389 5321 8401 5355
rect 8435 5352 8447 5355
rect 8570 5352 8576 5364
rect 8435 5324 8576 5352
rect 8435 5321 8447 5324
rect 8389 5315 8447 5321
rect 8570 5312 8576 5324
rect 8628 5312 8634 5364
rect 11790 5312 11796 5364
rect 11848 5352 11854 5364
rect 12170 5355 12228 5361
rect 12170 5352 12182 5355
rect 11848 5324 12182 5352
rect 11848 5312 11854 5324
rect 12170 5321 12182 5324
rect 12216 5321 12228 5355
rect 12170 5315 12228 5321
rect 4985 5287 5043 5293
rect 4985 5253 4997 5287
rect 5031 5253 5043 5287
rect 4985 5247 5043 5253
rect 5169 5287 5227 5293
rect 5169 5253 5181 5287
rect 5215 5284 5227 5287
rect 5442 5284 5448 5296
rect 5215 5256 5448 5284
rect 5215 5253 5227 5256
rect 5169 5247 5227 5253
rect 5442 5244 5448 5256
rect 5500 5244 5506 5296
rect 5902 5284 5908 5296
rect 5644 5256 5908 5284
rect 3697 5219 3832 5222
rect 3697 5206 3709 5219
rect 3528 5185 3709 5206
rect 3743 5194 3832 5219
rect 4062 5216 4068 5228
rect 3743 5185 3755 5194
rect 4023 5188 4068 5216
rect 3528 5179 3755 5185
rect 2961 5151 3019 5157
rect 2961 5117 2973 5151
rect 3007 5148 3019 5151
rect 3344 5148 3372 5179
rect 3528 5178 3740 5179
rect 4062 5176 4068 5188
rect 4120 5176 4126 5228
rect 4341 5219 4399 5225
rect 4341 5185 4353 5219
rect 4387 5185 4399 5219
rect 5350 5216 5356 5228
rect 5311 5188 5356 5216
rect 4341 5179 4399 5185
rect 4356 5148 4384 5179
rect 5350 5176 5356 5188
rect 5408 5176 5414 5228
rect 5644 5225 5672 5256
rect 5902 5244 5908 5256
rect 5960 5284 5966 5296
rect 8849 5287 8907 5293
rect 8849 5284 8861 5287
rect 5960 5256 6592 5284
rect 5960 5244 5966 5256
rect 5629 5219 5687 5225
rect 5629 5185 5641 5219
rect 5675 5185 5687 5219
rect 5994 5216 6000 5228
rect 5955 5188 6000 5216
rect 5629 5179 5687 5185
rect 5994 5176 6000 5188
rect 6052 5216 6058 5228
rect 6564 5225 6592 5256
rect 7576 5256 8861 5284
rect 7576 5225 7604 5256
rect 8849 5253 8861 5256
rect 8895 5253 8907 5287
rect 10042 5284 10048 5296
rect 8849 5247 8907 5253
rect 9508 5256 10048 5284
rect 6365 5219 6423 5225
rect 6365 5216 6377 5219
rect 6052 5188 6377 5216
rect 6052 5176 6058 5188
rect 6365 5185 6377 5188
rect 6411 5185 6423 5219
rect 6365 5179 6423 5185
rect 6549 5219 6607 5225
rect 6549 5185 6561 5219
rect 6595 5185 6607 5219
rect 7101 5219 7159 5225
rect 7101 5216 7113 5219
rect 6549 5179 6607 5185
rect 6656 5188 7113 5216
rect 4801 5151 4859 5157
rect 4801 5148 4813 5151
rect 3007 5120 3188 5148
rect 3344 5120 4813 5148
rect 3007 5117 3019 5120
rect 2961 5111 3019 5117
rect 2501 5083 2559 5089
rect 2501 5080 2513 5083
rect 2332 5052 2513 5080
rect 2332 5024 2360 5052
rect 2501 5049 2513 5052
rect 2547 5049 2559 5083
rect 2501 5043 2559 5049
rect 1762 4972 1768 5024
rect 1820 5012 1826 5024
rect 1949 5015 2007 5021
rect 1949 5012 1961 5015
rect 1820 4984 1961 5012
rect 1820 4972 1826 4984
rect 1949 4981 1961 4984
rect 1995 4981 2007 5015
rect 2314 5012 2320 5024
rect 2227 4984 2320 5012
rect 1949 4975 2007 4981
rect 2314 4972 2320 4984
rect 2372 4972 2378 5024
rect 3160 5021 3188 5120
rect 4801 5117 4813 5120
rect 4847 5117 4859 5151
rect 4801 5111 4859 5117
rect 3234 5040 3240 5092
rect 3292 5080 3298 5092
rect 6656 5080 6684 5188
rect 7101 5185 7113 5188
rect 7147 5185 7159 5219
rect 7101 5179 7159 5185
rect 7561 5219 7619 5225
rect 7561 5185 7573 5219
rect 7607 5185 7619 5219
rect 7561 5179 7619 5185
rect 6733 5151 6791 5157
rect 6733 5117 6745 5151
rect 6779 5117 6791 5151
rect 7116 5148 7144 5179
rect 8110 5176 8116 5228
rect 8168 5216 8174 5228
rect 8941 5219 8999 5225
rect 8941 5216 8953 5219
rect 8168 5188 8953 5216
rect 8168 5176 8174 5188
rect 8941 5185 8953 5188
rect 8987 5185 8999 5219
rect 8941 5179 8999 5185
rect 9030 5176 9036 5228
rect 9088 5216 9094 5228
rect 9125 5219 9183 5225
rect 9125 5216 9137 5219
rect 9088 5188 9137 5216
rect 9088 5176 9094 5188
rect 9125 5185 9137 5188
rect 9171 5185 9183 5219
rect 9125 5179 9183 5185
rect 7742 5148 7748 5160
rect 7116 5120 7748 5148
rect 6733 5111 6791 5117
rect 3292 5052 6684 5080
rect 6748 5080 6776 5111
rect 7742 5108 7748 5120
rect 7800 5108 7806 5160
rect 7929 5151 7987 5157
rect 7929 5117 7941 5151
rect 7975 5148 7987 5151
rect 8481 5151 8539 5157
rect 8481 5148 8493 5151
rect 7975 5120 8493 5148
rect 7975 5117 7987 5120
rect 7929 5111 7987 5117
rect 8481 5117 8493 5120
rect 8527 5117 8539 5151
rect 8481 5111 8539 5117
rect 8573 5151 8631 5157
rect 8573 5117 8585 5151
rect 8619 5117 8631 5151
rect 8573 5111 8631 5117
rect 7098 5080 7104 5092
rect 6748 5052 7104 5080
rect 3292 5040 3298 5052
rect 7098 5040 7104 5052
rect 7156 5040 7162 5092
rect 3145 5015 3203 5021
rect 3145 4981 3157 5015
rect 3191 5012 3203 5015
rect 3418 5012 3424 5024
rect 3191 4984 3424 5012
rect 3191 4981 3203 4984
rect 3145 4975 3203 4981
rect 3418 4972 3424 4984
rect 3476 4972 3482 5024
rect 3786 5012 3792 5024
rect 3747 4984 3792 5012
rect 3786 4972 3792 4984
rect 3844 4972 3850 5024
rect 5902 4972 5908 5024
rect 5960 5012 5966 5024
rect 5997 5015 6055 5021
rect 5997 5012 6009 5015
rect 5960 4984 6009 5012
rect 5960 4972 5966 4984
rect 5997 4981 6009 4984
rect 6043 4981 6055 5015
rect 5997 4975 6055 4981
rect 7650 4972 7656 5024
rect 7708 5012 7714 5024
rect 8021 5015 8079 5021
rect 8021 5012 8033 5015
rect 7708 4984 8033 5012
rect 7708 4972 7714 4984
rect 8021 4981 8033 4984
rect 8067 4981 8079 5015
rect 8588 5012 8616 5111
rect 8662 5108 8668 5160
rect 8720 5148 8726 5160
rect 9508 5157 9536 5256
rect 10042 5244 10048 5256
rect 10100 5244 10106 5296
rect 11146 5244 11152 5296
rect 11204 5284 11210 5296
rect 11701 5287 11759 5293
rect 11701 5284 11713 5287
rect 11204 5256 11713 5284
rect 11204 5244 11210 5256
rect 11701 5253 11713 5256
rect 11747 5284 11759 5287
rect 12066 5284 12072 5296
rect 11747 5256 12072 5284
rect 11747 5253 11759 5256
rect 11701 5247 11759 5253
rect 11606 5216 11612 5228
rect 10902 5188 11612 5216
rect 11606 5176 11612 5188
rect 11664 5176 11670 5228
rect 11808 5225 11836 5256
rect 12066 5244 12072 5256
rect 12124 5244 12130 5296
rect 13170 5244 13176 5296
rect 13228 5284 13234 5296
rect 13265 5287 13323 5293
rect 13265 5284 13277 5287
rect 13228 5256 13277 5284
rect 13228 5244 13234 5256
rect 13265 5253 13277 5256
rect 13311 5253 13323 5287
rect 13265 5247 13323 5253
rect 11793 5219 11851 5225
rect 11793 5185 11805 5219
rect 11839 5216 11851 5219
rect 12618 5216 12624 5228
rect 11839 5188 11873 5216
rect 12579 5188 12624 5216
rect 11839 5185 11851 5188
rect 11793 5179 11851 5185
rect 12618 5176 12624 5188
rect 12676 5176 12682 5228
rect 13538 5216 13544 5228
rect 13499 5188 13544 5216
rect 13538 5176 13544 5188
rect 13596 5176 13602 5228
rect 9493 5151 9551 5157
rect 9493 5148 9505 5151
rect 8720 5120 9505 5148
rect 8720 5108 8726 5120
rect 9493 5117 9505 5120
rect 9539 5117 9551 5151
rect 9766 5148 9772 5160
rect 9727 5120 9772 5148
rect 9493 5111 9551 5117
rect 9766 5108 9772 5120
rect 9824 5108 9830 5160
rect 11241 5083 11299 5089
rect 11241 5049 11253 5083
rect 11287 5049 11299 5083
rect 11241 5043 11299 5049
rect 9858 5012 9864 5024
rect 8588 4984 9864 5012
rect 8021 4975 8079 4981
rect 9858 4972 9864 4984
rect 9916 4972 9922 5024
rect 10410 4972 10416 5024
rect 10468 5012 10474 5024
rect 11256 5012 11284 5043
rect 12161 5015 12219 5021
rect 12161 5012 12173 5015
rect 10468 4984 12173 5012
rect 10468 4972 10474 4984
rect 12161 4981 12173 4984
rect 12207 4981 12219 5015
rect 12161 4975 12219 4981
rect 12345 5015 12403 5021
rect 12345 4981 12357 5015
rect 12391 5012 12403 5015
rect 12710 5012 12716 5024
rect 12391 4984 12716 5012
rect 12391 4981 12403 4984
rect 12345 4975 12403 4981
rect 12710 4972 12716 4984
rect 12768 4972 12774 5024
rect 1104 4922 13892 4944
rect 1104 4870 4214 4922
rect 4266 4870 4278 4922
rect 4330 4870 4342 4922
rect 4394 4870 4406 4922
rect 4458 4870 4470 4922
rect 4522 4870 12214 4922
rect 12266 4870 12278 4922
rect 12330 4870 12342 4922
rect 12394 4870 12406 4922
rect 12458 4870 12470 4922
rect 12522 4870 13892 4922
rect 1104 4848 13892 4870
rect 1394 4808 1400 4820
rect 1355 4780 1400 4808
rect 1394 4768 1400 4780
rect 1452 4808 1458 4820
rect 2774 4808 2780 4820
rect 1452 4780 2780 4808
rect 1452 4768 1458 4780
rect 2774 4768 2780 4780
rect 2832 4808 2838 4820
rect 3234 4808 3240 4820
rect 2832 4780 3240 4808
rect 2832 4768 2838 4780
rect 3234 4768 3240 4780
rect 3292 4768 3298 4820
rect 5626 4768 5632 4820
rect 5684 4808 5690 4820
rect 6638 4808 6644 4820
rect 5684 4780 6644 4808
rect 5684 4768 5690 4780
rect 6638 4768 6644 4780
rect 6696 4808 6702 4820
rect 6696 4780 6960 4808
rect 6696 4768 6702 4780
rect 6178 4740 6184 4752
rect 6012 4712 6184 4740
rect 2314 4672 2320 4684
rect 2275 4644 2320 4672
rect 2314 4632 2320 4644
rect 2372 4632 2378 4684
rect 3418 4672 3424 4684
rect 3379 4644 3424 4672
rect 3418 4632 3424 4644
rect 3476 4632 3482 4684
rect 5626 4672 5632 4684
rect 5587 4644 5632 4672
rect 5626 4632 5632 4644
rect 5684 4632 5690 4684
rect 1578 4604 1584 4616
rect 1539 4576 1584 4604
rect 1578 4564 1584 4576
rect 1636 4564 1642 4616
rect 1670 4564 1676 4616
rect 1728 4604 1734 4616
rect 1765 4607 1823 4613
rect 1765 4604 1777 4607
rect 1728 4576 1777 4604
rect 1728 4564 1734 4576
rect 1765 4573 1777 4576
rect 1811 4573 1823 4607
rect 2130 4604 2136 4616
rect 2091 4576 2136 4604
rect 1765 4567 1823 4573
rect 2130 4564 2136 4576
rect 2188 4564 2194 4616
rect 2406 4604 2412 4616
rect 2367 4576 2412 4604
rect 2406 4564 2412 4576
rect 2464 4564 2470 4616
rect 3125 4607 3183 4613
rect 3125 4573 3137 4607
rect 3171 4604 3183 4607
rect 3326 4604 3332 4616
rect 3171 4573 3188 4604
rect 3239 4576 3332 4604
rect 3125 4567 3188 4573
rect 2148 4536 2176 4564
rect 2682 4536 2688 4548
rect 2148 4508 2688 4536
rect 2682 4496 2688 4508
rect 2740 4496 2746 4548
rect 2774 4496 2780 4548
rect 2832 4536 2838 4548
rect 2869 4539 2927 4545
rect 2869 4536 2881 4539
rect 2832 4508 2881 4536
rect 2832 4496 2838 4508
rect 2869 4505 2881 4508
rect 2915 4505 2927 4539
rect 3160 4536 3188 4567
rect 3326 4564 3332 4576
rect 3384 4604 3390 4616
rect 3786 4604 3792 4616
rect 3384 4576 3792 4604
rect 3384 4564 3390 4576
rect 3786 4564 3792 4576
rect 3844 4564 3850 4616
rect 4246 4564 4252 4616
rect 4304 4564 4310 4616
rect 5718 4604 5724 4616
rect 5679 4576 5724 4604
rect 5718 4564 5724 4576
rect 5776 4564 5782 4616
rect 5902 4604 5908 4616
rect 5863 4576 5908 4604
rect 5902 4564 5908 4576
rect 5960 4564 5966 4616
rect 6012 4613 6040 4712
rect 6178 4700 6184 4712
rect 6236 4700 6242 4752
rect 6822 4672 6828 4684
rect 6564 4644 6828 4672
rect 5997 4607 6055 4613
rect 5997 4573 6009 4607
rect 6043 4573 6055 4607
rect 5997 4567 6055 4573
rect 6086 4564 6092 4616
rect 6144 4613 6150 4616
rect 6564 4613 6592 4644
rect 6822 4632 6828 4644
rect 6880 4632 6886 4684
rect 6932 4681 6960 4780
rect 8570 4768 8576 4820
rect 8628 4808 8634 4820
rect 8665 4811 8723 4817
rect 8665 4808 8677 4811
rect 8628 4780 8677 4808
rect 8628 4768 8634 4780
rect 8665 4777 8677 4780
rect 8711 4777 8723 4811
rect 8665 4771 8723 4777
rect 6917 4675 6975 4681
rect 6917 4641 6929 4675
rect 6963 4641 6975 4675
rect 6917 4635 6975 4641
rect 7193 4675 7251 4681
rect 7193 4641 7205 4675
rect 7239 4672 7251 4675
rect 7650 4672 7656 4684
rect 7239 4644 7656 4672
rect 7239 4641 7251 4644
rect 7193 4635 7251 4641
rect 7650 4632 7656 4644
rect 7708 4632 7714 4684
rect 7742 4632 7748 4684
rect 7800 4672 7806 4684
rect 8680 4672 8708 4771
rect 9398 4768 9404 4820
rect 9456 4808 9462 4820
rect 9493 4811 9551 4817
rect 9493 4808 9505 4811
rect 9456 4780 9505 4808
rect 9456 4768 9462 4780
rect 9493 4777 9505 4780
rect 9539 4777 9551 4811
rect 9493 4771 9551 4777
rect 10226 4768 10232 4820
rect 10284 4808 10290 4820
rect 11977 4811 12035 4817
rect 11977 4808 11989 4811
rect 10284 4780 11989 4808
rect 10284 4768 10290 4780
rect 11977 4777 11989 4780
rect 12023 4777 12035 4811
rect 11977 4771 12035 4777
rect 9674 4700 9680 4752
rect 9732 4740 9738 4752
rect 13170 4740 13176 4752
rect 9732 4712 10364 4740
rect 13131 4712 13176 4740
rect 9732 4700 9738 4712
rect 7800 4644 8432 4672
rect 8680 4644 9536 4672
rect 7800 4632 7806 4644
rect 6144 4607 6181 4613
rect 6169 4573 6181 4607
rect 6144 4567 6181 4573
rect 6549 4607 6607 4613
rect 6549 4573 6561 4607
rect 6595 4573 6607 4607
rect 6730 4604 6736 4616
rect 6691 4576 6736 4604
rect 6549 4567 6607 4573
rect 6144 4564 6150 4567
rect 6730 4564 6736 4576
rect 6788 4564 6794 4616
rect 8404 4604 8432 4644
rect 9033 4607 9091 4613
rect 9033 4604 9045 4607
rect 8404 4576 9045 4604
rect 9033 4573 9045 4576
rect 9079 4573 9091 4607
rect 9033 4567 9091 4573
rect 9122 4564 9128 4616
rect 9180 4604 9186 4616
rect 9508 4613 9536 4644
rect 10042 4632 10048 4684
rect 10100 4672 10106 4684
rect 10229 4675 10287 4681
rect 10229 4672 10241 4675
rect 10100 4644 10241 4672
rect 10100 4632 10106 4644
rect 10229 4641 10241 4644
rect 10275 4641 10287 4675
rect 10336 4672 10364 4712
rect 13170 4700 13176 4712
rect 13228 4700 13234 4752
rect 10505 4675 10563 4681
rect 10505 4672 10517 4675
rect 10336 4644 10517 4672
rect 10229 4635 10287 4641
rect 10505 4641 10517 4644
rect 10551 4641 10563 4675
rect 10505 4635 10563 4641
rect 9493 4607 9551 4613
rect 9180 4576 9225 4604
rect 9180 4564 9186 4576
rect 9493 4573 9505 4607
rect 9539 4573 9551 4607
rect 9493 4567 9551 4573
rect 12526 4564 12532 4616
rect 12584 4604 12590 4616
rect 12713 4607 12771 4613
rect 12713 4604 12725 4607
rect 12584 4576 12725 4604
rect 12584 4564 12590 4576
rect 12713 4573 12725 4576
rect 12759 4573 12771 4607
rect 13538 4604 13544 4616
rect 13499 4576 13544 4604
rect 12713 4567 12771 4573
rect 13538 4564 13544 4576
rect 13596 4564 13602 4616
rect 5353 4539 5411 4545
rect 3160 4508 3556 4536
rect 2869 4499 2927 4505
rect 3528 4480 3556 4508
rect 5353 4505 5365 4539
rect 5399 4505 5411 4539
rect 5353 4499 5411 4505
rect 6365 4539 6423 4545
rect 6365 4505 6377 4539
rect 6411 4536 6423 4539
rect 7190 4536 7196 4548
rect 6411 4508 7196 4536
rect 6411 4505 6423 4508
rect 6365 4499 6423 4505
rect 2225 4471 2283 4477
rect 2225 4437 2237 4471
rect 2271 4468 2283 4471
rect 2314 4468 2320 4480
rect 2271 4440 2320 4468
rect 2271 4437 2283 4440
rect 2225 4431 2283 4437
rect 2314 4428 2320 4440
rect 2372 4428 2378 4480
rect 3234 4468 3240 4480
rect 3195 4440 3240 4468
rect 3234 4428 3240 4440
rect 3292 4428 3298 4480
rect 3510 4468 3516 4480
rect 3471 4440 3516 4468
rect 3510 4428 3516 4440
rect 3568 4428 3574 4480
rect 3881 4471 3939 4477
rect 3881 4437 3893 4471
rect 3927 4468 3939 4471
rect 4522 4468 4528 4480
rect 3927 4440 4528 4468
rect 3927 4437 3939 4440
rect 3881 4431 3939 4437
rect 4522 4428 4528 4440
rect 4580 4428 4586 4480
rect 5368 4468 5396 4499
rect 7190 4496 7196 4508
rect 7248 4496 7254 4548
rect 11882 4536 11888 4548
rect 7300 4508 7682 4536
rect 11730 4508 11888 4536
rect 5534 4468 5540 4480
rect 5368 4440 5540 4468
rect 5534 4428 5540 4440
rect 5592 4428 5598 4480
rect 6733 4471 6791 4477
rect 6733 4437 6745 4471
rect 6779 4468 6791 4471
rect 7300 4468 7328 4508
rect 11882 4496 11888 4508
rect 11940 4496 11946 4548
rect 13265 4539 13323 4545
rect 13265 4505 13277 4539
rect 13311 4505 13323 4539
rect 13265 4499 13323 4505
rect 9674 4468 9680 4480
rect 6779 4440 7328 4468
rect 9635 4440 9680 4468
rect 6779 4437 6791 4440
rect 6733 4431 6791 4437
rect 9674 4428 9680 4440
rect 9732 4428 9738 4480
rect 13280 4468 13308 4499
rect 13357 4471 13415 4477
rect 13357 4468 13369 4471
rect 13280 4440 13369 4468
rect 13357 4437 13369 4440
rect 13403 4437 13415 4471
rect 13357 4431 13415 4437
rect 1104 4378 13892 4400
rect 1104 4326 8214 4378
rect 8266 4326 8278 4378
rect 8330 4326 8342 4378
rect 8394 4326 8406 4378
rect 8458 4326 8470 4378
rect 8522 4326 13892 4378
rect 1104 4304 13892 4326
rect 2406 4224 2412 4276
rect 2464 4264 2470 4276
rect 3329 4267 3387 4273
rect 3329 4264 3341 4267
rect 2464 4236 3341 4264
rect 2464 4224 2470 4236
rect 3329 4233 3341 4236
rect 3375 4233 3387 4267
rect 3329 4227 3387 4233
rect 4617 4267 4675 4273
rect 4617 4233 4629 4267
rect 4663 4233 4675 4267
rect 4617 4227 4675 4233
rect 2774 4156 2780 4208
rect 2832 4196 2838 4208
rect 2832 4168 3372 4196
rect 2832 4156 2838 4168
rect 1854 4128 1860 4140
rect 1815 4100 1860 4128
rect 1854 4088 1860 4100
rect 1912 4088 1918 4140
rect 2038 4128 2044 4140
rect 1999 4100 2044 4128
rect 2038 4088 2044 4100
rect 2096 4088 2102 4140
rect 2222 4128 2228 4140
rect 2183 4100 2228 4128
rect 2222 4088 2228 4100
rect 2280 4088 2286 4140
rect 2314 4088 2320 4140
rect 2372 4128 2378 4140
rect 2682 4128 2688 4140
rect 2372 4100 2417 4128
rect 2643 4100 2688 4128
rect 2372 4088 2378 4100
rect 2682 4088 2688 4100
rect 2740 4088 2746 4140
rect 2866 4128 2872 4140
rect 2827 4100 2872 4128
rect 2866 4088 2872 4100
rect 2924 4088 2930 4140
rect 3344 4137 3372 4168
rect 3694 4156 3700 4208
rect 3752 4196 3758 4208
rect 4632 4196 4660 4227
rect 4706 4224 4712 4276
rect 4764 4264 4770 4276
rect 5077 4267 5135 4273
rect 5077 4264 5089 4267
rect 4764 4236 5089 4264
rect 4764 4224 4770 4236
rect 5077 4233 5089 4236
rect 5123 4264 5135 4267
rect 5350 4264 5356 4276
rect 5123 4236 5356 4264
rect 5123 4233 5135 4236
rect 5077 4227 5135 4233
rect 5350 4224 5356 4236
rect 5408 4224 5414 4276
rect 5534 4264 5540 4276
rect 5495 4236 5540 4264
rect 5534 4224 5540 4236
rect 5592 4224 5598 4276
rect 6086 4224 6092 4276
rect 6144 4264 6150 4276
rect 6457 4267 6515 4273
rect 6457 4264 6469 4267
rect 6144 4236 6469 4264
rect 6144 4224 6150 4236
rect 6457 4233 6469 4236
rect 6503 4233 6515 4267
rect 6457 4227 6515 4233
rect 6638 4224 6644 4276
rect 6696 4264 6702 4276
rect 6696 4236 8248 4264
rect 6696 4224 6702 4236
rect 5718 4196 5724 4208
rect 3752 4168 4108 4196
rect 4632 4168 5724 4196
rect 3752 4156 3758 4168
rect 3329 4131 3387 4137
rect 3329 4097 3341 4131
rect 3375 4097 3387 4131
rect 3510 4128 3516 4140
rect 3471 4100 3516 4128
rect 3329 4091 3387 4097
rect 3510 4088 3516 4100
rect 3568 4088 3574 4140
rect 4080 4137 4108 4168
rect 5718 4156 5724 4168
rect 5776 4156 5782 4208
rect 6181 4199 6239 4205
rect 6181 4165 6193 4199
rect 6227 4196 6239 4199
rect 6227 4168 6762 4196
rect 6227 4165 6239 4168
rect 6181 4159 6239 4165
rect 3973 4131 4031 4137
rect 3973 4097 3985 4131
rect 4019 4097 4031 4131
rect 3973 4091 4031 4097
rect 4065 4131 4123 4137
rect 4065 4097 4077 4131
rect 4111 4097 4123 4131
rect 4246 4128 4252 4140
rect 4207 4100 4252 4128
rect 4065 4091 4123 4097
rect 1762 4060 1768 4072
rect 1723 4032 1768 4060
rect 1762 4020 1768 4032
rect 1820 4020 1826 4072
rect 2057 4032 3372 4060
rect 1489 3995 1547 4001
rect 1489 3961 1501 3995
rect 1535 3992 1547 3995
rect 2057 3992 2085 4032
rect 1535 3964 2085 3992
rect 2133 3995 2191 4001
rect 1535 3961 1547 3964
rect 1489 3955 1547 3961
rect 2133 3961 2145 3995
rect 2179 3992 2191 3995
rect 3053 3995 3111 4001
rect 3053 3992 3065 3995
rect 2179 3964 3065 3992
rect 2179 3961 2191 3964
rect 2133 3955 2191 3961
rect 3053 3961 3065 3964
rect 3099 3961 3111 3995
rect 3053 3955 3111 3961
rect 1857 3927 1915 3933
rect 1857 3893 1869 3927
rect 1903 3924 1915 3927
rect 2222 3924 2228 3936
rect 1903 3896 2228 3924
rect 1903 3893 1915 3896
rect 1857 3887 1915 3893
rect 2222 3884 2228 3896
rect 2280 3884 2286 3936
rect 2501 3927 2559 3933
rect 2501 3893 2513 3927
rect 2547 3924 2559 3927
rect 3142 3924 3148 3936
rect 2547 3896 3148 3924
rect 2547 3893 2559 3896
rect 2501 3887 2559 3893
rect 3142 3884 3148 3896
rect 3200 3884 3206 3936
rect 3344 3924 3372 4032
rect 3418 3952 3424 4004
rect 3476 3992 3482 4004
rect 3789 3995 3847 4001
rect 3789 3992 3801 3995
rect 3476 3964 3801 3992
rect 3476 3952 3482 3964
rect 3789 3961 3801 3964
rect 3835 3992 3847 3995
rect 3988 3992 4016 4091
rect 4246 4088 4252 4100
rect 4304 4088 4310 4140
rect 4522 4128 4528 4140
rect 4483 4100 4528 4128
rect 4522 4088 4528 4100
rect 4580 4088 4586 4140
rect 4709 4131 4767 4137
rect 4709 4097 4721 4131
rect 4755 4128 4767 4131
rect 5169 4131 5227 4137
rect 5169 4128 5181 4131
rect 4755 4100 5181 4128
rect 4755 4097 4767 4100
rect 4709 4091 4767 4097
rect 5169 4097 5181 4100
rect 5215 4128 5227 4131
rect 5442 4128 5448 4140
rect 5215 4100 5448 4128
rect 5215 4097 5227 4100
rect 5169 4091 5227 4097
rect 5442 4088 5448 4100
rect 5500 4088 5506 4140
rect 5813 4131 5871 4137
rect 5813 4097 5825 4131
rect 5859 4097 5871 4131
rect 5813 4091 5871 4097
rect 6089 4131 6147 4137
rect 6089 4097 6101 4131
rect 6135 4128 6147 4131
rect 6638 4128 6644 4140
rect 6135 4100 6644 4128
rect 6135 4097 6147 4100
rect 6089 4091 6147 4097
rect 4890 4060 4896 4072
rect 4851 4032 4896 4060
rect 4890 4020 4896 4032
rect 4948 4020 4954 4072
rect 4798 3992 4804 4004
rect 3835 3964 4804 3992
rect 3835 3961 3847 3964
rect 3789 3955 3847 3961
rect 4798 3952 4804 3964
rect 4856 3952 4862 4004
rect 4982 3952 4988 4004
rect 5040 3992 5046 4004
rect 5721 3995 5779 4001
rect 5721 3992 5733 3995
rect 5040 3964 5733 3992
rect 5040 3952 5046 3964
rect 5721 3961 5733 3964
rect 5767 3992 5779 3995
rect 5828 3992 5856 4091
rect 6638 4088 6644 4100
rect 6696 4088 6702 4140
rect 8220 4137 8248 4236
rect 8570 4224 8576 4276
rect 8628 4224 8634 4276
rect 9674 4264 9680 4276
rect 9635 4236 9680 4264
rect 9674 4224 9680 4236
rect 9732 4224 9738 4276
rect 9858 4224 9864 4276
rect 9916 4264 9922 4276
rect 11146 4264 11152 4276
rect 9916 4236 10824 4264
rect 11107 4236 11152 4264
rect 9916 4224 9922 4236
rect 8205 4131 8263 4137
rect 8205 4097 8217 4131
rect 8251 4128 8263 4131
rect 8478 4128 8484 4140
rect 8251 4100 8484 4128
rect 8251 4097 8263 4100
rect 8205 4091 8263 4097
rect 8478 4088 8484 4100
rect 8536 4088 8542 4140
rect 8588 4128 8616 4224
rect 9398 4196 9404 4208
rect 9048 4168 9404 4196
rect 9048 4137 9076 4168
rect 9398 4156 9404 4168
rect 9456 4196 9462 4208
rect 10796 4196 10824 4236
rect 11146 4224 11152 4236
rect 11204 4264 11210 4276
rect 11241 4267 11299 4273
rect 11241 4264 11253 4267
rect 11204 4236 11253 4264
rect 11204 4224 11210 4236
rect 11241 4233 11253 4236
rect 11287 4233 11299 4267
rect 11606 4264 11612 4276
rect 11567 4236 11612 4264
rect 11241 4227 11299 4233
rect 11256 4196 11284 4227
rect 11606 4224 11612 4236
rect 11664 4224 11670 4276
rect 11974 4196 11980 4208
rect 9456 4168 10456 4196
rect 10796 4168 10916 4196
rect 11256 4168 11980 4196
rect 9456 4156 9462 4168
rect 8757 4131 8815 4137
rect 8757 4128 8769 4131
rect 8588 4100 8769 4128
rect 8757 4097 8769 4100
rect 8803 4097 8815 4131
rect 8757 4091 8815 4097
rect 9033 4131 9091 4137
rect 9033 4097 9045 4131
rect 9079 4097 9091 4131
rect 9033 4091 9091 4097
rect 9493 4131 9551 4137
rect 9493 4097 9505 4131
rect 9539 4097 9551 4131
rect 9493 4091 9551 4097
rect 7190 4020 7196 4072
rect 7248 4060 7254 4072
rect 7929 4063 7987 4069
rect 7929 4060 7941 4063
rect 7248 4032 7941 4060
rect 7248 4020 7254 4032
rect 7929 4029 7941 4032
rect 7975 4029 7987 4063
rect 9508 4060 9536 4091
rect 9582 4088 9588 4140
rect 9640 4128 9646 4140
rect 9968 4137 9996 4168
rect 9953 4131 10011 4137
rect 9640 4100 9685 4128
rect 9640 4088 9646 4100
rect 9953 4097 9965 4131
rect 9999 4097 10011 4131
rect 9953 4091 10011 4097
rect 10045 4131 10103 4137
rect 10045 4097 10057 4131
rect 10091 4128 10103 4131
rect 10318 4128 10324 4140
rect 10091 4100 10324 4128
rect 10091 4097 10103 4100
rect 10045 4091 10103 4097
rect 10060 4060 10088 4091
rect 10318 4088 10324 4100
rect 10376 4088 10382 4140
rect 10428 4128 10456 4168
rect 10778 4128 10784 4140
rect 10428 4100 10784 4128
rect 10778 4088 10784 4100
rect 10836 4088 10842 4140
rect 10888 4137 10916 4168
rect 11808 4137 11836 4168
rect 11974 4156 11980 4168
rect 12032 4196 12038 4208
rect 12526 4196 12532 4208
rect 12032 4168 12296 4196
rect 12487 4168 12532 4196
rect 12032 4156 12038 4168
rect 10873 4131 10931 4137
rect 10873 4097 10885 4131
rect 10919 4097 10931 4131
rect 10873 4091 10931 4097
rect 11609 4131 11667 4137
rect 11609 4097 11621 4131
rect 11655 4097 11667 4131
rect 11609 4091 11667 4097
rect 11793 4131 11851 4137
rect 11793 4097 11805 4131
rect 11839 4097 11851 4131
rect 12066 4128 12072 4140
rect 12027 4100 12072 4128
rect 11793 4091 11851 4097
rect 7929 4023 7987 4029
rect 8266 4032 9536 4060
rect 9784 4032 10088 4060
rect 10229 4063 10287 4069
rect 6822 3992 6828 4004
rect 5767 3964 6828 3992
rect 5767 3961 5779 3964
rect 5721 3955 5779 3961
rect 6822 3952 6828 3964
rect 6880 3952 6886 4004
rect 8266 3924 8294 4032
rect 8573 3995 8631 4001
rect 8573 3961 8585 3995
rect 8619 3992 8631 3995
rect 9214 3992 9220 4004
rect 8619 3964 9220 3992
rect 8619 3961 8631 3964
rect 8573 3955 8631 3961
rect 9214 3952 9220 3964
rect 9272 3952 9278 4004
rect 9309 3995 9367 4001
rect 9309 3961 9321 3995
rect 9355 3992 9367 3995
rect 9784 3992 9812 4032
rect 10229 4029 10241 4063
rect 10275 4060 10287 4063
rect 10597 4063 10655 4069
rect 10597 4060 10609 4063
rect 10275 4032 10609 4060
rect 10275 4029 10287 4032
rect 10229 4023 10287 4029
rect 10597 4029 10609 4032
rect 10643 4029 10655 4063
rect 10597 4023 10655 4029
rect 9355 3964 9812 3992
rect 9861 3995 9919 4001
rect 9355 3961 9367 3964
rect 9309 3955 9367 3961
rect 9861 3961 9873 3995
rect 9907 3992 9919 3995
rect 9950 3992 9956 4004
rect 9907 3964 9956 3992
rect 9907 3961 9919 3964
rect 9861 3955 9919 3961
rect 9950 3952 9956 3964
rect 10008 3952 10014 4004
rect 11624 3992 11652 4091
rect 12066 4088 12072 4100
rect 12124 4088 12130 4140
rect 12268 4137 12296 4168
rect 12526 4156 12532 4168
rect 12584 4156 12590 4208
rect 12253 4131 12311 4137
rect 12253 4097 12265 4131
rect 12299 4128 12311 4131
rect 12710 4128 12716 4140
rect 12299 4100 12434 4128
rect 12671 4100 12716 4128
rect 12299 4097 12311 4100
rect 12253 4091 12311 4097
rect 11698 4020 11704 4072
rect 11756 4060 11762 4072
rect 11977 4063 12035 4069
rect 11977 4060 11989 4063
rect 11756 4032 11989 4060
rect 11756 4020 11762 4032
rect 11977 4029 11989 4032
rect 12023 4029 12035 4063
rect 11977 4023 12035 4029
rect 12084 3992 12112 4088
rect 12406 4060 12434 4100
rect 12710 4088 12716 4100
rect 12768 4088 12774 4140
rect 12897 4131 12955 4137
rect 12897 4097 12909 4131
rect 12943 4097 12955 4131
rect 12897 4091 12955 4097
rect 12989 4131 13047 4137
rect 12989 4097 13001 4131
rect 13035 4128 13047 4131
rect 13354 4128 13360 4140
rect 13035 4100 13360 4128
rect 13035 4097 13047 4100
rect 12989 4091 13047 4097
rect 12912 4060 12940 4091
rect 13354 4088 13360 4100
rect 13412 4088 13418 4140
rect 13081 4063 13139 4069
rect 13081 4060 13093 4063
rect 12406 4032 13093 4060
rect 13081 4029 13093 4032
rect 13127 4029 13139 4063
rect 13081 4023 13139 4029
rect 11624 3964 12112 3992
rect 3344 3896 8294 3924
rect 8941 3927 8999 3933
rect 8941 3893 8953 3927
rect 8987 3924 8999 3927
rect 9030 3924 9036 3936
rect 8987 3896 9036 3924
rect 8987 3893 8999 3896
rect 8941 3887 8999 3893
rect 9030 3884 9036 3896
rect 9088 3884 9094 3936
rect 10318 3884 10324 3936
rect 10376 3924 10382 3936
rect 10413 3927 10471 3933
rect 10413 3924 10425 3927
rect 10376 3896 10425 3924
rect 10376 3884 10382 3896
rect 10413 3893 10425 3896
rect 10459 3893 10471 3927
rect 13354 3924 13360 3936
rect 13315 3896 13360 3924
rect 10413 3887 10471 3893
rect 13354 3884 13360 3896
rect 13412 3884 13418 3936
rect 1104 3834 13892 3856
rect 1104 3782 4214 3834
rect 4266 3782 4278 3834
rect 4330 3782 4342 3834
rect 4394 3782 4406 3834
rect 4458 3782 4470 3834
rect 4522 3782 12214 3834
rect 12266 3782 12278 3834
rect 12330 3782 12342 3834
rect 12394 3782 12406 3834
rect 12458 3782 12470 3834
rect 12522 3782 13892 3834
rect 1104 3760 13892 3782
rect 1489 3723 1547 3729
rect 1489 3689 1501 3723
rect 1535 3720 1547 3723
rect 1670 3720 1676 3732
rect 1535 3692 1676 3720
rect 1535 3689 1547 3692
rect 1489 3683 1547 3689
rect 1670 3680 1676 3692
rect 1728 3720 1734 3732
rect 2225 3723 2283 3729
rect 2225 3720 2237 3723
rect 1728 3692 2237 3720
rect 1728 3680 1734 3692
rect 2225 3689 2237 3692
rect 2271 3689 2283 3723
rect 6457 3723 6515 3729
rect 6457 3720 6469 3723
rect 2225 3683 2283 3689
rect 3344 3692 6469 3720
rect 2130 3612 2136 3664
rect 2188 3652 2194 3664
rect 3344 3652 3372 3692
rect 6457 3689 6469 3692
rect 6503 3720 6515 3723
rect 6641 3723 6699 3729
rect 6641 3720 6653 3723
rect 6503 3692 6653 3720
rect 6503 3689 6515 3692
rect 6457 3683 6515 3689
rect 6641 3689 6653 3692
rect 6687 3689 6699 3723
rect 6641 3683 6699 3689
rect 6730 3680 6736 3732
rect 6788 3720 6794 3732
rect 9582 3720 9588 3732
rect 6788 3692 9076 3720
rect 9543 3692 9588 3720
rect 6788 3680 6794 3692
rect 5997 3655 6055 3661
rect 5997 3652 6009 3655
rect 2188 3624 3372 3652
rect 3436 3624 6009 3652
rect 2188 3612 2194 3624
rect 1857 3587 1915 3593
rect 1857 3553 1869 3587
rect 1903 3584 1915 3587
rect 2038 3584 2044 3596
rect 1903 3556 2044 3584
rect 1903 3553 1915 3556
rect 1857 3547 1915 3553
rect 2038 3544 2044 3556
rect 2096 3544 2102 3596
rect 2593 3587 2651 3593
rect 2593 3553 2605 3587
rect 2639 3584 2651 3587
rect 2774 3584 2780 3596
rect 2639 3556 2780 3584
rect 2639 3553 2651 3556
rect 2593 3547 2651 3553
rect 2774 3544 2780 3556
rect 2832 3544 2838 3596
rect 3436 3593 3464 3624
rect 5997 3621 6009 3624
rect 6043 3621 6055 3655
rect 5997 3615 6055 3621
rect 3421 3587 3479 3593
rect 3421 3553 3433 3587
rect 3467 3553 3479 3587
rect 3421 3547 3479 3553
rect 3510 3544 3516 3596
rect 3568 3584 3574 3596
rect 3789 3587 3847 3593
rect 3789 3584 3801 3587
rect 3568 3556 3801 3584
rect 3568 3544 3574 3556
rect 3789 3553 3801 3556
rect 3835 3553 3847 3587
rect 3789 3547 3847 3553
rect 4062 3544 4068 3596
rect 4120 3584 4126 3596
rect 4157 3587 4215 3593
rect 4157 3584 4169 3587
rect 4120 3556 4169 3584
rect 4120 3544 4126 3556
rect 4157 3553 4169 3556
rect 4203 3553 4215 3587
rect 5537 3587 5595 3593
rect 5537 3584 5549 3587
rect 4157 3547 4215 3553
rect 4632 3556 5549 3584
rect 1486 3516 1492 3528
rect 1447 3488 1492 3516
rect 1486 3476 1492 3488
rect 1544 3476 1550 3528
rect 1578 3476 1584 3528
rect 1636 3516 1642 3528
rect 2225 3519 2283 3525
rect 1636 3488 1681 3516
rect 1636 3476 1642 3488
rect 2225 3485 2237 3519
rect 2271 3516 2283 3519
rect 2314 3516 2320 3528
rect 2271 3488 2320 3516
rect 2271 3485 2283 3488
rect 2225 3479 2283 3485
rect 2314 3476 2320 3488
rect 2372 3476 2378 3528
rect 3326 3516 3332 3528
rect 3287 3488 3332 3516
rect 3326 3476 3332 3488
rect 3384 3476 3390 3528
rect 4338 3516 4344 3528
rect 4299 3488 4344 3516
rect 4338 3476 4344 3488
rect 4396 3476 4402 3528
rect 4430 3476 4436 3528
rect 4488 3516 4494 3528
rect 4632 3525 4660 3556
rect 5537 3553 5549 3556
rect 5583 3584 5595 3587
rect 6365 3587 6423 3593
rect 5583 3556 5948 3584
rect 5583 3553 5595 3556
rect 5537 3547 5595 3553
rect 4617 3519 4675 3525
rect 4488 3488 4533 3516
rect 4488 3476 4494 3488
rect 4617 3485 4629 3519
rect 4663 3485 4675 3519
rect 4617 3479 4675 3485
rect 4706 3476 4712 3528
rect 4764 3516 4770 3528
rect 5169 3519 5227 3525
rect 4764 3488 4809 3516
rect 4764 3476 4770 3488
rect 5169 3485 5181 3519
rect 5215 3485 5227 3519
rect 5350 3516 5356 3528
rect 5311 3488 5356 3516
rect 5169 3479 5227 3485
rect 2682 3408 2688 3460
rect 2740 3448 2746 3460
rect 4985 3451 5043 3457
rect 4985 3448 4997 3451
rect 2740 3420 4997 3448
rect 2740 3408 2746 3420
rect 4985 3417 4997 3420
rect 5031 3417 5043 3451
rect 5184 3448 5212 3479
rect 5350 3476 5356 3488
rect 5408 3476 5414 3528
rect 5718 3516 5724 3528
rect 5679 3488 5724 3516
rect 5718 3476 5724 3488
rect 5776 3476 5782 3528
rect 5920 3525 5948 3556
rect 6365 3553 6377 3587
rect 6411 3584 6423 3587
rect 6454 3584 6460 3596
rect 6411 3556 6460 3584
rect 6411 3553 6423 3556
rect 6365 3547 6423 3553
rect 6454 3544 6460 3556
rect 6512 3584 6518 3596
rect 6822 3584 6828 3596
rect 6512 3556 6828 3584
rect 6512 3544 6518 3556
rect 6822 3544 6828 3556
rect 6880 3544 6886 3596
rect 8478 3544 8484 3596
rect 8536 3584 8542 3596
rect 8757 3587 8815 3593
rect 8757 3584 8769 3587
rect 8536 3556 8769 3584
rect 8536 3544 8542 3556
rect 8757 3553 8769 3556
rect 8803 3584 8815 3587
rect 8846 3584 8852 3596
rect 8803 3556 8852 3584
rect 8803 3553 8815 3556
rect 8757 3547 8815 3553
rect 8846 3544 8852 3556
rect 8904 3544 8910 3596
rect 9048 3525 9076 3692
rect 9582 3680 9588 3692
rect 9640 3680 9646 3732
rect 9674 3680 9680 3732
rect 9732 3720 9738 3732
rect 9769 3723 9827 3729
rect 9769 3720 9781 3723
rect 9732 3692 9781 3720
rect 9732 3680 9738 3692
rect 9769 3689 9781 3692
rect 9815 3689 9827 3723
rect 9769 3683 9827 3689
rect 10778 3680 10784 3732
rect 10836 3720 10842 3732
rect 11793 3723 11851 3729
rect 11793 3720 11805 3723
rect 10836 3692 11805 3720
rect 10836 3680 10842 3692
rect 11793 3689 11805 3692
rect 11839 3689 11851 3723
rect 11793 3683 11851 3689
rect 9122 3544 9128 3596
rect 9180 3584 9186 3596
rect 10045 3587 10103 3593
rect 10045 3584 10057 3587
rect 9180 3556 10057 3584
rect 9180 3544 9186 3556
rect 10045 3553 10057 3556
rect 10091 3553 10103 3587
rect 10318 3584 10324 3596
rect 10279 3556 10324 3584
rect 10045 3547 10103 3553
rect 10318 3544 10324 3556
rect 10376 3544 10382 3596
rect 11974 3544 11980 3596
rect 12032 3584 12038 3596
rect 12897 3587 12955 3593
rect 12897 3584 12909 3587
rect 12032 3556 12909 3584
rect 12032 3544 12038 3556
rect 5905 3519 5963 3525
rect 5905 3485 5917 3519
rect 5951 3485 5963 3519
rect 5905 3479 5963 3485
rect 9033 3519 9091 3525
rect 9033 3485 9045 3519
rect 9079 3485 9091 3519
rect 9214 3516 9220 3528
rect 9175 3488 9220 3516
rect 9033 3479 9091 3485
rect 5442 3448 5448 3460
rect 5184 3420 5448 3448
rect 4985 3411 5043 3417
rect 5442 3408 5448 3420
rect 5500 3408 5506 3460
rect 8050 3420 8156 3448
rect 1854 3340 1860 3392
rect 1912 3380 1918 3392
rect 2041 3383 2099 3389
rect 2041 3380 2053 3383
rect 1912 3352 2053 3380
rect 1912 3340 1918 3352
rect 2041 3349 2053 3352
rect 2087 3349 2099 3383
rect 2041 3343 2099 3349
rect 3234 3340 3240 3392
rect 3292 3380 3298 3392
rect 4801 3383 4859 3389
rect 4801 3380 4813 3383
rect 3292 3352 4813 3380
rect 3292 3340 3298 3352
rect 4801 3349 4813 3352
rect 4847 3349 4859 3383
rect 4801 3343 4859 3349
rect 6914 3340 6920 3392
rect 6972 3380 6978 3392
rect 7009 3383 7067 3389
rect 7009 3380 7021 3383
rect 6972 3352 7021 3380
rect 6972 3340 6978 3352
rect 7009 3349 7021 3352
rect 7055 3349 7067 3383
rect 8128 3380 8156 3420
rect 8202 3408 8208 3460
rect 8260 3448 8266 3460
rect 8481 3451 8539 3457
rect 8481 3448 8493 3451
rect 8260 3420 8493 3448
rect 8260 3408 8266 3420
rect 8481 3417 8493 3420
rect 8527 3417 8539 3451
rect 9048 3448 9076 3479
rect 9214 3476 9220 3488
rect 9272 3516 9278 3528
rect 9490 3516 9496 3528
rect 9272 3488 9496 3516
rect 9272 3476 9278 3488
rect 9490 3476 9496 3488
rect 9548 3476 9554 3528
rect 12066 3516 12072 3528
rect 12027 3488 12072 3516
rect 12066 3476 12072 3488
rect 12124 3476 12130 3528
rect 12268 3525 12296 3556
rect 12897 3553 12909 3556
rect 12943 3584 12955 3587
rect 13081 3587 13139 3593
rect 13081 3584 13093 3587
rect 12943 3556 13093 3584
rect 12943 3553 12955 3556
rect 12897 3547 12955 3553
rect 13081 3553 13093 3556
rect 13127 3553 13139 3587
rect 13081 3547 13139 3553
rect 12253 3519 12311 3525
rect 12253 3485 12265 3519
rect 12299 3516 12311 3519
rect 12437 3519 12495 3525
rect 12437 3516 12449 3519
rect 12299 3488 12449 3516
rect 12299 3485 12311 3488
rect 12253 3479 12311 3485
rect 12437 3485 12449 3488
rect 12483 3485 12495 3519
rect 12437 3479 12495 3485
rect 12621 3519 12679 3525
rect 12621 3485 12633 3519
rect 12667 3485 12679 3519
rect 12621 3479 12679 3485
rect 9858 3448 9864 3460
rect 9048 3420 9864 3448
rect 8481 3411 8539 3417
rect 9858 3408 9864 3420
rect 9916 3408 9922 3460
rect 9953 3451 10011 3457
rect 9953 3417 9965 3451
rect 9999 3448 10011 3451
rect 10594 3448 10600 3460
rect 9999 3420 10600 3448
rect 9999 3417 10011 3420
rect 9953 3411 10011 3417
rect 10594 3408 10600 3420
rect 10652 3408 10658 3460
rect 11698 3448 11704 3460
rect 11546 3420 11704 3448
rect 11698 3408 11704 3420
rect 11756 3408 11762 3460
rect 11882 3408 11888 3460
rect 11940 3448 11946 3460
rect 11977 3451 12035 3457
rect 11977 3448 11989 3451
rect 11940 3420 11989 3448
rect 11940 3408 11946 3420
rect 11977 3417 11989 3420
rect 12023 3417 12035 3451
rect 12084 3448 12112 3476
rect 12636 3448 12664 3479
rect 12802 3448 12808 3460
rect 12084 3420 12664 3448
rect 12763 3420 12808 3448
rect 11977 3411 12035 3417
rect 12802 3408 12808 3420
rect 12860 3408 12866 3460
rect 9033 3383 9091 3389
rect 9033 3380 9045 3383
rect 8128 3352 9045 3380
rect 7009 3343 7067 3349
rect 9033 3349 9045 3352
rect 9079 3349 9091 3383
rect 9033 3343 9091 3349
rect 9582 3340 9588 3392
rect 9640 3380 9646 3392
rect 9769 3383 9827 3389
rect 9769 3380 9781 3383
rect 9640 3352 9781 3380
rect 9640 3340 9646 3352
rect 9769 3349 9781 3352
rect 9815 3349 9827 3383
rect 9769 3343 9827 3349
rect 1104 3290 13892 3312
rect 1104 3238 8214 3290
rect 8266 3238 8278 3290
rect 8330 3238 8342 3290
rect 8394 3238 8406 3290
rect 8458 3238 8470 3290
rect 8522 3238 13892 3290
rect 1104 3216 13892 3238
rect 1486 3136 1492 3188
rect 1544 3176 1550 3188
rect 1581 3179 1639 3185
rect 1581 3176 1593 3179
rect 1544 3148 1593 3176
rect 1544 3136 1550 3148
rect 1581 3145 1593 3148
rect 1627 3145 1639 3179
rect 2314 3176 2320 3188
rect 2275 3148 2320 3176
rect 1581 3139 1639 3145
rect 2314 3136 2320 3148
rect 2372 3136 2378 3188
rect 4706 3176 4712 3188
rect 3528 3148 4712 3176
rect 2777 3111 2835 3117
rect 2777 3108 2789 3111
rect 1780 3080 2789 3108
rect 1780 3049 1808 3080
rect 2516 3049 2544 3080
rect 2777 3077 2789 3080
rect 2823 3077 2835 3111
rect 3326 3108 3332 3120
rect 3287 3080 3332 3108
rect 2777 3071 2835 3077
rect 3326 3068 3332 3080
rect 3384 3068 3390 3120
rect 1765 3043 1823 3049
rect 1765 3009 1777 3043
rect 1811 3009 1823 3043
rect 1765 3003 1823 3009
rect 1857 3043 1915 3049
rect 1857 3009 1869 3043
rect 1903 3040 1915 3043
rect 2501 3043 2559 3049
rect 1903 3012 2268 3040
rect 1903 3009 1915 3012
rect 1857 3003 1915 3009
rect 1486 2932 1492 2984
rect 1544 2972 1550 2984
rect 1872 2972 1900 3003
rect 2130 2972 2136 2984
rect 1544 2944 1900 2972
rect 2091 2944 2136 2972
rect 1544 2932 1550 2944
rect 2130 2932 2136 2944
rect 2188 2932 2194 2984
rect 2240 2972 2268 3012
rect 2501 3009 2513 3043
rect 2547 3009 2559 3043
rect 2866 3040 2872 3052
rect 2827 3012 2872 3040
rect 2501 3003 2559 3009
rect 2866 3000 2872 3012
rect 2924 3000 2930 3052
rect 3145 3043 3203 3049
rect 3145 3009 3157 3043
rect 3191 3040 3203 3043
rect 3234 3040 3240 3052
rect 3191 3012 3240 3040
rect 3191 3009 3203 3012
rect 3145 3003 3203 3009
rect 3234 3000 3240 3012
rect 3292 3000 3298 3052
rect 3528 3049 3556 3148
rect 4706 3136 4712 3148
rect 4764 3176 4770 3188
rect 5169 3179 5227 3185
rect 5169 3176 5181 3179
rect 4764 3148 5181 3176
rect 4764 3136 4770 3148
rect 5169 3145 5181 3148
rect 5215 3145 5227 3179
rect 5169 3139 5227 3145
rect 5442 3136 5448 3188
rect 5500 3176 5506 3188
rect 6914 3176 6920 3188
rect 5500 3148 6920 3176
rect 5500 3136 5506 3148
rect 5736 3117 5764 3148
rect 6914 3136 6920 3148
rect 6972 3136 6978 3188
rect 7469 3179 7527 3185
rect 7469 3145 7481 3179
rect 7515 3176 7527 3179
rect 8110 3176 8116 3188
rect 7515 3148 8116 3176
rect 7515 3145 7527 3148
rect 7469 3139 7527 3145
rect 8110 3136 8116 3148
rect 8168 3136 8174 3188
rect 10594 3136 10600 3188
rect 10652 3176 10658 3188
rect 10781 3179 10839 3185
rect 10781 3176 10793 3179
rect 10652 3148 10793 3176
rect 10652 3136 10658 3148
rect 10781 3145 10793 3148
rect 10827 3176 10839 3179
rect 11054 3176 11060 3188
rect 10827 3148 11060 3176
rect 10827 3145 10839 3148
rect 10781 3139 10839 3145
rect 11054 3136 11060 3148
rect 11112 3136 11118 3188
rect 11330 3176 11336 3188
rect 11243 3148 11336 3176
rect 11330 3136 11336 3148
rect 11388 3176 11394 3188
rect 11974 3176 11980 3188
rect 11388 3148 11980 3176
rect 11388 3136 11394 3148
rect 3697 3111 3755 3117
rect 3697 3077 3709 3111
rect 3743 3108 3755 3111
rect 5721 3111 5779 3117
rect 3743 3080 4476 3108
rect 3743 3077 3755 3080
rect 3697 3071 3755 3077
rect 4448 3052 4476 3080
rect 5721 3077 5733 3111
rect 5767 3077 5779 3111
rect 5721 3071 5779 3077
rect 5905 3111 5963 3117
rect 5905 3077 5917 3111
rect 5951 3108 5963 3111
rect 8021 3111 8079 3117
rect 8021 3108 8033 3111
rect 5951 3080 6316 3108
rect 5951 3077 5963 3080
rect 5905 3071 5963 3077
rect 3513 3043 3571 3049
rect 3513 3009 3525 3043
rect 3559 3009 3571 3043
rect 3513 3003 3571 3009
rect 3789 3043 3847 3049
rect 3789 3009 3801 3043
rect 3835 3040 3847 3043
rect 3835 3012 4384 3040
rect 3835 3009 3847 3012
rect 3789 3003 3847 3009
rect 4356 2984 4384 3012
rect 4430 3000 4436 3052
rect 4488 3040 4494 3052
rect 4706 3040 4712 3052
rect 4488 3012 4712 3040
rect 4488 3000 4494 3012
rect 4706 3000 4712 3012
rect 4764 3000 4770 3052
rect 5350 3040 5356 3052
rect 5311 3012 5356 3040
rect 5350 3000 5356 3012
rect 5408 3000 5414 3052
rect 5442 3000 5448 3052
rect 5500 3040 5506 3052
rect 5537 3043 5595 3049
rect 5537 3040 5549 3043
rect 5500 3012 5549 3040
rect 5500 3000 5506 3012
rect 5537 3009 5549 3012
rect 5583 3040 5595 3043
rect 5583 3012 5948 3040
rect 5583 3009 5595 3012
rect 5537 3003 5595 3009
rect 2682 2972 2688 2984
rect 2240 2944 2688 2972
rect 2682 2932 2688 2944
rect 2740 2932 2746 2984
rect 3881 2975 3939 2981
rect 3881 2941 3893 2975
rect 3927 2941 3939 2975
rect 3881 2935 3939 2941
rect 2041 2907 2099 2913
rect 2041 2873 2053 2907
rect 2087 2904 2099 2907
rect 2314 2904 2320 2916
rect 2087 2876 2320 2904
rect 2087 2873 2099 2876
rect 2041 2867 2099 2873
rect 2314 2864 2320 2876
rect 2372 2904 2378 2916
rect 3896 2904 3924 2935
rect 4338 2932 4344 2984
rect 4396 2972 4402 2984
rect 4614 2972 4620 2984
rect 4396 2944 4620 2972
rect 4396 2932 4402 2944
rect 4614 2932 4620 2944
rect 4672 2932 4678 2984
rect 2372 2876 3924 2904
rect 5920 2904 5948 3012
rect 6288 2984 6316 3080
rect 7024 3080 8033 3108
rect 6546 3040 6552 3052
rect 6507 3012 6552 3040
rect 6546 3000 6552 3012
rect 6604 3000 6610 3052
rect 7024 3049 7052 3080
rect 8021 3077 8033 3080
rect 8067 3077 8079 3111
rect 8570 3108 8576 3120
rect 8021 3071 8079 3077
rect 8312 3080 8576 3108
rect 7009 3043 7067 3049
rect 7009 3009 7021 3043
rect 7055 3009 7067 3043
rect 7009 3003 7067 3009
rect 7098 3000 7104 3052
rect 7156 3040 7162 3052
rect 8312 3049 8340 3080
rect 8570 3068 8576 3080
rect 8628 3068 8634 3120
rect 9858 3108 9864 3120
rect 9798 3080 9864 3108
rect 9858 3068 9864 3080
rect 9916 3068 9922 3120
rect 11532 3049 11560 3148
rect 11974 3136 11980 3148
rect 12032 3136 12038 3188
rect 12066 3108 12072 3120
rect 11808 3080 12072 3108
rect 11808 3049 11836 3080
rect 12066 3068 12072 3080
rect 12124 3068 12130 3120
rect 7193 3043 7251 3049
rect 7193 3040 7205 3043
rect 7156 3012 7205 3040
rect 7156 3000 7162 3012
rect 7193 3009 7205 3012
rect 7239 3009 7251 3043
rect 7653 3043 7711 3049
rect 7653 3040 7665 3043
rect 7193 3003 7251 3009
rect 7300 3012 7665 3040
rect 6270 2932 6276 2984
rect 6328 2972 6334 2984
rect 6365 2975 6423 2981
rect 6365 2972 6377 2975
rect 6328 2944 6377 2972
rect 6328 2932 6334 2944
rect 6365 2941 6377 2944
rect 6411 2941 6423 2975
rect 6914 2972 6920 2984
rect 6875 2944 6920 2972
rect 6365 2935 6423 2941
rect 6914 2932 6920 2944
rect 6972 2932 6978 2984
rect 6546 2904 6552 2916
rect 5920 2876 6552 2904
rect 2372 2864 2378 2876
rect 5920 2845 5948 2876
rect 6546 2864 6552 2876
rect 6604 2864 6610 2916
rect 6825 2907 6883 2913
rect 6825 2873 6837 2907
rect 6871 2904 6883 2907
rect 7300 2904 7328 3012
rect 7653 3009 7665 3012
rect 7699 3009 7711 3043
rect 7653 3003 7711 3009
rect 7837 3043 7895 3049
rect 7837 3009 7849 3043
rect 7883 3009 7895 3043
rect 7837 3003 7895 3009
rect 8297 3043 8355 3049
rect 8297 3009 8309 3043
rect 8343 3009 8355 3043
rect 8297 3003 8355 3009
rect 10689 3043 10747 3049
rect 10689 3009 10701 3043
rect 10735 3009 10747 3043
rect 10689 3003 10747 3009
rect 11517 3043 11575 3049
rect 11517 3009 11529 3043
rect 11563 3009 11575 3043
rect 11517 3003 11575 3009
rect 11793 3043 11851 3049
rect 11793 3009 11805 3043
rect 11839 3009 11851 3043
rect 11793 3003 11851 3009
rect 12897 3043 12955 3049
rect 12897 3009 12909 3043
rect 12943 3009 12955 3043
rect 12897 3003 12955 3009
rect 13081 3043 13139 3049
rect 13081 3009 13093 3043
rect 13127 3040 13139 3043
rect 13170 3040 13176 3052
rect 13127 3012 13176 3040
rect 13127 3009 13139 3012
rect 13081 3003 13139 3009
rect 7561 2975 7619 2981
rect 7561 2941 7573 2975
rect 7607 2941 7619 2975
rect 7852 2972 7880 3003
rect 8573 2975 8631 2981
rect 7852 2944 7972 2972
rect 7561 2935 7619 2941
rect 6871 2876 7328 2904
rect 7576 2904 7604 2935
rect 7834 2904 7840 2916
rect 7576 2876 7840 2904
rect 6871 2873 6883 2876
rect 6825 2867 6883 2873
rect 7834 2864 7840 2876
rect 7892 2864 7898 2916
rect 5905 2839 5963 2845
rect 5905 2805 5917 2839
rect 5951 2805 5963 2839
rect 5905 2799 5963 2805
rect 6089 2839 6147 2845
rect 6089 2805 6101 2839
rect 6135 2836 6147 2839
rect 6178 2836 6184 2848
rect 6135 2808 6184 2836
rect 6135 2805 6147 2808
rect 6089 2799 6147 2805
rect 6178 2796 6184 2808
rect 6236 2836 6242 2848
rect 7944 2836 7972 2944
rect 8573 2941 8585 2975
rect 8619 2972 8631 2975
rect 8938 2972 8944 2984
rect 8619 2944 8944 2972
rect 8619 2941 8631 2944
rect 8573 2935 8631 2941
rect 8938 2932 8944 2944
rect 8996 2932 9002 2984
rect 9766 2932 9772 2984
rect 9824 2972 9830 2984
rect 10042 2972 10048 2984
rect 9824 2944 10048 2972
rect 9824 2932 9830 2944
rect 10042 2932 10048 2944
rect 10100 2972 10106 2984
rect 10704 2972 10732 3003
rect 10100 2944 10732 2972
rect 10965 2975 11023 2981
rect 10100 2932 10106 2944
rect 10965 2941 10977 2975
rect 11011 2972 11023 2975
rect 12069 2975 12127 2981
rect 12069 2972 12081 2975
rect 11011 2944 12081 2972
rect 11011 2941 11023 2944
rect 10965 2935 11023 2941
rect 12069 2941 12081 2944
rect 12115 2941 12127 2975
rect 12912 2972 12940 3003
rect 13170 3000 13176 3012
rect 13228 3000 13234 3052
rect 13262 2972 13268 2984
rect 12912 2944 13268 2972
rect 12069 2935 12127 2941
rect 10980 2904 11008 2935
rect 13262 2932 13268 2944
rect 13320 2932 13326 2984
rect 9600 2876 11008 2904
rect 11793 2907 11851 2913
rect 6236 2808 7972 2836
rect 6236 2796 6242 2808
rect 8018 2796 8024 2848
rect 8076 2836 8082 2848
rect 9600 2836 9628 2876
rect 11793 2873 11805 2907
rect 11839 2904 11851 2907
rect 12618 2904 12624 2916
rect 11839 2876 12624 2904
rect 11839 2873 11851 2876
rect 11793 2867 11851 2873
rect 12618 2864 12624 2876
rect 12676 2864 12682 2916
rect 8076 2808 9628 2836
rect 10321 2839 10379 2845
rect 8076 2796 8082 2808
rect 10321 2805 10333 2839
rect 10367 2836 10379 2839
rect 10594 2836 10600 2848
rect 10367 2808 10600 2836
rect 10367 2805 10379 2808
rect 10321 2799 10379 2805
rect 10594 2796 10600 2808
rect 10652 2796 10658 2848
rect 1104 2746 13892 2768
rect 1104 2694 4214 2746
rect 4266 2694 4278 2746
rect 4330 2694 4342 2746
rect 4394 2694 4406 2746
rect 4458 2694 4470 2746
rect 4522 2694 12214 2746
rect 12266 2694 12278 2746
rect 12330 2694 12342 2746
rect 12394 2694 12406 2746
rect 12458 2694 12470 2746
rect 12522 2694 13892 2746
rect 1104 2672 13892 2694
rect 2685 2635 2743 2641
rect 2685 2601 2697 2635
rect 2731 2632 2743 2635
rect 2866 2632 2872 2644
rect 2731 2604 2872 2632
rect 2731 2601 2743 2604
rect 2685 2595 2743 2601
rect 2866 2592 2872 2604
rect 2924 2592 2930 2644
rect 4157 2635 4215 2641
rect 4157 2601 4169 2635
rect 4203 2632 4215 2635
rect 4706 2632 4712 2644
rect 4203 2604 4712 2632
rect 4203 2601 4215 2604
rect 4157 2595 4215 2601
rect 4706 2592 4712 2604
rect 4764 2592 4770 2644
rect 8938 2632 8944 2644
rect 8899 2604 8944 2632
rect 8938 2592 8944 2604
rect 8996 2592 9002 2644
rect 11054 2592 11060 2644
rect 11112 2632 11118 2644
rect 12069 2635 12127 2641
rect 12069 2632 12081 2635
rect 11112 2604 12081 2632
rect 11112 2592 11118 2604
rect 12069 2601 12081 2604
rect 12115 2601 12127 2635
rect 12069 2595 12127 2601
rect 3418 2564 3424 2576
rect 1688 2536 3424 2564
rect 1688 2496 1716 2536
rect 3418 2524 3424 2536
rect 3476 2524 3482 2576
rect 3786 2524 3792 2576
rect 3844 2564 3850 2576
rect 9858 2564 9864 2576
rect 3844 2536 5672 2564
rect 9819 2536 9864 2564
rect 3844 2524 3850 2536
rect 1596 2468 1716 2496
rect 1596 2437 1624 2468
rect 1762 2456 1768 2508
rect 1820 2496 1826 2508
rect 1949 2499 2007 2505
rect 1949 2496 1961 2499
rect 1820 2468 1961 2496
rect 1820 2456 1826 2468
rect 1949 2465 1961 2468
rect 1995 2465 2007 2499
rect 1949 2459 2007 2465
rect 3513 2499 3571 2505
rect 3513 2465 3525 2499
rect 3559 2496 3571 2499
rect 3602 2496 3608 2508
rect 3559 2468 3608 2496
rect 3559 2465 3571 2468
rect 3513 2459 3571 2465
rect 3602 2456 3608 2468
rect 3660 2456 3666 2508
rect 4525 2499 4583 2505
rect 3896 2468 4108 2496
rect 1581 2431 1639 2437
rect 1581 2397 1593 2431
rect 1627 2397 1639 2431
rect 1581 2391 1639 2397
rect 1670 2388 1676 2440
rect 1728 2428 1734 2440
rect 2130 2428 2136 2440
rect 1728 2400 1773 2428
rect 2091 2400 2136 2428
rect 1728 2388 1734 2400
rect 2130 2388 2136 2400
rect 2188 2388 2194 2440
rect 2314 2428 2320 2440
rect 2275 2400 2320 2428
rect 2314 2388 2320 2400
rect 2372 2388 2378 2440
rect 2593 2431 2651 2437
rect 2593 2397 2605 2431
rect 2639 2397 2651 2431
rect 2593 2391 2651 2397
rect 2777 2431 2835 2437
rect 2777 2397 2789 2431
rect 2823 2428 2835 2431
rect 2866 2428 2872 2440
rect 2823 2400 2872 2428
rect 2823 2397 2835 2400
rect 2777 2391 2835 2397
rect 1854 2360 1860 2372
rect 1815 2332 1860 2360
rect 1854 2320 1860 2332
rect 1912 2320 1918 2372
rect 2608 2360 2636 2391
rect 2866 2388 2872 2400
rect 2924 2428 2930 2440
rect 3896 2437 3924 2468
rect 3329 2431 3387 2437
rect 3329 2428 3341 2431
rect 2924 2400 3341 2428
rect 2924 2388 2930 2400
rect 3329 2397 3341 2400
rect 3375 2397 3387 2431
rect 3329 2391 3387 2397
rect 3881 2431 3939 2437
rect 3881 2397 3893 2431
rect 3927 2397 3939 2431
rect 3881 2391 3939 2397
rect 3973 2431 4031 2437
rect 3973 2397 3985 2431
rect 4019 2397 4031 2431
rect 3973 2391 4031 2397
rect 3344 2360 3372 2391
rect 3694 2360 3700 2372
rect 2608 2332 3280 2360
rect 3344 2332 3700 2360
rect 2869 2295 2927 2301
rect 2869 2261 2881 2295
rect 2915 2292 2927 2295
rect 3142 2292 3148 2304
rect 2915 2264 3148 2292
rect 2915 2261 2927 2264
rect 2869 2255 2927 2261
rect 3142 2252 3148 2264
rect 3200 2252 3206 2304
rect 3252 2301 3280 2332
rect 3694 2320 3700 2332
rect 3752 2360 3758 2372
rect 3988 2360 4016 2391
rect 3752 2332 4016 2360
rect 3752 2320 3758 2332
rect 3237 2295 3295 2301
rect 3237 2261 3249 2295
rect 3283 2292 3295 2295
rect 3326 2292 3332 2304
rect 3283 2264 3332 2292
rect 3283 2261 3295 2264
rect 3237 2255 3295 2261
rect 3326 2252 3332 2264
rect 3384 2292 3390 2304
rect 4080 2292 4108 2468
rect 4525 2465 4537 2499
rect 4571 2496 4583 2499
rect 4614 2496 4620 2508
rect 4571 2468 4620 2496
rect 4571 2465 4583 2468
rect 4525 2459 4583 2465
rect 4614 2456 4620 2468
rect 4672 2456 4678 2508
rect 5644 2505 5672 2536
rect 9858 2524 9864 2536
rect 9916 2524 9922 2576
rect 5629 2499 5687 2505
rect 5629 2465 5641 2499
rect 5675 2496 5687 2499
rect 8570 2496 8576 2508
rect 5675 2468 8576 2496
rect 5675 2465 5687 2468
rect 5629 2459 5687 2465
rect 8570 2456 8576 2468
rect 8628 2456 8634 2508
rect 9582 2496 9588 2508
rect 9232 2468 9588 2496
rect 5356 2440 5408 2446
rect 5442 2388 5448 2440
rect 5500 2428 5506 2440
rect 7558 2428 7564 2440
rect 5500 2400 5545 2428
rect 7519 2400 7564 2428
rect 5500 2388 5506 2400
rect 7558 2388 7564 2400
rect 7616 2388 7622 2440
rect 7745 2431 7803 2437
rect 7745 2397 7757 2431
rect 7791 2397 7803 2431
rect 7745 2391 7803 2397
rect 5356 2382 5408 2388
rect 5902 2360 5908 2372
rect 5863 2332 5908 2360
rect 5902 2320 5908 2332
rect 5960 2320 5966 2372
rect 6362 2320 6368 2372
rect 6420 2320 6426 2372
rect 7190 2320 7196 2372
rect 7248 2360 7254 2372
rect 7760 2360 7788 2391
rect 7834 2388 7840 2440
rect 7892 2428 7898 2440
rect 8113 2431 8171 2437
rect 8113 2428 8125 2431
rect 7892 2400 8125 2428
rect 7892 2388 7898 2400
rect 8113 2397 8125 2400
rect 8159 2428 8171 2431
rect 9232 2428 9260 2468
rect 9582 2456 9588 2468
rect 9640 2496 9646 2508
rect 12253 2499 12311 2505
rect 12253 2496 12265 2499
rect 9640 2468 12265 2496
rect 9640 2456 9646 2468
rect 12253 2465 12265 2468
rect 12299 2465 12311 2499
rect 12253 2459 12311 2465
rect 13176 2440 13228 2446
rect 8159 2400 9260 2428
rect 9309 2431 9367 2437
rect 8159 2397 8171 2400
rect 8113 2391 8171 2397
rect 9309 2397 9321 2431
rect 9355 2428 9367 2431
rect 9766 2428 9772 2440
rect 9355 2400 9772 2428
rect 9355 2397 9367 2400
rect 9309 2391 9367 2397
rect 9766 2388 9772 2400
rect 9824 2388 9830 2440
rect 9950 2428 9956 2440
rect 9911 2400 9956 2428
rect 9950 2388 9956 2400
rect 10008 2388 10014 2440
rect 10045 2431 10103 2437
rect 10045 2397 10057 2431
rect 10091 2397 10103 2431
rect 10045 2391 10103 2397
rect 10321 2431 10379 2437
rect 10321 2397 10333 2431
rect 10367 2397 10379 2431
rect 10321 2391 10379 2397
rect 7248 2332 7788 2360
rect 7248 2320 7254 2332
rect 9122 2320 9128 2372
rect 9180 2360 9186 2372
rect 9401 2363 9459 2369
rect 9401 2360 9413 2363
rect 9180 2332 9413 2360
rect 9180 2320 9186 2332
rect 9401 2329 9413 2332
rect 9447 2360 9459 2363
rect 9674 2360 9680 2372
rect 9447 2332 9680 2360
rect 9447 2329 9459 2332
rect 9401 2323 9459 2329
rect 9674 2320 9680 2332
rect 9732 2320 9738 2372
rect 10060 2360 10088 2391
rect 9968 2332 10088 2360
rect 5626 2292 5632 2304
rect 3384 2264 5632 2292
rect 3384 2252 3390 2264
rect 5626 2252 5632 2264
rect 5684 2292 5690 2304
rect 6270 2292 6276 2304
rect 5684 2264 6276 2292
rect 5684 2252 5690 2264
rect 6270 2252 6276 2264
rect 6328 2292 6334 2304
rect 7282 2292 7288 2304
rect 6328 2264 7288 2292
rect 6328 2252 6334 2264
rect 7282 2252 7288 2264
rect 7340 2292 7346 2304
rect 7377 2295 7435 2301
rect 7377 2292 7389 2295
rect 7340 2264 7389 2292
rect 7340 2252 7346 2264
rect 7377 2261 7389 2264
rect 7423 2261 7435 2295
rect 7377 2255 7435 2261
rect 8021 2295 8079 2301
rect 8021 2261 8033 2295
rect 8067 2292 8079 2295
rect 8110 2292 8116 2304
rect 8067 2264 8116 2292
rect 8067 2261 8079 2264
rect 8021 2255 8079 2261
rect 8110 2252 8116 2264
rect 8168 2252 8174 2304
rect 8297 2295 8355 2301
rect 8297 2261 8309 2295
rect 8343 2292 8355 2295
rect 8662 2292 8668 2304
rect 8343 2264 8668 2292
rect 8343 2261 8355 2264
rect 8297 2255 8355 2261
rect 8662 2252 8668 2264
rect 8720 2292 8726 2304
rect 9490 2292 9496 2304
rect 8720 2264 9496 2292
rect 8720 2252 8726 2264
rect 9490 2252 9496 2264
rect 9548 2292 9554 2304
rect 9968 2292 9996 2332
rect 9548 2264 9996 2292
rect 10336 2292 10364 2391
rect 13262 2388 13268 2440
rect 13320 2428 13326 2440
rect 13320 2400 13365 2428
rect 13320 2388 13326 2400
rect 13176 2382 13228 2388
rect 10594 2360 10600 2372
rect 10555 2332 10600 2360
rect 10594 2320 10600 2332
rect 10652 2320 10658 2372
rect 11882 2360 11888 2372
rect 11822 2332 11888 2360
rect 11882 2320 11888 2332
rect 11940 2320 11946 2372
rect 11514 2292 11520 2304
rect 10336 2264 11520 2292
rect 9548 2252 9554 2264
rect 11514 2252 11520 2264
rect 11572 2252 11578 2304
rect 1104 2202 13892 2224
rect 1104 2150 8214 2202
rect 8266 2150 8278 2202
rect 8330 2150 8342 2202
rect 8394 2150 8406 2202
rect 8458 2150 8470 2202
rect 8522 2150 13892 2202
rect 1104 2128 13892 2150
rect 1578 2088 1584 2100
rect 1539 2060 1584 2088
rect 1578 2048 1584 2060
rect 1636 2048 1642 2100
rect 1765 2091 1823 2097
rect 1765 2057 1777 2091
rect 1811 2088 1823 2091
rect 2866 2088 2872 2100
rect 1811 2060 2872 2088
rect 1811 2057 1823 2060
rect 1765 2051 1823 2057
rect 2866 2048 2872 2060
rect 2924 2048 2930 2100
rect 3418 2048 3424 2100
rect 3476 2088 3482 2100
rect 3605 2091 3663 2097
rect 3605 2088 3617 2091
rect 3476 2060 3617 2088
rect 3476 2048 3482 2060
rect 3605 2057 3617 2060
rect 3651 2057 3663 2091
rect 3605 2051 3663 2057
rect 5350 2048 5356 2100
rect 5408 2088 5414 2100
rect 5537 2091 5595 2097
rect 5537 2088 5549 2091
rect 5408 2060 5549 2088
rect 5408 2048 5414 2060
rect 5537 2057 5549 2060
rect 5583 2057 5595 2091
rect 5537 2051 5595 2057
rect 6089 2091 6147 2097
rect 6089 2057 6101 2091
rect 6135 2088 6147 2091
rect 6362 2088 6368 2100
rect 6135 2060 6368 2088
rect 6135 2057 6147 2060
rect 6089 2051 6147 2057
rect 6362 2048 6368 2060
rect 6420 2048 6426 2100
rect 6454 2048 6460 2100
rect 6512 2088 6518 2100
rect 8662 2088 8668 2100
rect 6512 2060 8668 2088
rect 6512 2048 6518 2060
rect 8662 2048 8668 2060
rect 8720 2048 8726 2100
rect 9674 2048 9680 2100
rect 9732 2088 9738 2100
rect 10321 2091 10379 2097
rect 10321 2088 10333 2091
rect 9732 2060 10333 2088
rect 9732 2048 9738 2060
rect 10321 2057 10333 2060
rect 10367 2057 10379 2091
rect 10321 2051 10379 2057
rect 13170 2048 13176 2100
rect 13228 2088 13234 2100
rect 13265 2091 13323 2097
rect 13265 2088 13277 2091
rect 13228 2060 13277 2088
rect 13228 2048 13234 2060
rect 13265 2057 13277 2060
rect 13311 2057 13323 2091
rect 13265 2051 13323 2057
rect 1854 1980 1860 2032
rect 1912 2020 1918 2032
rect 1912 1992 2070 2020
rect 1912 1980 1918 1992
rect 3142 1980 3148 2032
rect 3200 2020 3206 2032
rect 3237 2023 3295 2029
rect 3237 2020 3249 2023
rect 3200 1992 3249 2020
rect 3200 1980 3206 1992
rect 3237 1989 3249 1992
rect 3283 1989 3295 2023
rect 3237 1983 3295 1989
rect 4614 1980 4620 2032
rect 4672 1980 4678 2032
rect 6472 2020 6500 2048
rect 7926 2020 7932 2032
rect 5920 1992 6500 2020
rect 7774 1992 7932 2020
rect 3510 1912 3516 1964
rect 3568 1952 3574 1964
rect 3786 1952 3792 1964
rect 3568 1924 3792 1952
rect 3568 1912 3574 1924
rect 3786 1912 3792 1924
rect 3844 1912 3850 1964
rect 5920 1961 5948 1992
rect 7926 1980 7932 1992
rect 7984 1980 7990 2032
rect 8110 1980 8116 2032
rect 8168 2020 8174 2032
rect 8205 2023 8263 2029
rect 8205 2020 8217 2023
rect 8168 1992 8217 2020
rect 8168 1980 8174 1992
rect 8205 1989 8217 1992
rect 8251 1989 8263 2023
rect 10505 2023 10563 2029
rect 10505 2020 10517 2023
rect 10074 1992 10517 2020
rect 8205 1983 8263 1989
rect 10505 1989 10517 1992
rect 10551 1989 10563 2023
rect 12066 2020 12072 2032
rect 10505 1983 10563 1989
rect 10704 1992 12072 2020
rect 5905 1955 5963 1961
rect 5905 1921 5917 1955
rect 5951 1921 5963 1955
rect 5905 1915 5963 1921
rect 6089 1955 6147 1961
rect 6089 1921 6101 1955
rect 6135 1952 6147 1955
rect 6730 1952 6736 1964
rect 6135 1924 6736 1952
rect 6135 1921 6147 1924
rect 6089 1915 6147 1921
rect 6730 1912 6736 1924
rect 6788 1912 6794 1964
rect 10134 1912 10140 1964
rect 10192 1952 10198 1964
rect 10704 1961 10732 1992
rect 11164 1961 11192 1992
rect 12066 1980 12072 1992
rect 12124 1980 12130 2032
rect 12526 1980 12532 2032
rect 12584 1980 12590 2032
rect 10689 1955 10747 1961
rect 10689 1952 10701 1955
rect 10192 1924 10701 1952
rect 10192 1912 10198 1924
rect 10689 1921 10701 1924
rect 10735 1921 10747 1955
rect 10689 1915 10747 1921
rect 10781 1955 10839 1961
rect 10781 1921 10793 1955
rect 10827 1921 10839 1955
rect 10781 1915 10839 1921
rect 11149 1955 11207 1961
rect 11149 1921 11161 1955
rect 11195 1921 11207 1955
rect 11149 1915 11207 1921
rect 11241 1955 11299 1961
rect 11241 1921 11253 1955
rect 11287 1952 11299 1955
rect 11330 1952 11336 1964
rect 11287 1924 11336 1952
rect 11287 1921 11299 1924
rect 11241 1915 11299 1921
rect 4062 1884 4068 1896
rect 4023 1856 4068 1884
rect 4062 1844 4068 1856
rect 4120 1844 4126 1896
rect 8481 1887 8539 1893
rect 8481 1853 8493 1887
rect 8527 1884 8539 1887
rect 8570 1884 8576 1896
rect 8527 1856 8576 1884
rect 8527 1853 8539 1856
rect 8481 1847 8539 1853
rect 8570 1844 8576 1856
rect 8628 1844 8634 1896
rect 8849 1887 8907 1893
rect 8849 1853 8861 1887
rect 8895 1884 8907 1887
rect 8938 1884 8944 1896
rect 8895 1856 8944 1884
rect 8895 1853 8907 1856
rect 8849 1847 8907 1853
rect 8938 1844 8944 1856
rect 8996 1844 9002 1896
rect 9490 1844 9496 1896
rect 9548 1884 9554 1896
rect 10796 1884 10824 1915
rect 11256 1884 11284 1915
rect 11330 1912 11336 1924
rect 11388 1912 11394 1964
rect 11514 1884 11520 1896
rect 9548 1856 11284 1884
rect 11475 1856 11520 1884
rect 9548 1844 9554 1856
rect 11054 1816 11060 1828
rect 11015 1788 11060 1816
rect 11054 1776 11060 1788
rect 11112 1776 11118 1828
rect 6546 1708 6552 1760
rect 6604 1748 6610 1760
rect 6733 1751 6791 1757
rect 6733 1748 6745 1751
rect 6604 1720 6745 1748
rect 6604 1708 6610 1720
rect 6733 1717 6745 1720
rect 6779 1748 6791 1751
rect 7006 1748 7012 1760
rect 6779 1720 7012 1748
rect 6779 1717 6791 1720
rect 6733 1711 6791 1717
rect 7006 1708 7012 1720
rect 7064 1708 7070 1760
rect 11256 1748 11284 1856
rect 11514 1844 11520 1856
rect 11572 1844 11578 1896
rect 11793 1887 11851 1893
rect 11793 1853 11805 1887
rect 11839 1884 11851 1887
rect 13262 1884 13268 1896
rect 11839 1856 13268 1884
rect 11839 1853 11851 1856
rect 11793 1847 11851 1853
rect 13262 1844 13268 1856
rect 13320 1844 13326 1896
rect 13449 1751 13507 1757
rect 13449 1748 13461 1751
rect 11256 1720 13461 1748
rect 13449 1717 13461 1720
rect 13495 1717 13507 1751
rect 13449 1711 13507 1717
rect 1104 1658 13892 1680
rect 1104 1606 4214 1658
rect 4266 1606 4278 1658
rect 4330 1606 4342 1658
rect 4394 1606 4406 1658
rect 4458 1606 4470 1658
rect 4522 1606 12214 1658
rect 12266 1606 12278 1658
rect 12330 1606 12342 1658
rect 12394 1606 12406 1658
rect 12458 1606 12470 1658
rect 12522 1606 13892 1658
rect 1104 1584 13892 1606
rect 1670 1504 1676 1556
rect 1728 1544 1734 1556
rect 4065 1547 4123 1553
rect 4065 1544 4077 1547
rect 1728 1516 4077 1544
rect 1728 1504 1734 1516
rect 4065 1513 4077 1516
rect 4111 1544 4123 1547
rect 4430 1544 4436 1556
rect 4111 1516 4436 1544
rect 4111 1513 4123 1516
rect 4065 1507 4123 1513
rect 4430 1504 4436 1516
rect 4488 1544 4494 1556
rect 6730 1544 6736 1556
rect 4488 1516 6736 1544
rect 4488 1504 4494 1516
rect 6730 1504 6736 1516
rect 6788 1504 6794 1556
rect 8481 1547 8539 1553
rect 8481 1513 8493 1547
rect 8527 1544 8539 1547
rect 8662 1544 8668 1556
rect 8527 1516 8668 1544
rect 8527 1513 8539 1516
rect 8481 1507 8539 1513
rect 3418 1436 3424 1488
rect 3476 1476 3482 1488
rect 4246 1476 4252 1488
rect 3476 1448 4252 1476
rect 3476 1436 3482 1448
rect 4246 1436 4252 1448
rect 4304 1436 4310 1488
rect 1394 1408 1400 1420
rect 1355 1380 1400 1408
rect 1394 1368 1400 1380
rect 1452 1368 1458 1420
rect 3694 1408 3700 1420
rect 3620 1380 3700 1408
rect 3145 1343 3203 1349
rect 3145 1309 3157 1343
rect 3191 1340 3203 1343
rect 3510 1340 3516 1352
rect 3191 1312 3516 1340
rect 3191 1309 3203 1312
rect 3145 1303 3203 1309
rect 3510 1300 3516 1312
rect 3568 1300 3574 1352
rect 3620 1349 3648 1380
rect 3694 1368 3700 1380
rect 3752 1368 3758 1420
rect 4080 1380 4752 1408
rect 3605 1343 3663 1349
rect 3605 1309 3617 1343
rect 3651 1309 3663 1343
rect 3605 1303 3663 1309
rect 3878 1300 3884 1352
rect 3936 1340 3942 1352
rect 4080 1349 4108 1380
rect 4065 1343 4123 1349
rect 3936 1312 3981 1340
rect 3936 1300 3942 1312
rect 4065 1309 4077 1343
rect 4111 1309 4123 1343
rect 4246 1340 4252 1352
rect 4207 1312 4252 1340
rect 4065 1303 4123 1309
rect 3234 1272 3240 1284
rect 3195 1244 3240 1272
rect 3234 1232 3240 1244
rect 3292 1232 3298 1284
rect 3326 1232 3332 1284
rect 3384 1272 3390 1284
rect 3421 1275 3479 1281
rect 3421 1272 3433 1275
rect 3384 1244 3433 1272
rect 3384 1232 3390 1244
rect 3421 1241 3433 1244
rect 3467 1241 3479 1275
rect 3421 1235 3479 1241
rect 3694 1164 3700 1216
rect 3752 1204 3758 1216
rect 4080 1204 4108 1303
rect 4246 1300 4252 1312
rect 4304 1300 4310 1352
rect 4430 1340 4436 1352
rect 4391 1312 4436 1340
rect 4430 1300 4436 1312
rect 4488 1300 4494 1352
rect 4614 1340 4620 1352
rect 4575 1312 4620 1340
rect 4614 1300 4620 1312
rect 4672 1300 4678 1352
rect 4724 1340 4752 1380
rect 4890 1368 4896 1420
rect 4948 1408 4954 1420
rect 5261 1411 5319 1417
rect 5261 1408 5273 1411
rect 4948 1380 5273 1408
rect 4948 1368 4954 1380
rect 5261 1377 5273 1380
rect 5307 1408 5319 1411
rect 5902 1408 5908 1420
rect 5307 1380 5764 1408
rect 5863 1380 5908 1408
rect 5307 1377 5319 1380
rect 5261 1371 5319 1377
rect 5169 1343 5227 1349
rect 4724 1312 4844 1340
rect 4522 1232 4528 1284
rect 4580 1272 4586 1284
rect 4816 1272 4844 1312
rect 5169 1309 5181 1343
rect 5215 1340 5227 1343
rect 5350 1340 5356 1352
rect 5215 1312 5356 1340
rect 5215 1309 5227 1312
rect 5169 1303 5227 1309
rect 5350 1300 5356 1312
rect 5408 1300 5414 1352
rect 5537 1343 5595 1349
rect 5537 1309 5549 1343
rect 5583 1340 5595 1343
rect 5626 1340 5632 1352
rect 5583 1312 5632 1340
rect 5583 1309 5595 1312
rect 5537 1303 5595 1309
rect 5626 1300 5632 1312
rect 5684 1300 5690 1352
rect 5736 1349 5764 1380
rect 5902 1368 5908 1380
rect 5960 1368 5966 1420
rect 6104 1380 6316 1408
rect 5721 1343 5779 1349
rect 5721 1309 5733 1343
rect 5767 1309 5779 1343
rect 5721 1303 5779 1309
rect 6104 1272 6132 1380
rect 6181 1343 6239 1349
rect 6181 1309 6193 1343
rect 6227 1309 6239 1343
rect 6288 1340 6316 1380
rect 6730 1368 6736 1420
rect 6788 1408 6794 1420
rect 7282 1408 7288 1420
rect 6788 1380 7144 1408
rect 7243 1380 7288 1408
rect 6788 1368 6794 1380
rect 6549 1343 6607 1349
rect 6549 1340 6561 1343
rect 6288 1312 6561 1340
rect 6181 1303 6239 1309
rect 6549 1309 6561 1312
rect 6595 1309 6607 1343
rect 7006 1340 7012 1352
rect 6967 1312 7012 1340
rect 6549 1303 6607 1309
rect 4580 1244 4752 1272
rect 4816 1244 6132 1272
rect 6196 1272 6224 1303
rect 7006 1300 7012 1312
rect 7064 1300 7070 1352
rect 7116 1340 7144 1380
rect 7282 1368 7288 1380
rect 7340 1368 7346 1420
rect 7558 1368 7564 1420
rect 7616 1408 7622 1420
rect 7745 1411 7803 1417
rect 7745 1408 7757 1411
rect 7616 1380 7757 1408
rect 7616 1368 7622 1380
rect 7745 1377 7757 1380
rect 7791 1377 7803 1411
rect 7926 1408 7932 1420
rect 7887 1380 7932 1408
rect 7745 1371 7803 1377
rect 7926 1368 7932 1380
rect 7984 1368 7990 1420
rect 8021 1343 8079 1349
rect 8021 1340 8033 1343
rect 7116 1312 8033 1340
rect 8021 1309 8033 1312
rect 8067 1309 8079 1343
rect 8021 1303 8079 1309
rect 8297 1343 8355 1349
rect 8297 1309 8309 1343
rect 8343 1340 8355 1343
rect 8496 1340 8524 1507
rect 8662 1504 8668 1516
rect 8720 1504 8726 1556
rect 9756 1547 9814 1553
rect 9756 1513 9768 1547
rect 9802 1544 9814 1547
rect 13262 1544 13268 1556
rect 9802 1516 11192 1544
rect 13223 1516 13268 1544
rect 9802 1513 9814 1516
rect 9756 1507 9814 1513
rect 11164 1488 11192 1516
rect 13262 1504 13268 1516
rect 13320 1504 13326 1556
rect 8938 1476 8944 1488
rect 8899 1448 8944 1476
rect 8938 1436 8944 1448
rect 8996 1436 9002 1488
rect 11146 1436 11152 1488
rect 11204 1476 11210 1488
rect 11204 1448 11652 1476
rect 11204 1436 11210 1448
rect 8570 1368 8576 1420
rect 8628 1408 8634 1420
rect 9493 1411 9551 1417
rect 9493 1408 9505 1411
rect 8628 1380 9505 1408
rect 8628 1368 8634 1380
rect 9493 1377 9505 1380
rect 9539 1408 9551 1411
rect 11514 1408 11520 1420
rect 9539 1380 11520 1408
rect 9539 1377 9551 1380
rect 9493 1371 9551 1377
rect 11514 1368 11520 1380
rect 11572 1368 11578 1420
rect 11624 1408 11652 1448
rect 11624 1380 13032 1408
rect 9122 1340 9128 1352
rect 8343 1312 8524 1340
rect 9083 1312 9128 1340
rect 8343 1309 8355 1312
rect 8297 1303 8355 1309
rect 9122 1300 9128 1312
rect 9180 1300 9186 1352
rect 13004 1340 13032 1380
rect 13449 1343 13507 1349
rect 13449 1340 13461 1343
rect 13004 1312 13461 1340
rect 13449 1309 13461 1312
rect 13495 1309 13507 1343
rect 13449 1303 13507 1309
rect 7098 1272 7104 1284
rect 6196 1244 7104 1272
rect 4580 1232 4586 1244
rect 4724 1213 4752 1244
rect 7098 1232 7104 1244
rect 7156 1232 7162 1284
rect 9309 1275 9367 1281
rect 9309 1241 9321 1275
rect 9355 1272 9367 1275
rect 9490 1272 9496 1284
rect 9355 1244 9496 1272
rect 9355 1241 9367 1244
rect 9309 1235 9367 1241
rect 9490 1232 9496 1244
rect 9548 1232 9554 1284
rect 11054 1272 11060 1284
rect 10994 1244 11060 1272
rect 11054 1232 11060 1244
rect 11112 1232 11118 1284
rect 11793 1275 11851 1281
rect 11793 1241 11805 1275
rect 11839 1241 11851 1275
rect 11793 1235 11851 1241
rect 3752 1176 4108 1204
rect 4709 1207 4767 1213
rect 3752 1164 3758 1176
rect 4709 1173 4721 1207
rect 4755 1173 4767 1207
rect 4709 1167 4767 1173
rect 5077 1207 5135 1213
rect 5077 1173 5089 1207
rect 5123 1204 5135 1207
rect 5442 1204 5448 1216
rect 5123 1176 5448 1204
rect 5123 1173 5135 1176
rect 5077 1167 5135 1173
rect 5442 1164 5448 1176
rect 5500 1164 5506 1216
rect 6362 1204 6368 1216
rect 6323 1176 6368 1204
rect 6362 1164 6368 1176
rect 6420 1164 6426 1216
rect 11241 1207 11299 1213
rect 11241 1173 11253 1207
rect 11287 1204 11299 1207
rect 11808 1204 11836 1235
rect 12802 1232 12808 1284
rect 12860 1232 12866 1284
rect 11287 1176 11836 1204
rect 11287 1173 11299 1176
rect 11241 1167 11299 1173
rect 1104 1114 13892 1136
rect 1104 1062 8214 1114
rect 8266 1062 8278 1114
rect 8330 1062 8342 1114
rect 8394 1062 8406 1114
rect 8458 1062 8470 1114
rect 8522 1062 13892 1114
rect 1104 1040 13892 1062
rect 3878 960 3884 1012
rect 3936 1000 3942 1012
rect 6362 1000 6368 1012
rect 3936 972 6368 1000
rect 3936 960 3942 972
rect 6362 960 6368 972
rect 6420 960 6426 1012
<< via1 >>
rect 2320 13744 2372 13796
rect 6644 13880 6696 13932
rect 1584 13676 1636 13728
rect 11244 13812 11296 13864
rect 5080 13676 5132 13728
rect 8116 13676 8168 13728
rect 4214 13574 4266 13626
rect 4278 13574 4330 13626
rect 4342 13574 4394 13626
rect 4406 13574 4458 13626
rect 4470 13574 4522 13626
rect 12214 13574 12266 13626
rect 12278 13574 12330 13626
rect 12342 13574 12394 13626
rect 12406 13574 12458 13626
rect 12470 13574 12522 13626
rect 1400 13515 1452 13524
rect 1400 13481 1409 13515
rect 1409 13481 1443 13515
rect 1443 13481 1452 13515
rect 1400 13472 1452 13481
rect 4068 13472 4120 13524
rect 1676 13404 1728 13456
rect 6920 13472 6972 13524
rect 848 13336 900 13388
rect 2320 13379 2372 13388
rect 2320 13345 2329 13379
rect 2329 13345 2363 13379
rect 2363 13345 2372 13379
rect 2320 13336 2372 13345
rect 5080 13379 5132 13388
rect 5080 13345 5089 13379
rect 5089 13345 5123 13379
rect 5123 13345 5132 13379
rect 5080 13336 5132 13345
rect 8116 13447 8168 13456
rect 8116 13413 8125 13447
rect 8125 13413 8159 13447
rect 8159 13413 8168 13447
rect 8668 13472 8720 13524
rect 8116 13404 8168 13413
rect 9036 13404 9088 13456
rect 7104 13336 7156 13388
rect 8208 13336 8260 13388
rect 14372 13472 14424 13524
rect 1584 13311 1636 13320
rect 1584 13277 1593 13311
rect 1593 13277 1627 13311
rect 1627 13277 1636 13311
rect 1584 13268 1636 13277
rect 2228 13268 2280 13320
rect 2688 13268 2740 13320
rect 2044 13243 2096 13252
rect 2044 13209 2053 13243
rect 2053 13209 2087 13243
rect 2087 13209 2096 13243
rect 2044 13200 2096 13209
rect 2136 13243 2188 13252
rect 2136 13209 2145 13243
rect 2145 13209 2179 13243
rect 2179 13209 2188 13243
rect 2872 13243 2924 13252
rect 2136 13200 2188 13209
rect 2872 13209 2881 13243
rect 2881 13209 2915 13243
rect 2915 13209 2924 13243
rect 2872 13200 2924 13209
rect 3424 13200 3476 13252
rect 3884 13268 3936 13320
rect 5724 13268 5776 13320
rect 6092 13268 6144 13320
rect 6644 13268 6696 13320
rect 7012 13311 7064 13320
rect 7012 13277 7021 13311
rect 7021 13277 7055 13311
rect 7055 13277 7064 13311
rect 7288 13311 7340 13320
rect 7012 13268 7064 13277
rect 7288 13277 7297 13311
rect 7297 13277 7331 13311
rect 7331 13277 7340 13311
rect 7288 13268 7340 13277
rect 7748 13268 7800 13320
rect 8668 13311 8720 13320
rect 8668 13277 8677 13311
rect 8677 13277 8711 13311
rect 8711 13277 8720 13311
rect 8668 13268 8720 13277
rect 8760 13268 8812 13320
rect 10600 13268 10652 13320
rect 11888 13336 11940 13388
rect 12072 13311 12124 13320
rect 5540 13243 5592 13252
rect 5540 13209 5549 13243
rect 5549 13209 5583 13243
rect 5583 13209 5592 13243
rect 5540 13200 5592 13209
rect 6000 13243 6052 13252
rect 6000 13209 6009 13243
rect 6009 13209 6043 13243
rect 6043 13209 6052 13243
rect 6000 13200 6052 13209
rect 6184 13200 6236 13252
rect 7104 13243 7156 13252
rect 7104 13209 7113 13243
rect 7113 13209 7147 13243
rect 7147 13209 7156 13243
rect 7104 13200 7156 13209
rect 7840 13243 7892 13252
rect 7840 13209 7849 13243
rect 7849 13209 7883 13243
rect 7883 13209 7892 13243
rect 7840 13200 7892 13209
rect 4252 13132 4304 13184
rect 5632 13132 5684 13184
rect 7656 13132 7708 13184
rect 8116 13200 8168 13252
rect 8484 13243 8536 13252
rect 8484 13209 8493 13243
rect 8493 13209 8527 13243
rect 8527 13209 8536 13243
rect 8484 13200 8536 13209
rect 10048 13200 10100 13252
rect 12072 13277 12081 13311
rect 12081 13277 12115 13311
rect 12115 13277 12124 13311
rect 12072 13268 12124 13277
rect 12164 13311 12216 13320
rect 12164 13277 12173 13311
rect 12173 13277 12207 13311
rect 12207 13277 12216 13311
rect 12164 13268 12216 13277
rect 12992 13268 13044 13320
rect 13176 13268 13228 13320
rect 9680 13175 9732 13184
rect 9680 13141 9689 13175
rect 9689 13141 9723 13175
rect 9723 13141 9732 13175
rect 9680 13132 9732 13141
rect 9864 13175 9916 13184
rect 9864 13141 9873 13175
rect 9873 13141 9907 13175
rect 9907 13141 9916 13175
rect 9864 13132 9916 13141
rect 9956 13175 10008 13184
rect 9956 13141 9965 13175
rect 9965 13141 9999 13175
rect 9999 13141 10008 13175
rect 10416 13175 10468 13184
rect 9956 13132 10008 13141
rect 10416 13141 10425 13175
rect 10425 13141 10459 13175
rect 10459 13141 10468 13175
rect 10416 13132 10468 13141
rect 11612 13243 11664 13252
rect 11612 13209 11621 13243
rect 11621 13209 11655 13243
rect 11655 13209 11664 13243
rect 12624 13243 12676 13252
rect 11612 13200 11664 13209
rect 12624 13209 12633 13243
rect 12633 13209 12667 13243
rect 12667 13209 12676 13243
rect 12624 13200 12676 13209
rect 13360 13243 13412 13252
rect 13360 13209 13369 13243
rect 13369 13209 13403 13243
rect 13403 13209 13412 13243
rect 13360 13200 13412 13209
rect 12900 13175 12952 13184
rect 12900 13141 12909 13175
rect 12909 13141 12943 13175
rect 12943 13141 12952 13175
rect 12900 13132 12952 13141
rect 13084 13132 13136 13184
rect 8214 13030 8266 13082
rect 8278 13030 8330 13082
rect 8342 13030 8394 13082
rect 8406 13030 8458 13082
rect 8470 13030 8522 13082
rect 3148 12928 3200 12980
rect 7104 12928 7156 12980
rect 7840 12928 7892 12980
rect 1492 12860 1544 12912
rect 3240 12860 3292 12912
rect 3700 12860 3752 12912
rect 4252 12903 4304 12912
rect 4252 12869 4261 12903
rect 4261 12869 4295 12903
rect 4295 12869 4304 12903
rect 4252 12860 4304 12869
rect 6644 12860 6696 12912
rect 7012 12860 7064 12912
rect 7288 12903 7340 12912
rect 7288 12869 7297 12903
rect 7297 12869 7331 12903
rect 7331 12869 7340 12903
rect 7288 12860 7340 12869
rect 8484 12860 8536 12912
rect 9680 12928 9732 12980
rect 10508 12928 10560 12980
rect 9864 12860 9916 12912
rect 10232 12860 10284 12912
rect 10876 12860 10928 12912
rect 1400 12792 1452 12844
rect 1860 12835 1912 12844
rect 1860 12801 1869 12835
rect 1869 12801 1903 12835
rect 1903 12801 1912 12835
rect 1860 12792 1912 12801
rect 2228 12835 2280 12844
rect 2228 12801 2237 12835
rect 2237 12801 2271 12835
rect 2271 12801 2280 12835
rect 2228 12792 2280 12801
rect 3884 12792 3936 12844
rect 4068 12835 4120 12844
rect 4068 12801 4117 12835
rect 4117 12801 4120 12835
rect 4068 12792 4120 12801
rect 4436 12792 4488 12844
rect 5724 12835 5776 12844
rect 2872 12656 2924 12708
rect 3792 12656 3844 12708
rect 5724 12801 5733 12835
rect 5733 12801 5767 12835
rect 5767 12801 5776 12835
rect 5724 12792 5776 12801
rect 6736 12835 6788 12844
rect 6460 12724 6512 12776
rect 6736 12801 6745 12835
rect 6745 12801 6779 12835
rect 6779 12801 6788 12835
rect 6736 12792 6788 12801
rect 6920 12835 6972 12844
rect 6920 12801 6934 12835
rect 6934 12801 6968 12835
rect 6968 12801 6972 12835
rect 6920 12792 6972 12801
rect 7380 12792 7432 12844
rect 7748 12792 7800 12844
rect 8760 12835 8812 12844
rect 8760 12801 8769 12835
rect 8769 12801 8803 12835
rect 8803 12801 8812 12835
rect 8760 12792 8812 12801
rect 8852 12835 8904 12844
rect 8852 12801 8861 12835
rect 8861 12801 8895 12835
rect 8895 12801 8904 12835
rect 9036 12835 9088 12844
rect 8852 12792 8904 12801
rect 9036 12801 9045 12835
rect 9045 12801 9079 12835
rect 9079 12801 9088 12835
rect 9036 12792 9088 12801
rect 7288 12724 7340 12776
rect 7656 12724 7708 12776
rect 10416 12792 10468 12844
rect 11888 12860 11940 12912
rect 10600 12767 10652 12776
rect 10600 12733 10609 12767
rect 10609 12733 10643 12767
rect 10643 12733 10652 12767
rect 10600 12724 10652 12733
rect 11796 12724 11848 12776
rect 6000 12656 6052 12708
rect 1400 12631 1452 12640
rect 1400 12597 1409 12631
rect 1409 12597 1443 12631
rect 1443 12597 1452 12631
rect 1400 12588 1452 12597
rect 4436 12588 4488 12640
rect 8484 12656 8536 12708
rect 8944 12656 8996 12708
rect 9864 12656 9916 12708
rect 12164 12792 12216 12844
rect 12624 12860 12676 12912
rect 12992 12656 13044 12708
rect 11244 12588 11296 12640
rect 4214 12486 4266 12538
rect 4278 12486 4330 12538
rect 4342 12486 4394 12538
rect 4406 12486 4458 12538
rect 4470 12486 4522 12538
rect 12214 12486 12266 12538
rect 12278 12486 12330 12538
rect 12342 12486 12394 12538
rect 12406 12486 12458 12538
rect 12470 12486 12522 12538
rect 2136 12384 2188 12436
rect 3884 12384 3936 12436
rect 7656 12427 7708 12436
rect 7656 12393 7665 12427
rect 7665 12393 7699 12427
rect 7699 12393 7708 12427
rect 7656 12384 7708 12393
rect 7748 12384 7800 12436
rect 8668 12384 8720 12436
rect 9496 12384 9548 12436
rect 10692 12384 10744 12436
rect 11980 12384 12032 12436
rect 1584 12180 1636 12232
rect 2044 12223 2096 12232
rect 2044 12189 2053 12223
rect 2053 12189 2087 12223
rect 2087 12189 2096 12223
rect 2044 12180 2096 12189
rect 2688 12223 2740 12232
rect 2688 12189 2697 12223
rect 2697 12189 2731 12223
rect 2731 12189 2740 12223
rect 3424 12223 3476 12232
rect 2688 12180 2740 12189
rect 3424 12189 3433 12223
rect 3433 12189 3467 12223
rect 3467 12189 3476 12223
rect 3424 12180 3476 12189
rect 6000 12359 6052 12368
rect 6000 12325 6009 12359
rect 6009 12325 6043 12359
rect 6043 12325 6052 12359
rect 6000 12316 6052 12325
rect 6644 12316 6696 12368
rect 6920 12316 6972 12368
rect 5632 12248 5684 12300
rect 6460 12291 6512 12300
rect 6460 12257 6469 12291
rect 6469 12257 6503 12291
rect 6503 12257 6512 12291
rect 6460 12248 6512 12257
rect 4068 12180 4120 12232
rect 4804 12223 4856 12232
rect 4804 12189 4813 12223
rect 4813 12189 4847 12223
rect 4847 12189 4856 12223
rect 4804 12180 4856 12189
rect 5080 12180 5132 12232
rect 5540 12223 5592 12232
rect 5540 12189 5549 12223
rect 5549 12189 5583 12223
rect 5583 12189 5592 12223
rect 5540 12180 5592 12189
rect 5816 12223 5868 12232
rect 5816 12189 5825 12223
rect 5825 12189 5859 12223
rect 5859 12189 5868 12223
rect 5816 12180 5868 12189
rect 6092 12180 6144 12232
rect 6276 12180 6328 12232
rect 6828 12180 6880 12232
rect 7104 12223 7156 12232
rect 7104 12189 7118 12223
rect 7118 12189 7152 12223
rect 7152 12189 7156 12223
rect 7104 12180 7156 12189
rect 2412 12112 2464 12164
rect 2872 12112 2924 12164
rect 6644 12112 6696 12164
rect 7012 12155 7064 12164
rect 7012 12121 7021 12155
rect 7021 12121 7055 12155
rect 7055 12121 7064 12155
rect 7012 12112 7064 12121
rect 8852 12248 8904 12300
rect 9036 12248 9088 12300
rect 9956 12291 10008 12300
rect 9956 12257 9965 12291
rect 9965 12257 9999 12291
rect 9999 12257 10008 12291
rect 9956 12248 10008 12257
rect 10692 12248 10744 12300
rect 11336 12248 11388 12300
rect 8668 12180 8720 12232
rect 9312 12223 9364 12232
rect 1860 12044 1912 12096
rect 5448 12044 5500 12096
rect 6552 12087 6604 12096
rect 6552 12053 6561 12087
rect 6561 12053 6595 12087
rect 6595 12053 6604 12087
rect 8116 12112 8168 12164
rect 6552 12044 6604 12053
rect 7748 12044 7800 12096
rect 8484 12044 8536 12096
rect 8668 12087 8720 12096
rect 8668 12053 8677 12087
rect 8677 12053 8711 12087
rect 8711 12053 8720 12087
rect 9312 12189 9321 12223
rect 9321 12189 9355 12223
rect 9355 12189 9364 12223
rect 9312 12180 9364 12189
rect 9864 12223 9916 12232
rect 9864 12189 9873 12223
rect 9873 12189 9907 12223
rect 9907 12189 9916 12223
rect 9864 12180 9916 12189
rect 10416 12180 10468 12232
rect 10876 12223 10928 12232
rect 10876 12189 10885 12223
rect 10885 12189 10919 12223
rect 10919 12189 10928 12223
rect 10876 12180 10928 12189
rect 11244 12180 11296 12232
rect 11612 12223 11664 12232
rect 9128 12155 9180 12164
rect 9128 12121 9137 12155
rect 9137 12121 9171 12155
rect 9171 12121 9180 12155
rect 9128 12112 9180 12121
rect 9220 12112 9272 12164
rect 11612 12189 11621 12223
rect 11621 12189 11655 12223
rect 11655 12189 11664 12223
rect 11612 12180 11664 12189
rect 11888 12223 11940 12232
rect 11888 12189 11897 12223
rect 11897 12189 11931 12223
rect 11931 12189 11940 12223
rect 11888 12180 11940 12189
rect 12808 12180 12860 12232
rect 12992 12223 13044 12232
rect 12992 12189 13001 12223
rect 13001 12189 13035 12223
rect 13035 12189 13044 12223
rect 12992 12180 13044 12189
rect 10692 12087 10744 12096
rect 8668 12044 8720 12053
rect 10692 12053 10701 12087
rect 10701 12053 10735 12087
rect 10735 12053 10744 12087
rect 10692 12044 10744 12053
rect 12072 12112 12124 12164
rect 13268 12112 13320 12164
rect 11428 12044 11480 12096
rect 8214 11942 8266 11994
rect 8278 11942 8330 11994
rect 8342 11942 8394 11994
rect 8406 11942 8458 11994
rect 8470 11942 8522 11994
rect 2044 11840 2096 11892
rect 4068 11840 4120 11892
rect 6552 11840 6604 11892
rect 6828 11883 6880 11892
rect 6828 11849 6837 11883
rect 6837 11849 6871 11883
rect 6871 11849 6880 11883
rect 6828 11840 6880 11849
rect 1400 11772 1452 11824
rect 3148 11772 3200 11824
rect 3792 11815 3844 11824
rect 3792 11781 3801 11815
rect 3801 11781 3835 11815
rect 3835 11781 3844 11815
rect 3792 11772 3844 11781
rect 5448 11772 5500 11824
rect 7840 11840 7892 11892
rect 8392 11883 8444 11892
rect 2504 11747 2556 11756
rect 2504 11713 2513 11747
rect 2513 11713 2547 11747
rect 2547 11713 2556 11747
rect 2504 11704 2556 11713
rect 2688 11704 2740 11756
rect 5080 11704 5132 11756
rect 2228 11636 2280 11688
rect 4712 11636 4764 11688
rect 4988 11636 5040 11688
rect 5632 11636 5684 11688
rect 2872 11568 2924 11620
rect 3148 11543 3200 11552
rect 3148 11509 3157 11543
rect 3157 11509 3191 11543
rect 3191 11509 3200 11543
rect 3700 11568 3752 11620
rect 3148 11500 3200 11509
rect 3884 11543 3936 11552
rect 3884 11509 3893 11543
rect 3893 11509 3927 11543
rect 3927 11509 3936 11543
rect 3884 11500 3936 11509
rect 4620 11568 4672 11620
rect 5540 11568 5592 11620
rect 6000 11747 6052 11756
rect 6000 11713 6009 11747
rect 6009 11713 6043 11747
rect 6043 11713 6052 11747
rect 6000 11704 6052 11713
rect 6184 11747 6236 11756
rect 6184 11713 6193 11747
rect 6193 11713 6227 11747
rect 6227 11713 6236 11747
rect 6184 11704 6236 11713
rect 6736 11704 6788 11756
rect 7288 11772 7340 11824
rect 7748 11772 7800 11824
rect 8392 11849 8401 11883
rect 8401 11849 8435 11883
rect 8435 11849 8444 11883
rect 8392 11840 8444 11849
rect 8668 11840 8720 11892
rect 7380 11747 7432 11756
rect 6460 11636 6512 11688
rect 6552 11568 6604 11620
rect 6736 11568 6788 11620
rect 7380 11713 7389 11747
rect 7389 11713 7423 11747
rect 7423 11713 7432 11747
rect 7656 11747 7708 11756
rect 7380 11704 7432 11713
rect 7656 11713 7665 11747
rect 7665 11713 7699 11747
rect 7699 11713 7708 11747
rect 7656 11704 7708 11713
rect 7840 11747 7892 11756
rect 7840 11713 7849 11747
rect 7849 11713 7883 11747
rect 7883 11713 7892 11747
rect 7840 11704 7892 11713
rect 8208 11747 8260 11756
rect 8208 11713 8217 11747
rect 8217 11713 8251 11747
rect 8251 11713 8260 11747
rect 8208 11704 8260 11713
rect 8760 11815 8812 11824
rect 7748 11636 7800 11688
rect 8760 11781 8769 11815
rect 8769 11781 8803 11815
rect 8803 11781 8812 11815
rect 8760 11772 8812 11781
rect 9588 11772 9640 11824
rect 10784 11840 10836 11892
rect 11980 11840 12032 11892
rect 13176 11840 13228 11892
rect 13452 11883 13504 11892
rect 13452 11849 13461 11883
rect 13461 11849 13495 11883
rect 13495 11849 13504 11883
rect 13452 11840 13504 11849
rect 10600 11772 10652 11824
rect 10692 11772 10744 11824
rect 12900 11772 12952 11824
rect 13360 11815 13412 11824
rect 13360 11781 13369 11815
rect 13369 11781 13403 11815
rect 13403 11781 13412 11815
rect 13360 11772 13412 11781
rect 9496 11747 9548 11756
rect 9496 11713 9505 11747
rect 9505 11713 9539 11747
rect 9539 11713 9548 11747
rect 9496 11704 9548 11713
rect 9680 11747 9732 11756
rect 9680 11713 9688 11747
rect 9688 11713 9722 11747
rect 9722 11713 9732 11747
rect 9864 11747 9916 11756
rect 9680 11704 9732 11713
rect 9864 11713 9873 11747
rect 9873 11713 9907 11747
rect 9907 11713 9916 11747
rect 9864 11704 9916 11713
rect 9956 11704 10008 11756
rect 9404 11636 9456 11688
rect 11152 11704 11204 11756
rect 11704 11747 11756 11756
rect 11704 11713 11713 11747
rect 11713 11713 11747 11747
rect 11747 11713 11756 11747
rect 11704 11704 11756 11713
rect 13084 11704 13136 11756
rect 13268 11747 13320 11756
rect 13268 11713 13277 11747
rect 13277 11713 13311 11747
rect 13311 11713 13320 11747
rect 13268 11704 13320 11713
rect 8208 11568 8260 11620
rect 9220 11568 9272 11620
rect 11336 11636 11388 11688
rect 12072 11636 12124 11688
rect 12808 11679 12860 11688
rect 12808 11645 12817 11679
rect 12817 11645 12851 11679
rect 12851 11645 12860 11679
rect 12808 11636 12860 11645
rect 10048 11568 10100 11620
rect 4804 11500 4856 11552
rect 6460 11500 6512 11552
rect 7380 11500 7432 11552
rect 8392 11500 8444 11552
rect 8668 11500 8720 11552
rect 9036 11500 9088 11552
rect 9496 11500 9548 11552
rect 10692 11543 10744 11552
rect 10692 11509 10701 11543
rect 10701 11509 10735 11543
rect 10735 11509 10744 11543
rect 10692 11500 10744 11509
rect 10876 11500 10928 11552
rect 11060 11500 11112 11552
rect 4214 11398 4266 11450
rect 4278 11398 4330 11450
rect 4342 11398 4394 11450
rect 4406 11398 4458 11450
rect 4470 11398 4522 11450
rect 12214 11398 12266 11450
rect 12278 11398 12330 11450
rect 12342 11398 12394 11450
rect 12406 11398 12458 11450
rect 12470 11398 12522 11450
rect 8668 11339 8720 11348
rect 8668 11305 8677 11339
rect 8677 11305 8711 11339
rect 8711 11305 8720 11339
rect 8668 11296 8720 11305
rect 8852 11296 8904 11348
rect 9128 11339 9180 11348
rect 9128 11305 9137 11339
rect 9137 11305 9171 11339
rect 9171 11305 9180 11339
rect 9128 11296 9180 11305
rect 2872 11271 2924 11280
rect 2872 11237 2881 11271
rect 2881 11237 2915 11271
rect 2915 11237 2924 11271
rect 2872 11228 2924 11237
rect 3516 11228 3568 11280
rect 5080 11271 5132 11280
rect 5080 11237 5089 11271
rect 5089 11237 5123 11271
rect 5123 11237 5132 11271
rect 5080 11228 5132 11237
rect 6092 11228 6144 11280
rect 4528 11160 4580 11212
rect 5172 11160 5224 11212
rect 2228 11092 2280 11144
rect 2412 11135 2464 11144
rect 2412 11101 2421 11135
rect 2421 11101 2455 11135
rect 2455 11101 2464 11135
rect 2412 11092 2464 11101
rect 3332 11092 3384 11144
rect 3884 11092 3936 11144
rect 4804 11092 4856 11144
rect 6552 11113 6604 11144
rect 6552 11092 6560 11113
rect 6560 11092 6594 11113
rect 6594 11092 6604 11113
rect 3516 11067 3568 11076
rect 3516 11033 3525 11067
rect 3525 11033 3559 11067
rect 3559 11033 3568 11067
rect 3516 11024 3568 11033
rect 3608 11067 3660 11076
rect 3608 11033 3617 11067
rect 3617 11033 3651 11067
rect 3651 11033 3660 11067
rect 3608 11024 3660 11033
rect 2688 10956 2740 11008
rect 5908 11024 5960 11076
rect 6092 11067 6144 11076
rect 6092 11033 6101 11067
rect 6101 11033 6135 11067
rect 6135 11033 6144 11067
rect 6092 11024 6144 11033
rect 6276 11067 6328 11076
rect 6276 11033 6285 11067
rect 6285 11033 6319 11067
rect 6319 11033 6328 11067
rect 6276 11024 6328 11033
rect 6000 10999 6052 11008
rect 6000 10965 6009 10999
rect 6009 10965 6043 10999
rect 6043 10965 6052 10999
rect 7012 11135 7064 11144
rect 7012 11101 7021 11135
rect 7021 11101 7055 11135
rect 7055 11101 7064 11135
rect 7748 11228 7800 11280
rect 7840 11228 7892 11280
rect 8576 11228 8628 11280
rect 7288 11160 7340 11212
rect 7564 11160 7616 11212
rect 8300 11160 8352 11212
rect 7012 11092 7064 11101
rect 8024 11092 8076 11144
rect 8668 11160 8720 11212
rect 9128 11160 9180 11212
rect 7288 11024 7340 11076
rect 7564 11024 7616 11076
rect 9036 11092 9088 11144
rect 9312 11296 9364 11348
rect 9772 11296 9824 11348
rect 11244 11296 11296 11348
rect 11980 11339 12032 11348
rect 11980 11305 11989 11339
rect 11989 11305 12023 11339
rect 12023 11305 12032 11339
rect 11980 11296 12032 11305
rect 10048 11228 10100 11280
rect 10692 11228 10744 11280
rect 9312 11203 9364 11212
rect 9312 11169 9321 11203
rect 9321 11169 9355 11203
rect 9355 11169 9364 11203
rect 11060 11203 11112 11212
rect 9312 11160 9364 11169
rect 11060 11169 11069 11203
rect 11069 11169 11103 11203
rect 11103 11169 11112 11203
rect 11060 11160 11112 11169
rect 11796 11228 11848 11280
rect 13452 11228 13504 11280
rect 13544 11203 13596 11212
rect 9588 11135 9640 11144
rect 9588 11101 9597 11135
rect 9597 11101 9631 11135
rect 9631 11101 9640 11135
rect 9588 11092 9640 11101
rect 9680 11135 9732 11144
rect 9680 11101 9689 11135
rect 9689 11101 9723 11135
rect 9723 11101 9732 11135
rect 9680 11092 9732 11101
rect 10048 11092 10100 11144
rect 10324 11135 10376 11144
rect 10324 11101 10333 11135
rect 10333 11101 10367 11135
rect 10367 11101 10376 11135
rect 10324 11092 10376 11101
rect 10600 11135 10652 11144
rect 10600 11101 10609 11135
rect 10609 11101 10643 11135
rect 10643 11101 10652 11135
rect 10600 11092 10652 11101
rect 13544 11169 13553 11203
rect 13553 11169 13587 11203
rect 13587 11169 13596 11203
rect 13544 11160 13596 11169
rect 6000 10956 6052 10965
rect 6736 10956 6788 11008
rect 7932 10956 7984 11008
rect 9956 11024 10008 11076
rect 10508 11067 10560 11076
rect 10508 11033 10517 11067
rect 10517 11033 10551 11067
rect 10551 11033 10560 11067
rect 10508 11024 10560 11033
rect 10968 11024 11020 11076
rect 12072 11135 12124 11144
rect 12072 11101 12081 11135
rect 12081 11101 12115 11135
rect 12115 11101 12124 11135
rect 12072 11092 12124 11101
rect 12992 11135 13044 11144
rect 12992 11101 13001 11135
rect 13001 11101 13035 11135
rect 13035 11101 13044 11135
rect 12992 11092 13044 11101
rect 13268 11135 13320 11144
rect 13268 11101 13277 11135
rect 13277 11101 13311 11135
rect 13311 11101 13320 11135
rect 13268 11092 13320 11101
rect 9036 10956 9088 11008
rect 10692 10956 10744 11008
rect 11336 10956 11388 11008
rect 11980 11024 12032 11076
rect 12256 11024 12308 11076
rect 13084 11024 13136 11076
rect 12532 10956 12584 11008
rect 12716 10956 12768 11008
rect 8214 10854 8266 10906
rect 8278 10854 8330 10906
rect 8342 10854 8394 10906
rect 8406 10854 8458 10906
rect 8470 10854 8522 10906
rect 2412 10795 2464 10804
rect 2412 10761 2421 10795
rect 2421 10761 2455 10795
rect 2455 10761 2464 10795
rect 2412 10752 2464 10761
rect 2780 10752 2832 10804
rect 1584 10659 1636 10668
rect 2688 10684 2740 10736
rect 4528 10752 4580 10804
rect 4712 10752 4764 10804
rect 5816 10795 5868 10804
rect 5816 10761 5825 10795
rect 5825 10761 5859 10795
rect 5859 10761 5868 10795
rect 5816 10752 5868 10761
rect 5908 10752 5960 10804
rect 6276 10752 6328 10804
rect 3332 10727 3384 10736
rect 3332 10693 3341 10727
rect 3341 10693 3375 10727
rect 3375 10693 3384 10727
rect 3332 10684 3384 10693
rect 3608 10684 3660 10736
rect 4620 10684 4672 10736
rect 6460 10684 6512 10736
rect 7012 10727 7064 10736
rect 7012 10693 7021 10727
rect 7021 10693 7055 10727
rect 7055 10693 7064 10727
rect 7012 10684 7064 10693
rect 7380 10727 7432 10736
rect 7380 10693 7389 10727
rect 7389 10693 7423 10727
rect 7423 10693 7432 10727
rect 7380 10684 7432 10693
rect 7932 10727 7984 10736
rect 7932 10693 7941 10727
rect 7941 10693 7975 10727
rect 7975 10693 7984 10727
rect 7932 10684 7984 10693
rect 8392 10752 8444 10804
rect 8944 10752 8996 10804
rect 1584 10625 1633 10659
rect 1633 10625 1636 10659
rect 1584 10616 1636 10625
rect 1400 10480 1452 10532
rect 2780 10616 2832 10668
rect 2688 10548 2740 10600
rect 3884 10616 3936 10668
rect 4988 10659 5040 10668
rect 4988 10625 4997 10659
rect 4997 10625 5031 10659
rect 5031 10625 5040 10659
rect 4988 10616 5040 10625
rect 5264 10659 5316 10668
rect 5264 10625 5273 10659
rect 5273 10625 5307 10659
rect 5307 10625 5316 10659
rect 5264 10616 5316 10625
rect 6736 10616 6788 10668
rect 7656 10616 7708 10668
rect 7840 10659 7892 10668
rect 7840 10625 7844 10659
rect 7844 10625 7878 10659
rect 7878 10625 7892 10659
rect 7840 10616 7892 10625
rect 8208 10659 8260 10668
rect 8208 10625 8217 10659
rect 8217 10625 8251 10659
rect 8251 10625 8260 10659
rect 8208 10616 8260 10625
rect 8760 10684 8812 10736
rect 9220 10684 9272 10736
rect 9680 10684 9732 10736
rect 10324 10752 10376 10804
rect 9128 10659 9180 10668
rect 5908 10548 5960 10600
rect 1492 10455 1544 10464
rect 1492 10421 1501 10455
rect 1501 10421 1535 10455
rect 1535 10421 1544 10455
rect 1492 10412 1544 10421
rect 2136 10455 2188 10464
rect 2136 10421 2145 10455
rect 2145 10421 2179 10455
rect 2179 10421 2188 10455
rect 2136 10412 2188 10421
rect 6276 10480 6328 10532
rect 3148 10412 3200 10464
rect 4620 10412 4672 10464
rect 5356 10412 5408 10464
rect 6000 10455 6052 10464
rect 6000 10421 6009 10455
rect 6009 10421 6043 10455
rect 6043 10421 6052 10455
rect 6000 10412 6052 10421
rect 6184 10412 6236 10464
rect 6828 10548 6880 10600
rect 7104 10548 7156 10600
rect 7288 10548 7340 10600
rect 9128 10625 9137 10659
rect 9137 10625 9171 10659
rect 9171 10625 9180 10659
rect 9128 10616 9180 10625
rect 9404 10616 9456 10668
rect 9588 10659 9640 10668
rect 9588 10625 9597 10659
rect 9597 10625 9631 10659
rect 9631 10625 9640 10659
rect 9588 10616 9640 10625
rect 10692 10684 10744 10736
rect 11336 10659 11388 10668
rect 8944 10591 8996 10600
rect 8944 10557 8953 10591
rect 8953 10557 8987 10591
rect 8987 10557 8996 10591
rect 8944 10548 8996 10557
rect 7380 10480 7432 10532
rect 8392 10480 8444 10532
rect 8576 10480 8628 10532
rect 11336 10625 11345 10659
rect 11345 10625 11379 10659
rect 11379 10625 11388 10659
rect 11336 10616 11388 10625
rect 11796 10659 11848 10668
rect 11796 10625 11800 10659
rect 11800 10625 11834 10659
rect 11834 10625 11848 10659
rect 11796 10616 11848 10625
rect 12256 10684 12308 10736
rect 12164 10659 12216 10668
rect 9864 10548 9916 10600
rect 11244 10548 11296 10600
rect 12164 10625 12173 10659
rect 12173 10625 12207 10659
rect 12207 10625 12216 10659
rect 12164 10616 12216 10625
rect 12624 10616 12676 10668
rect 12072 10548 12124 10600
rect 12348 10548 12400 10600
rect 12900 10591 12952 10600
rect 12900 10557 12909 10591
rect 12909 10557 12943 10591
rect 12943 10557 12952 10591
rect 12900 10548 12952 10557
rect 13360 10523 13412 10532
rect 13360 10489 13369 10523
rect 13369 10489 13403 10523
rect 13403 10489 13412 10523
rect 13360 10480 13412 10489
rect 9956 10412 10008 10464
rect 10600 10412 10652 10464
rect 10876 10455 10928 10464
rect 10876 10421 10885 10455
rect 10885 10421 10919 10455
rect 10919 10421 10928 10455
rect 10876 10412 10928 10421
rect 11704 10412 11756 10464
rect 11980 10412 12032 10464
rect 12256 10412 12308 10464
rect 4214 10310 4266 10362
rect 4278 10310 4330 10362
rect 4342 10310 4394 10362
rect 4406 10310 4458 10362
rect 4470 10310 4522 10362
rect 12214 10310 12266 10362
rect 12278 10310 12330 10362
rect 12342 10310 12394 10362
rect 12406 10310 12458 10362
rect 12470 10310 12522 10362
rect 1400 10251 1452 10260
rect 1400 10217 1409 10251
rect 1409 10217 1443 10251
rect 1443 10217 1452 10251
rect 1400 10208 1452 10217
rect 2872 10208 2924 10260
rect 3332 10208 3384 10260
rect 5816 10208 5868 10260
rect 7196 10208 7248 10260
rect 8484 10208 8536 10260
rect 9496 10208 9548 10260
rect 1492 10072 1544 10124
rect 2688 10140 2740 10192
rect 8208 10183 8260 10192
rect 4620 10115 4672 10124
rect 4620 10081 4629 10115
rect 4629 10081 4663 10115
rect 4663 10081 4672 10115
rect 4620 10072 4672 10081
rect 2412 10047 2464 10056
rect 2412 10013 2421 10047
rect 2421 10013 2455 10047
rect 2455 10013 2464 10047
rect 2872 10047 2924 10056
rect 2412 10004 2464 10013
rect 2872 10013 2881 10047
rect 2881 10013 2915 10047
rect 2915 10013 2924 10047
rect 2872 10004 2924 10013
rect 2780 9936 2832 9988
rect 2964 9979 3016 9988
rect 2964 9945 2973 9979
rect 2973 9945 3007 9979
rect 3007 9945 3016 9979
rect 2964 9936 3016 9945
rect 3332 10047 3384 10056
rect 3332 10013 3341 10047
rect 3341 10013 3375 10047
rect 3375 10013 3384 10047
rect 3332 10004 3384 10013
rect 3700 10004 3752 10056
rect 5356 10047 5408 10056
rect 5356 10013 5365 10047
rect 5365 10013 5399 10047
rect 5399 10013 5408 10047
rect 5356 10004 5408 10013
rect 5540 10047 5592 10056
rect 5540 10013 5549 10047
rect 5549 10013 5583 10047
rect 5583 10013 5592 10047
rect 5540 10004 5592 10013
rect 7656 10072 7708 10124
rect 7840 10072 7892 10124
rect 8208 10149 8217 10183
rect 8217 10149 8251 10183
rect 8251 10149 8260 10183
rect 8208 10140 8260 10149
rect 8484 10072 8536 10124
rect 6368 10004 6420 10056
rect 6644 10047 6696 10056
rect 6644 10013 6653 10047
rect 6653 10013 6687 10047
rect 6687 10013 6696 10047
rect 6644 10004 6696 10013
rect 6828 10047 6880 10056
rect 6828 10013 6837 10047
rect 6837 10013 6871 10047
rect 6871 10013 6880 10047
rect 6828 10004 6880 10013
rect 4528 9979 4580 9988
rect 2136 9868 2188 9920
rect 4528 9945 4537 9979
rect 4537 9945 4571 9979
rect 4571 9945 4580 9979
rect 4528 9936 4580 9945
rect 4988 9979 5040 9988
rect 4988 9945 4997 9979
rect 4997 9945 5031 9979
rect 5031 9945 5040 9979
rect 4988 9936 5040 9945
rect 5172 9979 5224 9988
rect 5172 9945 5181 9979
rect 5181 9945 5215 9979
rect 5215 9945 5224 9979
rect 5172 9936 5224 9945
rect 3148 9911 3200 9920
rect 3148 9877 3157 9911
rect 3157 9877 3191 9911
rect 3191 9877 3200 9911
rect 3148 9868 3200 9877
rect 3976 9868 4028 9920
rect 6736 9936 6788 9988
rect 7104 10004 7156 10056
rect 7564 10047 7616 10056
rect 7564 10013 7573 10047
rect 7573 10013 7607 10047
rect 7607 10013 7616 10047
rect 7564 10004 7616 10013
rect 7748 10047 7800 10056
rect 7748 10013 7757 10047
rect 7757 10013 7791 10047
rect 7791 10013 7800 10047
rect 7748 10004 7800 10013
rect 8576 10047 8628 10056
rect 8576 10013 8585 10047
rect 8585 10013 8619 10047
rect 8619 10013 8628 10047
rect 8576 10004 8628 10013
rect 8944 10072 8996 10124
rect 10968 10208 11020 10260
rect 9864 10183 9916 10192
rect 9864 10149 9873 10183
rect 9873 10149 9907 10183
rect 9907 10149 9916 10183
rect 9864 10140 9916 10149
rect 11060 10140 11112 10192
rect 9772 10072 9824 10124
rect 10416 10072 10468 10124
rect 10692 10072 10744 10124
rect 9588 10004 9640 10056
rect 10600 10047 10652 10056
rect 10600 10013 10609 10047
rect 10609 10013 10643 10047
rect 10643 10013 10652 10047
rect 10600 10004 10652 10013
rect 10784 10047 10836 10056
rect 10784 10013 10793 10047
rect 10793 10013 10827 10047
rect 10827 10013 10836 10047
rect 10784 10004 10836 10013
rect 6184 9868 6236 9920
rect 7196 9868 7248 9920
rect 7840 9868 7892 9920
rect 9772 9936 9824 9988
rect 10140 9936 10192 9988
rect 10324 9979 10376 9988
rect 10324 9945 10343 9979
rect 10343 9945 10376 9979
rect 10324 9936 10376 9945
rect 11796 10072 11848 10124
rect 11060 10047 11112 10056
rect 11060 10013 11069 10047
rect 11069 10013 11103 10047
rect 11103 10013 11112 10047
rect 11060 10004 11112 10013
rect 11152 10004 11204 10056
rect 12900 10140 12952 10192
rect 13360 10183 13412 10192
rect 13360 10149 13369 10183
rect 13369 10149 13403 10183
rect 13403 10149 13412 10183
rect 13360 10140 13412 10149
rect 12716 10004 12768 10056
rect 11244 9936 11296 9988
rect 11796 9936 11848 9988
rect 8392 9868 8444 9920
rect 9312 9868 9364 9920
rect 9496 9868 9548 9920
rect 10600 9868 10652 9920
rect 8214 9766 8266 9818
rect 8278 9766 8330 9818
rect 8342 9766 8394 9818
rect 8406 9766 8458 9818
rect 8470 9766 8522 9818
rect 6460 9664 6512 9716
rect 7012 9664 7064 9716
rect 7472 9664 7524 9716
rect 7748 9664 7800 9716
rect 1768 9596 1820 9648
rect 4528 9596 4580 9648
rect 5264 9596 5316 9648
rect 8392 9664 8444 9716
rect 8852 9707 8904 9716
rect 8852 9673 8861 9707
rect 8861 9673 8895 9707
rect 8895 9673 8904 9707
rect 8852 9664 8904 9673
rect 9220 9664 9272 9716
rect 1492 9528 1544 9580
rect 3240 9528 3292 9580
rect 3700 9571 3752 9580
rect 3700 9537 3709 9571
rect 3709 9537 3743 9571
rect 3743 9537 3752 9571
rect 3700 9528 3752 9537
rect 5172 9571 5224 9580
rect 5172 9537 5181 9571
rect 5181 9537 5215 9571
rect 5215 9537 5224 9571
rect 5172 9528 5224 9537
rect 6644 9571 6696 9580
rect 6644 9537 6648 9571
rect 6648 9537 6682 9571
rect 6682 9537 6696 9571
rect 6644 9528 6696 9537
rect 6736 9571 6788 9580
rect 6736 9537 6748 9571
rect 6748 9537 6782 9571
rect 6782 9537 6788 9571
rect 6736 9528 6788 9537
rect 5908 9503 5960 9512
rect 2780 9392 2832 9444
rect 4528 9392 4580 9444
rect 5908 9469 5917 9503
rect 5917 9469 5951 9503
rect 5951 9469 5960 9503
rect 5908 9460 5960 9469
rect 6828 9392 6880 9444
rect 7656 9528 7708 9580
rect 8116 9528 8168 9580
rect 8484 9571 8536 9580
rect 8484 9537 8492 9571
rect 8492 9537 8526 9571
rect 8526 9537 8536 9571
rect 8484 9528 8536 9537
rect 8760 9571 8812 9580
rect 8760 9537 8764 9571
rect 8764 9537 8798 9571
rect 8798 9537 8812 9571
rect 9772 9664 9824 9716
rect 10140 9664 10192 9716
rect 10784 9707 10836 9716
rect 10784 9673 10793 9707
rect 10793 9673 10827 9707
rect 10827 9673 10836 9707
rect 10784 9664 10836 9673
rect 11244 9664 11296 9716
rect 9864 9596 9916 9648
rect 10692 9639 10744 9648
rect 10692 9605 10701 9639
rect 10701 9605 10735 9639
rect 10735 9605 10744 9639
rect 10692 9596 10744 9605
rect 8760 9528 8812 9537
rect 7196 9460 7248 9512
rect 7840 9460 7892 9512
rect 7564 9435 7616 9444
rect 7564 9401 7573 9435
rect 7573 9401 7607 9435
rect 7607 9401 7616 9435
rect 7564 9392 7616 9401
rect 9312 9460 9364 9512
rect 9680 9460 9732 9512
rect 9956 9460 10008 9512
rect 10232 9460 10284 9512
rect 6184 9324 6236 9376
rect 6644 9324 6696 9376
rect 8024 9392 8076 9444
rect 9864 9392 9916 9444
rect 10048 9392 10100 9444
rect 10416 9528 10468 9580
rect 11152 9571 11204 9580
rect 11152 9537 11161 9571
rect 11161 9537 11195 9571
rect 11195 9537 11204 9571
rect 11152 9528 11204 9537
rect 12808 9639 12860 9648
rect 12808 9605 12817 9639
rect 12817 9605 12851 9639
rect 12851 9605 12860 9639
rect 12808 9596 12860 9605
rect 13360 9596 13412 9648
rect 11612 9460 11664 9512
rect 11428 9392 11480 9444
rect 7932 9324 7984 9376
rect 8852 9324 8904 9376
rect 9404 9367 9456 9376
rect 9404 9333 9413 9367
rect 9413 9333 9447 9367
rect 9447 9333 9456 9367
rect 9404 9324 9456 9333
rect 10140 9324 10192 9376
rect 11336 9324 11388 9376
rect 12072 9528 12124 9580
rect 12716 9528 12768 9580
rect 13452 9435 13504 9444
rect 13452 9401 13461 9435
rect 13461 9401 13495 9435
rect 13495 9401 13504 9435
rect 13452 9392 13504 9401
rect 4214 9222 4266 9274
rect 4278 9222 4330 9274
rect 4342 9222 4394 9274
rect 4406 9222 4458 9274
rect 4470 9222 4522 9274
rect 12214 9222 12266 9274
rect 12278 9222 12330 9274
rect 12342 9222 12394 9274
rect 12406 9222 12458 9274
rect 12470 9222 12522 9274
rect 1584 9120 1636 9172
rect 2964 9120 3016 9172
rect 6552 9120 6604 9172
rect 3516 9052 3568 9104
rect 5724 9052 5776 9104
rect 7104 9120 7156 9172
rect 8024 9120 8076 9172
rect 8392 9120 8444 9172
rect 8944 9120 8996 9172
rect 9128 9163 9180 9172
rect 9128 9129 9137 9163
rect 9137 9129 9171 9163
rect 9171 9129 9180 9163
rect 9680 9163 9732 9172
rect 9128 9120 9180 9129
rect 9680 9129 9689 9163
rect 9689 9129 9723 9163
rect 9723 9129 9732 9163
rect 9680 9120 9732 9129
rect 9956 9120 10008 9172
rect 11244 9120 11296 9172
rect 12072 9163 12124 9172
rect 2596 8916 2648 8968
rect 1768 8823 1820 8832
rect 1768 8789 1777 8823
rect 1777 8789 1811 8823
rect 1811 8789 1820 8823
rect 1768 8780 1820 8789
rect 2136 8823 2188 8832
rect 2136 8789 2145 8823
rect 2145 8789 2179 8823
rect 2179 8789 2188 8823
rect 2872 8916 2924 8968
rect 3240 8959 3292 8968
rect 3240 8925 3249 8959
rect 3249 8925 3283 8959
rect 3283 8925 3292 8959
rect 3240 8916 3292 8925
rect 4620 8916 4672 8968
rect 5264 8916 5316 8968
rect 3976 8848 4028 8900
rect 4252 8891 4304 8900
rect 4252 8857 4261 8891
rect 4261 8857 4295 8891
rect 4295 8857 4304 8891
rect 4252 8848 4304 8857
rect 5172 8848 5224 8900
rect 5908 8916 5960 8968
rect 6460 8984 6512 9036
rect 6552 8959 6604 8968
rect 6552 8925 6561 8959
rect 6561 8925 6595 8959
rect 6595 8925 6604 8959
rect 6552 8916 6604 8925
rect 7012 8984 7064 9036
rect 7104 8959 7156 8968
rect 6828 8891 6880 8900
rect 6828 8857 6837 8891
rect 6837 8857 6871 8891
rect 6871 8857 6880 8891
rect 6828 8848 6880 8857
rect 7104 8925 7113 8959
rect 7113 8925 7147 8959
rect 7147 8925 7156 8959
rect 7104 8916 7156 8925
rect 7840 8959 7892 8968
rect 7840 8925 7849 8959
rect 7849 8925 7883 8959
rect 7883 8925 7892 8959
rect 7840 8916 7892 8925
rect 8208 8916 8260 8968
rect 2136 8780 2188 8789
rect 5448 8780 5500 8832
rect 5724 8823 5776 8832
rect 5724 8789 5733 8823
rect 5733 8789 5767 8823
rect 5767 8789 5776 8823
rect 5724 8780 5776 8789
rect 7564 8848 7616 8900
rect 8668 9052 8720 9104
rect 8852 9052 8904 9104
rect 9404 9052 9456 9104
rect 9772 9052 9824 9104
rect 11612 9052 11664 9104
rect 9036 9027 9088 9036
rect 9036 8993 9045 9027
rect 9045 8993 9079 9027
rect 9079 8993 9088 9027
rect 9036 8984 9088 8993
rect 9312 8984 9364 9036
rect 9588 8984 9640 9036
rect 8576 8916 8628 8968
rect 8760 8916 8812 8968
rect 10048 8984 10100 9036
rect 10876 8984 10928 9036
rect 10140 8959 10192 8968
rect 10140 8925 10149 8959
rect 10149 8925 10183 8959
rect 10183 8925 10192 8959
rect 10140 8916 10192 8925
rect 11336 8916 11388 8968
rect 10232 8848 10284 8900
rect 9128 8780 9180 8832
rect 10692 8780 10744 8832
rect 10876 8848 10928 8900
rect 12072 9129 12081 9163
rect 12081 9129 12115 9163
rect 12115 9129 12124 9163
rect 12072 9120 12124 9129
rect 12348 9052 12400 9104
rect 11888 8916 11940 8968
rect 13268 8916 13320 8968
rect 12900 8848 12952 8900
rect 13084 8891 13136 8900
rect 13084 8857 13093 8891
rect 13093 8857 13127 8891
rect 13127 8857 13136 8891
rect 13084 8848 13136 8857
rect 11336 8780 11388 8832
rect 8214 8678 8266 8730
rect 8278 8678 8330 8730
rect 8342 8678 8394 8730
rect 8406 8678 8458 8730
rect 8470 8678 8522 8730
rect 5540 8576 5592 8628
rect 6552 8576 6604 8628
rect 4988 8508 5040 8560
rect 5448 8551 5500 8560
rect 5448 8517 5457 8551
rect 5457 8517 5491 8551
rect 5491 8517 5500 8551
rect 5448 8508 5500 8517
rect 6828 8508 6880 8560
rect 7564 8576 7616 8628
rect 9312 8576 9364 8628
rect 9496 8619 9548 8628
rect 9496 8585 9505 8619
rect 9505 8585 9539 8619
rect 9539 8585 9548 8619
rect 9496 8576 9548 8585
rect 9588 8576 9640 8628
rect 8116 8508 8168 8560
rect 1492 8483 1544 8492
rect 1492 8449 1501 8483
rect 1501 8449 1535 8483
rect 1535 8449 1544 8483
rect 1492 8440 1544 8449
rect 4252 8440 4304 8492
rect 5264 8483 5316 8492
rect 5264 8449 5273 8483
rect 5273 8449 5307 8483
rect 5307 8449 5316 8483
rect 5264 8440 5316 8449
rect 6184 8483 6236 8492
rect 6184 8449 6193 8483
rect 6193 8449 6227 8483
rect 6227 8449 6236 8483
rect 6184 8440 6236 8449
rect 6552 8483 6604 8492
rect 6552 8449 6561 8483
rect 6561 8449 6595 8483
rect 6595 8449 6604 8483
rect 6552 8440 6604 8449
rect 7012 8483 7064 8492
rect 2964 8347 3016 8356
rect 2964 8313 2973 8347
rect 2973 8313 3007 8347
rect 3007 8313 3016 8347
rect 2964 8304 3016 8313
rect 7012 8449 7021 8483
rect 7021 8449 7055 8483
rect 7055 8449 7064 8483
rect 7012 8440 7064 8449
rect 7840 8440 7892 8492
rect 9956 8508 10008 8560
rect 11152 8576 11204 8628
rect 11704 8576 11756 8628
rect 11612 8508 11664 8560
rect 11980 8576 12032 8628
rect 6920 8415 6972 8424
rect 6920 8381 6929 8415
rect 6929 8381 6963 8415
rect 6963 8381 6972 8415
rect 6920 8372 6972 8381
rect 8024 8415 8076 8424
rect 8024 8381 8033 8415
rect 8033 8381 8067 8415
rect 8067 8381 8076 8415
rect 8024 8372 8076 8381
rect 9496 8372 9548 8424
rect 9864 8440 9916 8492
rect 10416 8440 10468 8492
rect 12716 8508 12768 8560
rect 13084 8551 13136 8560
rect 13084 8517 13093 8551
rect 13093 8517 13127 8551
rect 13127 8517 13136 8551
rect 13084 8508 13136 8517
rect 12348 8483 12400 8492
rect 12348 8449 12357 8483
rect 12357 8449 12391 8483
rect 12391 8449 12400 8483
rect 12348 8440 12400 8449
rect 13268 8483 13320 8492
rect 13268 8449 13277 8483
rect 13277 8449 13311 8483
rect 13311 8449 13320 8483
rect 13268 8440 13320 8449
rect 9220 8304 9272 8356
rect 10048 8372 10100 8424
rect 10232 8415 10284 8424
rect 10232 8381 10241 8415
rect 10241 8381 10275 8415
rect 10275 8381 10284 8415
rect 10232 8372 10284 8381
rect 10600 8372 10652 8424
rect 11244 8372 11296 8424
rect 12072 8304 12124 8356
rect 3056 8236 3108 8288
rect 7656 8236 7708 8288
rect 8944 8279 8996 8288
rect 8944 8245 8953 8279
rect 8953 8245 8987 8279
rect 8987 8245 8996 8279
rect 8944 8236 8996 8245
rect 9680 8236 9732 8288
rect 4214 8134 4266 8186
rect 4278 8134 4330 8186
rect 4342 8134 4394 8186
rect 4406 8134 4458 8186
rect 4470 8134 4522 8186
rect 12214 8134 12266 8186
rect 12278 8134 12330 8186
rect 12342 8134 12394 8186
rect 12406 8134 12458 8186
rect 12470 8134 12522 8186
rect 1492 8075 1544 8084
rect 1492 8041 1501 8075
rect 1501 8041 1535 8075
rect 1535 8041 1544 8075
rect 1492 8032 1544 8041
rect 1768 7871 1820 7880
rect 1768 7837 1777 7871
rect 1777 7837 1811 7871
rect 1811 7837 1820 7871
rect 1768 7828 1820 7837
rect 3792 7896 3844 7948
rect 4068 7896 4120 7948
rect 4620 7896 4672 7948
rect 3056 7871 3108 7880
rect 3056 7837 3065 7871
rect 3065 7837 3099 7871
rect 3099 7837 3108 7871
rect 3056 7828 3108 7837
rect 3976 7871 4028 7880
rect 3976 7837 3985 7871
rect 3985 7837 4019 7871
rect 4019 7837 4028 7871
rect 3976 7828 4028 7837
rect 5264 8032 5316 8084
rect 7840 8075 7892 8084
rect 7840 8041 7849 8075
rect 7849 8041 7883 8075
rect 7883 8041 7892 8075
rect 7840 8032 7892 8041
rect 12900 8032 12952 8084
rect 13544 8032 13596 8084
rect 5448 7964 5500 8016
rect 10232 8007 10284 8016
rect 6092 7896 6144 7948
rect 4988 7828 5040 7880
rect 10232 7973 10241 8007
rect 10241 7973 10275 8007
rect 10275 7973 10284 8007
rect 10232 7964 10284 7973
rect 7196 7896 7248 7948
rect 7748 7896 7800 7948
rect 8024 7896 8076 7948
rect 9680 7896 9732 7948
rect 6828 7828 6880 7880
rect 7656 7871 7708 7880
rect 7656 7837 7665 7871
rect 7665 7837 7699 7871
rect 7699 7837 7708 7871
rect 8116 7871 8168 7880
rect 7656 7828 7708 7837
rect 8116 7837 8125 7871
rect 8125 7837 8159 7871
rect 8159 7837 8168 7871
rect 8116 7828 8168 7837
rect 9036 7828 9088 7880
rect 9496 7871 9548 7880
rect 9496 7837 9505 7871
rect 9505 7837 9539 7871
rect 9539 7837 9548 7871
rect 9496 7828 9548 7837
rect 9956 7828 10008 7880
rect 10692 7871 10744 7880
rect 10692 7837 10701 7871
rect 10701 7837 10735 7871
rect 10735 7837 10744 7871
rect 10692 7828 10744 7837
rect 10876 7871 10928 7880
rect 10876 7837 10885 7871
rect 10885 7837 10919 7871
rect 10919 7837 10928 7871
rect 10876 7828 10928 7837
rect 11060 7828 11112 7880
rect 13268 7871 13320 7880
rect 13268 7837 13277 7871
rect 13277 7837 13311 7871
rect 13311 7837 13320 7871
rect 13268 7828 13320 7837
rect 1676 7760 1728 7812
rect 3516 7803 3568 7812
rect 2872 7692 2924 7744
rect 3056 7692 3108 7744
rect 3516 7769 3525 7803
rect 3525 7769 3559 7803
rect 3559 7769 3568 7803
rect 3516 7760 3568 7769
rect 3700 7692 3752 7744
rect 5448 7760 5500 7812
rect 6276 7692 6328 7744
rect 7380 7735 7432 7744
rect 7380 7701 7389 7735
rect 7389 7701 7423 7735
rect 7423 7701 7432 7735
rect 7380 7692 7432 7701
rect 10140 7735 10192 7744
rect 10140 7701 10149 7735
rect 10149 7701 10183 7735
rect 10183 7701 10192 7735
rect 10140 7692 10192 7701
rect 11980 7760 12032 7812
rect 12256 7692 12308 7744
rect 8214 7590 8266 7642
rect 8278 7590 8330 7642
rect 8342 7590 8394 7642
rect 8406 7590 8458 7642
rect 8470 7590 8522 7642
rect 3424 7488 3476 7540
rect 3700 7488 3752 7540
rect 3056 7420 3108 7472
rect 1676 7395 1728 7404
rect 1676 7361 1685 7395
rect 1685 7361 1719 7395
rect 1719 7361 1728 7395
rect 1676 7352 1728 7361
rect 1768 7395 1820 7404
rect 1768 7361 1777 7395
rect 1777 7361 1811 7395
rect 1811 7361 1820 7395
rect 1768 7352 1820 7361
rect 4160 7352 4212 7404
rect 6828 7488 6880 7540
rect 7472 7531 7524 7540
rect 7472 7497 7481 7531
rect 7481 7497 7515 7531
rect 7515 7497 7524 7531
rect 7472 7488 7524 7497
rect 8116 7488 8168 7540
rect 5448 7395 5500 7404
rect 2596 7327 2648 7336
rect 2596 7293 2605 7327
rect 2605 7293 2639 7327
rect 2639 7293 2648 7327
rect 2596 7284 2648 7293
rect 2780 7327 2832 7336
rect 2780 7293 2789 7327
rect 2789 7293 2823 7327
rect 2823 7293 2832 7327
rect 3056 7327 3108 7336
rect 2780 7284 2832 7293
rect 3056 7293 3065 7327
rect 3065 7293 3099 7327
rect 3099 7293 3108 7327
rect 3056 7284 3108 7293
rect 3516 7284 3568 7336
rect 5448 7361 5457 7395
rect 5457 7361 5491 7395
rect 5491 7361 5500 7395
rect 5448 7352 5500 7361
rect 5540 7352 5592 7404
rect 6736 7420 6788 7472
rect 6920 7463 6972 7472
rect 5724 7352 5776 7404
rect 6276 7352 6328 7404
rect 6920 7429 6929 7463
rect 6929 7429 6963 7463
rect 6963 7429 6972 7463
rect 6920 7420 6972 7429
rect 7564 7420 7616 7472
rect 6092 7284 6144 7336
rect 7196 7352 7248 7404
rect 7012 7284 7064 7336
rect 1768 7216 1820 7268
rect 1492 7191 1544 7200
rect 1492 7157 1501 7191
rect 1501 7157 1535 7191
rect 1535 7157 1544 7191
rect 1492 7148 1544 7157
rect 1952 7191 2004 7200
rect 1952 7157 1961 7191
rect 1961 7157 1995 7191
rect 1995 7157 2004 7191
rect 1952 7148 2004 7157
rect 5724 7216 5776 7268
rect 8392 7284 8444 7336
rect 8300 7216 8352 7268
rect 8944 7352 8996 7404
rect 10692 7488 10744 7540
rect 12256 7488 12308 7540
rect 12072 7420 12124 7472
rect 10232 7395 10284 7404
rect 8852 7327 8904 7336
rect 8852 7293 8861 7327
rect 8861 7293 8895 7327
rect 8895 7293 8904 7327
rect 8852 7284 8904 7293
rect 4620 7148 4672 7200
rect 5264 7191 5316 7200
rect 5264 7157 5273 7191
rect 5273 7157 5307 7191
rect 5307 7157 5316 7191
rect 5264 7148 5316 7157
rect 8024 7148 8076 7200
rect 10232 7361 10241 7395
rect 10241 7361 10275 7395
rect 10275 7361 10284 7395
rect 10232 7352 10284 7361
rect 11060 7352 11112 7404
rect 12256 7395 12308 7404
rect 12256 7361 12265 7395
rect 12265 7361 12299 7395
rect 12299 7361 12308 7395
rect 12256 7352 12308 7361
rect 10508 7284 10560 7336
rect 12072 7284 12124 7336
rect 4214 7046 4266 7098
rect 4278 7046 4330 7098
rect 4342 7046 4394 7098
rect 4406 7046 4458 7098
rect 4470 7046 4522 7098
rect 12214 7046 12266 7098
rect 12278 7046 12330 7098
rect 12342 7046 12394 7098
rect 12406 7046 12458 7098
rect 12470 7046 12522 7098
rect 1952 6944 2004 6996
rect 3516 6944 3568 6996
rect 3976 6944 4028 6996
rect 4160 6944 4212 6996
rect 5632 6944 5684 6996
rect 7380 6944 7432 6996
rect 2780 6808 2832 6860
rect 3976 6808 4028 6860
rect 5632 6851 5684 6860
rect 5632 6817 5641 6851
rect 5641 6817 5675 6851
rect 5675 6817 5684 6851
rect 5632 6808 5684 6817
rect 7840 6876 7892 6928
rect 6460 6808 6512 6860
rect 6920 6808 6972 6860
rect 7656 6808 7708 6860
rect 8576 6808 8628 6860
rect 9680 6876 9732 6928
rect 13268 6919 13320 6928
rect 13268 6885 13277 6919
rect 13277 6885 13311 6919
rect 13311 6885 13320 6919
rect 13268 6876 13320 6885
rect 2872 6740 2924 6792
rect 3332 6740 3384 6792
rect 3792 6740 3844 6792
rect 4160 6783 4212 6792
rect 4160 6749 4169 6783
rect 4169 6749 4203 6783
rect 4203 6749 4212 6783
rect 4160 6740 4212 6749
rect 5264 6783 5316 6792
rect 5264 6749 5273 6783
rect 5273 6749 5307 6783
rect 5307 6749 5316 6783
rect 5264 6740 5316 6749
rect 7196 6740 7248 6792
rect 8024 6740 8076 6792
rect 6552 6672 6604 6724
rect 7748 6672 7800 6724
rect 8300 6740 8352 6792
rect 8392 6783 8444 6792
rect 8392 6749 8401 6783
rect 8401 6749 8435 6783
rect 8435 6749 8444 6783
rect 8392 6740 8444 6749
rect 8852 6740 8904 6792
rect 11612 6808 11664 6860
rect 10048 6783 10100 6792
rect 8668 6715 8720 6724
rect 1492 6604 1544 6656
rect 2504 6604 2556 6656
rect 4068 6647 4120 6656
rect 4068 6613 4077 6647
rect 4077 6613 4111 6647
rect 4111 6613 4120 6647
rect 4068 6604 4120 6613
rect 8668 6681 8677 6715
rect 8677 6681 8711 6715
rect 8711 6681 8720 6715
rect 8668 6672 8720 6681
rect 8760 6672 8812 6724
rect 9312 6604 9364 6656
rect 10048 6749 10057 6783
rect 10057 6749 10091 6783
rect 10091 6749 10100 6783
rect 10048 6740 10100 6749
rect 11704 6740 11756 6792
rect 12348 6740 12400 6792
rect 13452 6783 13504 6792
rect 13452 6749 13461 6783
rect 13461 6749 13495 6783
rect 13495 6749 13504 6783
rect 13452 6740 13504 6749
rect 11888 6672 11940 6724
rect 8214 6502 8266 6554
rect 8278 6502 8330 6554
rect 8342 6502 8394 6554
rect 8406 6502 8458 6554
rect 8470 6502 8522 6554
rect 2044 6400 2096 6452
rect 3056 6400 3108 6452
rect 1768 6307 1820 6316
rect 1768 6273 1777 6307
rect 1777 6273 1811 6307
rect 1811 6273 1820 6307
rect 1768 6264 1820 6273
rect 1952 6307 2004 6316
rect 1952 6273 1977 6307
rect 1977 6273 2004 6307
rect 1952 6264 2004 6273
rect 2504 6307 2556 6316
rect 2504 6273 2513 6307
rect 2513 6273 2547 6307
rect 2547 6273 2556 6307
rect 2504 6264 2556 6273
rect 2688 6307 2740 6316
rect 2688 6273 2697 6307
rect 2697 6273 2731 6307
rect 2731 6273 2740 6307
rect 2688 6264 2740 6273
rect 5540 6400 5592 6452
rect 6092 6443 6144 6452
rect 6092 6409 6101 6443
rect 6101 6409 6135 6443
rect 6135 6409 6144 6443
rect 6092 6400 6144 6409
rect 6552 6443 6604 6452
rect 6552 6409 6561 6443
rect 6561 6409 6595 6443
rect 6595 6409 6604 6443
rect 6552 6400 6604 6409
rect 10416 6400 10468 6452
rect 10876 6400 10928 6452
rect 3976 6332 4028 6384
rect 6920 6375 6972 6384
rect 6920 6341 6929 6375
rect 6929 6341 6963 6375
rect 6963 6341 6972 6375
rect 6920 6332 6972 6341
rect 7472 6332 7524 6384
rect 1400 6103 1452 6112
rect 1400 6069 1409 6103
rect 1409 6069 1443 6103
rect 1443 6069 1452 6103
rect 1400 6060 1452 6069
rect 5724 6264 5776 6316
rect 6460 6264 6512 6316
rect 7932 6307 7984 6316
rect 2228 6128 2280 6180
rect 3148 6171 3200 6180
rect 3148 6137 3157 6171
rect 3157 6137 3191 6171
rect 3191 6137 3200 6171
rect 3148 6128 3200 6137
rect 2320 6060 2372 6112
rect 4068 6239 4120 6248
rect 4068 6205 4077 6239
rect 4077 6205 4111 6239
rect 4111 6205 4120 6239
rect 4068 6196 4120 6205
rect 5356 6196 5408 6248
rect 7932 6273 7941 6307
rect 7941 6273 7975 6307
rect 7975 6273 7984 6307
rect 7932 6264 7984 6273
rect 8668 6307 8720 6316
rect 8668 6273 8677 6307
rect 8677 6273 8711 6307
rect 8711 6273 8720 6307
rect 8668 6264 8720 6273
rect 9680 6332 9732 6384
rect 12072 6400 12124 6452
rect 10692 6307 10744 6316
rect 6736 6196 6788 6248
rect 7748 6239 7800 6248
rect 7748 6205 7757 6239
rect 7757 6205 7791 6239
rect 7791 6205 7800 6239
rect 7748 6196 7800 6205
rect 10692 6273 10701 6307
rect 10701 6273 10735 6307
rect 10735 6273 10744 6307
rect 10692 6264 10744 6273
rect 10784 6307 10836 6316
rect 10784 6273 10793 6307
rect 10793 6273 10827 6307
rect 10827 6273 10836 6307
rect 11888 6332 11940 6384
rect 13268 6332 13320 6384
rect 10784 6264 10836 6273
rect 12072 6307 12124 6316
rect 10508 6196 10560 6248
rect 11152 6196 11204 6248
rect 12072 6273 12081 6307
rect 12081 6273 12115 6307
rect 12115 6273 12124 6307
rect 12072 6264 12124 6273
rect 12348 6264 12400 6316
rect 13268 6239 13320 6248
rect 11612 6171 11664 6180
rect 11612 6137 11621 6171
rect 11621 6137 11655 6171
rect 11655 6137 11664 6171
rect 11612 6128 11664 6137
rect 4620 6060 4672 6112
rect 9772 6103 9824 6112
rect 9772 6069 9781 6103
rect 9781 6069 9815 6103
rect 9815 6069 9824 6103
rect 9772 6060 9824 6069
rect 12072 6060 12124 6112
rect 13268 6205 13277 6239
rect 13277 6205 13311 6239
rect 13311 6205 13320 6239
rect 13268 6196 13320 6205
rect 4214 5958 4266 6010
rect 4278 5958 4330 6010
rect 4342 5958 4394 6010
rect 4406 5958 4458 6010
rect 4470 5958 4522 6010
rect 12214 5958 12266 6010
rect 12278 5958 12330 6010
rect 12342 5958 12394 6010
rect 12406 5958 12458 6010
rect 12470 5958 12522 6010
rect 1584 5856 1636 5908
rect 2688 5856 2740 5908
rect 5356 5899 5408 5908
rect 2320 5831 2372 5840
rect 2320 5797 2329 5831
rect 2329 5797 2363 5831
rect 2363 5797 2372 5831
rect 2320 5788 2372 5797
rect 5356 5865 5365 5899
rect 5365 5865 5399 5899
rect 5399 5865 5408 5899
rect 5356 5856 5408 5865
rect 4068 5788 4120 5840
rect 5724 5856 5776 5908
rect 8116 5856 8168 5908
rect 10324 5856 10376 5908
rect 10692 5856 10744 5908
rect 13268 5899 13320 5908
rect 13268 5865 13277 5899
rect 13277 5865 13311 5899
rect 13311 5865 13320 5899
rect 13268 5856 13320 5865
rect 1400 5720 1452 5772
rect 2780 5720 2832 5772
rect 3148 5720 3200 5772
rect 1492 5695 1544 5704
rect 1492 5661 1501 5695
rect 1501 5661 1535 5695
rect 1535 5661 1544 5695
rect 1492 5652 1544 5661
rect 1584 5695 1636 5704
rect 1584 5661 1593 5695
rect 1593 5661 1627 5695
rect 1627 5661 1636 5695
rect 1584 5652 1636 5661
rect 2044 5652 2096 5704
rect 4620 5720 4672 5772
rect 8760 5788 8812 5840
rect 6000 5763 6052 5772
rect 6000 5729 6009 5763
rect 6009 5729 6043 5763
rect 6043 5729 6052 5763
rect 6000 5720 6052 5729
rect 7748 5720 7800 5772
rect 4712 5695 4764 5704
rect 2872 5584 2924 5636
rect 3608 5584 3660 5636
rect 3976 5627 4028 5636
rect 3976 5593 3985 5627
rect 3985 5593 4019 5627
rect 4019 5593 4028 5627
rect 3976 5584 4028 5593
rect 2228 5516 2280 5568
rect 3332 5516 3384 5568
rect 3424 5516 3476 5568
rect 4068 5559 4120 5568
rect 4068 5525 4077 5559
rect 4077 5525 4111 5559
rect 4111 5525 4120 5559
rect 4068 5516 4120 5525
rect 4712 5661 4721 5695
rect 4721 5661 4755 5695
rect 4755 5661 4764 5695
rect 4712 5652 4764 5661
rect 4436 5584 4488 5636
rect 5908 5652 5960 5704
rect 6184 5695 6236 5704
rect 6184 5661 6193 5695
rect 6193 5661 6227 5695
rect 6227 5661 6236 5695
rect 6184 5652 6236 5661
rect 8576 5695 8628 5704
rect 6092 5584 6144 5636
rect 8576 5661 8585 5695
rect 8585 5661 8619 5695
rect 8619 5661 8628 5695
rect 8576 5652 8628 5661
rect 10048 5720 10100 5772
rect 10600 5763 10652 5772
rect 10600 5729 10609 5763
rect 10609 5729 10643 5763
rect 10643 5729 10652 5763
rect 10600 5720 10652 5729
rect 9312 5695 9364 5704
rect 9312 5661 9321 5695
rect 9321 5661 9355 5695
rect 9355 5661 9364 5695
rect 9312 5652 9364 5661
rect 9680 5695 9732 5704
rect 9680 5661 9719 5695
rect 9719 5661 9732 5695
rect 9680 5652 9732 5661
rect 9864 5652 9916 5704
rect 10232 5695 10284 5704
rect 10232 5661 10241 5695
rect 10241 5661 10275 5695
rect 10275 5661 10284 5695
rect 10232 5652 10284 5661
rect 11980 5652 12032 5704
rect 5540 5516 5592 5568
rect 9404 5584 9456 5636
rect 11612 5584 11664 5636
rect 11888 5584 11940 5636
rect 8576 5516 8628 5568
rect 9680 5516 9732 5568
rect 10140 5516 10192 5568
rect 11428 5516 11480 5568
rect 12164 5516 12216 5568
rect 13176 5559 13228 5568
rect 13176 5525 13185 5559
rect 13185 5525 13219 5559
rect 13219 5525 13228 5559
rect 13176 5516 13228 5525
rect 8214 5414 8266 5466
rect 8278 5414 8330 5466
rect 8342 5414 8394 5466
rect 8406 5414 8458 5466
rect 8470 5414 8522 5466
rect 2780 5312 2832 5364
rect 4068 5312 4120 5364
rect 1952 5244 2004 5296
rect 1492 5219 1544 5228
rect 1492 5185 1501 5219
rect 1501 5185 1535 5219
rect 1535 5185 1544 5219
rect 1492 5176 1544 5185
rect 1584 5176 1636 5228
rect 2136 5219 2188 5228
rect 2136 5185 2145 5219
rect 2145 5185 2179 5219
rect 2179 5185 2188 5219
rect 2136 5176 2188 5185
rect 2320 5219 2372 5228
rect 2320 5185 2329 5219
rect 2329 5185 2363 5219
rect 2363 5185 2372 5219
rect 2320 5176 2372 5185
rect 3240 5176 3292 5228
rect 3608 5287 3660 5296
rect 3608 5253 3617 5287
rect 3617 5253 3651 5287
rect 3651 5253 3660 5287
rect 4436 5287 4488 5296
rect 3608 5244 3660 5253
rect 4436 5253 4445 5287
rect 4445 5253 4479 5287
rect 4479 5253 4488 5287
rect 4436 5244 4488 5253
rect 4620 5287 4672 5296
rect 4620 5253 4629 5287
rect 4629 5253 4663 5287
rect 4663 5253 4672 5287
rect 4620 5244 4672 5253
rect 8576 5312 8628 5364
rect 11796 5312 11848 5364
rect 5448 5244 5500 5296
rect 4068 5219 4120 5228
rect 4068 5185 4077 5219
rect 4077 5185 4111 5219
rect 4111 5185 4120 5219
rect 4068 5176 4120 5185
rect 5356 5219 5408 5228
rect 5356 5185 5365 5219
rect 5365 5185 5399 5219
rect 5399 5185 5408 5219
rect 5356 5176 5408 5185
rect 5908 5244 5960 5296
rect 6000 5219 6052 5228
rect 6000 5185 6009 5219
rect 6009 5185 6043 5219
rect 6043 5185 6052 5219
rect 6000 5176 6052 5185
rect 1768 4972 1820 5024
rect 2320 5015 2372 5024
rect 2320 4981 2329 5015
rect 2329 4981 2363 5015
rect 2363 4981 2372 5015
rect 2320 4972 2372 4981
rect 3240 5040 3292 5092
rect 8116 5176 8168 5228
rect 9036 5176 9088 5228
rect 7748 5108 7800 5160
rect 7104 5040 7156 5092
rect 3424 4972 3476 5024
rect 3792 5015 3844 5024
rect 3792 4981 3801 5015
rect 3801 4981 3835 5015
rect 3835 4981 3844 5015
rect 3792 4972 3844 4981
rect 5908 4972 5960 5024
rect 7656 4972 7708 5024
rect 8668 5108 8720 5160
rect 10048 5244 10100 5296
rect 11152 5244 11204 5296
rect 11612 5176 11664 5228
rect 12072 5244 12124 5296
rect 13176 5244 13228 5296
rect 12624 5219 12676 5228
rect 12624 5185 12633 5219
rect 12633 5185 12667 5219
rect 12667 5185 12676 5219
rect 12624 5176 12676 5185
rect 13544 5219 13596 5228
rect 13544 5185 13553 5219
rect 13553 5185 13587 5219
rect 13587 5185 13596 5219
rect 13544 5176 13596 5185
rect 9772 5151 9824 5160
rect 9772 5117 9781 5151
rect 9781 5117 9815 5151
rect 9815 5117 9824 5151
rect 9772 5108 9824 5117
rect 9864 4972 9916 5024
rect 10416 4972 10468 5024
rect 12716 4972 12768 5024
rect 4214 4870 4266 4922
rect 4278 4870 4330 4922
rect 4342 4870 4394 4922
rect 4406 4870 4458 4922
rect 4470 4870 4522 4922
rect 12214 4870 12266 4922
rect 12278 4870 12330 4922
rect 12342 4870 12394 4922
rect 12406 4870 12458 4922
rect 12470 4870 12522 4922
rect 1400 4811 1452 4820
rect 1400 4777 1409 4811
rect 1409 4777 1443 4811
rect 1443 4777 1452 4811
rect 1400 4768 1452 4777
rect 2780 4768 2832 4820
rect 3240 4768 3292 4820
rect 5632 4768 5684 4820
rect 6644 4768 6696 4820
rect 2320 4675 2372 4684
rect 2320 4641 2329 4675
rect 2329 4641 2363 4675
rect 2363 4641 2372 4675
rect 2320 4632 2372 4641
rect 3424 4675 3476 4684
rect 3424 4641 3433 4675
rect 3433 4641 3467 4675
rect 3467 4641 3476 4675
rect 3424 4632 3476 4641
rect 5632 4675 5684 4684
rect 5632 4641 5641 4675
rect 5641 4641 5675 4675
rect 5675 4641 5684 4675
rect 5632 4632 5684 4641
rect 1584 4607 1636 4616
rect 1584 4573 1593 4607
rect 1593 4573 1627 4607
rect 1627 4573 1636 4607
rect 1584 4564 1636 4573
rect 1676 4564 1728 4616
rect 2136 4607 2188 4616
rect 2136 4573 2145 4607
rect 2145 4573 2179 4607
rect 2179 4573 2188 4607
rect 2136 4564 2188 4573
rect 2412 4607 2464 4616
rect 2412 4573 2421 4607
rect 2421 4573 2455 4607
rect 2455 4573 2464 4607
rect 2412 4564 2464 4573
rect 3332 4607 3384 4616
rect 2688 4539 2740 4548
rect 2688 4505 2697 4539
rect 2697 4505 2731 4539
rect 2731 4505 2740 4539
rect 2688 4496 2740 4505
rect 2780 4496 2832 4548
rect 3332 4573 3341 4607
rect 3341 4573 3375 4607
rect 3375 4573 3384 4607
rect 3332 4564 3384 4573
rect 3792 4564 3844 4616
rect 4252 4564 4304 4616
rect 5724 4607 5776 4616
rect 5724 4573 5733 4607
rect 5733 4573 5767 4607
rect 5767 4573 5776 4607
rect 5724 4564 5776 4573
rect 5908 4607 5960 4616
rect 5908 4573 5917 4607
rect 5917 4573 5951 4607
rect 5951 4573 5960 4607
rect 5908 4564 5960 4573
rect 6184 4700 6236 4752
rect 6092 4607 6144 4616
rect 6828 4632 6880 4684
rect 8576 4768 8628 4820
rect 7656 4632 7708 4684
rect 7748 4632 7800 4684
rect 9404 4768 9456 4820
rect 10232 4768 10284 4820
rect 9680 4700 9732 4752
rect 13176 4743 13228 4752
rect 6092 4573 6135 4607
rect 6135 4573 6144 4607
rect 6092 4564 6144 4573
rect 6736 4607 6788 4616
rect 6736 4573 6745 4607
rect 6745 4573 6779 4607
rect 6779 4573 6788 4607
rect 6736 4564 6788 4573
rect 9128 4607 9180 4616
rect 9128 4573 9137 4607
rect 9137 4573 9171 4607
rect 9171 4573 9180 4607
rect 10048 4632 10100 4684
rect 13176 4709 13185 4743
rect 13185 4709 13219 4743
rect 13219 4709 13228 4743
rect 13176 4700 13228 4709
rect 9128 4564 9180 4573
rect 12532 4564 12584 4616
rect 13544 4607 13596 4616
rect 13544 4573 13553 4607
rect 13553 4573 13587 4607
rect 13587 4573 13596 4607
rect 13544 4564 13596 4573
rect 2320 4428 2372 4480
rect 3240 4471 3292 4480
rect 3240 4437 3249 4471
rect 3249 4437 3283 4471
rect 3283 4437 3292 4471
rect 3240 4428 3292 4437
rect 3516 4471 3568 4480
rect 3516 4437 3525 4471
rect 3525 4437 3559 4471
rect 3559 4437 3568 4471
rect 3516 4428 3568 4437
rect 4528 4428 4580 4480
rect 7196 4496 7248 4548
rect 5540 4428 5592 4480
rect 11888 4496 11940 4548
rect 9680 4471 9732 4480
rect 9680 4437 9689 4471
rect 9689 4437 9723 4471
rect 9723 4437 9732 4471
rect 9680 4428 9732 4437
rect 8214 4326 8266 4378
rect 8278 4326 8330 4378
rect 8342 4326 8394 4378
rect 8406 4326 8458 4378
rect 8470 4326 8522 4378
rect 2412 4224 2464 4276
rect 2780 4156 2832 4208
rect 1860 4131 1912 4140
rect 1860 4097 1869 4131
rect 1869 4097 1903 4131
rect 1903 4097 1912 4131
rect 1860 4088 1912 4097
rect 2044 4131 2096 4140
rect 2044 4097 2053 4131
rect 2053 4097 2087 4131
rect 2087 4097 2096 4131
rect 2044 4088 2096 4097
rect 2228 4131 2280 4140
rect 2228 4097 2237 4131
rect 2237 4097 2271 4131
rect 2271 4097 2280 4131
rect 2228 4088 2280 4097
rect 2320 4131 2372 4140
rect 2320 4097 2329 4131
rect 2329 4097 2363 4131
rect 2363 4097 2372 4131
rect 2688 4131 2740 4140
rect 2320 4088 2372 4097
rect 2688 4097 2697 4131
rect 2697 4097 2731 4131
rect 2731 4097 2740 4131
rect 2688 4088 2740 4097
rect 2872 4131 2924 4140
rect 2872 4097 2881 4131
rect 2881 4097 2915 4131
rect 2915 4097 2924 4131
rect 2872 4088 2924 4097
rect 3700 4156 3752 4208
rect 4712 4224 4764 4276
rect 5356 4224 5408 4276
rect 5540 4267 5592 4276
rect 5540 4233 5549 4267
rect 5549 4233 5583 4267
rect 5583 4233 5592 4267
rect 5540 4224 5592 4233
rect 6092 4224 6144 4276
rect 6644 4224 6696 4276
rect 3516 4131 3568 4140
rect 3516 4097 3525 4131
rect 3525 4097 3559 4131
rect 3559 4097 3568 4131
rect 3516 4088 3568 4097
rect 5724 4156 5776 4208
rect 4252 4131 4304 4140
rect 1768 4063 1820 4072
rect 1768 4029 1777 4063
rect 1777 4029 1811 4063
rect 1811 4029 1820 4063
rect 1768 4020 1820 4029
rect 2228 3884 2280 3936
rect 3148 3884 3200 3936
rect 3424 3952 3476 4004
rect 4252 4097 4261 4131
rect 4261 4097 4295 4131
rect 4295 4097 4304 4131
rect 4252 4088 4304 4097
rect 4528 4131 4580 4140
rect 4528 4097 4537 4131
rect 4537 4097 4571 4131
rect 4571 4097 4580 4131
rect 4528 4088 4580 4097
rect 5448 4088 5500 4140
rect 4896 4063 4948 4072
rect 4896 4029 4905 4063
rect 4905 4029 4939 4063
rect 4939 4029 4948 4063
rect 4896 4020 4948 4029
rect 4804 3952 4856 4004
rect 4988 3952 5040 4004
rect 6644 4088 6696 4140
rect 8576 4224 8628 4276
rect 9680 4267 9732 4276
rect 9680 4233 9689 4267
rect 9689 4233 9723 4267
rect 9723 4233 9732 4267
rect 9680 4224 9732 4233
rect 9864 4224 9916 4276
rect 11152 4267 11204 4276
rect 8484 4088 8536 4140
rect 9404 4156 9456 4208
rect 11152 4233 11161 4267
rect 11161 4233 11195 4267
rect 11195 4233 11204 4267
rect 11152 4224 11204 4233
rect 11612 4267 11664 4276
rect 11612 4233 11621 4267
rect 11621 4233 11655 4267
rect 11655 4233 11664 4267
rect 11612 4224 11664 4233
rect 7196 4020 7248 4072
rect 9588 4131 9640 4140
rect 9588 4097 9597 4131
rect 9597 4097 9631 4131
rect 9631 4097 9640 4131
rect 9588 4088 9640 4097
rect 10324 4088 10376 4140
rect 10784 4131 10836 4140
rect 10784 4097 10793 4131
rect 10793 4097 10827 4131
rect 10827 4097 10836 4131
rect 10784 4088 10836 4097
rect 11980 4156 12032 4208
rect 12532 4199 12584 4208
rect 12072 4131 12124 4140
rect 6828 3952 6880 4004
rect 9220 3952 9272 4004
rect 9956 3952 10008 4004
rect 12072 4097 12081 4131
rect 12081 4097 12115 4131
rect 12115 4097 12124 4131
rect 12072 4088 12124 4097
rect 12532 4165 12541 4199
rect 12541 4165 12575 4199
rect 12575 4165 12584 4199
rect 12532 4156 12584 4165
rect 12716 4131 12768 4140
rect 11704 4020 11756 4072
rect 12716 4097 12725 4131
rect 12725 4097 12759 4131
rect 12759 4097 12768 4131
rect 12716 4088 12768 4097
rect 13360 4088 13412 4140
rect 9036 3884 9088 3936
rect 10324 3884 10376 3936
rect 13360 3927 13412 3936
rect 13360 3893 13369 3927
rect 13369 3893 13403 3927
rect 13403 3893 13412 3927
rect 13360 3884 13412 3893
rect 4214 3782 4266 3834
rect 4278 3782 4330 3834
rect 4342 3782 4394 3834
rect 4406 3782 4458 3834
rect 4470 3782 4522 3834
rect 12214 3782 12266 3834
rect 12278 3782 12330 3834
rect 12342 3782 12394 3834
rect 12406 3782 12458 3834
rect 12470 3782 12522 3834
rect 1676 3680 1728 3732
rect 2136 3612 2188 3664
rect 6736 3680 6788 3732
rect 9588 3723 9640 3732
rect 2044 3544 2096 3596
rect 2780 3544 2832 3596
rect 3516 3544 3568 3596
rect 4068 3544 4120 3596
rect 1492 3519 1544 3528
rect 1492 3485 1501 3519
rect 1501 3485 1535 3519
rect 1535 3485 1544 3519
rect 1492 3476 1544 3485
rect 1584 3519 1636 3528
rect 1584 3485 1593 3519
rect 1593 3485 1627 3519
rect 1627 3485 1636 3519
rect 1584 3476 1636 3485
rect 2320 3476 2372 3528
rect 3332 3519 3384 3528
rect 3332 3485 3341 3519
rect 3341 3485 3375 3519
rect 3375 3485 3384 3519
rect 3332 3476 3384 3485
rect 4344 3519 4396 3528
rect 4344 3485 4353 3519
rect 4353 3485 4387 3519
rect 4387 3485 4396 3519
rect 4344 3476 4396 3485
rect 4436 3519 4488 3528
rect 4436 3485 4445 3519
rect 4445 3485 4479 3519
rect 4479 3485 4488 3519
rect 4436 3476 4488 3485
rect 4712 3519 4764 3528
rect 4712 3485 4721 3519
rect 4721 3485 4755 3519
rect 4755 3485 4764 3519
rect 4712 3476 4764 3485
rect 5356 3519 5408 3528
rect 2688 3408 2740 3460
rect 5356 3485 5365 3519
rect 5365 3485 5399 3519
rect 5399 3485 5408 3519
rect 5356 3476 5408 3485
rect 5724 3519 5776 3528
rect 5724 3485 5733 3519
rect 5733 3485 5767 3519
rect 5767 3485 5776 3519
rect 5724 3476 5776 3485
rect 6460 3544 6512 3596
rect 6828 3544 6880 3596
rect 8484 3544 8536 3596
rect 8852 3544 8904 3596
rect 9588 3689 9597 3723
rect 9597 3689 9631 3723
rect 9631 3689 9640 3723
rect 9588 3680 9640 3689
rect 9680 3680 9732 3732
rect 10784 3680 10836 3732
rect 9128 3544 9180 3596
rect 10324 3587 10376 3596
rect 10324 3553 10333 3587
rect 10333 3553 10367 3587
rect 10367 3553 10376 3587
rect 10324 3544 10376 3553
rect 11980 3544 12032 3596
rect 9220 3519 9272 3528
rect 5448 3408 5500 3460
rect 1860 3340 1912 3392
rect 3240 3340 3292 3392
rect 6920 3340 6972 3392
rect 8208 3408 8260 3460
rect 9220 3485 9229 3519
rect 9229 3485 9263 3519
rect 9263 3485 9272 3519
rect 9220 3476 9272 3485
rect 9496 3476 9548 3528
rect 12072 3519 12124 3528
rect 12072 3485 12081 3519
rect 12081 3485 12115 3519
rect 12115 3485 12124 3519
rect 12072 3476 12124 3485
rect 9864 3408 9916 3460
rect 10600 3408 10652 3460
rect 11704 3408 11756 3460
rect 11888 3408 11940 3460
rect 12808 3451 12860 3460
rect 12808 3417 12817 3451
rect 12817 3417 12851 3451
rect 12851 3417 12860 3451
rect 12808 3408 12860 3417
rect 9588 3340 9640 3392
rect 8214 3238 8266 3290
rect 8278 3238 8330 3290
rect 8342 3238 8394 3290
rect 8406 3238 8458 3290
rect 8470 3238 8522 3290
rect 1492 3136 1544 3188
rect 2320 3179 2372 3188
rect 2320 3145 2329 3179
rect 2329 3145 2363 3179
rect 2363 3145 2372 3179
rect 2320 3136 2372 3145
rect 3332 3111 3384 3120
rect 3332 3077 3341 3111
rect 3341 3077 3375 3111
rect 3375 3077 3384 3111
rect 3332 3068 3384 3077
rect 1492 2932 1544 2984
rect 2136 2975 2188 2984
rect 2136 2941 2145 2975
rect 2145 2941 2179 2975
rect 2179 2941 2188 2975
rect 2136 2932 2188 2941
rect 2872 3043 2924 3052
rect 2872 3009 2881 3043
rect 2881 3009 2915 3043
rect 2915 3009 2924 3043
rect 2872 3000 2924 3009
rect 3240 3000 3292 3052
rect 4712 3136 4764 3188
rect 5448 3136 5500 3188
rect 6920 3136 6972 3188
rect 8116 3136 8168 3188
rect 10600 3136 10652 3188
rect 11060 3136 11112 3188
rect 11336 3179 11388 3188
rect 11336 3145 11345 3179
rect 11345 3145 11379 3179
rect 11379 3145 11388 3179
rect 11336 3136 11388 3145
rect 4436 3000 4488 3052
rect 4712 3043 4764 3052
rect 4712 3009 4721 3043
rect 4721 3009 4755 3043
rect 4755 3009 4764 3043
rect 4712 3000 4764 3009
rect 5356 3043 5408 3052
rect 5356 3009 5365 3043
rect 5365 3009 5399 3043
rect 5399 3009 5408 3043
rect 5356 3000 5408 3009
rect 5448 3000 5500 3052
rect 2688 2975 2740 2984
rect 2688 2941 2697 2975
rect 2697 2941 2731 2975
rect 2731 2941 2740 2975
rect 2688 2932 2740 2941
rect 2320 2864 2372 2916
rect 4344 2932 4396 2984
rect 4620 2975 4672 2984
rect 4620 2941 4629 2975
rect 4629 2941 4663 2975
rect 4663 2941 4672 2975
rect 4620 2932 4672 2941
rect 6552 3043 6604 3052
rect 6552 3009 6561 3043
rect 6561 3009 6595 3043
rect 6595 3009 6604 3043
rect 6552 3000 6604 3009
rect 7104 3000 7156 3052
rect 8576 3068 8628 3120
rect 9864 3068 9916 3120
rect 11980 3136 12032 3188
rect 12072 3068 12124 3120
rect 6276 2932 6328 2984
rect 6920 2975 6972 2984
rect 6920 2941 6929 2975
rect 6929 2941 6963 2975
rect 6963 2941 6972 2975
rect 6920 2932 6972 2941
rect 6552 2864 6604 2916
rect 7840 2864 7892 2916
rect 6184 2796 6236 2848
rect 8944 2932 8996 2984
rect 9772 2932 9824 2984
rect 10048 2975 10100 2984
rect 10048 2941 10057 2975
rect 10057 2941 10091 2975
rect 10091 2941 10100 2975
rect 10048 2932 10100 2941
rect 13176 3000 13228 3052
rect 13268 2932 13320 2984
rect 8024 2796 8076 2848
rect 12624 2864 12676 2916
rect 10600 2796 10652 2848
rect 4214 2694 4266 2746
rect 4278 2694 4330 2746
rect 4342 2694 4394 2746
rect 4406 2694 4458 2746
rect 4470 2694 4522 2746
rect 12214 2694 12266 2746
rect 12278 2694 12330 2746
rect 12342 2694 12394 2746
rect 12406 2694 12458 2746
rect 12470 2694 12522 2746
rect 2872 2592 2924 2644
rect 4712 2592 4764 2644
rect 8944 2635 8996 2644
rect 8944 2601 8953 2635
rect 8953 2601 8987 2635
rect 8987 2601 8996 2635
rect 8944 2592 8996 2601
rect 11060 2592 11112 2644
rect 3424 2524 3476 2576
rect 3792 2524 3844 2576
rect 9864 2567 9916 2576
rect 1768 2456 1820 2508
rect 3608 2456 3660 2508
rect 1676 2431 1728 2440
rect 1676 2397 1685 2431
rect 1685 2397 1719 2431
rect 1719 2397 1728 2431
rect 2136 2431 2188 2440
rect 1676 2388 1728 2397
rect 2136 2397 2145 2431
rect 2145 2397 2179 2431
rect 2179 2397 2188 2431
rect 2136 2388 2188 2397
rect 2320 2431 2372 2440
rect 2320 2397 2329 2431
rect 2329 2397 2363 2431
rect 2363 2397 2372 2431
rect 2320 2388 2372 2397
rect 1860 2363 1912 2372
rect 1860 2329 1869 2363
rect 1869 2329 1903 2363
rect 1903 2329 1912 2363
rect 1860 2320 1912 2329
rect 2872 2388 2924 2440
rect 3148 2252 3200 2304
rect 3700 2320 3752 2372
rect 3332 2252 3384 2304
rect 4620 2456 4672 2508
rect 9864 2533 9873 2567
rect 9873 2533 9907 2567
rect 9907 2533 9916 2567
rect 9864 2524 9916 2533
rect 8576 2456 8628 2508
rect 9588 2499 9640 2508
rect 5356 2388 5408 2440
rect 5448 2431 5500 2440
rect 5448 2397 5457 2431
rect 5457 2397 5491 2431
rect 5491 2397 5500 2431
rect 7564 2431 7616 2440
rect 5448 2388 5500 2397
rect 7564 2397 7573 2431
rect 7573 2397 7607 2431
rect 7607 2397 7616 2431
rect 7564 2388 7616 2397
rect 5908 2363 5960 2372
rect 5908 2329 5917 2363
rect 5917 2329 5951 2363
rect 5951 2329 5960 2363
rect 5908 2320 5960 2329
rect 6368 2320 6420 2372
rect 7196 2320 7248 2372
rect 7840 2388 7892 2440
rect 9588 2465 9597 2499
rect 9597 2465 9631 2499
rect 9631 2465 9640 2499
rect 9588 2456 9640 2465
rect 9772 2388 9824 2440
rect 9956 2431 10008 2440
rect 9956 2397 9965 2431
rect 9965 2397 9999 2431
rect 9999 2397 10008 2431
rect 9956 2388 10008 2397
rect 9128 2320 9180 2372
rect 9680 2320 9732 2372
rect 5632 2252 5684 2304
rect 6276 2252 6328 2304
rect 7288 2252 7340 2304
rect 8116 2252 8168 2304
rect 8668 2295 8720 2304
rect 8668 2261 8677 2295
rect 8677 2261 8711 2295
rect 8711 2261 8720 2295
rect 8668 2252 8720 2261
rect 9496 2252 9548 2304
rect 13176 2388 13228 2440
rect 13268 2431 13320 2440
rect 13268 2397 13277 2431
rect 13277 2397 13311 2431
rect 13311 2397 13320 2431
rect 13268 2388 13320 2397
rect 10600 2363 10652 2372
rect 10600 2329 10609 2363
rect 10609 2329 10643 2363
rect 10643 2329 10652 2363
rect 10600 2320 10652 2329
rect 11888 2320 11940 2372
rect 11520 2252 11572 2304
rect 8214 2150 8266 2202
rect 8278 2150 8330 2202
rect 8342 2150 8394 2202
rect 8406 2150 8458 2202
rect 8470 2150 8522 2202
rect 1584 2091 1636 2100
rect 1584 2057 1593 2091
rect 1593 2057 1627 2091
rect 1627 2057 1636 2091
rect 1584 2048 1636 2057
rect 2872 2048 2924 2100
rect 3424 2048 3476 2100
rect 5356 2048 5408 2100
rect 6368 2048 6420 2100
rect 6460 2091 6512 2100
rect 6460 2057 6469 2091
rect 6469 2057 6503 2091
rect 6503 2057 6512 2091
rect 6460 2048 6512 2057
rect 8668 2048 8720 2100
rect 9680 2048 9732 2100
rect 13176 2048 13228 2100
rect 1860 1980 1912 2032
rect 3148 1980 3200 2032
rect 4620 1980 4672 2032
rect 3516 1955 3568 1964
rect 3516 1921 3525 1955
rect 3525 1921 3559 1955
rect 3559 1921 3568 1955
rect 3792 1955 3844 1964
rect 3516 1912 3568 1921
rect 3792 1921 3801 1955
rect 3801 1921 3835 1955
rect 3835 1921 3844 1955
rect 3792 1912 3844 1921
rect 7932 1980 7984 2032
rect 8116 1980 8168 2032
rect 6736 1912 6788 1964
rect 10140 1912 10192 1964
rect 12072 1980 12124 2032
rect 12532 1980 12584 2032
rect 4068 1887 4120 1896
rect 4068 1853 4077 1887
rect 4077 1853 4111 1887
rect 4111 1853 4120 1887
rect 4068 1844 4120 1853
rect 8576 1887 8628 1896
rect 8576 1853 8585 1887
rect 8585 1853 8619 1887
rect 8619 1853 8628 1887
rect 8576 1844 8628 1853
rect 8944 1844 8996 1896
rect 9496 1844 9548 1896
rect 11336 1912 11388 1964
rect 11520 1887 11572 1896
rect 11060 1819 11112 1828
rect 11060 1785 11069 1819
rect 11069 1785 11103 1819
rect 11103 1785 11112 1819
rect 11060 1776 11112 1785
rect 6552 1708 6604 1760
rect 7012 1708 7064 1760
rect 11520 1853 11529 1887
rect 11529 1853 11563 1887
rect 11563 1853 11572 1887
rect 11520 1844 11572 1853
rect 13268 1844 13320 1896
rect 4214 1606 4266 1658
rect 4278 1606 4330 1658
rect 4342 1606 4394 1658
rect 4406 1606 4458 1658
rect 4470 1606 4522 1658
rect 12214 1606 12266 1658
rect 12278 1606 12330 1658
rect 12342 1606 12394 1658
rect 12406 1606 12458 1658
rect 12470 1606 12522 1658
rect 1676 1504 1728 1556
rect 4436 1504 4488 1556
rect 6736 1504 6788 1556
rect 8668 1547 8720 1556
rect 3424 1436 3476 1488
rect 4252 1436 4304 1488
rect 1400 1411 1452 1420
rect 1400 1377 1409 1411
rect 1409 1377 1443 1411
rect 1443 1377 1452 1411
rect 1400 1368 1452 1377
rect 3516 1300 3568 1352
rect 3700 1368 3752 1420
rect 3884 1343 3936 1352
rect 3884 1309 3893 1343
rect 3893 1309 3927 1343
rect 3927 1309 3936 1343
rect 3884 1300 3936 1309
rect 4252 1343 4304 1352
rect 3240 1275 3292 1284
rect 3240 1241 3249 1275
rect 3249 1241 3283 1275
rect 3283 1241 3292 1275
rect 3240 1232 3292 1241
rect 3332 1232 3384 1284
rect 3700 1164 3752 1216
rect 4252 1309 4261 1343
rect 4261 1309 4295 1343
rect 4295 1309 4304 1343
rect 4252 1300 4304 1309
rect 4436 1343 4488 1352
rect 4436 1309 4445 1343
rect 4445 1309 4479 1343
rect 4479 1309 4488 1343
rect 4436 1300 4488 1309
rect 4620 1343 4672 1352
rect 4620 1309 4629 1343
rect 4629 1309 4663 1343
rect 4663 1309 4672 1343
rect 4620 1300 4672 1309
rect 4896 1368 4948 1420
rect 5908 1411 5960 1420
rect 4528 1232 4580 1284
rect 5356 1300 5408 1352
rect 5632 1300 5684 1352
rect 5908 1377 5917 1411
rect 5917 1377 5951 1411
rect 5951 1377 5960 1411
rect 5908 1368 5960 1377
rect 6736 1368 6788 1420
rect 7288 1411 7340 1420
rect 7012 1343 7064 1352
rect 7012 1309 7021 1343
rect 7021 1309 7055 1343
rect 7055 1309 7064 1343
rect 7012 1300 7064 1309
rect 7288 1377 7297 1411
rect 7297 1377 7331 1411
rect 7331 1377 7340 1411
rect 7288 1368 7340 1377
rect 7564 1368 7616 1420
rect 7932 1411 7984 1420
rect 7932 1377 7941 1411
rect 7941 1377 7975 1411
rect 7975 1377 7984 1411
rect 7932 1368 7984 1377
rect 8668 1513 8677 1547
rect 8677 1513 8711 1547
rect 8711 1513 8720 1547
rect 8668 1504 8720 1513
rect 13268 1547 13320 1556
rect 13268 1513 13277 1547
rect 13277 1513 13311 1547
rect 13311 1513 13320 1547
rect 13268 1504 13320 1513
rect 8944 1479 8996 1488
rect 8944 1445 8953 1479
rect 8953 1445 8987 1479
rect 8987 1445 8996 1479
rect 8944 1436 8996 1445
rect 11152 1436 11204 1488
rect 8576 1368 8628 1420
rect 11520 1411 11572 1420
rect 11520 1377 11529 1411
rect 11529 1377 11563 1411
rect 11563 1377 11572 1411
rect 11520 1368 11572 1377
rect 9128 1343 9180 1352
rect 9128 1309 9137 1343
rect 9137 1309 9171 1343
rect 9171 1309 9180 1343
rect 9128 1300 9180 1309
rect 7104 1232 7156 1284
rect 9496 1232 9548 1284
rect 11060 1232 11112 1284
rect 5448 1164 5500 1216
rect 6368 1207 6420 1216
rect 6368 1173 6377 1207
rect 6377 1173 6411 1207
rect 6411 1173 6420 1207
rect 6368 1164 6420 1173
rect 12808 1232 12860 1284
rect 8214 1062 8266 1114
rect 8278 1062 8330 1114
rect 8342 1062 8394 1114
rect 8406 1062 8458 1114
rect 8470 1062 8522 1114
rect 3884 960 3936 1012
rect 6368 960 6420 1012
<< metal2 >>
rect 570 14362 626 15000
rect 1398 14512 1454 14521
rect 1398 14447 1454 14456
rect 570 14334 888 14362
rect 570 14200 626 14334
rect 860 13394 888 14334
rect 1412 13530 1440 14447
rect 1674 14200 1730 15000
rect 2870 14362 2926 15000
rect 2870 14334 3188 14362
rect 2870 14200 2926 14334
rect 1584 13728 1636 13734
rect 1584 13670 1636 13676
rect 1400 13524 1452 13530
rect 1400 13466 1452 13472
rect 848 13388 900 13394
rect 848 13330 900 13336
rect 1596 13326 1624 13670
rect 1688 13462 1716 14200
rect 2320 13796 2372 13802
rect 2320 13738 2372 13744
rect 1676 13456 1728 13462
rect 1676 13398 1728 13404
rect 2332 13394 2360 13738
rect 2778 13560 2834 13569
rect 2778 13495 2834 13504
rect 2320 13388 2372 13394
rect 2320 13330 2372 13336
rect 1584 13320 1636 13326
rect 1584 13262 1636 13268
rect 2228 13320 2280 13326
rect 2228 13262 2280 13268
rect 2688 13320 2740 13326
rect 2688 13262 2740 13268
rect 1492 12912 1544 12918
rect 1492 12854 1544 12860
rect 1400 12844 1452 12850
rect 1400 12786 1452 12792
rect 1412 12646 1440 12786
rect 1400 12640 1452 12646
rect 1504 12617 1532 12854
rect 1400 12582 1452 12588
rect 1490 12608 1546 12617
rect 1412 11830 1440 12582
rect 1490 12543 1546 12552
rect 1596 12238 1624 13262
rect 2044 13252 2096 13258
rect 2044 13194 2096 13200
rect 2136 13252 2188 13258
rect 2136 13194 2188 13200
rect 1860 12844 1912 12850
rect 1860 12786 1912 12792
rect 1584 12232 1636 12238
rect 1584 12174 1636 12180
rect 1872 12102 1900 12786
rect 2056 12238 2084 13194
rect 2148 12442 2176 13194
rect 2240 12850 2268 13262
rect 2228 12844 2280 12850
rect 2228 12786 2280 12792
rect 2136 12436 2188 12442
rect 2136 12378 2188 12384
rect 2700 12345 2728 13262
rect 2686 12336 2742 12345
rect 2686 12271 2742 12280
rect 2700 12238 2728 12271
rect 2044 12232 2096 12238
rect 2044 12174 2096 12180
rect 2688 12232 2740 12238
rect 2688 12174 2740 12180
rect 1860 12096 1912 12102
rect 1860 12038 1912 12044
rect 2056 11898 2084 12174
rect 2412 12164 2464 12170
rect 2412 12106 2464 12112
rect 2044 11892 2096 11898
rect 2044 11834 2096 11840
rect 1400 11824 1452 11830
rect 1400 11766 1452 11772
rect 2228 11688 2280 11694
rect 1766 11656 1822 11665
rect 2228 11630 2280 11636
rect 1766 11591 1822 11600
rect 1582 10704 1638 10713
rect 1582 10639 1584 10648
rect 1636 10639 1638 10648
rect 1584 10610 1636 10616
rect 1400 10532 1452 10538
rect 1400 10474 1452 10480
rect 1412 10266 1440 10474
rect 1492 10464 1544 10470
rect 1492 10406 1544 10412
rect 1400 10260 1452 10266
rect 1400 10202 1452 10208
rect 1504 10130 1532 10406
rect 1492 10124 1544 10130
rect 1492 10066 1544 10072
rect 1504 9586 1532 10066
rect 1492 9580 1544 9586
rect 1492 9522 1544 9528
rect 1596 9178 1624 10610
rect 1780 9654 1808 11591
rect 2240 11150 2268 11630
rect 2424 11150 2452 12106
rect 2504 11756 2556 11762
rect 2504 11698 2556 11704
rect 2688 11756 2740 11762
rect 2688 11698 2740 11704
rect 2516 11665 2544 11698
rect 2502 11656 2558 11665
rect 2502 11591 2558 11600
rect 2228 11144 2280 11150
rect 2228 11086 2280 11092
rect 2412 11144 2464 11150
rect 2412 11086 2464 11092
rect 2424 10810 2452 11086
rect 2700 11014 2728 11698
rect 2688 11008 2740 11014
rect 2688 10950 2740 10956
rect 2412 10804 2464 10810
rect 2412 10746 2464 10752
rect 2700 10742 2728 10950
rect 2792 10810 2820 13495
rect 2872 13252 2924 13258
rect 2872 13194 2924 13200
rect 2884 12714 2912 13194
rect 3160 12986 3188 14334
rect 3974 14200 4030 15000
rect 5170 14200 5226 15000
rect 6274 14362 6330 15000
rect 6274 14334 6408 14362
rect 6274 14200 6330 14334
rect 3884 13320 3936 13326
rect 3884 13262 3936 13268
rect 3424 13252 3476 13258
rect 3424 13194 3476 13200
rect 3148 12980 3200 12986
rect 3148 12922 3200 12928
rect 3240 12912 3292 12918
rect 3240 12854 3292 12860
rect 2872 12708 2924 12714
rect 2872 12650 2924 12656
rect 2872 12164 2924 12170
rect 2872 12106 2924 12112
rect 2884 11626 2912 12106
rect 3148 11824 3200 11830
rect 3148 11766 3200 11772
rect 2872 11620 2924 11626
rect 2872 11562 2924 11568
rect 2884 11286 2912 11562
rect 3160 11558 3188 11766
rect 3148 11552 3200 11558
rect 3148 11494 3200 11500
rect 2872 11280 2924 11286
rect 2872 11222 2924 11228
rect 2780 10804 2832 10810
rect 2832 10764 2912 10792
rect 2780 10746 2832 10752
rect 2688 10736 2740 10742
rect 2688 10678 2740 10684
rect 2780 10668 2832 10674
rect 2780 10610 2832 10616
rect 2688 10600 2740 10606
rect 2688 10542 2740 10548
rect 2136 10464 2188 10470
rect 2136 10406 2188 10412
rect 2148 9926 2176 10406
rect 2700 10198 2728 10542
rect 2688 10192 2740 10198
rect 2410 10160 2466 10169
rect 2688 10134 2740 10140
rect 2410 10095 2466 10104
rect 2424 10062 2452 10095
rect 2412 10056 2464 10062
rect 2412 9998 2464 10004
rect 2136 9920 2188 9926
rect 2136 9862 2188 9868
rect 2148 9761 2176 9862
rect 2134 9752 2190 9761
rect 2134 9687 2190 9696
rect 2424 9674 2452 9998
rect 2792 9994 2820 10610
rect 2884 10266 2912 10764
rect 3160 10470 3188 11494
rect 3148 10464 3200 10470
rect 3148 10406 3200 10412
rect 2872 10260 2924 10266
rect 2872 10202 2924 10208
rect 2872 10056 2924 10062
rect 2872 9998 2924 10004
rect 2780 9988 2832 9994
rect 2780 9930 2832 9936
rect 1768 9648 1820 9654
rect 2424 9646 2636 9674
rect 1768 9590 1820 9596
rect 1584 9172 1636 9178
rect 1584 9114 1636 9120
rect 2608 8974 2636 9646
rect 2792 9450 2820 9930
rect 2780 9444 2832 9450
rect 2780 9386 2832 9392
rect 2884 8974 2912 9998
rect 2964 9988 3016 9994
rect 2964 9930 3016 9936
rect 2976 9178 3004 9930
rect 3160 9926 3188 10406
rect 3148 9920 3200 9926
rect 3148 9862 3200 9868
rect 3252 9738 3280 12854
rect 3436 12238 3464 13194
rect 3700 12912 3752 12918
rect 3700 12854 3752 12860
rect 3424 12232 3476 12238
rect 3424 12174 3476 12180
rect 3712 11626 3740 12854
rect 3896 12850 3924 13262
rect 3884 12844 3936 12850
rect 3884 12786 3936 12792
rect 3792 12708 3844 12714
rect 3792 12650 3844 12656
rect 3804 11830 3832 12650
rect 3896 12442 3924 12786
rect 3988 12730 4016 14200
rect 5080 13728 5132 13734
rect 5080 13670 5132 13676
rect 4214 13628 4522 13637
rect 4214 13626 4220 13628
rect 4276 13626 4300 13628
rect 4356 13626 4380 13628
rect 4436 13626 4460 13628
rect 4516 13626 4522 13628
rect 4276 13574 4278 13626
rect 4458 13574 4460 13626
rect 4214 13572 4220 13574
rect 4276 13572 4300 13574
rect 4356 13572 4380 13574
rect 4436 13572 4460 13574
rect 4516 13572 4522 13574
rect 4214 13563 4522 13572
rect 4068 13524 4120 13530
rect 4068 13466 4120 13472
rect 4080 12850 4108 13466
rect 5092 13394 5120 13670
rect 5080 13388 5132 13394
rect 5080 13330 5132 13336
rect 4252 13184 4304 13190
rect 4252 13126 4304 13132
rect 4264 12918 4292 13126
rect 4252 12912 4304 12918
rect 4252 12854 4304 12860
rect 4068 12844 4120 12850
rect 4068 12786 4120 12792
rect 4436 12844 4488 12850
rect 4436 12786 4488 12792
rect 3988 12702 4108 12730
rect 3884 12436 3936 12442
rect 3884 12378 3936 12384
rect 4080 12238 4108 12702
rect 4448 12646 4476 12786
rect 4436 12640 4488 12646
rect 4436 12582 4488 12588
rect 4214 12540 4522 12549
rect 4214 12538 4220 12540
rect 4276 12538 4300 12540
rect 4356 12538 4380 12540
rect 4436 12538 4460 12540
rect 4516 12538 4522 12540
rect 4276 12486 4278 12538
rect 4458 12486 4460 12538
rect 4214 12484 4220 12486
rect 4276 12484 4300 12486
rect 4356 12484 4380 12486
rect 4436 12484 4460 12486
rect 4516 12484 4522 12486
rect 4214 12475 4522 12484
rect 5092 12238 5120 13330
rect 4068 12232 4120 12238
rect 4068 12174 4120 12180
rect 4804 12232 4856 12238
rect 4804 12174 4856 12180
rect 5080 12232 5132 12238
rect 5080 12174 5132 12180
rect 4080 11898 4108 12174
rect 4068 11892 4120 11898
rect 4068 11834 4120 11840
rect 3792 11824 3844 11830
rect 3792 11766 3844 11772
rect 4712 11688 4764 11694
rect 4712 11630 4764 11636
rect 3700 11620 3752 11626
rect 3700 11562 3752 11568
rect 4620 11620 4672 11626
rect 4620 11562 4672 11568
rect 3884 11552 3936 11558
rect 3884 11494 3936 11500
rect 3516 11280 3568 11286
rect 3516 11222 3568 11228
rect 3332 11144 3384 11150
rect 3332 11086 3384 11092
rect 3344 10742 3372 11086
rect 3528 11082 3556 11222
rect 3896 11150 3924 11494
rect 4214 11452 4522 11461
rect 4214 11450 4220 11452
rect 4276 11450 4300 11452
rect 4356 11450 4380 11452
rect 4436 11450 4460 11452
rect 4516 11450 4522 11452
rect 4276 11398 4278 11450
rect 4458 11398 4460 11450
rect 4214 11396 4220 11398
rect 4276 11396 4300 11398
rect 4356 11396 4380 11398
rect 4436 11396 4460 11398
rect 4516 11396 4522 11398
rect 4214 11387 4522 11396
rect 4528 11212 4580 11218
rect 4528 11154 4580 11160
rect 3884 11144 3936 11150
rect 3884 11086 3936 11092
rect 3516 11076 3568 11082
rect 3516 11018 3568 11024
rect 3608 11076 3660 11082
rect 3608 11018 3660 11024
rect 3332 10736 3384 10742
rect 3332 10678 3384 10684
rect 3332 10260 3384 10266
rect 3332 10202 3384 10208
rect 3344 10062 3372 10202
rect 3332 10056 3384 10062
rect 3332 9998 3384 10004
rect 3252 9710 3372 9738
rect 3240 9580 3292 9586
rect 3240 9522 3292 9528
rect 2964 9172 3016 9178
rect 2964 9114 3016 9120
rect 3252 8974 3280 9522
rect 2596 8968 2648 8974
rect 2596 8910 2648 8916
rect 2872 8968 2924 8974
rect 2872 8910 2924 8916
rect 3240 8968 3292 8974
rect 3240 8910 3292 8916
rect 1768 8832 1820 8838
rect 2136 8832 2188 8838
rect 1768 8774 1820 8780
rect 2134 8800 2136 8809
rect 2188 8800 2190 8809
rect 1492 8492 1544 8498
rect 1492 8434 1544 8440
rect 1504 8090 1532 8434
rect 1492 8084 1544 8090
rect 1492 8026 1544 8032
rect 1780 7886 1808 8774
rect 2134 8735 2190 8744
rect 2964 8356 3016 8362
rect 2964 8298 3016 8304
rect 1768 7880 1820 7886
rect 1768 7822 1820 7828
rect 1676 7812 1728 7818
rect 1676 7754 1728 7760
rect 1688 7410 1716 7754
rect 2872 7744 2924 7750
rect 2872 7686 2924 7692
rect 1676 7404 1728 7410
rect 1676 7346 1728 7352
rect 1768 7404 1820 7410
rect 1768 7346 1820 7352
rect 1780 7274 1808 7346
rect 2596 7336 2648 7342
rect 2596 7278 2648 7284
rect 2780 7336 2832 7342
rect 2780 7278 2832 7284
rect 1768 7268 1820 7274
rect 1768 7210 1820 7216
rect 1492 7200 1544 7206
rect 1492 7142 1544 7148
rect 1504 6662 1532 7142
rect 1492 6656 1544 6662
rect 1492 6598 1544 6604
rect 1400 6112 1452 6118
rect 1398 6080 1400 6089
rect 1452 6080 1454 6089
rect 1398 6015 1454 6024
rect 1412 5778 1440 6015
rect 1400 5772 1452 5778
rect 1400 5714 1452 5720
rect 1504 5710 1532 6598
rect 1780 6322 1808 7210
rect 1952 7200 2004 7206
rect 1952 7142 2004 7148
rect 1964 7002 1992 7142
rect 1952 6996 2004 7002
rect 1952 6938 2004 6944
rect 2504 6656 2556 6662
rect 2504 6598 2556 6604
rect 2044 6452 2096 6458
rect 2044 6394 2096 6400
rect 1768 6316 1820 6322
rect 1768 6258 1820 6264
rect 1952 6316 2004 6322
rect 1952 6258 2004 6264
rect 1584 5908 1636 5914
rect 1584 5850 1636 5856
rect 1596 5710 1624 5850
rect 1492 5704 1544 5710
rect 1492 5646 1544 5652
rect 1584 5704 1636 5710
rect 1584 5646 1636 5652
rect 1504 5234 1532 5646
rect 1596 5234 1624 5646
rect 1964 5302 1992 6258
rect 2056 5710 2084 6394
rect 2516 6322 2544 6598
rect 2608 6361 2636 7278
rect 2792 6866 2820 7278
rect 2780 6860 2832 6866
rect 2780 6802 2832 6808
rect 2884 6798 2912 7686
rect 2872 6792 2924 6798
rect 2872 6734 2924 6740
rect 2594 6352 2650 6361
rect 2504 6316 2556 6322
rect 2594 6287 2650 6296
rect 2688 6316 2740 6322
rect 2504 6258 2556 6264
rect 2688 6258 2740 6264
rect 2228 6180 2280 6186
rect 2228 6122 2280 6128
rect 2044 5704 2096 5710
rect 2240 5658 2268 6122
rect 2320 6112 2372 6118
rect 2320 6054 2372 6060
rect 2332 5846 2360 6054
rect 2700 5914 2728 6258
rect 2688 5908 2740 5914
rect 2688 5850 2740 5856
rect 2320 5840 2372 5846
rect 2320 5782 2372 5788
rect 2780 5772 2832 5778
rect 2780 5714 2832 5720
rect 2044 5646 2096 5652
rect 2148 5630 2268 5658
rect 2148 5386 2176 5630
rect 2228 5568 2280 5574
rect 2228 5510 2280 5516
rect 2056 5358 2176 5386
rect 1952 5296 2004 5302
rect 1952 5238 2004 5244
rect 1492 5228 1544 5234
rect 1492 5170 1544 5176
rect 1584 5228 1636 5234
rect 1584 5170 1636 5176
rect 1398 5128 1454 5137
rect 1398 5063 1454 5072
rect 1412 4826 1440 5063
rect 1768 5024 1820 5030
rect 1768 4966 1820 4972
rect 1400 4820 1452 4826
rect 1400 4762 1452 4768
rect 1584 4616 1636 4622
rect 1584 4558 1636 4564
rect 1676 4616 1728 4622
rect 1676 4558 1728 4564
rect 1596 3534 1624 4558
rect 1688 3738 1716 4558
rect 1780 4078 1808 4966
rect 2056 4146 2084 5358
rect 2136 5228 2188 5234
rect 2136 5170 2188 5176
rect 2148 4622 2176 5170
rect 2136 4616 2188 4622
rect 2136 4558 2188 4564
rect 2240 4146 2268 5510
rect 2792 5370 2820 5714
rect 2872 5636 2924 5642
rect 2872 5578 2924 5584
rect 2780 5364 2832 5370
rect 2780 5306 2832 5312
rect 2320 5228 2372 5234
rect 2372 5188 2452 5216
rect 2320 5170 2372 5176
rect 2320 5024 2372 5030
rect 2320 4966 2372 4972
rect 2332 4690 2360 4966
rect 2320 4684 2372 4690
rect 2320 4626 2372 4632
rect 2424 4622 2452 5188
rect 2792 4826 2820 5306
rect 2780 4820 2832 4826
rect 2780 4762 2832 4768
rect 2412 4616 2464 4622
rect 2412 4558 2464 4564
rect 2320 4480 2372 4486
rect 2320 4422 2372 4428
rect 2332 4146 2360 4422
rect 2424 4282 2452 4558
rect 2688 4548 2740 4554
rect 2688 4490 2740 4496
rect 2780 4548 2832 4554
rect 2780 4490 2832 4496
rect 2412 4276 2464 4282
rect 2412 4218 2464 4224
rect 2700 4146 2728 4490
rect 2792 4214 2820 4490
rect 2780 4208 2832 4214
rect 2780 4150 2832 4156
rect 1860 4140 1912 4146
rect 1860 4082 1912 4088
rect 2044 4140 2096 4146
rect 2044 4082 2096 4088
rect 2228 4140 2280 4146
rect 2228 4082 2280 4088
rect 2320 4140 2372 4146
rect 2320 4082 2372 4088
rect 2688 4140 2740 4146
rect 2688 4082 2740 4088
rect 1768 4072 1820 4078
rect 1768 4014 1820 4020
rect 1676 3732 1728 3738
rect 1676 3674 1728 3680
rect 1492 3528 1544 3534
rect 1492 3470 1544 3476
rect 1584 3528 1636 3534
rect 1584 3470 1636 3476
rect 1504 3194 1532 3470
rect 1492 3188 1544 3194
rect 1492 3130 1544 3136
rect 1492 2984 1544 2990
rect 1492 2926 1544 2932
rect 1504 2774 1532 2926
rect 1596 2836 1624 3470
rect 1872 3398 1900 4082
rect 2056 3602 2084 4082
rect 2240 3942 2268 4082
rect 2228 3936 2280 3942
rect 2228 3878 2280 3884
rect 2136 3664 2188 3670
rect 2136 3606 2188 3612
rect 2044 3596 2096 3602
rect 2044 3538 2096 3544
rect 1860 3392 1912 3398
rect 1860 3334 1912 3340
rect 2148 3233 2176 3606
rect 2792 3602 2820 4150
rect 2884 4146 2912 5578
rect 2872 4140 2924 4146
rect 2872 4082 2924 4088
rect 2780 3596 2832 3602
rect 2780 3538 2832 3544
rect 2320 3528 2372 3534
rect 2320 3470 2372 3476
rect 2134 3224 2190 3233
rect 2332 3194 2360 3470
rect 2688 3460 2740 3466
rect 2688 3402 2740 3408
rect 2134 3159 2190 3168
rect 2320 3188 2372 3194
rect 2148 2990 2176 3159
rect 2320 3130 2372 3136
rect 2700 2990 2728 3402
rect 2872 3052 2924 3058
rect 2872 2994 2924 3000
rect 2136 2984 2188 2990
rect 2136 2926 2188 2932
rect 2688 2984 2740 2990
rect 2688 2926 2740 2932
rect 1596 2808 1808 2836
rect 1504 2746 1624 2774
rect 1596 2281 1624 2746
rect 1780 2514 1808 2808
rect 1768 2508 1820 2514
rect 1768 2450 1820 2456
rect 2148 2446 2176 2926
rect 2320 2916 2372 2922
rect 2320 2858 2372 2864
rect 2332 2446 2360 2858
rect 2884 2650 2912 2994
rect 2872 2644 2924 2650
rect 2872 2586 2924 2592
rect 1676 2440 1728 2446
rect 1676 2382 1728 2388
rect 2136 2440 2188 2446
rect 2136 2382 2188 2388
rect 2320 2440 2372 2446
rect 2320 2382 2372 2388
rect 2872 2440 2924 2446
rect 2872 2382 2924 2388
rect 1582 2272 1638 2281
rect 1582 2207 1638 2216
rect 1596 2106 1624 2207
rect 1584 2100 1636 2106
rect 1584 2042 1636 2048
rect 1688 1562 1716 2382
rect 1860 2372 1912 2378
rect 1860 2314 1912 2320
rect 1872 2038 1900 2314
rect 2884 2106 2912 2382
rect 2872 2100 2924 2106
rect 2872 2042 2924 2048
rect 1860 2032 1912 2038
rect 1860 1974 1912 1980
rect 1676 1556 1728 1562
rect 1676 1498 1728 1504
rect 1400 1420 1452 1426
rect 1400 1362 1452 1368
rect 1412 513 1440 1362
rect 2976 1329 3004 8298
rect 3056 8288 3108 8294
rect 3056 8230 3108 8236
rect 3068 7993 3096 8230
rect 3054 7984 3110 7993
rect 3054 7919 3110 7928
rect 3068 7886 3096 7919
rect 3056 7880 3108 7886
rect 3056 7822 3108 7828
rect 3056 7744 3108 7750
rect 3056 7686 3108 7692
rect 3068 7478 3096 7686
rect 3056 7472 3108 7478
rect 3056 7414 3108 7420
rect 3056 7336 3108 7342
rect 3056 7278 3108 7284
rect 3068 6458 3096 7278
rect 3344 6798 3372 9710
rect 3528 9110 3556 11018
rect 3620 10742 3648 11018
rect 3608 10736 3660 10742
rect 3608 10678 3660 10684
rect 3896 10674 3924 11086
rect 4540 10810 4568 11154
rect 4528 10804 4580 10810
rect 4528 10746 4580 10752
rect 4632 10742 4660 11562
rect 4724 10810 4752 11630
rect 4816 11558 4844 12174
rect 5080 11756 5132 11762
rect 5080 11698 5132 11704
rect 4988 11688 5040 11694
rect 4988 11630 5040 11636
rect 4804 11552 4856 11558
rect 4804 11494 4856 11500
rect 4816 11150 4844 11494
rect 4804 11144 4856 11150
rect 4804 11086 4856 11092
rect 4712 10804 4764 10810
rect 4712 10746 4764 10752
rect 4620 10736 4672 10742
rect 4620 10678 4672 10684
rect 5000 10674 5028 11630
rect 5092 11286 5120 11698
rect 5080 11280 5132 11286
rect 5080 11222 5132 11228
rect 5184 11218 5212 14200
rect 5724 13320 5776 13326
rect 5724 13262 5776 13268
rect 6092 13320 6144 13326
rect 6092 13262 6144 13268
rect 5540 13252 5592 13258
rect 5540 13194 5592 13200
rect 5552 12238 5580 13194
rect 5632 13184 5684 13190
rect 5632 13126 5684 13132
rect 5644 12306 5672 13126
rect 5736 12850 5764 13262
rect 6000 13252 6052 13258
rect 6000 13194 6052 13200
rect 5724 12844 5776 12850
rect 5724 12786 5776 12792
rect 6012 12714 6040 13194
rect 6000 12708 6052 12714
rect 6000 12650 6052 12656
rect 6012 12374 6040 12650
rect 6000 12368 6052 12374
rect 6000 12310 6052 12316
rect 5632 12300 5684 12306
rect 5632 12242 5684 12248
rect 6104 12238 6132 13262
rect 6184 13252 6236 13258
rect 6184 13194 6236 13200
rect 5540 12232 5592 12238
rect 5446 12200 5502 12209
rect 5540 12174 5592 12180
rect 5816 12232 5868 12238
rect 5816 12174 5868 12180
rect 6092 12232 6144 12238
rect 6092 12174 6144 12180
rect 5446 12135 5502 12144
rect 5460 12102 5488 12135
rect 5448 12096 5500 12102
rect 5448 12038 5500 12044
rect 5460 11830 5488 12038
rect 5448 11824 5500 11830
rect 5448 11766 5500 11772
rect 5632 11688 5684 11694
rect 5828 11642 5856 12174
rect 6196 11880 6224 13194
rect 6276 12232 6328 12238
rect 6276 12174 6328 12180
rect 5684 11636 5856 11642
rect 5632 11630 5856 11636
rect 5540 11620 5592 11626
rect 5644 11614 5856 11630
rect 5920 11852 6224 11880
rect 5540 11562 5592 11568
rect 5172 11212 5224 11218
rect 5172 11154 5224 11160
rect 3884 10668 3936 10674
rect 3884 10610 3936 10616
rect 4988 10668 5040 10674
rect 4988 10610 5040 10616
rect 5264 10668 5316 10674
rect 5264 10610 5316 10616
rect 5000 10577 5028 10610
rect 4986 10568 5042 10577
rect 4986 10503 5042 10512
rect 4620 10464 4672 10470
rect 4620 10406 4672 10412
rect 4214 10364 4522 10373
rect 4214 10362 4220 10364
rect 4276 10362 4300 10364
rect 4356 10362 4380 10364
rect 4436 10362 4460 10364
rect 4516 10362 4522 10364
rect 4276 10310 4278 10362
rect 4458 10310 4460 10362
rect 4214 10308 4220 10310
rect 4276 10308 4300 10310
rect 4356 10308 4380 10310
rect 4436 10308 4460 10310
rect 4516 10308 4522 10310
rect 4214 10299 4522 10308
rect 4632 10130 4660 10406
rect 4620 10124 4672 10130
rect 4620 10066 4672 10072
rect 3700 10056 3752 10062
rect 3700 9998 3752 10004
rect 3712 9586 3740 9998
rect 4528 9988 4580 9994
rect 4528 9930 4580 9936
rect 4988 9988 5040 9994
rect 4988 9930 5040 9936
rect 5172 9988 5224 9994
rect 5172 9930 5224 9936
rect 3976 9920 4028 9926
rect 3976 9862 4028 9868
rect 3700 9580 3752 9586
rect 3700 9522 3752 9528
rect 3516 9104 3568 9110
rect 3516 9046 3568 9052
rect 3988 8906 4016 9862
rect 4540 9654 4568 9930
rect 4528 9648 4580 9654
rect 4528 9590 4580 9596
rect 4540 9450 4568 9590
rect 4528 9444 4580 9450
rect 4528 9386 4580 9392
rect 4214 9276 4522 9285
rect 4214 9274 4220 9276
rect 4276 9274 4300 9276
rect 4356 9274 4380 9276
rect 4436 9274 4460 9276
rect 4516 9274 4522 9276
rect 4276 9222 4278 9274
rect 4458 9222 4460 9274
rect 4214 9220 4220 9222
rect 4276 9220 4300 9222
rect 4356 9220 4380 9222
rect 4436 9220 4460 9222
rect 4516 9220 4522 9222
rect 4214 9211 4522 9220
rect 4620 8968 4672 8974
rect 4620 8910 4672 8916
rect 3976 8900 4028 8906
rect 3976 8842 4028 8848
rect 4252 8900 4304 8906
rect 4252 8842 4304 8848
rect 3792 7948 3844 7954
rect 3792 7890 3844 7896
rect 3516 7812 3568 7818
rect 3516 7754 3568 7760
rect 3528 7562 3556 7754
rect 3700 7744 3752 7750
rect 3700 7686 3752 7692
rect 3436 7546 3556 7562
rect 3712 7546 3740 7686
rect 3424 7540 3556 7546
rect 3476 7534 3556 7540
rect 3424 7482 3476 7488
rect 3528 7342 3556 7534
rect 3700 7540 3752 7546
rect 3700 7482 3752 7488
rect 3804 7449 3832 7890
rect 3988 7886 4016 8842
rect 4264 8498 4292 8842
rect 4252 8492 4304 8498
rect 4252 8434 4304 8440
rect 4264 8378 4292 8434
rect 4080 8350 4292 8378
rect 4080 7954 4108 8350
rect 4214 8188 4522 8197
rect 4214 8186 4220 8188
rect 4276 8186 4300 8188
rect 4356 8186 4380 8188
rect 4436 8186 4460 8188
rect 4516 8186 4522 8188
rect 4276 8134 4278 8186
rect 4458 8134 4460 8186
rect 4214 8132 4220 8134
rect 4276 8132 4300 8134
rect 4356 8132 4380 8134
rect 4436 8132 4460 8134
rect 4516 8132 4522 8134
rect 4214 8123 4522 8132
rect 4632 7954 4660 8910
rect 5000 8566 5028 9930
rect 5184 9586 5212 9930
rect 5276 9654 5304 10610
rect 5356 10464 5408 10470
rect 5356 10406 5408 10412
rect 5368 10062 5396 10406
rect 5552 10062 5580 11562
rect 5920 11336 5948 11852
rect 6000 11756 6052 11762
rect 6000 11698 6052 11704
rect 6184 11756 6236 11762
rect 6184 11698 6236 11704
rect 5828 11308 5948 11336
rect 5828 10810 5856 11308
rect 5908 11076 5960 11082
rect 5908 11018 5960 11024
rect 5920 10810 5948 11018
rect 6012 11014 6040 11698
rect 6092 11280 6144 11286
rect 6090 11248 6092 11257
rect 6144 11248 6146 11257
rect 6090 11183 6146 11192
rect 6092 11076 6144 11082
rect 6196 11064 6224 11698
rect 6288 11082 6316 12174
rect 6144 11036 6224 11064
rect 6092 11018 6144 11024
rect 6000 11008 6052 11014
rect 6000 10950 6052 10956
rect 5816 10804 5868 10810
rect 5816 10746 5868 10752
rect 5908 10804 5960 10810
rect 5908 10746 5960 10752
rect 5828 10266 5856 10746
rect 5908 10600 5960 10606
rect 5908 10542 5960 10548
rect 5816 10260 5868 10266
rect 5816 10202 5868 10208
rect 5356 10056 5408 10062
rect 5356 9998 5408 10004
rect 5540 10056 5592 10062
rect 5540 9998 5592 10004
rect 5264 9648 5316 9654
rect 5264 9590 5316 9596
rect 5172 9580 5224 9586
rect 5172 9522 5224 9528
rect 5184 8906 5212 9522
rect 5276 8974 5304 9590
rect 5264 8968 5316 8974
rect 5264 8910 5316 8916
rect 5172 8900 5224 8906
rect 5172 8842 5224 8848
rect 5448 8832 5500 8838
rect 5448 8774 5500 8780
rect 5460 8566 5488 8774
rect 5552 8634 5580 9998
rect 5828 9489 5856 10202
rect 5920 9518 5948 10542
rect 6012 10470 6040 10950
rect 6196 10470 6224 11036
rect 6276 11076 6328 11082
rect 6276 11018 6328 11024
rect 6288 10810 6316 11018
rect 6276 10804 6328 10810
rect 6276 10746 6328 10752
rect 6288 10538 6316 10746
rect 6276 10532 6328 10538
rect 6276 10474 6328 10480
rect 6000 10464 6052 10470
rect 6000 10406 6052 10412
rect 6184 10464 6236 10470
rect 6184 10406 6236 10412
rect 6196 9926 6224 10406
rect 6380 10062 6408 14334
rect 7470 14200 7526 15000
rect 8574 14200 8630 15000
rect 9770 14200 9826 15000
rect 10874 14200 10930 15000
rect 12070 14200 12126 15000
rect 13174 14362 13230 15000
rect 13174 14334 13492 14362
rect 13174 14200 13230 14334
rect 6644 13932 6696 13938
rect 6644 13874 6696 13880
rect 6656 13326 6684 13874
rect 6920 13524 6972 13530
rect 6920 13466 6972 13472
rect 6644 13320 6696 13326
rect 6644 13262 6696 13268
rect 6644 12912 6696 12918
rect 6644 12854 6696 12860
rect 6460 12776 6512 12782
rect 6460 12718 6512 12724
rect 6472 12306 6500 12718
rect 6656 12374 6684 12854
rect 6932 12850 6960 13466
rect 7104 13388 7156 13394
rect 7104 13330 7156 13336
rect 7012 13320 7064 13326
rect 7012 13262 7064 13268
rect 7024 12918 7052 13262
rect 7116 13258 7144 13330
rect 7288 13320 7340 13326
rect 7288 13262 7340 13268
rect 7104 13252 7156 13258
rect 7104 13194 7156 13200
rect 7104 12980 7156 12986
rect 7104 12922 7156 12928
rect 7012 12912 7064 12918
rect 7012 12854 7064 12860
rect 6736 12844 6788 12850
rect 6736 12786 6788 12792
rect 6920 12844 6972 12850
rect 6920 12786 6972 12792
rect 6644 12368 6696 12374
rect 6644 12310 6696 12316
rect 6460 12300 6512 12306
rect 6460 12242 6512 12248
rect 6644 12164 6696 12170
rect 6644 12106 6696 12112
rect 6552 12096 6604 12102
rect 6552 12038 6604 12044
rect 6564 11898 6592 12038
rect 6552 11892 6604 11898
rect 6552 11834 6604 11840
rect 6460 11688 6512 11694
rect 6460 11630 6512 11636
rect 6472 11558 6500 11630
rect 6564 11626 6592 11834
rect 6552 11620 6604 11626
rect 6552 11562 6604 11568
rect 6460 11552 6512 11558
rect 6460 11494 6512 11500
rect 6472 10742 6500 11494
rect 6552 11144 6604 11150
rect 6550 11112 6552 11121
rect 6604 11112 6606 11121
rect 6550 11047 6606 11056
rect 6460 10736 6512 10742
rect 6460 10678 6512 10684
rect 6368 10056 6420 10062
rect 6368 9998 6420 10004
rect 6184 9920 6236 9926
rect 6184 9862 6236 9868
rect 6460 9716 6512 9722
rect 6460 9658 6512 9664
rect 5908 9512 5960 9518
rect 5814 9480 5870 9489
rect 5908 9454 5960 9460
rect 5814 9415 5870 9424
rect 5724 9104 5776 9110
rect 5724 9046 5776 9052
rect 5736 8838 5764 9046
rect 5920 8974 5948 9454
rect 6184 9376 6236 9382
rect 6184 9318 6236 9324
rect 5908 8968 5960 8974
rect 5908 8910 5960 8916
rect 5724 8832 5776 8838
rect 5724 8774 5776 8780
rect 5540 8628 5592 8634
rect 5540 8570 5592 8576
rect 4988 8560 5040 8566
rect 4988 8502 5040 8508
rect 5448 8560 5500 8566
rect 5448 8502 5500 8508
rect 4068 7948 4120 7954
rect 4068 7890 4120 7896
rect 4620 7948 4672 7954
rect 4620 7890 4672 7896
rect 5000 7886 5028 8502
rect 5264 8492 5316 8498
rect 5264 8434 5316 8440
rect 5276 8090 5304 8434
rect 5264 8084 5316 8090
rect 5264 8026 5316 8032
rect 5460 8022 5488 8502
rect 5448 8016 5500 8022
rect 5448 7958 5500 7964
rect 3976 7880 4028 7886
rect 3976 7822 4028 7828
rect 4988 7880 5040 7886
rect 4988 7822 5040 7828
rect 3790 7440 3846 7449
rect 3790 7375 3846 7384
rect 3516 7336 3568 7342
rect 3516 7278 3568 7284
rect 3528 7002 3556 7278
rect 3516 6996 3568 7002
rect 3516 6938 3568 6944
rect 3804 6798 3832 7375
rect 3882 7032 3938 7041
rect 3988 7002 4016 7822
rect 5448 7812 5500 7818
rect 5448 7754 5500 7760
rect 5460 7410 5488 7754
rect 5538 7440 5594 7449
rect 4160 7404 4212 7410
rect 4160 7346 4212 7352
rect 5448 7404 5500 7410
rect 5736 7410 5764 8774
rect 6196 8498 6224 9318
rect 6472 9042 6500 9658
rect 6564 9178 6592 11047
rect 6656 10062 6684 12106
rect 6748 11762 6776 12786
rect 6920 12368 6972 12374
rect 6920 12310 6972 12316
rect 6828 12232 6880 12238
rect 6828 12174 6880 12180
rect 6840 11898 6868 12174
rect 6828 11892 6880 11898
rect 6828 11834 6880 11840
rect 6736 11756 6788 11762
rect 6736 11698 6788 11704
rect 6736 11620 6788 11626
rect 6736 11562 6788 11568
rect 6748 11014 6776 11562
rect 6736 11008 6788 11014
rect 6736 10950 6788 10956
rect 6748 10674 6776 10950
rect 6736 10668 6788 10674
rect 6736 10610 6788 10616
rect 6644 10056 6696 10062
rect 6644 9998 6696 10004
rect 6748 9994 6776 10610
rect 6828 10600 6880 10606
rect 6828 10542 6880 10548
rect 6840 10062 6868 10542
rect 6828 10056 6880 10062
rect 6828 9998 6880 10004
rect 6736 9988 6788 9994
rect 6736 9930 6788 9936
rect 6642 9752 6698 9761
rect 6642 9687 6698 9696
rect 6656 9586 6684 9687
rect 6748 9586 6776 9930
rect 6644 9580 6696 9586
rect 6644 9522 6696 9528
rect 6736 9580 6788 9586
rect 6736 9522 6788 9528
rect 6826 9480 6882 9489
rect 6826 9415 6828 9424
rect 6880 9415 6882 9424
rect 6828 9386 6880 9392
rect 6644 9376 6696 9382
rect 6644 9318 6696 9324
rect 6552 9172 6604 9178
rect 6552 9114 6604 9120
rect 6460 9036 6512 9042
rect 6460 8978 6512 8984
rect 6552 8968 6604 8974
rect 6656 8956 6684 9318
rect 6604 8928 6684 8956
rect 6552 8910 6604 8916
rect 6828 8900 6880 8906
rect 6932 8888 6960 12310
rect 7024 12170 7052 12854
rect 7116 12238 7144 12922
rect 7300 12918 7328 13262
rect 7288 12912 7340 12918
rect 7288 12854 7340 12860
rect 7380 12844 7432 12850
rect 7380 12786 7432 12792
rect 7288 12776 7340 12782
rect 7288 12718 7340 12724
rect 7104 12232 7156 12238
rect 7104 12174 7156 12180
rect 7012 12164 7064 12170
rect 7012 12106 7064 12112
rect 7300 11830 7328 12718
rect 7288 11824 7340 11830
rect 7288 11766 7340 11772
rect 7300 11218 7328 11766
rect 7392 11762 7420 12786
rect 7380 11756 7432 11762
rect 7380 11698 7432 11704
rect 7380 11552 7432 11558
rect 7380 11494 7432 11500
rect 7288 11212 7340 11218
rect 7288 11154 7340 11160
rect 7012 11144 7064 11150
rect 7012 11086 7064 11092
rect 7024 10742 7052 11086
rect 7288 11076 7340 11082
rect 7288 11018 7340 11024
rect 7012 10736 7064 10742
rect 7012 10678 7064 10684
rect 7300 10606 7328 11018
rect 7392 10742 7420 11494
rect 7380 10736 7432 10742
rect 7380 10678 7432 10684
rect 7104 10600 7156 10606
rect 7024 10560 7104 10588
rect 7024 9722 7052 10560
rect 7104 10542 7156 10548
rect 7288 10600 7340 10606
rect 7288 10542 7340 10548
rect 7392 10538 7420 10678
rect 7380 10532 7432 10538
rect 7380 10474 7432 10480
rect 7194 10432 7250 10441
rect 7194 10367 7250 10376
rect 7208 10266 7236 10367
rect 7196 10260 7248 10266
rect 7196 10202 7248 10208
rect 7104 10056 7156 10062
rect 7104 9998 7156 10004
rect 7012 9716 7064 9722
rect 7012 9658 7064 9664
rect 7024 9042 7052 9658
rect 7116 9178 7144 9998
rect 7196 9920 7248 9926
rect 7196 9862 7248 9868
rect 7208 9625 7236 9862
rect 7484 9761 7512 14200
rect 8116 13728 8168 13734
rect 8116 13670 8168 13676
rect 8128 13462 8156 13670
rect 8116 13456 8168 13462
rect 8116 13398 8168 13404
rect 8208 13388 8260 13394
rect 8208 13330 8260 13336
rect 7748 13320 7800 13326
rect 7748 13262 7800 13268
rect 7656 13184 7708 13190
rect 7656 13126 7708 13132
rect 7668 12782 7696 13126
rect 7760 12850 7788 13262
rect 7840 13252 7892 13258
rect 7840 13194 7892 13200
rect 8116 13252 8168 13258
rect 8220 13240 8248 13330
rect 8484 13252 8536 13258
rect 8220 13212 8484 13240
rect 8116 13194 8168 13200
rect 8484 13194 8536 13200
rect 7852 12986 7880 13194
rect 7840 12980 7892 12986
rect 7840 12922 7892 12928
rect 7748 12844 7800 12850
rect 7748 12786 7800 12792
rect 7656 12776 7708 12782
rect 7656 12718 7708 12724
rect 7654 12472 7710 12481
rect 7760 12442 7788 12786
rect 7654 12407 7656 12416
rect 7708 12407 7710 12416
rect 7748 12436 7800 12442
rect 7656 12378 7708 12384
rect 7748 12378 7800 12384
rect 8128 12170 8156 13194
rect 8214 13084 8522 13093
rect 8214 13082 8220 13084
rect 8276 13082 8300 13084
rect 8356 13082 8380 13084
rect 8436 13082 8460 13084
rect 8516 13082 8522 13084
rect 8276 13030 8278 13082
rect 8458 13030 8460 13082
rect 8214 13028 8220 13030
rect 8276 13028 8300 13030
rect 8356 13028 8380 13030
rect 8436 13028 8460 13030
rect 8516 13028 8522 13030
rect 8214 13019 8522 13028
rect 8484 12912 8536 12918
rect 8482 12880 8484 12889
rect 8536 12880 8538 12889
rect 8482 12815 8538 12824
rect 8484 12708 8536 12714
rect 8484 12650 8536 12656
rect 8116 12164 8168 12170
rect 8116 12106 8168 12112
rect 8496 12102 8524 12650
rect 7748 12096 7800 12102
rect 7748 12038 7800 12044
rect 8484 12096 8536 12102
rect 8484 12038 8536 12044
rect 7760 11830 7788 12038
rect 8214 11996 8522 12005
rect 8214 11994 8220 11996
rect 8276 11994 8300 11996
rect 8356 11994 8380 11996
rect 8436 11994 8460 11996
rect 8516 11994 8522 11996
rect 8276 11942 8278 11994
rect 8458 11942 8460 11994
rect 8214 11940 8220 11942
rect 8276 11940 8300 11942
rect 8356 11940 8380 11942
rect 8436 11940 8460 11942
rect 8516 11940 8522 11942
rect 8214 11931 8522 11940
rect 7840 11892 7892 11898
rect 7840 11834 7892 11840
rect 8392 11892 8444 11898
rect 8392 11834 8444 11840
rect 7748 11824 7800 11830
rect 7748 11766 7800 11772
rect 7852 11762 7880 11834
rect 8404 11801 8432 11834
rect 8390 11792 8446 11801
rect 7656 11756 7708 11762
rect 7656 11698 7708 11704
rect 7840 11756 7892 11762
rect 7840 11698 7892 11704
rect 8208 11756 8260 11762
rect 8390 11727 8446 11736
rect 8208 11698 8260 11704
rect 7668 11529 7696 11698
rect 7748 11688 7800 11694
rect 7748 11630 7800 11636
rect 7654 11520 7710 11529
rect 7654 11455 7710 11464
rect 7654 11384 7710 11393
rect 7654 11319 7710 11328
rect 7564 11212 7616 11218
rect 7564 11154 7616 11160
rect 7576 11121 7604 11154
rect 7562 11112 7618 11121
rect 7562 11047 7564 11056
rect 7616 11047 7618 11056
rect 7564 11018 7616 11024
rect 7576 10987 7604 11018
rect 7668 10674 7696 11319
rect 7760 11286 7788 11630
rect 7852 11286 7880 11698
rect 8220 11626 8248 11698
rect 8208 11620 8260 11626
rect 8260 11580 8340 11608
rect 8208 11562 8260 11568
rect 8114 11520 8170 11529
rect 8114 11455 8170 11464
rect 7748 11280 7800 11286
rect 7748 11222 7800 11228
rect 7840 11280 7892 11286
rect 7840 11222 7892 11228
rect 8024 11144 8076 11150
rect 7838 11112 7894 11121
rect 8024 11086 8076 11092
rect 7838 11047 7894 11056
rect 7852 10674 7880 11047
rect 7932 11008 7984 11014
rect 7932 10950 7984 10956
rect 7944 10742 7972 10950
rect 7932 10736 7984 10742
rect 7932 10678 7984 10684
rect 7656 10668 7708 10674
rect 7656 10610 7708 10616
rect 7840 10668 7892 10674
rect 7840 10610 7892 10616
rect 7668 10130 7696 10610
rect 7656 10124 7708 10130
rect 7656 10066 7708 10072
rect 7840 10124 7892 10130
rect 7892 10084 7972 10112
rect 7840 10066 7892 10072
rect 7564 10056 7616 10062
rect 7564 9998 7616 10004
rect 7470 9752 7526 9761
rect 7470 9687 7472 9696
rect 7524 9687 7526 9696
rect 7472 9658 7524 9664
rect 7484 9627 7512 9658
rect 7194 9616 7250 9625
rect 7194 9551 7250 9560
rect 7196 9512 7248 9518
rect 7196 9454 7248 9460
rect 7104 9172 7156 9178
rect 7104 9114 7156 9120
rect 7012 9036 7064 9042
rect 7012 8978 7064 8984
rect 7116 8974 7144 9114
rect 7104 8968 7156 8974
rect 7104 8910 7156 8916
rect 6880 8860 6960 8888
rect 6828 8842 6880 8848
rect 6552 8628 6604 8634
rect 7208 8616 7236 9454
rect 7576 9450 7604 9998
rect 7668 9586 7696 10066
rect 7748 10056 7800 10062
rect 7748 9998 7800 10004
rect 7760 9722 7788 9998
rect 7840 9920 7892 9926
rect 7840 9862 7892 9868
rect 7748 9716 7800 9722
rect 7748 9658 7800 9664
rect 7656 9580 7708 9586
rect 7656 9522 7708 9528
rect 7852 9518 7880 9862
rect 7840 9512 7892 9518
rect 7840 9454 7892 9460
rect 7564 9444 7616 9450
rect 7564 9386 7616 9392
rect 7852 8974 7880 9454
rect 7944 9382 7972 10084
rect 8036 9450 8064 11086
rect 8128 9586 8156 11455
rect 8312 11218 8340 11580
rect 8404 11558 8432 11727
rect 8588 11642 8616 14200
rect 8668 13524 8720 13530
rect 8668 13466 8720 13472
rect 8680 13326 8708 13466
rect 9036 13456 9088 13462
rect 8850 13424 8906 13433
rect 9036 13398 9088 13404
rect 8850 13359 8906 13368
rect 8668 13320 8720 13326
rect 8668 13262 8720 13268
rect 8760 13320 8812 13326
rect 8760 13262 8812 13268
rect 8680 12481 8708 13262
rect 8772 12850 8800 13262
rect 8864 12850 8892 13359
rect 9048 12850 9076 13398
rect 9680 13184 9732 13190
rect 9680 13126 9732 13132
rect 9692 12986 9720 13126
rect 9680 12980 9732 12986
rect 9680 12922 9732 12928
rect 9310 12880 9366 12889
rect 8760 12844 8812 12850
rect 8760 12786 8812 12792
rect 8852 12844 8904 12850
rect 8852 12786 8904 12792
rect 9036 12844 9088 12850
rect 9310 12815 9366 12824
rect 9036 12786 9088 12792
rect 8666 12472 8722 12481
rect 8666 12407 8668 12416
rect 8720 12407 8722 12416
rect 8668 12378 8720 12384
rect 8680 12347 8708 12378
rect 8864 12306 8892 12786
rect 8944 12708 8996 12714
rect 8944 12650 8996 12656
rect 8852 12300 8904 12306
rect 8852 12242 8904 12248
rect 8668 12232 8720 12238
rect 8720 12180 8800 12186
rect 8668 12174 8800 12180
rect 8680 12158 8800 12174
rect 8668 12096 8720 12102
rect 8668 12038 8720 12044
rect 8680 11898 8708 12038
rect 8668 11892 8720 11898
rect 8668 11834 8720 11840
rect 8772 11830 8800 12158
rect 8850 11928 8906 11937
rect 8850 11863 8906 11872
rect 8760 11824 8812 11830
rect 8760 11766 8812 11772
rect 8588 11614 8800 11642
rect 8392 11552 8444 11558
rect 8392 11494 8444 11500
rect 8668 11552 8720 11558
rect 8668 11494 8720 11500
rect 8680 11354 8708 11494
rect 8668 11348 8720 11354
rect 8668 11290 8720 11296
rect 8576 11280 8628 11286
rect 8576 11222 8628 11228
rect 8300 11212 8352 11218
rect 8300 11154 8352 11160
rect 8214 10908 8522 10917
rect 8214 10906 8220 10908
rect 8276 10906 8300 10908
rect 8356 10906 8380 10908
rect 8436 10906 8460 10908
rect 8516 10906 8522 10908
rect 8276 10854 8278 10906
rect 8458 10854 8460 10906
rect 8214 10852 8220 10854
rect 8276 10852 8300 10854
rect 8356 10852 8380 10854
rect 8436 10852 8460 10854
rect 8516 10852 8522 10854
rect 8214 10843 8522 10852
rect 8392 10804 8444 10810
rect 8588 10792 8616 11222
rect 8668 11212 8720 11218
rect 8668 11154 8720 11160
rect 8392 10746 8444 10752
rect 8496 10764 8616 10792
rect 8404 10713 8432 10746
rect 8390 10704 8446 10713
rect 8208 10668 8260 10674
rect 8390 10639 8446 10648
rect 8208 10610 8260 10616
rect 8220 10198 8248 10610
rect 8392 10532 8444 10538
rect 8392 10474 8444 10480
rect 8208 10192 8260 10198
rect 8208 10134 8260 10140
rect 8404 9926 8432 10474
rect 8496 10266 8524 10764
rect 8576 10532 8628 10538
rect 8576 10474 8628 10480
rect 8484 10260 8536 10266
rect 8484 10202 8536 10208
rect 8484 10124 8536 10130
rect 8484 10066 8536 10072
rect 8496 10033 8524 10066
rect 8588 10062 8616 10474
rect 8576 10056 8628 10062
rect 8482 10024 8538 10033
rect 8576 9998 8628 10004
rect 8482 9959 8538 9968
rect 8392 9920 8444 9926
rect 8392 9862 8444 9868
rect 8214 9820 8522 9829
rect 8214 9818 8220 9820
rect 8276 9818 8300 9820
rect 8356 9818 8380 9820
rect 8436 9818 8460 9820
rect 8516 9818 8522 9820
rect 8276 9766 8278 9818
rect 8458 9766 8460 9818
rect 8214 9764 8220 9766
rect 8276 9764 8300 9766
rect 8356 9764 8380 9766
rect 8436 9764 8460 9766
rect 8516 9764 8522 9766
rect 8214 9755 8522 9764
rect 8392 9716 8444 9722
rect 8392 9658 8444 9664
rect 8116 9580 8168 9586
rect 8116 9522 8168 9528
rect 8024 9444 8076 9450
rect 8024 9386 8076 9392
rect 7932 9376 7984 9382
rect 7932 9318 7984 9324
rect 7840 8968 7892 8974
rect 7760 8928 7840 8956
rect 7564 8900 7616 8906
rect 7564 8842 7616 8848
rect 7576 8634 7604 8842
rect 6552 8570 6604 8576
rect 6932 8588 7236 8616
rect 7564 8628 7616 8634
rect 6564 8498 6592 8570
rect 6828 8560 6880 8566
rect 6932 8548 6960 8588
rect 7564 8570 7616 8576
rect 6880 8520 6960 8548
rect 6828 8502 6880 8508
rect 6184 8492 6236 8498
rect 6184 8434 6236 8440
rect 6552 8492 6604 8498
rect 6552 8434 6604 8440
rect 7012 8492 7064 8498
rect 7012 8434 7064 8440
rect 6196 7970 6224 8434
rect 6920 8424 6972 8430
rect 6920 8366 6972 8372
rect 6104 7954 6224 7970
rect 6092 7948 6224 7954
rect 6144 7942 6224 7948
rect 6092 7890 6144 7896
rect 6828 7880 6880 7886
rect 6828 7822 6880 7828
rect 6276 7744 6328 7750
rect 6276 7686 6328 7692
rect 6288 7410 6316 7686
rect 6840 7546 6868 7822
rect 6828 7540 6880 7546
rect 6828 7482 6880 7488
rect 6932 7478 6960 8366
rect 6736 7472 6788 7478
rect 6736 7414 6788 7420
rect 6920 7472 6972 7478
rect 6920 7414 6972 7420
rect 5724 7404 5776 7410
rect 5538 7375 5540 7384
rect 5448 7346 5500 7352
rect 5592 7375 5594 7384
rect 5540 7346 5592 7352
rect 5644 7364 5724 7392
rect 4172 7256 4200 7346
rect 4080 7228 4200 7256
rect 3882 6967 3938 6976
rect 3976 6996 4028 7002
rect 3332 6792 3384 6798
rect 3792 6792 3844 6798
rect 3332 6734 3384 6740
rect 3712 6752 3792 6780
rect 3056 6452 3108 6458
rect 3056 6394 3108 6400
rect 3148 6180 3200 6186
rect 3148 6122 3200 6128
rect 3160 5778 3188 6122
rect 3148 5772 3200 5778
rect 3148 5714 3200 5720
rect 3608 5636 3660 5642
rect 3608 5578 3660 5584
rect 3332 5568 3384 5574
rect 3332 5510 3384 5516
rect 3424 5568 3476 5574
rect 3424 5510 3476 5516
rect 3240 5228 3292 5234
rect 3344 5216 3372 5510
rect 3292 5188 3372 5216
rect 3240 5170 3292 5176
rect 3240 5092 3292 5098
rect 3160 5052 3240 5080
rect 3160 3942 3188 5052
rect 3240 5034 3292 5040
rect 3240 4820 3292 4826
rect 3240 4762 3292 4768
rect 3252 4486 3280 4762
rect 3344 4622 3372 5188
rect 3436 5030 3464 5510
rect 3620 5302 3648 5578
rect 3608 5296 3660 5302
rect 3608 5238 3660 5244
rect 3424 5024 3476 5030
rect 3424 4966 3476 4972
rect 3436 4690 3464 4966
rect 3424 4684 3476 4690
rect 3424 4626 3476 4632
rect 3332 4616 3384 4622
rect 3332 4558 3384 4564
rect 3240 4480 3292 4486
rect 3240 4422 3292 4428
rect 3516 4480 3568 4486
rect 3516 4422 3568 4428
rect 3148 3936 3200 3942
rect 3148 3878 3200 3884
rect 3252 3398 3280 4422
rect 3528 4185 3556 4422
rect 3712 4214 3740 6752
rect 3792 6734 3844 6740
rect 3792 5024 3844 5030
rect 3792 4966 3844 4972
rect 3804 4622 3832 4966
rect 3792 4616 3844 4622
rect 3792 4558 3844 4564
rect 3700 4208 3752 4214
rect 3514 4176 3570 4185
rect 3700 4150 3752 4156
rect 3514 4111 3516 4120
rect 3568 4111 3570 4120
rect 3516 4082 3568 4088
rect 3424 4004 3476 4010
rect 3424 3946 3476 3952
rect 3332 3528 3384 3534
rect 3332 3470 3384 3476
rect 3240 3392 3292 3398
rect 3240 3334 3292 3340
rect 3344 3126 3372 3470
rect 3332 3120 3384 3126
rect 3332 3062 3384 3068
rect 3240 3052 3292 3058
rect 3240 2994 3292 3000
rect 3148 2304 3200 2310
rect 3148 2246 3200 2252
rect 3160 2038 3188 2246
rect 3148 2032 3200 2038
rect 3148 1974 3200 1980
rect 2962 1320 3018 1329
rect 3252 1290 3280 2994
rect 3436 2582 3464 3946
rect 3528 3602 3556 4082
rect 3606 4040 3662 4049
rect 3606 3975 3662 3984
rect 3516 3596 3568 3602
rect 3516 3538 3568 3544
rect 3424 2576 3476 2582
rect 3424 2518 3476 2524
rect 3332 2304 3384 2310
rect 3332 2246 3384 2252
rect 3344 1290 3372 2246
rect 3436 2106 3464 2518
rect 3620 2514 3648 3975
rect 3792 2576 3844 2582
rect 3792 2518 3844 2524
rect 3608 2508 3660 2514
rect 3608 2450 3660 2456
rect 3700 2372 3752 2378
rect 3700 2314 3752 2320
rect 3424 2100 3476 2106
rect 3424 2042 3476 2048
rect 3436 1494 3464 2042
rect 3516 1964 3568 1970
rect 3516 1906 3568 1912
rect 3424 1488 3476 1494
rect 3424 1430 3476 1436
rect 3528 1358 3556 1906
rect 3712 1426 3740 2314
rect 3804 1970 3832 2518
rect 3792 1964 3844 1970
rect 3792 1906 3844 1912
rect 3700 1420 3752 1426
rect 3700 1362 3752 1368
rect 3896 1358 3924 6967
rect 3976 6938 4028 6944
rect 3976 6860 4028 6866
rect 3976 6802 4028 6808
rect 3988 6390 4016 6802
rect 4080 6662 4108 7228
rect 4620 7200 4672 7206
rect 4620 7142 4672 7148
rect 5264 7200 5316 7206
rect 5264 7142 5316 7148
rect 4214 7100 4522 7109
rect 4214 7098 4220 7100
rect 4276 7098 4300 7100
rect 4356 7098 4380 7100
rect 4436 7098 4460 7100
rect 4516 7098 4522 7100
rect 4276 7046 4278 7098
rect 4458 7046 4460 7098
rect 4214 7044 4220 7046
rect 4276 7044 4300 7046
rect 4356 7044 4380 7046
rect 4436 7044 4460 7046
rect 4516 7044 4522 7046
rect 4214 7035 4522 7044
rect 4160 6996 4212 7002
rect 4160 6938 4212 6944
rect 4172 6798 4200 6938
rect 4160 6792 4212 6798
rect 4160 6734 4212 6740
rect 4068 6656 4120 6662
rect 4068 6598 4120 6604
rect 3976 6384 4028 6390
rect 3976 6326 4028 6332
rect 4066 6352 4122 6361
rect 4066 6287 4122 6296
rect 4080 6254 4108 6287
rect 4068 6248 4120 6254
rect 4068 6190 4120 6196
rect 4080 5846 4108 6190
rect 4632 6118 4660 7142
rect 5276 6798 5304 7142
rect 5644 7002 5672 7364
rect 5724 7346 5776 7352
rect 6276 7404 6328 7410
rect 6276 7346 6328 7352
rect 6092 7336 6144 7342
rect 6092 7278 6144 7284
rect 5724 7268 5776 7274
rect 5724 7210 5776 7216
rect 5632 6996 5684 7002
rect 5632 6938 5684 6944
rect 5632 6860 5684 6866
rect 5632 6802 5684 6808
rect 5264 6792 5316 6798
rect 5264 6734 5316 6740
rect 5540 6452 5592 6458
rect 5540 6394 5592 6400
rect 5356 6248 5408 6254
rect 5356 6190 5408 6196
rect 4620 6112 4672 6118
rect 4672 6072 4752 6100
rect 4620 6054 4672 6060
rect 4214 6012 4522 6021
rect 4214 6010 4220 6012
rect 4276 6010 4300 6012
rect 4356 6010 4380 6012
rect 4436 6010 4460 6012
rect 4516 6010 4522 6012
rect 4276 5958 4278 6010
rect 4458 5958 4460 6010
rect 4214 5956 4220 5958
rect 4276 5956 4300 5958
rect 4356 5956 4380 5958
rect 4436 5956 4460 5958
rect 4516 5956 4522 5958
rect 4214 5947 4522 5956
rect 4068 5840 4120 5846
rect 4068 5782 4120 5788
rect 4620 5772 4672 5778
rect 4620 5714 4672 5720
rect 3976 5636 4028 5642
rect 3976 5578 4028 5584
rect 4436 5636 4488 5642
rect 4436 5578 4488 5584
rect 3988 5250 4016 5578
rect 4068 5568 4120 5574
rect 4068 5510 4120 5516
rect 4080 5370 4108 5510
rect 4068 5364 4120 5370
rect 4068 5306 4120 5312
rect 4448 5302 4476 5578
rect 4632 5302 4660 5714
rect 4724 5710 4752 6072
rect 5368 5914 5396 6190
rect 5356 5908 5408 5914
rect 5356 5850 5408 5856
rect 4712 5704 4764 5710
rect 4712 5646 4764 5652
rect 5552 5574 5580 6394
rect 5540 5568 5592 5574
rect 5540 5510 5592 5516
rect 4436 5296 4488 5302
rect 3988 5234 4108 5250
rect 4436 5238 4488 5244
rect 4620 5296 4672 5302
rect 4620 5238 4672 5244
rect 5448 5296 5500 5302
rect 5448 5238 5500 5244
rect 3988 5228 4120 5234
rect 3988 5222 4068 5228
rect 4068 5170 4120 5176
rect 5356 5228 5408 5234
rect 5356 5170 5408 5176
rect 4080 3602 4108 5170
rect 4214 4924 4522 4933
rect 4214 4922 4220 4924
rect 4276 4922 4300 4924
rect 4356 4922 4380 4924
rect 4436 4922 4460 4924
rect 4516 4922 4522 4924
rect 4276 4870 4278 4922
rect 4458 4870 4460 4922
rect 4214 4868 4220 4870
rect 4276 4868 4300 4870
rect 4356 4868 4380 4870
rect 4436 4868 4460 4870
rect 4516 4868 4522 4870
rect 4214 4859 4522 4868
rect 4252 4616 4304 4622
rect 4252 4558 4304 4564
rect 4264 4146 4292 4558
rect 4528 4480 4580 4486
rect 4528 4422 4580 4428
rect 4540 4146 4568 4422
rect 5368 4282 5396 5170
rect 4712 4276 4764 4282
rect 4712 4218 4764 4224
rect 5356 4276 5408 4282
rect 5356 4218 5408 4224
rect 4252 4140 4304 4146
rect 4252 4082 4304 4088
rect 4528 4140 4580 4146
rect 4724 4128 4752 4218
rect 4580 4100 4752 4128
rect 4816 4134 5028 4162
rect 4528 4082 4580 4088
rect 4816 4010 4844 4134
rect 4896 4072 4948 4078
rect 4894 4040 4896 4049
rect 4948 4040 4950 4049
rect 4804 4004 4856 4010
rect 5000 4010 5028 4134
rect 4894 3975 4950 3984
rect 4988 4004 5040 4010
rect 4804 3946 4856 3952
rect 4214 3836 4522 3845
rect 4214 3834 4220 3836
rect 4276 3834 4300 3836
rect 4356 3834 4380 3836
rect 4436 3834 4460 3836
rect 4516 3834 4522 3836
rect 4276 3782 4278 3834
rect 4458 3782 4460 3834
rect 4214 3780 4220 3782
rect 4276 3780 4300 3782
rect 4356 3780 4380 3782
rect 4436 3780 4460 3782
rect 4516 3780 4522 3782
rect 4214 3771 4522 3780
rect 4068 3596 4120 3602
rect 4068 3538 4120 3544
rect 4344 3528 4396 3534
rect 4344 3470 4396 3476
rect 4436 3528 4488 3534
rect 4436 3470 4488 3476
rect 4712 3528 4764 3534
rect 4712 3470 4764 3476
rect 4356 2990 4384 3470
rect 4448 3058 4476 3470
rect 4724 3194 4752 3470
rect 4712 3188 4764 3194
rect 4712 3130 4764 3136
rect 4436 3052 4488 3058
rect 4436 2994 4488 3000
rect 4712 3052 4764 3058
rect 4712 2994 4764 3000
rect 4344 2984 4396 2990
rect 4344 2926 4396 2932
rect 4620 2984 4672 2990
rect 4620 2926 4672 2932
rect 4214 2748 4522 2757
rect 4214 2746 4220 2748
rect 4276 2746 4300 2748
rect 4356 2746 4380 2748
rect 4436 2746 4460 2748
rect 4516 2746 4522 2748
rect 4276 2694 4278 2746
rect 4458 2694 4460 2746
rect 4214 2692 4220 2694
rect 4276 2692 4300 2694
rect 4356 2692 4380 2694
rect 4436 2692 4460 2694
rect 4516 2692 4522 2694
rect 4214 2683 4522 2692
rect 4632 2514 4660 2926
rect 4724 2650 4752 2994
rect 4712 2644 4764 2650
rect 4712 2586 4764 2592
rect 4620 2508 4672 2514
rect 4620 2450 4672 2456
rect 4620 2032 4672 2038
rect 4620 1974 4672 1980
rect 4068 1896 4120 1902
rect 4068 1838 4120 1844
rect 3516 1352 3568 1358
rect 3516 1294 3568 1300
rect 3884 1352 3936 1358
rect 3884 1294 3936 1300
rect 2962 1255 3018 1264
rect 3240 1284 3292 1290
rect 3240 1226 3292 1232
rect 3332 1284 3384 1290
rect 3332 1226 3384 1232
rect 3700 1216 3752 1222
rect 3700 1158 3752 1164
rect 3712 800 3740 1158
rect 3896 1018 3924 1294
rect 4080 1170 4108 1838
rect 4214 1660 4522 1669
rect 4214 1658 4220 1660
rect 4276 1658 4300 1660
rect 4356 1658 4380 1660
rect 4436 1658 4460 1660
rect 4516 1658 4522 1660
rect 4276 1606 4278 1658
rect 4458 1606 4460 1658
rect 4214 1604 4220 1606
rect 4276 1604 4300 1606
rect 4356 1604 4380 1606
rect 4436 1604 4460 1606
rect 4516 1604 4522 1606
rect 4214 1595 4522 1604
rect 4436 1556 4488 1562
rect 4436 1498 4488 1504
rect 4252 1488 4304 1494
rect 4252 1430 4304 1436
rect 4264 1358 4292 1430
rect 4448 1358 4476 1498
rect 4632 1358 4660 1974
rect 4908 1426 4936 3975
rect 4988 3946 5040 3952
rect 5368 3534 5396 4218
rect 5460 4146 5488 5238
rect 5644 4826 5672 6802
rect 5736 6322 5764 7210
rect 6104 6458 6132 7278
rect 6460 6860 6512 6866
rect 6460 6802 6512 6808
rect 6092 6452 6144 6458
rect 6092 6394 6144 6400
rect 5724 6316 5776 6322
rect 5724 6258 5776 6264
rect 5724 5908 5776 5914
rect 6104 5896 6132 6394
rect 6472 6322 6500 6802
rect 6552 6724 6604 6730
rect 6552 6666 6604 6672
rect 6564 6458 6592 6666
rect 6552 6452 6604 6458
rect 6552 6394 6604 6400
rect 6460 6316 6512 6322
rect 6460 6258 6512 6264
rect 6748 6254 6776 7414
rect 7024 7342 7052 8434
rect 7196 7948 7248 7954
rect 7196 7890 7248 7896
rect 7208 7410 7236 7890
rect 7380 7744 7432 7750
rect 7380 7686 7432 7692
rect 7196 7404 7248 7410
rect 7196 7346 7248 7352
rect 7012 7336 7064 7342
rect 7012 7278 7064 7284
rect 6920 6860 6972 6866
rect 6920 6802 6972 6808
rect 6932 6390 6960 6802
rect 7208 6798 7236 7346
rect 7392 7002 7420 7686
rect 7472 7540 7524 7546
rect 7472 7482 7524 7488
rect 7380 6996 7432 7002
rect 7380 6938 7432 6944
rect 7196 6792 7248 6798
rect 7196 6734 7248 6740
rect 7484 6390 7512 7482
rect 7576 7478 7604 8570
rect 7656 8288 7708 8294
rect 7656 8230 7708 8236
rect 7668 7886 7696 8230
rect 7760 7954 7788 8928
rect 7840 8910 7892 8916
rect 7840 8492 7892 8498
rect 7840 8434 7892 8440
rect 7852 8090 7880 8434
rect 7840 8084 7892 8090
rect 7840 8026 7892 8032
rect 7748 7948 7800 7954
rect 7748 7890 7800 7896
rect 7656 7880 7708 7886
rect 7656 7822 7708 7828
rect 7564 7472 7616 7478
rect 7564 7414 7616 7420
rect 7760 6882 7788 7890
rect 7852 6934 7880 8026
rect 7668 6866 7788 6882
rect 7840 6928 7892 6934
rect 7840 6870 7892 6876
rect 7656 6860 7788 6866
rect 7708 6854 7788 6860
rect 7656 6802 7708 6808
rect 7748 6724 7800 6730
rect 7748 6666 7800 6672
rect 6920 6384 6972 6390
rect 6920 6326 6972 6332
rect 7472 6384 7524 6390
rect 7472 6326 7524 6332
rect 6736 6248 6788 6254
rect 6736 6190 6788 6196
rect 5724 5850 5776 5856
rect 5920 5868 6132 5896
rect 5632 4820 5684 4826
rect 5632 4762 5684 4768
rect 5644 4690 5672 4762
rect 5632 4684 5684 4690
rect 5632 4626 5684 4632
rect 5736 4622 5764 5850
rect 5920 5710 5948 5868
rect 6000 5772 6052 5778
rect 6000 5714 6052 5720
rect 5908 5704 5960 5710
rect 5908 5646 5960 5652
rect 5920 5302 5948 5646
rect 5908 5296 5960 5302
rect 5908 5238 5960 5244
rect 6012 5234 6040 5714
rect 6184 5704 6236 5710
rect 6184 5646 6236 5652
rect 6092 5636 6144 5642
rect 6092 5578 6144 5584
rect 6000 5228 6052 5234
rect 6000 5170 6052 5176
rect 5908 5024 5960 5030
rect 5908 4966 5960 4972
rect 5920 4622 5948 4966
rect 6104 4622 6132 5578
rect 6196 4758 6224 5646
rect 6644 4820 6696 4826
rect 6644 4762 6696 4768
rect 6184 4752 6236 4758
rect 6184 4694 6236 4700
rect 5724 4616 5776 4622
rect 5724 4558 5776 4564
rect 5908 4616 5960 4622
rect 5908 4558 5960 4564
rect 6092 4616 6144 4622
rect 6092 4558 6144 4564
rect 5540 4480 5592 4486
rect 5540 4422 5592 4428
rect 5552 4282 5580 4422
rect 5736 4298 5764 4558
rect 5540 4276 5592 4282
rect 5540 4218 5592 4224
rect 5644 4270 5764 4298
rect 6104 4282 6132 4558
rect 6092 4276 6144 4282
rect 5448 4140 5500 4146
rect 5448 4082 5500 4088
rect 5356 3528 5408 3534
rect 5356 3470 5408 3476
rect 5460 3466 5488 4082
rect 5644 4049 5672 4270
rect 6092 4218 6144 4224
rect 5724 4208 5776 4214
rect 5724 4150 5776 4156
rect 5630 4040 5686 4049
rect 5630 3975 5686 3984
rect 5736 3534 5764 4150
rect 5724 3528 5776 3534
rect 5724 3470 5776 3476
rect 5448 3460 5500 3466
rect 5448 3402 5500 3408
rect 5460 3194 5488 3402
rect 5448 3188 5500 3194
rect 5448 3130 5500 3136
rect 5356 3052 5408 3058
rect 5356 2994 5408 3000
rect 5448 3052 5500 3058
rect 5448 2994 5500 3000
rect 5368 2446 5396 2994
rect 5460 2446 5488 2994
rect 6196 2854 6224 4694
rect 6656 4282 6684 4762
rect 6748 4622 6776 6190
rect 6828 4684 6880 4690
rect 6932 4672 6960 6326
rect 7760 6254 7788 6666
rect 7944 6322 7972 9318
rect 8036 9178 8064 9386
rect 8404 9178 8432 9658
rect 8484 9580 8536 9586
rect 8484 9522 8536 9528
rect 8496 9353 8524 9522
rect 8482 9344 8538 9353
rect 8482 9279 8538 9288
rect 8024 9172 8076 9178
rect 8024 9114 8076 9120
rect 8392 9172 8444 9178
rect 8392 9114 8444 9120
rect 8588 8974 8616 9998
rect 8680 9110 8708 11154
rect 8772 11121 8800 11614
rect 8864 11354 8892 11863
rect 8852 11348 8904 11354
rect 8852 11290 8904 11296
rect 8758 11112 8814 11121
rect 8758 11047 8814 11056
rect 8772 10742 8800 11047
rect 8850 10976 8906 10985
rect 8850 10911 8906 10920
rect 8760 10736 8812 10742
rect 8760 10678 8812 10684
rect 8864 9722 8892 10911
rect 8956 10810 8984 12650
rect 9048 12306 9076 12786
rect 9218 12336 9274 12345
rect 9036 12300 9088 12306
rect 9218 12271 9274 12280
rect 9036 12242 9088 12248
rect 9232 12170 9260 12271
rect 9324 12238 9352 12815
rect 9496 12436 9548 12442
rect 9496 12378 9548 12384
rect 9312 12232 9364 12238
rect 9312 12174 9364 12180
rect 9128 12164 9180 12170
rect 9128 12106 9180 12112
rect 9220 12164 9272 12170
rect 9220 12106 9272 12112
rect 9140 11744 9168 12106
rect 9140 11716 9260 11744
rect 9232 11626 9260 11716
rect 9220 11620 9272 11626
rect 9220 11562 9272 11568
rect 9036 11552 9088 11558
rect 9036 11494 9088 11500
rect 9048 11336 9076 11494
rect 9232 11393 9260 11562
rect 9218 11384 9274 11393
rect 9128 11348 9180 11354
rect 9048 11308 9128 11336
rect 9324 11354 9352 12174
rect 9508 11762 9536 12378
rect 9586 12200 9642 12209
rect 9586 12135 9642 12144
rect 9600 11830 9628 12135
rect 9588 11824 9640 11830
rect 9588 11766 9640 11772
rect 9496 11756 9548 11762
rect 9496 11698 9548 11704
rect 9680 11756 9732 11762
rect 9680 11698 9732 11704
rect 9404 11688 9456 11694
rect 9404 11630 9456 11636
rect 9494 11656 9550 11665
rect 9218 11319 9274 11328
rect 9312 11348 9364 11354
rect 9128 11290 9180 11296
rect 9312 11290 9364 11296
rect 9128 11212 9180 11218
rect 9312 11212 9364 11218
rect 9180 11172 9312 11200
rect 9128 11154 9180 11160
rect 9416 11200 9444 11630
rect 9494 11591 9550 11600
rect 9508 11558 9536 11591
rect 9496 11552 9548 11558
rect 9496 11494 9548 11500
rect 9586 11520 9642 11529
rect 9586 11455 9642 11464
rect 9364 11172 9444 11200
rect 9312 11154 9364 11160
rect 9600 11150 9628 11455
rect 9692 11150 9720 11698
rect 9784 11354 9812 14200
rect 10600 13320 10652 13326
rect 10600 13262 10652 13268
rect 10048 13252 10100 13258
rect 10048 13194 10100 13200
rect 9864 13184 9916 13190
rect 9864 13126 9916 13132
rect 9956 13184 10008 13190
rect 9956 13126 10008 13132
rect 9876 12918 9904 13126
rect 9864 12912 9916 12918
rect 9864 12854 9916 12860
rect 9864 12708 9916 12714
rect 9864 12650 9916 12656
rect 9876 12238 9904 12650
rect 9968 12306 9996 13126
rect 9956 12300 10008 12306
rect 9956 12242 10008 12248
rect 9864 12232 9916 12238
rect 9864 12174 9916 12180
rect 9862 11792 9918 11801
rect 9862 11727 9864 11736
rect 9916 11727 9918 11736
rect 9956 11756 10008 11762
rect 9864 11698 9916 11704
rect 9956 11698 10008 11704
rect 9772 11348 9824 11354
rect 9772 11290 9824 11296
rect 9036 11144 9088 11150
rect 9588 11144 9640 11150
rect 9088 11092 9352 11098
rect 9036 11086 9352 11092
rect 9588 11086 9640 11092
rect 9680 11144 9732 11150
rect 9680 11086 9732 11092
rect 9048 11070 9352 11086
rect 9036 11008 9088 11014
rect 9036 10950 9088 10956
rect 8944 10804 8996 10810
rect 8944 10746 8996 10752
rect 8944 10600 8996 10606
rect 8944 10542 8996 10548
rect 8956 10130 8984 10542
rect 8944 10124 8996 10130
rect 8944 10066 8996 10072
rect 8852 9716 8904 9722
rect 8852 9658 8904 9664
rect 8760 9580 8812 9586
rect 8760 9522 8812 9528
rect 8668 9104 8720 9110
rect 8668 9046 8720 9052
rect 8772 8974 8800 9522
rect 8852 9376 8904 9382
rect 8852 9318 8904 9324
rect 8864 9110 8892 9318
rect 8956 9178 8984 10066
rect 9048 9217 9076 10950
rect 9220 10736 9272 10742
rect 9220 10678 9272 10684
rect 9128 10668 9180 10674
rect 9128 10610 9180 10616
rect 9034 9208 9090 9217
rect 8944 9172 8996 9178
rect 9140 9178 9168 10610
rect 9232 10577 9260 10678
rect 9218 10568 9274 10577
rect 9218 10503 9274 10512
rect 9324 10452 9352 11070
rect 9692 10742 9720 11086
rect 9680 10736 9732 10742
rect 9680 10678 9732 10684
rect 9404 10668 9456 10674
rect 9404 10610 9456 10616
rect 9588 10668 9640 10674
rect 9588 10610 9640 10616
rect 9232 10424 9352 10452
rect 9232 9722 9260 10424
rect 9416 10305 9444 10610
rect 9600 10418 9628 10610
rect 9678 10432 9734 10441
rect 9600 10390 9678 10418
rect 9678 10367 9734 10376
rect 9402 10296 9458 10305
rect 9586 10296 9642 10305
rect 9402 10231 9458 10240
rect 9496 10260 9548 10266
rect 9586 10231 9642 10240
rect 9496 10202 9548 10208
rect 9508 9926 9536 10202
rect 9600 10062 9628 10231
rect 9784 10130 9812 11290
rect 9968 11082 9996 11698
rect 10060 11626 10088 13194
rect 10416 13184 10468 13190
rect 10416 13126 10468 13132
rect 10232 12912 10284 12918
rect 10232 12854 10284 12860
rect 10048 11620 10100 11626
rect 10048 11562 10100 11568
rect 10060 11286 10088 11562
rect 10048 11280 10100 11286
rect 10048 11222 10100 11228
rect 10048 11144 10100 11150
rect 10048 11086 10100 11092
rect 9956 11076 10008 11082
rect 9956 11018 10008 11024
rect 9862 10704 9918 10713
rect 9862 10639 9918 10648
rect 9876 10606 9904 10639
rect 9864 10600 9916 10606
rect 9864 10542 9916 10548
rect 9956 10464 10008 10470
rect 9956 10406 10008 10412
rect 9864 10192 9916 10198
rect 9862 10160 9864 10169
rect 9916 10160 9918 10169
rect 9772 10124 9824 10130
rect 9862 10095 9918 10104
rect 9772 10066 9824 10072
rect 9588 10056 9640 10062
rect 9588 9998 9640 10004
rect 9772 9988 9824 9994
rect 9772 9930 9824 9936
rect 9312 9920 9364 9926
rect 9310 9888 9312 9897
rect 9496 9920 9548 9926
rect 9364 9888 9366 9897
rect 9496 9862 9548 9868
rect 9310 9823 9366 9832
rect 9220 9716 9272 9722
rect 9220 9658 9272 9664
rect 9034 9143 9090 9152
rect 9128 9172 9180 9178
rect 8944 9114 8996 9120
rect 9128 9114 9180 9120
rect 8852 9104 8904 9110
rect 8852 9046 8904 9052
rect 9036 9036 9088 9042
rect 9036 8978 9088 8984
rect 8208 8968 8260 8974
rect 8206 8936 8208 8945
rect 8576 8968 8628 8974
rect 8260 8936 8262 8945
rect 8128 8894 8206 8922
rect 8128 8566 8156 8894
rect 8576 8910 8628 8916
rect 8760 8968 8812 8974
rect 8760 8910 8812 8916
rect 8206 8871 8262 8880
rect 8214 8732 8522 8741
rect 8214 8730 8220 8732
rect 8276 8730 8300 8732
rect 8356 8730 8380 8732
rect 8436 8730 8460 8732
rect 8516 8730 8522 8732
rect 8276 8678 8278 8730
rect 8458 8678 8460 8730
rect 8214 8676 8220 8678
rect 8276 8676 8300 8678
rect 8356 8676 8380 8678
rect 8436 8676 8460 8678
rect 8516 8676 8522 8678
rect 8214 8667 8522 8676
rect 8116 8560 8168 8566
rect 8116 8502 8168 8508
rect 8024 8424 8076 8430
rect 8024 8366 8076 8372
rect 8036 7954 8064 8366
rect 8944 8288 8996 8294
rect 8944 8230 8996 8236
rect 8024 7948 8076 7954
rect 8024 7890 8076 7896
rect 8036 7206 8064 7890
rect 8116 7880 8168 7886
rect 8116 7822 8168 7828
rect 8128 7546 8156 7822
rect 8214 7644 8522 7653
rect 8214 7642 8220 7644
rect 8276 7642 8300 7644
rect 8356 7642 8380 7644
rect 8436 7642 8460 7644
rect 8516 7642 8522 7644
rect 8276 7590 8278 7642
rect 8458 7590 8460 7642
rect 8214 7588 8220 7590
rect 8276 7588 8300 7590
rect 8356 7588 8380 7590
rect 8436 7588 8460 7590
rect 8516 7588 8522 7590
rect 8214 7579 8522 7588
rect 8116 7540 8168 7546
rect 8116 7482 8168 7488
rect 8024 7200 8076 7206
rect 8024 7142 8076 7148
rect 8036 6798 8064 7142
rect 8024 6792 8076 6798
rect 8024 6734 8076 6740
rect 7932 6316 7984 6322
rect 7932 6258 7984 6264
rect 7748 6248 7800 6254
rect 7748 6190 7800 6196
rect 7760 5778 7788 6190
rect 8128 5914 8156 7482
rect 8956 7410 8984 8230
rect 9048 7886 9076 8978
rect 9128 8832 9180 8838
rect 9128 8774 9180 8780
rect 9036 7880 9088 7886
rect 9036 7822 9088 7828
rect 8944 7404 8996 7410
rect 8944 7346 8996 7352
rect 8392 7336 8444 7342
rect 8392 7278 8444 7284
rect 8852 7336 8904 7342
rect 8852 7278 8904 7284
rect 8300 7268 8352 7274
rect 8300 7210 8352 7216
rect 8312 6798 8340 7210
rect 8404 6798 8432 7278
rect 8576 6860 8628 6866
rect 8576 6802 8628 6808
rect 8300 6792 8352 6798
rect 8300 6734 8352 6740
rect 8392 6792 8444 6798
rect 8392 6734 8444 6740
rect 8214 6556 8522 6565
rect 8214 6554 8220 6556
rect 8276 6554 8300 6556
rect 8356 6554 8380 6556
rect 8436 6554 8460 6556
rect 8516 6554 8522 6556
rect 8276 6502 8278 6554
rect 8458 6502 8460 6554
rect 8214 6500 8220 6502
rect 8276 6500 8300 6502
rect 8356 6500 8380 6502
rect 8436 6500 8460 6502
rect 8516 6500 8522 6502
rect 8214 6491 8522 6500
rect 8116 5908 8168 5914
rect 8116 5850 8168 5856
rect 7748 5772 7800 5778
rect 7748 5714 7800 5720
rect 7760 5166 7788 5714
rect 8128 5234 8156 5850
rect 8588 5710 8616 6802
rect 8864 6798 8892 7278
rect 8852 6792 8904 6798
rect 8852 6734 8904 6740
rect 8668 6724 8720 6730
rect 8668 6666 8720 6672
rect 8760 6724 8812 6730
rect 8760 6666 8812 6672
rect 8680 6322 8708 6666
rect 8668 6316 8720 6322
rect 8668 6258 8720 6264
rect 8772 5846 8800 6666
rect 8760 5840 8812 5846
rect 8760 5782 8812 5788
rect 8576 5704 8628 5710
rect 8576 5646 8628 5652
rect 8576 5568 8628 5574
rect 8576 5510 8628 5516
rect 8214 5468 8522 5477
rect 8214 5466 8220 5468
rect 8276 5466 8300 5468
rect 8356 5466 8380 5468
rect 8436 5466 8460 5468
rect 8516 5466 8522 5468
rect 8276 5414 8278 5466
rect 8458 5414 8460 5466
rect 8214 5412 8220 5414
rect 8276 5412 8300 5414
rect 8356 5412 8380 5414
rect 8436 5412 8460 5414
rect 8516 5412 8522 5414
rect 8214 5403 8522 5412
rect 8588 5370 8616 5510
rect 8576 5364 8628 5370
rect 8576 5306 8628 5312
rect 8116 5228 8168 5234
rect 8116 5170 8168 5176
rect 7748 5160 7800 5166
rect 7748 5102 7800 5108
rect 7104 5092 7156 5098
rect 7104 5034 7156 5040
rect 6880 4644 6960 4672
rect 6828 4626 6880 4632
rect 6736 4616 6788 4622
rect 6736 4558 6788 4564
rect 6644 4276 6696 4282
rect 6644 4218 6696 4224
rect 6644 4140 6696 4146
rect 6748 4128 6776 4558
rect 6696 4100 6776 4128
rect 6644 4082 6696 4088
rect 6748 3738 6776 4100
rect 6840 4010 6868 4626
rect 6828 4004 6880 4010
rect 6828 3946 6880 3952
rect 6736 3732 6788 3738
rect 6736 3674 6788 3680
rect 6460 3596 6512 3602
rect 6460 3538 6512 3544
rect 6276 2984 6328 2990
rect 6276 2926 6328 2932
rect 6184 2848 6236 2854
rect 6184 2790 6236 2796
rect 5356 2440 5408 2446
rect 5356 2382 5408 2388
rect 5448 2440 5500 2446
rect 5448 2382 5500 2388
rect 5368 2106 5396 2382
rect 5356 2100 5408 2106
rect 5356 2042 5408 2048
rect 4896 1420 4948 1426
rect 4896 1362 4948 1368
rect 5368 1358 5396 2042
rect 4252 1352 4304 1358
rect 4252 1294 4304 1300
rect 4436 1352 4488 1358
rect 4436 1294 4488 1300
rect 4620 1352 4672 1358
rect 4620 1294 4672 1300
rect 5356 1352 5408 1358
rect 5356 1294 5408 1300
rect 4528 1284 4580 1290
rect 4528 1226 4580 1232
rect 4540 1170 4568 1226
rect 5460 1222 5488 2382
rect 5908 2372 5960 2378
rect 5908 2314 5960 2320
rect 5632 2304 5684 2310
rect 5632 2246 5684 2252
rect 5644 1358 5672 2246
rect 5920 1426 5948 2314
rect 6288 2310 6316 2926
rect 6368 2372 6420 2378
rect 6368 2314 6420 2320
rect 6276 2304 6328 2310
rect 6276 2246 6328 2252
rect 6380 2106 6408 2314
rect 6472 2106 6500 3538
rect 6552 3052 6604 3058
rect 6552 2994 6604 3000
rect 6564 2922 6592 2994
rect 6552 2916 6604 2922
rect 6552 2858 6604 2864
rect 6368 2100 6420 2106
rect 6368 2042 6420 2048
rect 6460 2100 6512 2106
rect 6460 2042 6512 2048
rect 6564 1766 6592 2858
rect 6748 1970 6776 3674
rect 6840 3602 6868 3946
rect 6828 3596 6880 3602
rect 6828 3538 6880 3544
rect 6920 3392 6972 3398
rect 6920 3334 6972 3340
rect 6932 3194 6960 3334
rect 6920 3188 6972 3194
rect 6920 3130 6972 3136
rect 6932 2990 6960 3130
rect 7116 3058 7144 5034
rect 7656 5024 7708 5030
rect 7656 4966 7708 4972
rect 7668 4690 7696 4966
rect 7760 4690 7788 5102
rect 8588 4826 8616 5306
rect 9048 5234 9076 7822
rect 9036 5228 9088 5234
rect 9036 5170 9088 5176
rect 8668 5160 8720 5166
rect 8668 5102 8720 5108
rect 8576 4820 8628 4826
rect 8576 4762 8628 4768
rect 7656 4684 7708 4690
rect 7656 4626 7708 4632
rect 7748 4684 7800 4690
rect 7748 4626 7800 4632
rect 7196 4548 7248 4554
rect 7196 4490 7248 4496
rect 7208 4078 7236 4490
rect 8214 4380 8522 4389
rect 8214 4378 8220 4380
rect 8276 4378 8300 4380
rect 8356 4378 8380 4380
rect 8436 4378 8460 4380
rect 8516 4378 8522 4380
rect 8276 4326 8278 4378
rect 8458 4326 8460 4378
rect 8214 4324 8220 4326
rect 8276 4324 8300 4326
rect 8356 4324 8380 4326
rect 8436 4324 8460 4326
rect 8516 4324 8522 4326
rect 8214 4315 8522 4324
rect 8588 4282 8616 4762
rect 8576 4276 8628 4282
rect 8576 4218 8628 4224
rect 8484 4140 8536 4146
rect 8680 4128 8708 5102
rect 8536 4100 8708 4128
rect 8484 4082 8536 4088
rect 7196 4072 7248 4078
rect 7196 4014 7248 4020
rect 8022 4040 8078 4049
rect 8022 3975 8078 3984
rect 7104 3052 7156 3058
rect 7104 2994 7156 3000
rect 6920 2984 6972 2990
rect 6920 2926 6972 2932
rect 7116 2394 7144 2994
rect 7840 2916 7892 2922
rect 7840 2858 7892 2864
rect 7852 2446 7880 2858
rect 8036 2854 8064 3975
rect 8496 3602 8524 4082
rect 9048 3942 9076 5170
rect 9140 4622 9168 8774
rect 9232 8362 9260 9658
rect 9324 9518 9352 9823
rect 9312 9512 9364 9518
rect 9312 9454 9364 9460
rect 9404 9376 9456 9382
rect 9508 9364 9536 9862
rect 9678 9752 9734 9761
rect 9784 9722 9812 9930
rect 9678 9687 9734 9696
rect 9772 9716 9824 9722
rect 9692 9602 9720 9687
rect 9772 9658 9824 9664
rect 9456 9336 9536 9364
rect 9600 9574 9720 9602
rect 9404 9318 9456 9324
rect 9416 9110 9444 9318
rect 9494 9208 9550 9217
rect 9494 9143 9550 9152
rect 9404 9104 9456 9110
rect 9404 9046 9456 9052
rect 9312 9036 9364 9042
rect 9312 8978 9364 8984
rect 9324 8634 9352 8978
rect 9508 8634 9536 9143
rect 9600 9042 9628 9574
rect 9680 9512 9732 9518
rect 9680 9454 9732 9460
rect 9692 9178 9720 9454
rect 9680 9172 9732 9178
rect 9680 9114 9732 9120
rect 9784 9110 9812 9658
rect 9864 9648 9916 9654
rect 9864 9590 9916 9596
rect 9876 9450 9904 9590
rect 9968 9518 9996 10406
rect 9956 9512 10008 9518
rect 9956 9454 10008 9460
rect 9864 9444 9916 9450
rect 9864 9386 9916 9392
rect 9772 9104 9824 9110
rect 9772 9046 9824 9052
rect 9588 9036 9640 9042
rect 9588 8978 9640 8984
rect 9600 8634 9628 8978
rect 9312 8628 9364 8634
rect 9312 8570 9364 8576
rect 9496 8628 9548 8634
rect 9496 8570 9548 8576
rect 9588 8628 9640 8634
rect 9588 8570 9640 8576
rect 9876 8498 9904 9386
rect 9968 9178 9996 9454
rect 10060 9450 10088 11086
rect 10244 10985 10272 12854
rect 10428 12850 10456 13126
rect 10508 12980 10560 12986
rect 10508 12922 10560 12928
rect 10416 12844 10468 12850
rect 10416 12786 10468 12792
rect 10428 12238 10456 12786
rect 10416 12232 10468 12238
rect 10416 12174 10468 12180
rect 10428 11665 10456 12174
rect 10414 11656 10470 11665
rect 10414 11591 10470 11600
rect 10324 11144 10376 11150
rect 10324 11086 10376 11092
rect 10230 10976 10286 10985
rect 10230 10911 10286 10920
rect 10336 10810 10364 11086
rect 10520 11082 10548 12922
rect 10612 12782 10640 13262
rect 10888 12918 10916 14200
rect 11244 13864 11296 13870
rect 11244 13806 11296 13812
rect 10876 12912 10928 12918
rect 10876 12854 10928 12860
rect 10600 12776 10652 12782
rect 10600 12718 10652 12724
rect 11256 12646 11284 13806
rect 12084 13410 12112 14200
rect 12214 13628 12522 13637
rect 12214 13626 12220 13628
rect 12276 13626 12300 13628
rect 12356 13626 12380 13628
rect 12436 13626 12460 13628
rect 12516 13626 12522 13628
rect 12276 13574 12278 13626
rect 12458 13574 12460 13626
rect 12214 13572 12220 13574
rect 12276 13572 12300 13574
rect 12356 13572 12380 13574
rect 12436 13572 12460 13574
rect 12516 13572 12522 13574
rect 12214 13563 12522 13572
rect 11888 13388 11940 13394
rect 11888 13330 11940 13336
rect 11992 13382 12112 13410
rect 11612 13252 11664 13258
rect 11612 13194 11664 13200
rect 11244 12640 11296 12646
rect 11244 12582 11296 12588
rect 10692 12436 10744 12442
rect 10692 12378 10744 12384
rect 10704 12306 10732 12378
rect 10692 12300 10744 12306
rect 10692 12242 10744 12248
rect 11336 12300 11388 12306
rect 11336 12242 11388 12248
rect 10704 12186 10732 12242
rect 10612 12158 10732 12186
rect 10876 12232 10928 12238
rect 10876 12174 10928 12180
rect 11244 12232 11296 12238
rect 11244 12174 11296 12180
rect 10612 11830 10640 12158
rect 10692 12096 10744 12102
rect 10692 12038 10744 12044
rect 10704 11830 10732 12038
rect 10784 11892 10836 11898
rect 10784 11834 10836 11840
rect 10600 11824 10652 11830
rect 10600 11766 10652 11772
rect 10692 11824 10744 11830
rect 10692 11766 10744 11772
rect 10692 11552 10744 11558
rect 10692 11494 10744 11500
rect 10704 11286 10732 11494
rect 10692 11280 10744 11286
rect 10692 11222 10744 11228
rect 10600 11144 10652 11150
rect 10598 11112 10600 11121
rect 10652 11112 10654 11121
rect 10508 11076 10560 11082
rect 10598 11047 10654 11056
rect 10508 11018 10560 11024
rect 10324 10804 10376 10810
rect 10324 10746 10376 10752
rect 10322 10432 10378 10441
rect 10322 10367 10378 10376
rect 10336 9994 10364 10367
rect 10416 10124 10468 10130
rect 10416 10066 10468 10072
rect 10140 9988 10192 9994
rect 10140 9930 10192 9936
rect 10324 9988 10376 9994
rect 10324 9930 10376 9936
rect 10152 9722 10180 9930
rect 10336 9761 10364 9930
rect 10322 9752 10378 9761
rect 10140 9716 10192 9722
rect 10322 9687 10378 9696
rect 10140 9658 10192 9664
rect 10048 9444 10100 9450
rect 10048 9386 10100 9392
rect 9956 9172 10008 9178
rect 9956 9114 10008 9120
rect 9968 8566 9996 9114
rect 10060 9042 10088 9386
rect 10152 9382 10180 9658
rect 10428 9586 10456 10066
rect 10416 9580 10468 9586
rect 10416 9522 10468 9528
rect 10232 9512 10284 9518
rect 10230 9480 10232 9489
rect 10284 9480 10286 9489
rect 10230 9415 10286 9424
rect 10140 9376 10192 9382
rect 10428 9353 10456 9522
rect 10520 9466 10548 11018
rect 10612 10588 10640 11047
rect 10692 11008 10744 11014
rect 10692 10950 10744 10956
rect 10704 10742 10732 10950
rect 10692 10736 10744 10742
rect 10692 10678 10744 10684
rect 10612 10560 10732 10588
rect 10600 10464 10652 10470
rect 10600 10406 10652 10412
rect 10612 10062 10640 10406
rect 10704 10282 10732 10560
rect 10796 10452 10824 11834
rect 10888 11558 10916 12174
rect 10966 11928 11022 11937
rect 10966 11863 11022 11872
rect 10876 11552 10928 11558
rect 10876 11494 10928 11500
rect 10980 11082 11008 11863
rect 11152 11756 11204 11762
rect 11152 11698 11204 11704
rect 11060 11552 11112 11558
rect 11060 11494 11112 11500
rect 11072 11218 11100 11494
rect 11060 11212 11112 11218
rect 11060 11154 11112 11160
rect 10968 11076 11020 11082
rect 10968 11018 11020 11024
rect 11058 10568 11114 10577
rect 11058 10503 11114 10512
rect 10876 10464 10928 10470
rect 10796 10424 10876 10452
rect 10876 10406 10928 10412
rect 10704 10254 10824 10282
rect 10692 10124 10744 10130
rect 10692 10066 10744 10072
rect 10600 10056 10652 10062
rect 10600 9998 10652 10004
rect 10612 9926 10640 9998
rect 10600 9920 10652 9926
rect 10600 9862 10652 9868
rect 10704 9654 10732 10066
rect 10796 10062 10824 10254
rect 10784 10056 10836 10062
rect 10784 9998 10836 10004
rect 10796 9722 10824 9998
rect 10784 9716 10836 9722
rect 10784 9658 10836 9664
rect 10692 9648 10744 9654
rect 10692 9590 10744 9596
rect 10520 9438 10732 9466
rect 10140 9318 10192 9324
rect 10414 9344 10470 9353
rect 10414 9279 10470 9288
rect 10048 9036 10100 9042
rect 10048 8978 10100 8984
rect 9956 8560 10008 8566
rect 9956 8502 10008 8508
rect 9864 8492 9916 8498
rect 9864 8434 9916 8440
rect 9496 8424 9548 8430
rect 9496 8366 9548 8372
rect 9220 8356 9272 8362
rect 9220 8298 9272 8304
rect 9508 7886 9536 8366
rect 9680 8288 9732 8294
rect 9680 8230 9732 8236
rect 9692 7954 9720 8230
rect 9680 7948 9732 7954
rect 9680 7890 9732 7896
rect 9968 7886 9996 8502
rect 10060 8430 10088 8978
rect 10140 8968 10192 8974
rect 10140 8910 10192 8916
rect 10230 8936 10286 8945
rect 10048 8424 10100 8430
rect 10048 8366 10100 8372
rect 9496 7880 9548 7886
rect 9496 7822 9548 7828
rect 9956 7880 10008 7886
rect 9956 7822 10008 7828
rect 10152 7834 10180 8910
rect 10230 8871 10232 8880
rect 10284 8871 10286 8880
rect 10232 8842 10284 8848
rect 10428 8498 10456 9279
rect 10704 8922 10732 9438
rect 10888 9042 10916 10406
rect 10968 10260 11020 10266
rect 10968 10202 11020 10208
rect 10980 10044 11008 10202
rect 11072 10198 11100 10503
rect 11164 10452 11192 11698
rect 11256 11354 11284 12174
rect 11348 11694 11376 12242
rect 11624 12238 11652 13194
rect 11900 12918 11928 13330
rect 11888 12912 11940 12918
rect 11888 12854 11940 12860
rect 11796 12776 11848 12782
rect 11796 12718 11848 12724
rect 11612 12232 11664 12238
rect 11612 12174 11664 12180
rect 11428 12096 11480 12102
rect 11428 12038 11480 12044
rect 11336 11688 11388 11694
rect 11336 11630 11388 11636
rect 11244 11348 11296 11354
rect 11244 11290 11296 11296
rect 11348 11014 11376 11630
rect 11336 11008 11388 11014
rect 11336 10950 11388 10956
rect 11334 10704 11390 10713
rect 11334 10639 11336 10648
rect 11388 10639 11390 10648
rect 11336 10610 11388 10616
rect 11244 10600 11296 10606
rect 11334 10568 11390 10577
rect 11296 10548 11334 10554
rect 11244 10542 11334 10548
rect 11256 10526 11334 10542
rect 11334 10503 11390 10512
rect 11164 10424 11284 10452
rect 11060 10192 11112 10198
rect 11060 10134 11112 10140
rect 11060 10056 11112 10062
rect 10980 10016 11060 10044
rect 11060 9998 11112 10004
rect 11152 10056 11204 10062
rect 11152 9998 11204 10004
rect 11164 9897 11192 9998
rect 11256 9994 11284 10424
rect 11244 9988 11296 9994
rect 11244 9930 11296 9936
rect 11150 9888 11206 9897
rect 11150 9823 11206 9832
rect 11058 9616 11114 9625
rect 11164 9586 11192 9823
rect 11244 9716 11296 9722
rect 11244 9658 11296 9664
rect 11058 9551 11114 9560
rect 11152 9580 11204 9586
rect 10876 9036 10928 9042
rect 10876 8978 10928 8984
rect 10704 8906 10916 8922
rect 10704 8900 10928 8906
rect 10704 8894 10876 8900
rect 10876 8842 10928 8848
rect 10692 8832 10744 8838
rect 10692 8774 10744 8780
rect 10416 8492 10468 8498
rect 10416 8434 10468 8440
rect 10232 8424 10284 8430
rect 10232 8366 10284 8372
rect 10244 8022 10272 8366
rect 10232 8016 10284 8022
rect 10232 7958 10284 7964
rect 10152 7806 10272 7834
rect 10140 7744 10192 7750
rect 10140 7686 10192 7692
rect 9680 6928 9732 6934
rect 9680 6870 9732 6876
rect 9312 6656 9364 6662
rect 9312 6598 9364 6604
rect 9324 5710 9352 6598
rect 9692 6390 9720 6870
rect 10048 6792 10100 6798
rect 10048 6734 10100 6740
rect 9680 6384 9732 6390
rect 9680 6326 9732 6332
rect 9692 5710 9720 6326
rect 9772 6112 9824 6118
rect 9772 6054 9824 6060
rect 9312 5704 9364 5710
rect 9312 5646 9364 5652
rect 9680 5704 9732 5710
rect 9680 5646 9732 5652
rect 9404 5636 9456 5642
rect 9404 5578 9456 5584
rect 9416 4826 9444 5578
rect 9680 5568 9732 5574
rect 9680 5510 9732 5516
rect 9404 4820 9456 4826
rect 9404 4762 9456 4768
rect 9128 4616 9180 4622
rect 9128 4558 9180 4564
rect 9416 4214 9444 4762
rect 9692 4758 9720 5510
rect 9784 5166 9812 6054
rect 10060 5778 10088 6734
rect 10048 5772 10100 5778
rect 10048 5714 10100 5720
rect 9864 5704 9916 5710
rect 9864 5646 9916 5652
rect 9772 5160 9824 5166
rect 9772 5102 9824 5108
rect 9876 5030 9904 5646
rect 10060 5302 10088 5714
rect 10152 5574 10180 7686
rect 10244 7410 10272 7806
rect 10232 7404 10284 7410
rect 10232 7346 10284 7352
rect 10244 5710 10272 7346
rect 10428 6458 10456 8434
rect 10600 8424 10652 8430
rect 10600 8366 10652 8372
rect 10508 7336 10560 7342
rect 10508 7278 10560 7284
rect 10416 6452 10468 6458
rect 10416 6394 10468 6400
rect 10324 5908 10376 5914
rect 10324 5850 10376 5856
rect 10232 5704 10284 5710
rect 10232 5646 10284 5652
rect 10140 5568 10192 5574
rect 10140 5510 10192 5516
rect 10048 5296 10100 5302
rect 10048 5238 10100 5244
rect 9864 5024 9916 5030
rect 9864 4966 9916 4972
rect 9680 4752 9732 4758
rect 9680 4694 9732 4700
rect 9680 4480 9732 4486
rect 9680 4422 9732 4428
rect 9692 4282 9720 4422
rect 9876 4282 9904 4966
rect 10060 4690 10088 5238
rect 10244 4826 10272 5646
rect 10232 4820 10284 4826
rect 10232 4762 10284 4768
rect 10048 4684 10100 4690
rect 10048 4626 10100 4632
rect 9680 4276 9732 4282
rect 9680 4218 9732 4224
rect 9864 4276 9916 4282
rect 9864 4218 9916 4224
rect 9404 4208 9456 4214
rect 9404 4150 9456 4156
rect 10336 4146 10364 5850
rect 10428 5030 10456 6394
rect 10520 6254 10548 7278
rect 10508 6248 10560 6254
rect 10508 6190 10560 6196
rect 10612 5778 10640 8366
rect 10704 7970 10732 8774
rect 10704 7942 10824 7970
rect 10692 7880 10744 7886
rect 10692 7822 10744 7828
rect 10704 7546 10732 7822
rect 10692 7540 10744 7546
rect 10692 7482 10744 7488
rect 10796 6322 10824 7942
rect 11072 7886 11100 9551
rect 11152 9522 11204 9528
rect 11256 9178 11284 9658
rect 11348 9382 11376 10503
rect 11440 9450 11468 12038
rect 11808 11880 11836 12718
rect 11900 12238 11928 12854
rect 11992 12442 12020 13382
rect 12072 13320 12124 13326
rect 12072 13262 12124 13268
rect 12164 13320 12216 13326
rect 12164 13262 12216 13268
rect 12992 13320 13044 13326
rect 12992 13262 13044 13268
rect 13176 13320 13228 13326
rect 13176 13262 13228 13268
rect 11980 12436 12032 12442
rect 11980 12378 12032 12384
rect 11888 12232 11940 12238
rect 11888 12174 11940 12180
rect 12084 12170 12112 13262
rect 12176 12850 12204 13262
rect 12624 13252 12676 13258
rect 12624 13194 12676 13200
rect 12636 12918 12664 13194
rect 12900 13184 12952 13190
rect 12900 13126 12952 13132
rect 12624 12912 12676 12918
rect 12624 12854 12676 12860
rect 12164 12844 12216 12850
rect 12164 12786 12216 12792
rect 12214 12540 12522 12549
rect 12214 12538 12220 12540
rect 12276 12538 12300 12540
rect 12356 12538 12380 12540
rect 12436 12538 12460 12540
rect 12516 12538 12522 12540
rect 12276 12486 12278 12538
rect 12458 12486 12460 12538
rect 12214 12484 12220 12486
rect 12276 12484 12300 12486
rect 12356 12484 12380 12486
rect 12436 12484 12460 12486
rect 12516 12484 12522 12486
rect 12214 12475 12522 12484
rect 12808 12232 12860 12238
rect 12808 12174 12860 12180
rect 12072 12164 12124 12170
rect 12072 12106 12124 12112
rect 11980 11892 12032 11898
rect 11808 11852 11980 11880
rect 11980 11834 12032 11840
rect 11704 11756 11756 11762
rect 11704 11698 11756 11704
rect 11518 11248 11574 11257
rect 11518 11183 11574 11192
rect 11428 9444 11480 9450
rect 11428 9386 11480 9392
rect 11336 9376 11388 9382
rect 11388 9324 11468 9330
rect 11336 9318 11468 9324
rect 11348 9302 11468 9318
rect 11244 9172 11296 9178
rect 11244 9114 11296 9120
rect 11256 9058 11284 9114
rect 11164 9030 11284 9058
rect 11164 8634 11192 9030
rect 11336 8968 11388 8974
rect 11256 8928 11336 8956
rect 11152 8628 11204 8634
rect 11152 8570 11204 8576
rect 10876 7880 10928 7886
rect 10876 7822 10928 7828
rect 11060 7880 11112 7886
rect 11060 7822 11112 7828
rect 10888 6458 10916 7822
rect 11072 7410 11100 7822
rect 11060 7404 11112 7410
rect 11060 7346 11112 7352
rect 10876 6452 10928 6458
rect 10876 6394 10928 6400
rect 10692 6316 10744 6322
rect 10692 6258 10744 6264
rect 10784 6316 10836 6322
rect 10784 6258 10836 6264
rect 10704 5914 10732 6258
rect 11164 6254 11192 8570
rect 11256 8430 11284 8928
rect 11336 8910 11388 8916
rect 11336 8832 11388 8838
rect 11440 8786 11468 9302
rect 11388 8780 11468 8786
rect 11336 8774 11468 8780
rect 11348 8758 11468 8774
rect 11244 8424 11296 8430
rect 11244 8366 11296 8372
rect 11152 6248 11204 6254
rect 11152 6190 11204 6196
rect 10692 5908 10744 5914
rect 10692 5850 10744 5856
rect 10600 5772 10652 5778
rect 10600 5714 10652 5720
rect 11152 5296 11204 5302
rect 11152 5238 11204 5244
rect 10416 5024 10468 5030
rect 10416 4966 10468 4972
rect 11164 4282 11192 5238
rect 11152 4276 11204 4282
rect 11152 4218 11204 4224
rect 9588 4140 9640 4146
rect 9588 4082 9640 4088
rect 10324 4140 10376 4146
rect 10324 4082 10376 4088
rect 10784 4140 10836 4146
rect 10784 4082 10836 4088
rect 9220 4004 9272 4010
rect 9220 3946 9272 3952
rect 9036 3936 9088 3942
rect 9036 3878 9088 3884
rect 8864 3602 9168 3618
rect 8484 3596 8536 3602
rect 8484 3538 8536 3544
rect 8852 3596 9180 3602
rect 8904 3590 9128 3596
rect 8852 3538 8904 3544
rect 9128 3538 9180 3544
rect 8208 3460 8260 3466
rect 8128 3420 8208 3448
rect 8128 3194 8156 3420
rect 8496 3448 8524 3538
rect 9232 3534 9260 3946
rect 9600 3738 9628 4082
rect 9956 4004 10008 4010
rect 9956 3946 10008 3952
rect 9588 3732 9640 3738
rect 9588 3674 9640 3680
rect 9680 3732 9732 3738
rect 9680 3674 9732 3680
rect 9220 3528 9272 3534
rect 9220 3470 9272 3476
rect 9496 3528 9548 3534
rect 9496 3470 9548 3476
rect 8496 3420 8616 3448
rect 8208 3402 8260 3408
rect 8214 3292 8522 3301
rect 8214 3290 8220 3292
rect 8276 3290 8300 3292
rect 8356 3290 8380 3292
rect 8436 3290 8460 3292
rect 8516 3290 8522 3292
rect 8276 3238 8278 3290
rect 8458 3238 8460 3290
rect 8214 3236 8220 3238
rect 8276 3236 8300 3238
rect 8356 3236 8380 3238
rect 8436 3236 8460 3238
rect 8516 3236 8522 3238
rect 8214 3227 8522 3236
rect 8116 3188 8168 3194
rect 8116 3130 8168 3136
rect 8588 3126 8616 3420
rect 8576 3120 8628 3126
rect 8576 3062 8628 3068
rect 8024 2848 8076 2854
rect 8024 2790 8076 2796
rect 8588 2514 8616 3062
rect 8944 2984 8996 2990
rect 8944 2926 8996 2932
rect 8956 2650 8984 2926
rect 8944 2644 8996 2650
rect 8944 2586 8996 2592
rect 8576 2508 8628 2514
rect 8576 2450 8628 2456
rect 7564 2440 7616 2446
rect 7116 2378 7236 2394
rect 7564 2382 7616 2388
rect 7840 2440 7892 2446
rect 7840 2382 7892 2388
rect 7116 2372 7248 2378
rect 7116 2366 7196 2372
rect 6736 1964 6788 1970
rect 6736 1906 6788 1912
rect 6552 1760 6604 1766
rect 6552 1702 6604 1708
rect 6748 1562 6776 1906
rect 7012 1760 7064 1766
rect 7012 1702 7064 1708
rect 6736 1556 6788 1562
rect 6736 1498 6788 1504
rect 6748 1426 6776 1498
rect 5908 1420 5960 1426
rect 5908 1362 5960 1368
rect 6736 1420 6788 1426
rect 6736 1362 6788 1368
rect 7024 1358 7052 1702
rect 5632 1352 5684 1358
rect 5632 1294 5684 1300
rect 7012 1352 7064 1358
rect 7012 1294 7064 1300
rect 7116 1290 7144 2366
rect 7196 2314 7248 2320
rect 7288 2304 7340 2310
rect 7288 2246 7340 2252
rect 7300 1426 7328 2246
rect 7576 1426 7604 2382
rect 8116 2304 8168 2310
rect 8116 2246 8168 2252
rect 8128 2038 8156 2246
rect 8214 2204 8522 2213
rect 8214 2202 8220 2204
rect 8276 2202 8300 2204
rect 8356 2202 8380 2204
rect 8436 2202 8460 2204
rect 8516 2202 8522 2204
rect 8276 2150 8278 2202
rect 8458 2150 8460 2202
rect 8214 2148 8220 2150
rect 8276 2148 8300 2150
rect 8356 2148 8380 2150
rect 8436 2148 8460 2150
rect 8516 2148 8522 2150
rect 8214 2139 8522 2148
rect 7932 2032 7984 2038
rect 7932 1974 7984 1980
rect 8116 2032 8168 2038
rect 8116 1974 8168 1980
rect 7944 1426 7972 1974
rect 8588 1902 8616 2450
rect 9128 2372 9180 2378
rect 9128 2314 9180 2320
rect 8668 2304 8720 2310
rect 8668 2246 8720 2252
rect 8680 2106 8708 2246
rect 8668 2100 8720 2106
rect 8668 2042 8720 2048
rect 8576 1896 8628 1902
rect 8576 1838 8628 1844
rect 8588 1426 8616 1838
rect 8680 1562 8708 2042
rect 8944 1896 8996 1902
rect 8944 1838 8996 1844
rect 8668 1556 8720 1562
rect 8668 1498 8720 1504
rect 8956 1494 8984 1838
rect 8944 1488 8996 1494
rect 8944 1430 8996 1436
rect 7288 1420 7340 1426
rect 7288 1362 7340 1368
rect 7564 1420 7616 1426
rect 7564 1362 7616 1368
rect 7932 1420 7984 1426
rect 7932 1362 7984 1368
rect 8576 1420 8628 1426
rect 8576 1362 8628 1368
rect 9140 1358 9168 2314
rect 9508 2310 9536 3470
rect 9588 3392 9640 3398
rect 9588 3334 9640 3340
rect 9600 2514 9628 3334
rect 9588 2508 9640 2514
rect 9588 2450 9640 2456
rect 9496 2304 9548 2310
rect 9496 2246 9548 2252
rect 9508 1902 9536 2246
rect 9496 1896 9548 1902
rect 9496 1838 9548 1844
rect 9128 1352 9180 1358
rect 9600 1306 9628 2450
rect 9692 2378 9720 3674
rect 9968 3618 9996 3946
rect 10324 3936 10376 3942
rect 10324 3878 10376 3884
rect 9968 3590 10088 3618
rect 10336 3602 10364 3878
rect 10796 3738 10824 4082
rect 10784 3732 10836 3738
rect 10784 3674 10836 3680
rect 9864 3460 9916 3466
rect 9916 3420 9996 3448
rect 9864 3402 9916 3408
rect 9864 3120 9916 3126
rect 9864 3062 9916 3068
rect 9772 2984 9824 2990
rect 9772 2926 9824 2932
rect 9784 2446 9812 2926
rect 9876 2582 9904 3062
rect 9864 2576 9916 2582
rect 9864 2518 9916 2524
rect 9968 2446 9996 3420
rect 10060 2990 10088 3590
rect 10324 3596 10376 3602
rect 10324 3538 10376 3544
rect 10600 3460 10652 3466
rect 10600 3402 10652 3408
rect 10612 3194 10640 3402
rect 10600 3188 10652 3194
rect 10600 3130 10652 3136
rect 11060 3188 11112 3194
rect 11060 3130 11112 3136
rect 10048 2984 10100 2990
rect 10048 2926 10100 2932
rect 10600 2848 10652 2854
rect 10600 2790 10652 2796
rect 9772 2440 9824 2446
rect 9772 2382 9824 2388
rect 9956 2440 10008 2446
rect 10008 2400 10180 2428
rect 9956 2382 10008 2388
rect 9680 2372 9732 2378
rect 9680 2314 9732 2320
rect 9692 2106 9720 2314
rect 9680 2100 9732 2106
rect 9680 2042 9732 2048
rect 10152 1970 10180 2400
rect 10612 2378 10640 2790
rect 11072 2650 11100 3130
rect 11060 2644 11112 2650
rect 11060 2586 11112 2592
rect 10600 2372 10652 2378
rect 10600 2314 10652 2320
rect 10140 1964 10192 1970
rect 10140 1906 10192 1912
rect 11060 1828 11112 1834
rect 11060 1770 11112 1776
rect 9128 1294 9180 1300
rect 9508 1290 9628 1306
rect 11072 1290 11100 1770
rect 11152 1488 11204 1494
rect 11152 1430 11204 1436
rect 7104 1284 7156 1290
rect 7104 1226 7156 1232
rect 9496 1284 9628 1290
rect 9548 1278 9628 1284
rect 11060 1284 11112 1290
rect 9496 1226 9548 1232
rect 11060 1226 11112 1232
rect 4080 1142 4568 1170
rect 5448 1216 5500 1222
rect 5448 1158 5500 1164
rect 6368 1216 6420 1222
rect 6368 1158 6420 1164
rect 6380 1018 6408 1158
rect 8214 1116 8522 1125
rect 8214 1114 8220 1116
rect 8276 1114 8300 1116
rect 8356 1114 8380 1116
rect 8436 1114 8460 1116
rect 8516 1114 8522 1116
rect 8276 1062 8278 1114
rect 8458 1062 8460 1114
rect 8214 1060 8220 1062
rect 8276 1060 8300 1062
rect 8356 1060 8380 1062
rect 8436 1060 8460 1062
rect 8516 1060 8522 1062
rect 8214 1051 8522 1060
rect 3884 1012 3936 1018
rect 3884 954 3936 960
rect 6368 1012 6420 1018
rect 6368 954 6420 960
rect 11164 800 11192 1430
rect 11256 1329 11284 8366
rect 11440 5574 11468 8758
rect 11532 6746 11560 11183
rect 11716 10577 11744 11698
rect 11992 11354 12020 11834
rect 12820 11694 12848 12174
rect 12912 11830 12940 13126
rect 13004 12714 13032 13262
rect 13084 13184 13136 13190
rect 13084 13126 13136 13132
rect 12992 12708 13044 12714
rect 12992 12650 13044 12656
rect 13004 12238 13032 12650
rect 12992 12232 13044 12238
rect 12992 12174 13044 12180
rect 12900 11824 12952 11830
rect 12900 11766 12952 11772
rect 12072 11688 12124 11694
rect 12072 11630 12124 11636
rect 12808 11688 12860 11694
rect 12808 11630 12860 11636
rect 11980 11348 12032 11354
rect 11980 11290 12032 11296
rect 11796 11280 11848 11286
rect 11796 11222 11848 11228
rect 11808 10674 11836 11222
rect 11992 11121 12020 11290
rect 12084 11150 12112 11630
rect 12214 11452 12522 11461
rect 12214 11450 12220 11452
rect 12276 11450 12300 11452
rect 12356 11450 12380 11452
rect 12436 11450 12460 11452
rect 12516 11450 12522 11452
rect 12276 11398 12278 11450
rect 12458 11398 12460 11450
rect 12214 11396 12220 11398
rect 12276 11396 12300 11398
rect 12356 11396 12380 11398
rect 12436 11396 12460 11398
rect 12516 11396 12522 11398
rect 12214 11387 12522 11396
rect 13004 11150 13032 12174
rect 13096 11762 13124 13126
rect 13188 11898 13216 13262
rect 13360 13252 13412 13258
rect 13360 13194 13412 13200
rect 13268 12164 13320 12170
rect 13268 12106 13320 12112
rect 13176 11892 13228 11898
rect 13176 11834 13228 11840
rect 13280 11762 13308 12106
rect 13372 11830 13400 13194
rect 13464 11898 13492 14334
rect 14370 14200 14426 15000
rect 14384 13530 14412 14200
rect 14372 13524 14424 13530
rect 14372 13466 14424 13472
rect 13452 11892 13504 11898
rect 13452 11834 13504 11840
rect 13360 11824 13412 11830
rect 13360 11766 13412 11772
rect 13084 11756 13136 11762
rect 13084 11698 13136 11704
rect 13268 11756 13320 11762
rect 13268 11698 13320 11704
rect 12072 11144 12124 11150
rect 11978 11112 12034 11121
rect 12072 11086 12124 11092
rect 12992 11144 13044 11150
rect 12992 11086 13044 11092
rect 13096 11082 13124 11698
rect 13280 11150 13308 11698
rect 13464 11286 13492 11834
rect 13452 11280 13504 11286
rect 13452 11222 13504 11228
rect 13542 11248 13598 11257
rect 13542 11183 13544 11192
rect 13596 11183 13598 11192
rect 13544 11154 13596 11160
rect 13268 11144 13320 11150
rect 13268 11086 13320 11092
rect 11978 11047 11980 11056
rect 12032 11047 12034 11056
rect 12256 11076 12308 11082
rect 11980 11018 12032 11024
rect 12256 11018 12308 11024
rect 13084 11076 13136 11082
rect 13084 11018 13136 11024
rect 11992 10987 12020 11018
rect 12268 10742 12296 11018
rect 12532 11008 12584 11014
rect 12532 10950 12584 10956
rect 12716 11008 12768 11014
rect 12716 10950 12768 10956
rect 12256 10736 12308 10742
rect 11900 10674 12204 10690
rect 12256 10678 12308 10684
rect 11796 10668 11848 10674
rect 11796 10610 11848 10616
rect 11900 10668 12216 10674
rect 11900 10662 12164 10668
rect 11702 10568 11758 10577
rect 11702 10503 11758 10512
rect 11704 10464 11756 10470
rect 11704 10406 11756 10412
rect 11612 9512 11664 9518
rect 11612 9454 11664 9460
rect 11624 9110 11652 9454
rect 11612 9104 11664 9110
rect 11612 9046 11664 9052
rect 11624 8566 11652 9046
rect 11716 8634 11744 10406
rect 11796 10124 11848 10130
rect 11900 10112 11928 10662
rect 12164 10610 12216 10616
rect 12072 10600 12124 10606
rect 12072 10542 12124 10548
rect 12348 10600 12400 10606
rect 12348 10542 12400 10548
rect 11980 10464 12032 10470
rect 11980 10406 12032 10412
rect 11848 10084 11928 10112
rect 11796 10066 11848 10072
rect 11796 9988 11848 9994
rect 11796 9930 11848 9936
rect 11704 8628 11756 8634
rect 11704 8570 11756 8576
rect 11612 8560 11664 8566
rect 11612 8502 11664 8508
rect 11624 6866 11652 8502
rect 11612 6860 11664 6866
rect 11612 6802 11664 6808
rect 11704 6792 11756 6798
rect 11532 6740 11704 6746
rect 11532 6734 11756 6740
rect 11532 6718 11744 6734
rect 11612 6180 11664 6186
rect 11612 6122 11664 6128
rect 11624 5642 11652 6122
rect 11612 5636 11664 5642
rect 11612 5578 11664 5584
rect 11428 5568 11480 5574
rect 11428 5510 11480 5516
rect 11808 5370 11836 9930
rect 11900 8974 11928 10084
rect 11888 8968 11940 8974
rect 11888 8910 11940 8916
rect 11992 8634 12020 10406
rect 12084 9586 12112 10542
rect 12256 10464 12308 10470
rect 12360 10452 12388 10542
rect 12544 10520 12572 10950
rect 12622 10704 12678 10713
rect 12622 10639 12624 10648
rect 12676 10639 12678 10648
rect 12624 10610 12676 10616
rect 12544 10492 12664 10520
rect 12308 10424 12388 10452
rect 12256 10406 12308 10412
rect 12214 10364 12522 10373
rect 12214 10362 12220 10364
rect 12276 10362 12300 10364
rect 12356 10362 12380 10364
rect 12436 10362 12460 10364
rect 12516 10362 12522 10364
rect 12276 10310 12278 10362
rect 12458 10310 12460 10362
rect 12214 10308 12220 10310
rect 12276 10308 12300 10310
rect 12356 10308 12380 10310
rect 12436 10308 12460 10310
rect 12516 10308 12522 10310
rect 12214 10299 12522 10308
rect 12072 9580 12124 9586
rect 12072 9522 12124 9528
rect 12084 9178 12112 9522
rect 12214 9276 12522 9285
rect 12214 9274 12220 9276
rect 12276 9274 12300 9276
rect 12356 9274 12380 9276
rect 12436 9274 12460 9276
rect 12516 9274 12522 9276
rect 12276 9222 12278 9274
rect 12458 9222 12460 9274
rect 12214 9220 12220 9222
rect 12276 9220 12300 9222
rect 12356 9220 12380 9222
rect 12436 9220 12460 9222
rect 12516 9220 12522 9222
rect 12214 9211 12522 9220
rect 12072 9172 12124 9178
rect 12072 9114 12124 9120
rect 12348 9104 12400 9110
rect 12348 9046 12400 9052
rect 11980 8628 12032 8634
rect 11980 8570 12032 8576
rect 12360 8498 12388 9046
rect 12636 8809 12664 10492
rect 12728 10062 12756 10950
rect 12806 10704 12862 10713
rect 12806 10639 12862 10648
rect 12716 10056 12768 10062
rect 12716 9998 12768 10004
rect 12728 9586 12756 9998
rect 12820 9654 12848 10639
rect 12900 10600 12952 10606
rect 12900 10542 12952 10548
rect 12912 10198 12940 10542
rect 13360 10532 13412 10538
rect 13360 10474 13412 10480
rect 13372 10198 13400 10474
rect 12900 10192 12952 10198
rect 12900 10134 12952 10140
rect 13360 10192 13412 10198
rect 13360 10134 13412 10140
rect 13372 9654 13400 10134
rect 12808 9648 12860 9654
rect 12808 9590 12860 9596
rect 13360 9648 13412 9654
rect 13360 9590 13412 9596
rect 12716 9580 12768 9586
rect 12716 9522 12768 9528
rect 12622 8800 12678 8809
rect 12622 8735 12678 8744
rect 12728 8566 12756 9522
rect 13452 9444 13504 9450
rect 13452 9386 13504 9392
rect 13268 8968 13320 8974
rect 13268 8910 13320 8916
rect 12900 8900 12952 8906
rect 12900 8842 12952 8848
rect 13084 8900 13136 8906
rect 13084 8842 13136 8848
rect 12716 8560 12768 8566
rect 12716 8502 12768 8508
rect 12348 8492 12400 8498
rect 12348 8434 12400 8440
rect 12072 8356 12124 8362
rect 12072 8298 12124 8304
rect 11980 7812 12032 7818
rect 11980 7754 12032 7760
rect 11992 7324 12020 7754
rect 12084 7478 12112 8298
rect 12214 8188 12522 8197
rect 12214 8186 12220 8188
rect 12276 8186 12300 8188
rect 12356 8186 12380 8188
rect 12436 8186 12460 8188
rect 12516 8186 12522 8188
rect 12276 8134 12278 8186
rect 12458 8134 12460 8186
rect 12214 8132 12220 8134
rect 12276 8132 12300 8134
rect 12356 8132 12380 8134
rect 12436 8132 12460 8134
rect 12516 8132 12522 8134
rect 12214 8123 12522 8132
rect 12912 8090 12940 8842
rect 13096 8566 13124 8842
rect 13084 8560 13136 8566
rect 13084 8502 13136 8508
rect 13280 8498 13308 8910
rect 13268 8492 13320 8498
rect 13268 8434 13320 8440
rect 12900 8084 12952 8090
rect 12900 8026 12952 8032
rect 13280 7886 13308 8434
rect 13268 7880 13320 7886
rect 13268 7822 13320 7828
rect 12256 7744 12308 7750
rect 12256 7686 12308 7692
rect 12268 7546 12296 7686
rect 12256 7540 12308 7546
rect 12256 7482 12308 7488
rect 12072 7472 12124 7478
rect 12072 7414 12124 7420
rect 12268 7410 12296 7482
rect 12256 7404 12308 7410
rect 12256 7346 12308 7352
rect 12072 7336 12124 7342
rect 11992 7296 12072 7324
rect 12072 7278 12124 7284
rect 11888 6724 11940 6730
rect 11888 6666 11940 6672
rect 11900 6390 11928 6666
rect 12084 6458 12112 7278
rect 12214 7100 12522 7109
rect 12214 7098 12220 7100
rect 12276 7098 12300 7100
rect 12356 7098 12380 7100
rect 12436 7098 12460 7100
rect 12516 7098 12522 7100
rect 12276 7046 12278 7098
rect 12458 7046 12460 7098
rect 12214 7044 12220 7046
rect 12276 7044 12300 7046
rect 12356 7044 12380 7046
rect 12436 7044 12460 7046
rect 12516 7044 12522 7046
rect 12214 7035 12522 7044
rect 13280 6934 13308 7822
rect 13268 6928 13320 6934
rect 13268 6870 13320 6876
rect 12348 6792 12400 6798
rect 12348 6734 12400 6740
rect 12072 6452 12124 6458
rect 12072 6394 12124 6400
rect 11888 6384 11940 6390
rect 11888 6326 11940 6332
rect 12084 6322 12112 6394
rect 12360 6322 12388 6734
rect 13280 6390 13308 6870
rect 13464 6798 13492 9386
rect 13544 8084 13596 8090
rect 13544 8026 13596 8032
rect 13452 6792 13504 6798
rect 13452 6734 13504 6740
rect 13268 6384 13320 6390
rect 13268 6326 13320 6332
rect 12072 6316 12124 6322
rect 11992 6276 12072 6304
rect 11992 5710 12020 6276
rect 12072 6258 12124 6264
rect 12348 6316 12400 6322
rect 12348 6258 12400 6264
rect 13268 6248 13320 6254
rect 13268 6190 13320 6196
rect 12072 6112 12124 6118
rect 12072 6054 12124 6060
rect 11980 5704 12032 5710
rect 11980 5646 12032 5652
rect 12084 5658 12112 6054
rect 12214 6012 12522 6021
rect 12214 6010 12220 6012
rect 12276 6010 12300 6012
rect 12356 6010 12380 6012
rect 12436 6010 12460 6012
rect 12516 6010 12522 6012
rect 12276 5958 12278 6010
rect 12458 5958 12460 6010
rect 12214 5956 12220 5958
rect 12276 5956 12300 5958
rect 12356 5956 12380 5958
rect 12436 5956 12460 5958
rect 12516 5956 12522 5958
rect 12214 5947 12522 5956
rect 13280 5914 13308 6190
rect 13464 5930 13492 6734
rect 13556 6225 13584 8026
rect 13542 6216 13598 6225
rect 13542 6151 13598 6160
rect 13268 5908 13320 5914
rect 13464 5902 13584 5930
rect 13268 5850 13320 5856
rect 11888 5636 11940 5642
rect 11888 5578 11940 5584
rect 11796 5364 11848 5370
rect 11796 5306 11848 5312
rect 11612 5228 11664 5234
rect 11612 5170 11664 5176
rect 11624 4282 11652 5170
rect 11900 4554 11928 5578
rect 11888 4548 11940 4554
rect 11888 4490 11940 4496
rect 11992 4298 12020 5646
rect 12084 5630 12204 5658
rect 12084 5302 12112 5630
rect 12176 5574 12204 5630
rect 12164 5568 12216 5574
rect 12164 5510 12216 5516
rect 13176 5568 13228 5574
rect 13176 5510 13228 5516
rect 13188 5302 13216 5510
rect 12072 5296 12124 5302
rect 12072 5238 12124 5244
rect 13176 5296 13228 5302
rect 13176 5238 13228 5244
rect 12624 5228 12676 5234
rect 12624 5170 12676 5176
rect 12214 4924 12522 4933
rect 12214 4922 12220 4924
rect 12276 4922 12300 4924
rect 12356 4922 12380 4924
rect 12436 4922 12460 4924
rect 12516 4922 12522 4924
rect 12276 4870 12278 4922
rect 12458 4870 12460 4922
rect 12214 4868 12220 4870
rect 12276 4868 12300 4870
rect 12356 4868 12380 4870
rect 12436 4868 12460 4870
rect 12516 4868 12522 4870
rect 12214 4859 12522 4868
rect 12636 4706 12664 5170
rect 12716 5024 12768 5030
rect 12716 4966 12768 4972
rect 12544 4678 12664 4706
rect 12544 4622 12572 4678
rect 12532 4616 12584 4622
rect 12532 4558 12584 4564
rect 11612 4276 11664 4282
rect 11992 4270 12112 4298
rect 11612 4218 11664 4224
rect 11980 4208 12032 4214
rect 11980 4150 12032 4156
rect 11704 4072 11756 4078
rect 11704 4014 11756 4020
rect 11716 3466 11744 4014
rect 11992 3602 12020 4150
rect 12084 4146 12112 4270
rect 12544 4214 12572 4558
rect 12532 4208 12584 4214
rect 12532 4150 12584 4156
rect 12728 4146 12756 4966
rect 13188 4758 13216 5238
rect 13556 5234 13584 5902
rect 13544 5228 13596 5234
rect 13544 5170 13596 5176
rect 13176 4752 13228 4758
rect 13176 4694 13228 4700
rect 13556 4622 13584 5170
rect 13544 4616 13596 4622
rect 13544 4558 13596 4564
rect 12072 4140 12124 4146
rect 12072 4082 12124 4088
rect 12716 4140 12768 4146
rect 12716 4082 12768 4088
rect 13360 4140 13412 4146
rect 13360 4082 13412 4088
rect 11980 3596 12032 3602
rect 11980 3538 12032 3544
rect 11704 3460 11756 3466
rect 11704 3402 11756 3408
rect 11888 3460 11940 3466
rect 11888 3402 11940 3408
rect 11336 3188 11388 3194
rect 11336 3130 11388 3136
rect 11348 1970 11376 3130
rect 11900 2378 11928 3402
rect 11992 3194 12020 3538
rect 12084 3534 12112 4082
rect 13372 3942 13400 4082
rect 13360 3936 13412 3942
rect 13360 3878 13412 3884
rect 12214 3836 12522 3845
rect 12214 3834 12220 3836
rect 12276 3834 12300 3836
rect 12356 3834 12380 3836
rect 12436 3834 12460 3836
rect 12516 3834 12522 3836
rect 12276 3782 12278 3834
rect 12458 3782 12460 3834
rect 12214 3780 12220 3782
rect 12276 3780 12300 3782
rect 12356 3780 12380 3782
rect 12436 3780 12460 3782
rect 12516 3780 12522 3782
rect 12214 3771 12522 3780
rect 13372 3777 13400 3878
rect 13358 3768 13414 3777
rect 13358 3703 13414 3712
rect 12072 3528 12124 3534
rect 12072 3470 12124 3476
rect 11980 3188 12032 3194
rect 11980 3130 12032 3136
rect 12084 3126 12112 3470
rect 12808 3460 12860 3466
rect 12808 3402 12860 3408
rect 12072 3120 12124 3126
rect 12072 3062 12124 3068
rect 11888 2372 11940 2378
rect 11888 2314 11940 2320
rect 11520 2304 11572 2310
rect 11520 2246 11572 2252
rect 11336 1964 11388 1970
rect 11336 1906 11388 1912
rect 11532 1902 11560 2246
rect 12084 2038 12112 3062
rect 12624 2916 12676 2922
rect 12624 2858 12676 2864
rect 12214 2748 12522 2757
rect 12214 2746 12220 2748
rect 12276 2746 12300 2748
rect 12356 2746 12380 2748
rect 12436 2746 12460 2748
rect 12516 2746 12522 2748
rect 12276 2694 12278 2746
rect 12458 2694 12460 2746
rect 12214 2692 12220 2694
rect 12276 2692 12300 2694
rect 12356 2692 12380 2694
rect 12436 2692 12460 2694
rect 12516 2692 12522 2694
rect 12214 2683 12522 2692
rect 12636 2394 12664 2858
rect 12544 2366 12664 2394
rect 12544 2038 12572 2366
rect 12072 2032 12124 2038
rect 12072 1974 12124 1980
rect 12532 2032 12584 2038
rect 12532 1974 12584 1980
rect 11520 1896 11572 1902
rect 11520 1838 11572 1844
rect 11532 1426 11560 1838
rect 12214 1660 12522 1669
rect 12214 1658 12220 1660
rect 12276 1658 12300 1660
rect 12356 1658 12380 1660
rect 12436 1658 12460 1660
rect 12516 1658 12522 1660
rect 12276 1606 12278 1658
rect 12458 1606 12460 1658
rect 12214 1604 12220 1606
rect 12276 1604 12300 1606
rect 12356 1604 12380 1606
rect 12436 1604 12460 1606
rect 12516 1604 12522 1606
rect 12214 1595 12522 1604
rect 11520 1420 11572 1426
rect 11520 1362 11572 1368
rect 11242 1320 11298 1329
rect 12820 1290 12848 3402
rect 13176 3052 13228 3058
rect 13176 2994 13228 3000
rect 13188 2446 13216 2994
rect 13268 2984 13320 2990
rect 13268 2926 13320 2932
rect 13280 2446 13308 2926
rect 13176 2440 13228 2446
rect 13176 2382 13228 2388
rect 13268 2440 13320 2446
rect 13268 2382 13320 2388
rect 13188 2106 13216 2382
rect 13176 2100 13228 2106
rect 13176 2042 13228 2048
rect 13280 1902 13308 2382
rect 13268 1896 13320 1902
rect 13268 1838 13320 1844
rect 13280 1562 13308 1838
rect 13268 1556 13320 1562
rect 13268 1498 13320 1504
rect 11242 1255 11298 1264
rect 12808 1284 12860 1290
rect 12808 1226 12860 1232
rect 1398 504 1454 513
rect 1398 439 1454 448
rect 3698 0 3754 800
rect 11150 0 11206 800
<< via2 >>
rect 1398 14456 1454 14512
rect 2778 13504 2834 13560
rect 1490 12552 1546 12608
rect 2686 12280 2742 12336
rect 1766 11600 1822 11656
rect 1582 10668 1638 10704
rect 1582 10648 1584 10668
rect 1584 10648 1636 10668
rect 1636 10648 1638 10668
rect 2502 11600 2558 11656
rect 2410 10104 2466 10160
rect 2134 9696 2190 9752
rect 4220 13626 4276 13628
rect 4300 13626 4356 13628
rect 4380 13626 4436 13628
rect 4460 13626 4516 13628
rect 4220 13574 4266 13626
rect 4266 13574 4276 13626
rect 4300 13574 4330 13626
rect 4330 13574 4342 13626
rect 4342 13574 4356 13626
rect 4380 13574 4394 13626
rect 4394 13574 4406 13626
rect 4406 13574 4436 13626
rect 4460 13574 4470 13626
rect 4470 13574 4516 13626
rect 4220 13572 4276 13574
rect 4300 13572 4356 13574
rect 4380 13572 4436 13574
rect 4460 13572 4516 13574
rect 4220 12538 4276 12540
rect 4300 12538 4356 12540
rect 4380 12538 4436 12540
rect 4460 12538 4516 12540
rect 4220 12486 4266 12538
rect 4266 12486 4276 12538
rect 4300 12486 4330 12538
rect 4330 12486 4342 12538
rect 4342 12486 4356 12538
rect 4380 12486 4394 12538
rect 4394 12486 4406 12538
rect 4406 12486 4436 12538
rect 4460 12486 4470 12538
rect 4470 12486 4516 12538
rect 4220 12484 4276 12486
rect 4300 12484 4356 12486
rect 4380 12484 4436 12486
rect 4460 12484 4516 12486
rect 4220 11450 4276 11452
rect 4300 11450 4356 11452
rect 4380 11450 4436 11452
rect 4460 11450 4516 11452
rect 4220 11398 4266 11450
rect 4266 11398 4276 11450
rect 4300 11398 4330 11450
rect 4330 11398 4342 11450
rect 4342 11398 4356 11450
rect 4380 11398 4394 11450
rect 4394 11398 4406 11450
rect 4406 11398 4436 11450
rect 4460 11398 4470 11450
rect 4470 11398 4516 11450
rect 4220 11396 4276 11398
rect 4300 11396 4356 11398
rect 4380 11396 4436 11398
rect 4460 11396 4516 11398
rect 2134 8780 2136 8800
rect 2136 8780 2188 8800
rect 2188 8780 2190 8800
rect 2134 8744 2190 8780
rect 1398 6060 1400 6080
rect 1400 6060 1452 6080
rect 1452 6060 1454 6080
rect 1398 6024 1454 6060
rect 2594 6296 2650 6352
rect 1398 5072 1454 5128
rect 2134 3168 2190 3224
rect 1582 2216 1638 2272
rect 3054 7928 3110 7984
rect 5446 12144 5502 12200
rect 4986 10512 5042 10568
rect 4220 10362 4276 10364
rect 4300 10362 4356 10364
rect 4380 10362 4436 10364
rect 4460 10362 4516 10364
rect 4220 10310 4266 10362
rect 4266 10310 4276 10362
rect 4300 10310 4330 10362
rect 4330 10310 4342 10362
rect 4342 10310 4356 10362
rect 4380 10310 4394 10362
rect 4394 10310 4406 10362
rect 4406 10310 4436 10362
rect 4460 10310 4470 10362
rect 4470 10310 4516 10362
rect 4220 10308 4276 10310
rect 4300 10308 4356 10310
rect 4380 10308 4436 10310
rect 4460 10308 4516 10310
rect 4220 9274 4276 9276
rect 4300 9274 4356 9276
rect 4380 9274 4436 9276
rect 4460 9274 4516 9276
rect 4220 9222 4266 9274
rect 4266 9222 4276 9274
rect 4300 9222 4330 9274
rect 4330 9222 4342 9274
rect 4342 9222 4356 9274
rect 4380 9222 4394 9274
rect 4394 9222 4406 9274
rect 4406 9222 4436 9274
rect 4460 9222 4470 9274
rect 4470 9222 4516 9274
rect 4220 9220 4276 9222
rect 4300 9220 4356 9222
rect 4380 9220 4436 9222
rect 4460 9220 4516 9222
rect 4220 8186 4276 8188
rect 4300 8186 4356 8188
rect 4380 8186 4436 8188
rect 4460 8186 4516 8188
rect 4220 8134 4266 8186
rect 4266 8134 4276 8186
rect 4300 8134 4330 8186
rect 4330 8134 4342 8186
rect 4342 8134 4356 8186
rect 4380 8134 4394 8186
rect 4394 8134 4406 8186
rect 4406 8134 4436 8186
rect 4460 8134 4470 8186
rect 4470 8134 4516 8186
rect 4220 8132 4276 8134
rect 4300 8132 4356 8134
rect 4380 8132 4436 8134
rect 4460 8132 4516 8134
rect 6090 11228 6092 11248
rect 6092 11228 6144 11248
rect 6144 11228 6146 11248
rect 6090 11192 6146 11228
rect 6550 11092 6552 11112
rect 6552 11092 6604 11112
rect 6604 11092 6606 11112
rect 6550 11056 6606 11092
rect 5814 9424 5870 9480
rect 3790 7384 3846 7440
rect 3882 6976 3938 7032
rect 5538 7404 5594 7440
rect 6642 9696 6698 9752
rect 6826 9444 6882 9480
rect 6826 9424 6828 9444
rect 6828 9424 6880 9444
rect 6880 9424 6882 9444
rect 7194 10376 7250 10432
rect 7654 12436 7710 12472
rect 7654 12416 7656 12436
rect 7656 12416 7708 12436
rect 7708 12416 7710 12436
rect 8220 13082 8276 13084
rect 8300 13082 8356 13084
rect 8380 13082 8436 13084
rect 8460 13082 8516 13084
rect 8220 13030 8266 13082
rect 8266 13030 8276 13082
rect 8300 13030 8330 13082
rect 8330 13030 8342 13082
rect 8342 13030 8356 13082
rect 8380 13030 8394 13082
rect 8394 13030 8406 13082
rect 8406 13030 8436 13082
rect 8460 13030 8470 13082
rect 8470 13030 8516 13082
rect 8220 13028 8276 13030
rect 8300 13028 8356 13030
rect 8380 13028 8436 13030
rect 8460 13028 8516 13030
rect 8482 12860 8484 12880
rect 8484 12860 8536 12880
rect 8536 12860 8538 12880
rect 8482 12824 8538 12860
rect 8220 11994 8276 11996
rect 8300 11994 8356 11996
rect 8380 11994 8436 11996
rect 8460 11994 8516 11996
rect 8220 11942 8266 11994
rect 8266 11942 8276 11994
rect 8300 11942 8330 11994
rect 8330 11942 8342 11994
rect 8342 11942 8356 11994
rect 8380 11942 8394 11994
rect 8394 11942 8406 11994
rect 8406 11942 8436 11994
rect 8460 11942 8470 11994
rect 8470 11942 8516 11994
rect 8220 11940 8276 11942
rect 8300 11940 8356 11942
rect 8380 11940 8436 11942
rect 8460 11940 8516 11942
rect 8390 11736 8446 11792
rect 7654 11464 7710 11520
rect 7654 11328 7710 11384
rect 7562 11076 7618 11112
rect 7562 11056 7564 11076
rect 7564 11056 7616 11076
rect 7616 11056 7618 11076
rect 8114 11464 8170 11520
rect 7838 11056 7894 11112
rect 7470 9716 7526 9752
rect 7470 9696 7472 9716
rect 7472 9696 7524 9716
rect 7524 9696 7526 9716
rect 7194 9560 7250 9616
rect 8850 13368 8906 13424
rect 9310 12824 9366 12880
rect 8666 12436 8722 12472
rect 8666 12416 8668 12436
rect 8668 12416 8720 12436
rect 8720 12416 8722 12436
rect 8850 11872 8906 11928
rect 8220 10906 8276 10908
rect 8300 10906 8356 10908
rect 8380 10906 8436 10908
rect 8460 10906 8516 10908
rect 8220 10854 8266 10906
rect 8266 10854 8276 10906
rect 8300 10854 8330 10906
rect 8330 10854 8342 10906
rect 8342 10854 8356 10906
rect 8380 10854 8394 10906
rect 8394 10854 8406 10906
rect 8406 10854 8436 10906
rect 8460 10854 8470 10906
rect 8470 10854 8516 10906
rect 8220 10852 8276 10854
rect 8300 10852 8356 10854
rect 8380 10852 8436 10854
rect 8460 10852 8516 10854
rect 8390 10648 8446 10704
rect 8482 9968 8538 10024
rect 8220 9818 8276 9820
rect 8300 9818 8356 9820
rect 8380 9818 8436 9820
rect 8460 9818 8516 9820
rect 8220 9766 8266 9818
rect 8266 9766 8276 9818
rect 8300 9766 8330 9818
rect 8330 9766 8342 9818
rect 8342 9766 8356 9818
rect 8380 9766 8394 9818
rect 8394 9766 8406 9818
rect 8406 9766 8436 9818
rect 8460 9766 8470 9818
rect 8470 9766 8516 9818
rect 8220 9764 8276 9766
rect 8300 9764 8356 9766
rect 8380 9764 8436 9766
rect 8460 9764 8516 9766
rect 5538 7384 5540 7404
rect 5540 7384 5592 7404
rect 5592 7384 5594 7404
rect 3514 4140 3570 4176
rect 3514 4120 3516 4140
rect 3516 4120 3568 4140
rect 3568 4120 3570 4140
rect 2962 1264 3018 1320
rect 3606 3984 3662 4040
rect 4220 7098 4276 7100
rect 4300 7098 4356 7100
rect 4380 7098 4436 7100
rect 4460 7098 4516 7100
rect 4220 7046 4266 7098
rect 4266 7046 4276 7098
rect 4300 7046 4330 7098
rect 4330 7046 4342 7098
rect 4342 7046 4356 7098
rect 4380 7046 4394 7098
rect 4394 7046 4406 7098
rect 4406 7046 4436 7098
rect 4460 7046 4470 7098
rect 4470 7046 4516 7098
rect 4220 7044 4276 7046
rect 4300 7044 4356 7046
rect 4380 7044 4436 7046
rect 4460 7044 4516 7046
rect 4066 6296 4122 6352
rect 4220 6010 4276 6012
rect 4300 6010 4356 6012
rect 4380 6010 4436 6012
rect 4460 6010 4516 6012
rect 4220 5958 4266 6010
rect 4266 5958 4276 6010
rect 4300 5958 4330 6010
rect 4330 5958 4342 6010
rect 4342 5958 4356 6010
rect 4380 5958 4394 6010
rect 4394 5958 4406 6010
rect 4406 5958 4436 6010
rect 4460 5958 4470 6010
rect 4470 5958 4516 6010
rect 4220 5956 4276 5958
rect 4300 5956 4356 5958
rect 4380 5956 4436 5958
rect 4460 5956 4516 5958
rect 4220 4922 4276 4924
rect 4300 4922 4356 4924
rect 4380 4922 4436 4924
rect 4460 4922 4516 4924
rect 4220 4870 4266 4922
rect 4266 4870 4276 4922
rect 4300 4870 4330 4922
rect 4330 4870 4342 4922
rect 4342 4870 4356 4922
rect 4380 4870 4394 4922
rect 4394 4870 4406 4922
rect 4406 4870 4436 4922
rect 4460 4870 4470 4922
rect 4470 4870 4516 4922
rect 4220 4868 4276 4870
rect 4300 4868 4356 4870
rect 4380 4868 4436 4870
rect 4460 4868 4516 4870
rect 4894 4020 4896 4040
rect 4896 4020 4948 4040
rect 4948 4020 4950 4040
rect 4894 3984 4950 4020
rect 4220 3834 4276 3836
rect 4300 3834 4356 3836
rect 4380 3834 4436 3836
rect 4460 3834 4516 3836
rect 4220 3782 4266 3834
rect 4266 3782 4276 3834
rect 4300 3782 4330 3834
rect 4330 3782 4342 3834
rect 4342 3782 4356 3834
rect 4380 3782 4394 3834
rect 4394 3782 4406 3834
rect 4406 3782 4436 3834
rect 4460 3782 4470 3834
rect 4470 3782 4516 3834
rect 4220 3780 4276 3782
rect 4300 3780 4356 3782
rect 4380 3780 4436 3782
rect 4460 3780 4516 3782
rect 4220 2746 4276 2748
rect 4300 2746 4356 2748
rect 4380 2746 4436 2748
rect 4460 2746 4516 2748
rect 4220 2694 4266 2746
rect 4266 2694 4276 2746
rect 4300 2694 4330 2746
rect 4330 2694 4342 2746
rect 4342 2694 4356 2746
rect 4380 2694 4394 2746
rect 4394 2694 4406 2746
rect 4406 2694 4436 2746
rect 4460 2694 4470 2746
rect 4470 2694 4516 2746
rect 4220 2692 4276 2694
rect 4300 2692 4356 2694
rect 4380 2692 4436 2694
rect 4460 2692 4516 2694
rect 4220 1658 4276 1660
rect 4300 1658 4356 1660
rect 4380 1658 4436 1660
rect 4460 1658 4516 1660
rect 4220 1606 4266 1658
rect 4266 1606 4276 1658
rect 4300 1606 4330 1658
rect 4330 1606 4342 1658
rect 4342 1606 4356 1658
rect 4380 1606 4394 1658
rect 4394 1606 4406 1658
rect 4406 1606 4436 1658
rect 4460 1606 4470 1658
rect 4470 1606 4516 1658
rect 4220 1604 4276 1606
rect 4300 1604 4356 1606
rect 4380 1604 4436 1606
rect 4460 1604 4516 1606
rect 5630 3984 5686 4040
rect 8482 9288 8538 9344
rect 8758 11056 8814 11112
rect 8850 10920 8906 10976
rect 9218 12280 9274 12336
rect 9218 11328 9274 11384
rect 9586 12144 9642 12200
rect 9494 11600 9550 11656
rect 9586 11464 9642 11520
rect 9862 11756 9918 11792
rect 9862 11736 9864 11756
rect 9864 11736 9916 11756
rect 9916 11736 9918 11756
rect 9034 9152 9090 9208
rect 9218 10512 9274 10568
rect 9678 10376 9734 10432
rect 9402 10240 9458 10296
rect 9586 10240 9642 10296
rect 9862 10648 9918 10704
rect 9862 10140 9864 10160
rect 9864 10140 9916 10160
rect 9916 10140 9918 10160
rect 9862 10104 9918 10140
rect 9310 9868 9312 9888
rect 9312 9868 9364 9888
rect 9364 9868 9366 9888
rect 9310 9832 9366 9868
rect 8206 8916 8208 8936
rect 8208 8916 8260 8936
rect 8260 8916 8262 8936
rect 8206 8880 8262 8916
rect 8220 8730 8276 8732
rect 8300 8730 8356 8732
rect 8380 8730 8436 8732
rect 8460 8730 8516 8732
rect 8220 8678 8266 8730
rect 8266 8678 8276 8730
rect 8300 8678 8330 8730
rect 8330 8678 8342 8730
rect 8342 8678 8356 8730
rect 8380 8678 8394 8730
rect 8394 8678 8406 8730
rect 8406 8678 8436 8730
rect 8460 8678 8470 8730
rect 8470 8678 8516 8730
rect 8220 8676 8276 8678
rect 8300 8676 8356 8678
rect 8380 8676 8436 8678
rect 8460 8676 8516 8678
rect 8220 7642 8276 7644
rect 8300 7642 8356 7644
rect 8380 7642 8436 7644
rect 8460 7642 8516 7644
rect 8220 7590 8266 7642
rect 8266 7590 8276 7642
rect 8300 7590 8330 7642
rect 8330 7590 8342 7642
rect 8342 7590 8356 7642
rect 8380 7590 8394 7642
rect 8394 7590 8406 7642
rect 8406 7590 8436 7642
rect 8460 7590 8470 7642
rect 8470 7590 8516 7642
rect 8220 7588 8276 7590
rect 8300 7588 8356 7590
rect 8380 7588 8436 7590
rect 8460 7588 8516 7590
rect 8220 6554 8276 6556
rect 8300 6554 8356 6556
rect 8380 6554 8436 6556
rect 8460 6554 8516 6556
rect 8220 6502 8266 6554
rect 8266 6502 8276 6554
rect 8300 6502 8330 6554
rect 8330 6502 8342 6554
rect 8342 6502 8356 6554
rect 8380 6502 8394 6554
rect 8394 6502 8406 6554
rect 8406 6502 8436 6554
rect 8460 6502 8470 6554
rect 8470 6502 8516 6554
rect 8220 6500 8276 6502
rect 8300 6500 8356 6502
rect 8380 6500 8436 6502
rect 8460 6500 8516 6502
rect 8220 5466 8276 5468
rect 8300 5466 8356 5468
rect 8380 5466 8436 5468
rect 8460 5466 8516 5468
rect 8220 5414 8266 5466
rect 8266 5414 8276 5466
rect 8300 5414 8330 5466
rect 8330 5414 8342 5466
rect 8342 5414 8356 5466
rect 8380 5414 8394 5466
rect 8394 5414 8406 5466
rect 8406 5414 8436 5466
rect 8460 5414 8470 5466
rect 8470 5414 8516 5466
rect 8220 5412 8276 5414
rect 8300 5412 8356 5414
rect 8380 5412 8436 5414
rect 8460 5412 8516 5414
rect 8220 4378 8276 4380
rect 8300 4378 8356 4380
rect 8380 4378 8436 4380
rect 8460 4378 8516 4380
rect 8220 4326 8266 4378
rect 8266 4326 8276 4378
rect 8300 4326 8330 4378
rect 8330 4326 8342 4378
rect 8342 4326 8356 4378
rect 8380 4326 8394 4378
rect 8394 4326 8406 4378
rect 8406 4326 8436 4378
rect 8460 4326 8470 4378
rect 8470 4326 8516 4378
rect 8220 4324 8276 4326
rect 8300 4324 8356 4326
rect 8380 4324 8436 4326
rect 8460 4324 8516 4326
rect 8022 3984 8078 4040
rect 9678 9696 9734 9752
rect 9494 9152 9550 9208
rect 10414 11600 10470 11656
rect 10230 10920 10286 10976
rect 12220 13626 12276 13628
rect 12300 13626 12356 13628
rect 12380 13626 12436 13628
rect 12460 13626 12516 13628
rect 12220 13574 12266 13626
rect 12266 13574 12276 13626
rect 12300 13574 12330 13626
rect 12330 13574 12342 13626
rect 12342 13574 12356 13626
rect 12380 13574 12394 13626
rect 12394 13574 12406 13626
rect 12406 13574 12436 13626
rect 12460 13574 12470 13626
rect 12470 13574 12516 13626
rect 12220 13572 12276 13574
rect 12300 13572 12356 13574
rect 12380 13572 12436 13574
rect 12460 13572 12516 13574
rect 10598 11092 10600 11112
rect 10600 11092 10652 11112
rect 10652 11092 10654 11112
rect 10598 11056 10654 11092
rect 10322 10376 10378 10432
rect 10322 9696 10378 9752
rect 10230 9460 10232 9480
rect 10232 9460 10284 9480
rect 10284 9460 10286 9480
rect 10230 9424 10286 9460
rect 10966 11872 11022 11928
rect 11058 10512 11114 10568
rect 10414 9288 10470 9344
rect 10230 8900 10286 8936
rect 10230 8880 10232 8900
rect 10232 8880 10284 8900
rect 10284 8880 10286 8900
rect 11334 10668 11390 10704
rect 11334 10648 11336 10668
rect 11336 10648 11388 10668
rect 11388 10648 11390 10668
rect 11334 10512 11390 10568
rect 11150 9832 11206 9888
rect 11058 9560 11114 9616
rect 12220 12538 12276 12540
rect 12300 12538 12356 12540
rect 12380 12538 12436 12540
rect 12460 12538 12516 12540
rect 12220 12486 12266 12538
rect 12266 12486 12276 12538
rect 12300 12486 12330 12538
rect 12330 12486 12342 12538
rect 12342 12486 12356 12538
rect 12380 12486 12394 12538
rect 12394 12486 12406 12538
rect 12406 12486 12436 12538
rect 12460 12486 12470 12538
rect 12470 12486 12516 12538
rect 12220 12484 12276 12486
rect 12300 12484 12356 12486
rect 12380 12484 12436 12486
rect 12460 12484 12516 12486
rect 11518 11192 11574 11248
rect 8220 3290 8276 3292
rect 8300 3290 8356 3292
rect 8380 3290 8436 3292
rect 8460 3290 8516 3292
rect 8220 3238 8266 3290
rect 8266 3238 8276 3290
rect 8300 3238 8330 3290
rect 8330 3238 8342 3290
rect 8342 3238 8356 3290
rect 8380 3238 8394 3290
rect 8394 3238 8406 3290
rect 8406 3238 8436 3290
rect 8460 3238 8470 3290
rect 8470 3238 8516 3290
rect 8220 3236 8276 3238
rect 8300 3236 8356 3238
rect 8380 3236 8436 3238
rect 8460 3236 8516 3238
rect 8220 2202 8276 2204
rect 8300 2202 8356 2204
rect 8380 2202 8436 2204
rect 8460 2202 8516 2204
rect 8220 2150 8266 2202
rect 8266 2150 8276 2202
rect 8300 2150 8330 2202
rect 8330 2150 8342 2202
rect 8342 2150 8356 2202
rect 8380 2150 8394 2202
rect 8394 2150 8406 2202
rect 8406 2150 8436 2202
rect 8460 2150 8470 2202
rect 8470 2150 8516 2202
rect 8220 2148 8276 2150
rect 8300 2148 8356 2150
rect 8380 2148 8436 2150
rect 8460 2148 8516 2150
rect 8220 1114 8276 1116
rect 8300 1114 8356 1116
rect 8380 1114 8436 1116
rect 8460 1114 8516 1116
rect 8220 1062 8266 1114
rect 8266 1062 8276 1114
rect 8300 1062 8330 1114
rect 8330 1062 8342 1114
rect 8342 1062 8356 1114
rect 8380 1062 8394 1114
rect 8394 1062 8406 1114
rect 8406 1062 8436 1114
rect 8460 1062 8470 1114
rect 8470 1062 8516 1114
rect 8220 1060 8276 1062
rect 8300 1060 8356 1062
rect 8380 1060 8436 1062
rect 8460 1060 8516 1062
rect 12220 11450 12276 11452
rect 12300 11450 12356 11452
rect 12380 11450 12436 11452
rect 12460 11450 12516 11452
rect 12220 11398 12266 11450
rect 12266 11398 12276 11450
rect 12300 11398 12330 11450
rect 12330 11398 12342 11450
rect 12342 11398 12356 11450
rect 12380 11398 12394 11450
rect 12394 11398 12406 11450
rect 12406 11398 12436 11450
rect 12460 11398 12470 11450
rect 12470 11398 12516 11450
rect 12220 11396 12276 11398
rect 12300 11396 12356 11398
rect 12380 11396 12436 11398
rect 12460 11396 12516 11398
rect 11978 11076 12034 11112
rect 13542 11212 13598 11248
rect 13542 11192 13544 11212
rect 13544 11192 13596 11212
rect 13596 11192 13598 11212
rect 11978 11056 11980 11076
rect 11980 11056 12032 11076
rect 12032 11056 12034 11076
rect 11702 10512 11758 10568
rect 12622 10668 12678 10704
rect 12622 10648 12624 10668
rect 12624 10648 12676 10668
rect 12676 10648 12678 10668
rect 12220 10362 12276 10364
rect 12300 10362 12356 10364
rect 12380 10362 12436 10364
rect 12460 10362 12516 10364
rect 12220 10310 12266 10362
rect 12266 10310 12276 10362
rect 12300 10310 12330 10362
rect 12330 10310 12342 10362
rect 12342 10310 12356 10362
rect 12380 10310 12394 10362
rect 12394 10310 12406 10362
rect 12406 10310 12436 10362
rect 12460 10310 12470 10362
rect 12470 10310 12516 10362
rect 12220 10308 12276 10310
rect 12300 10308 12356 10310
rect 12380 10308 12436 10310
rect 12460 10308 12516 10310
rect 12220 9274 12276 9276
rect 12300 9274 12356 9276
rect 12380 9274 12436 9276
rect 12460 9274 12516 9276
rect 12220 9222 12266 9274
rect 12266 9222 12276 9274
rect 12300 9222 12330 9274
rect 12330 9222 12342 9274
rect 12342 9222 12356 9274
rect 12380 9222 12394 9274
rect 12394 9222 12406 9274
rect 12406 9222 12436 9274
rect 12460 9222 12470 9274
rect 12470 9222 12516 9274
rect 12220 9220 12276 9222
rect 12300 9220 12356 9222
rect 12380 9220 12436 9222
rect 12460 9220 12516 9222
rect 12806 10648 12862 10704
rect 12622 8744 12678 8800
rect 12220 8186 12276 8188
rect 12300 8186 12356 8188
rect 12380 8186 12436 8188
rect 12460 8186 12516 8188
rect 12220 8134 12266 8186
rect 12266 8134 12276 8186
rect 12300 8134 12330 8186
rect 12330 8134 12342 8186
rect 12342 8134 12356 8186
rect 12380 8134 12394 8186
rect 12394 8134 12406 8186
rect 12406 8134 12436 8186
rect 12460 8134 12470 8186
rect 12470 8134 12516 8186
rect 12220 8132 12276 8134
rect 12300 8132 12356 8134
rect 12380 8132 12436 8134
rect 12460 8132 12516 8134
rect 12220 7098 12276 7100
rect 12300 7098 12356 7100
rect 12380 7098 12436 7100
rect 12460 7098 12516 7100
rect 12220 7046 12266 7098
rect 12266 7046 12276 7098
rect 12300 7046 12330 7098
rect 12330 7046 12342 7098
rect 12342 7046 12356 7098
rect 12380 7046 12394 7098
rect 12394 7046 12406 7098
rect 12406 7046 12436 7098
rect 12460 7046 12470 7098
rect 12470 7046 12516 7098
rect 12220 7044 12276 7046
rect 12300 7044 12356 7046
rect 12380 7044 12436 7046
rect 12460 7044 12516 7046
rect 12220 6010 12276 6012
rect 12300 6010 12356 6012
rect 12380 6010 12436 6012
rect 12460 6010 12516 6012
rect 12220 5958 12266 6010
rect 12266 5958 12276 6010
rect 12300 5958 12330 6010
rect 12330 5958 12342 6010
rect 12342 5958 12356 6010
rect 12380 5958 12394 6010
rect 12394 5958 12406 6010
rect 12406 5958 12436 6010
rect 12460 5958 12470 6010
rect 12470 5958 12516 6010
rect 12220 5956 12276 5958
rect 12300 5956 12356 5958
rect 12380 5956 12436 5958
rect 12460 5956 12516 5958
rect 13542 6160 13598 6216
rect 12220 4922 12276 4924
rect 12300 4922 12356 4924
rect 12380 4922 12436 4924
rect 12460 4922 12516 4924
rect 12220 4870 12266 4922
rect 12266 4870 12276 4922
rect 12300 4870 12330 4922
rect 12330 4870 12342 4922
rect 12342 4870 12356 4922
rect 12380 4870 12394 4922
rect 12394 4870 12406 4922
rect 12406 4870 12436 4922
rect 12460 4870 12470 4922
rect 12470 4870 12516 4922
rect 12220 4868 12276 4870
rect 12300 4868 12356 4870
rect 12380 4868 12436 4870
rect 12460 4868 12516 4870
rect 12220 3834 12276 3836
rect 12300 3834 12356 3836
rect 12380 3834 12436 3836
rect 12460 3834 12516 3836
rect 12220 3782 12266 3834
rect 12266 3782 12276 3834
rect 12300 3782 12330 3834
rect 12330 3782 12342 3834
rect 12342 3782 12356 3834
rect 12380 3782 12394 3834
rect 12394 3782 12406 3834
rect 12406 3782 12436 3834
rect 12460 3782 12470 3834
rect 12470 3782 12516 3834
rect 12220 3780 12276 3782
rect 12300 3780 12356 3782
rect 12380 3780 12436 3782
rect 12460 3780 12516 3782
rect 13358 3712 13414 3768
rect 12220 2746 12276 2748
rect 12300 2746 12356 2748
rect 12380 2746 12436 2748
rect 12460 2746 12516 2748
rect 12220 2694 12266 2746
rect 12266 2694 12276 2746
rect 12300 2694 12330 2746
rect 12330 2694 12342 2746
rect 12342 2694 12356 2746
rect 12380 2694 12394 2746
rect 12394 2694 12406 2746
rect 12406 2694 12436 2746
rect 12460 2694 12470 2746
rect 12470 2694 12516 2746
rect 12220 2692 12276 2694
rect 12300 2692 12356 2694
rect 12380 2692 12436 2694
rect 12460 2692 12516 2694
rect 12220 1658 12276 1660
rect 12300 1658 12356 1660
rect 12380 1658 12436 1660
rect 12460 1658 12516 1660
rect 12220 1606 12266 1658
rect 12266 1606 12276 1658
rect 12300 1606 12330 1658
rect 12330 1606 12342 1658
rect 12342 1606 12356 1658
rect 12380 1606 12394 1658
rect 12394 1606 12406 1658
rect 12406 1606 12436 1658
rect 12460 1606 12470 1658
rect 12470 1606 12516 1658
rect 12220 1604 12276 1606
rect 12300 1604 12356 1606
rect 12380 1604 12436 1606
rect 12460 1604 12516 1606
rect 11242 1264 11298 1320
rect 1398 448 1454 504
<< metal3 >>
rect 0 14514 800 14544
rect 1393 14514 1459 14517
rect 0 14512 1459 14514
rect 0 14456 1398 14512
rect 1454 14456 1459 14512
rect 0 14454 1459 14456
rect 0 14424 800 14454
rect 1393 14451 1459 14454
rect 14200 13698 15000 13728
rect 12758 13638 15000 13698
rect 4210 13632 4526 13633
rect 0 13562 800 13592
rect 4210 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4526 13632
rect 4210 13567 4526 13568
rect 12210 13632 12526 13633
rect 12210 13568 12216 13632
rect 12280 13568 12296 13632
rect 12360 13568 12376 13632
rect 12440 13568 12456 13632
rect 12520 13568 12526 13632
rect 12210 13567 12526 13568
rect 2773 13562 2839 13565
rect 0 13560 2839 13562
rect 0 13504 2778 13560
rect 2834 13504 2839 13560
rect 0 13502 2839 13504
rect 0 13472 800 13502
rect 2773 13499 2839 13502
rect 8845 13426 8911 13429
rect 12758 13426 12818 13638
rect 14200 13608 15000 13638
rect 8845 13424 12818 13426
rect 8845 13368 8850 13424
rect 8906 13368 12818 13424
rect 8845 13366 12818 13368
rect 8845 13363 8911 13366
rect 8210 13088 8526 13089
rect 8210 13024 8216 13088
rect 8280 13024 8296 13088
rect 8360 13024 8376 13088
rect 8440 13024 8456 13088
rect 8520 13024 8526 13088
rect 8210 13023 8526 13024
rect 8477 12882 8543 12885
rect 9305 12882 9371 12885
rect 8477 12880 9371 12882
rect 8477 12824 8482 12880
rect 8538 12824 9310 12880
rect 9366 12824 9371 12880
rect 8477 12822 9371 12824
rect 8477 12819 8543 12822
rect 9305 12819 9371 12822
rect 0 12610 800 12640
rect 1485 12610 1551 12613
rect 0 12608 1551 12610
rect 0 12552 1490 12608
rect 1546 12552 1551 12608
rect 0 12550 1551 12552
rect 0 12520 800 12550
rect 1485 12547 1551 12550
rect 4210 12544 4526 12545
rect 4210 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4526 12544
rect 4210 12479 4526 12480
rect 12210 12544 12526 12545
rect 12210 12480 12216 12544
rect 12280 12480 12296 12544
rect 12360 12480 12376 12544
rect 12440 12480 12456 12544
rect 12520 12480 12526 12544
rect 12210 12479 12526 12480
rect 7649 12474 7715 12477
rect 8661 12474 8727 12477
rect 7649 12472 8727 12474
rect 7649 12416 7654 12472
rect 7710 12416 8666 12472
rect 8722 12416 8727 12472
rect 7649 12414 8727 12416
rect 7649 12411 7715 12414
rect 8661 12411 8727 12414
rect 2681 12338 2747 12341
rect 9213 12338 9279 12341
rect 2681 12336 9279 12338
rect 2681 12280 2686 12336
rect 2742 12280 9218 12336
rect 9274 12280 9279 12336
rect 2681 12278 9279 12280
rect 2681 12275 2747 12278
rect 9213 12275 9279 12278
rect 5441 12202 5507 12205
rect 9581 12202 9647 12205
rect 5441 12200 9647 12202
rect 5441 12144 5446 12200
rect 5502 12144 9586 12200
rect 9642 12144 9647 12200
rect 5441 12142 9647 12144
rect 5441 12139 5507 12142
rect 9581 12139 9647 12142
rect 8210 12000 8526 12001
rect 8210 11936 8216 12000
rect 8280 11936 8296 12000
rect 8360 11936 8376 12000
rect 8440 11936 8456 12000
rect 8520 11936 8526 12000
rect 8210 11935 8526 11936
rect 8845 11930 8911 11933
rect 10961 11930 11027 11933
rect 8845 11928 11027 11930
rect 8845 11872 8850 11928
rect 8906 11872 10966 11928
rect 11022 11872 11027 11928
rect 8845 11870 11027 11872
rect 8845 11867 8911 11870
rect 10961 11867 11027 11870
rect 8385 11794 8451 11797
rect 9857 11794 9923 11797
rect 8385 11792 9923 11794
rect 8385 11736 8390 11792
rect 8446 11736 9862 11792
rect 9918 11736 9923 11792
rect 8385 11734 9923 11736
rect 8385 11731 8451 11734
rect 9857 11731 9923 11734
rect 0 11658 800 11688
rect 1761 11658 1827 11661
rect 2497 11658 2563 11661
rect 0 11656 2563 11658
rect 0 11600 1766 11656
rect 1822 11600 2502 11656
rect 2558 11600 2563 11656
rect 0 11598 2563 11600
rect 0 11568 800 11598
rect 1761 11595 1827 11598
rect 2497 11595 2563 11598
rect 9489 11658 9555 11661
rect 10409 11658 10475 11661
rect 9489 11656 10475 11658
rect 9489 11600 9494 11656
rect 9550 11600 10414 11656
rect 10470 11600 10475 11656
rect 9489 11598 10475 11600
rect 9489 11595 9555 11598
rect 10409 11595 10475 11598
rect 7649 11522 7715 11525
rect 8109 11522 8175 11525
rect 9581 11522 9647 11525
rect 7649 11520 9647 11522
rect 7649 11464 7654 11520
rect 7710 11464 8114 11520
rect 8170 11464 9586 11520
rect 9642 11464 9647 11520
rect 7649 11462 9647 11464
rect 7649 11459 7715 11462
rect 8109 11459 8175 11462
rect 9581 11459 9647 11462
rect 4210 11456 4526 11457
rect 4210 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4526 11456
rect 4210 11391 4526 11392
rect 12210 11456 12526 11457
rect 12210 11392 12216 11456
rect 12280 11392 12296 11456
rect 12360 11392 12376 11456
rect 12440 11392 12456 11456
rect 12520 11392 12526 11456
rect 12210 11391 12526 11392
rect 7649 11386 7715 11389
rect 9213 11386 9279 11389
rect 7649 11384 9279 11386
rect 7649 11328 7654 11384
rect 7710 11328 9218 11384
rect 9274 11328 9279 11384
rect 7649 11326 9279 11328
rect 7649 11323 7715 11326
rect 9213 11323 9279 11326
rect 6085 11250 6151 11253
rect 11513 11250 11579 11253
rect 6085 11248 11579 11250
rect 6085 11192 6090 11248
rect 6146 11192 11518 11248
rect 11574 11192 11579 11248
rect 6085 11190 11579 11192
rect 6085 11187 6151 11190
rect 11513 11187 11579 11190
rect 13537 11250 13603 11253
rect 14200 11250 15000 11280
rect 13537 11248 15000 11250
rect 13537 11192 13542 11248
rect 13598 11192 15000 11248
rect 13537 11190 15000 11192
rect 13537 11187 13603 11190
rect 14200 11160 15000 11190
rect 6545 11114 6611 11117
rect 7557 11114 7623 11117
rect 6545 11112 7623 11114
rect 6545 11056 6550 11112
rect 6606 11056 7562 11112
rect 7618 11056 7623 11112
rect 6545 11054 7623 11056
rect 6545 11051 6611 11054
rect 7557 11051 7623 11054
rect 7833 11114 7899 11117
rect 8753 11114 8819 11117
rect 7833 11112 8819 11114
rect 7833 11056 7838 11112
rect 7894 11056 8758 11112
rect 8814 11056 8819 11112
rect 7833 11054 8819 11056
rect 7833 11051 7899 11054
rect 8753 11051 8819 11054
rect 10593 11114 10659 11117
rect 11973 11114 12039 11117
rect 10593 11112 12039 11114
rect 10593 11056 10598 11112
rect 10654 11056 11978 11112
rect 12034 11056 12039 11112
rect 10593 11054 12039 11056
rect 10593 11051 10659 11054
rect 11973 11051 12039 11054
rect 8845 10978 8911 10981
rect 10225 10978 10291 10981
rect 8845 10976 10291 10978
rect 8845 10920 8850 10976
rect 8906 10920 10230 10976
rect 10286 10920 10291 10976
rect 8845 10918 10291 10920
rect 8845 10915 8911 10918
rect 10225 10915 10291 10918
rect 8210 10912 8526 10913
rect 8210 10848 8216 10912
rect 8280 10848 8296 10912
rect 8360 10848 8376 10912
rect 8440 10848 8456 10912
rect 8520 10848 8526 10912
rect 8210 10847 8526 10848
rect 0 10706 800 10736
rect 1577 10706 1643 10709
rect 0 10704 1643 10706
rect 0 10648 1582 10704
rect 1638 10648 1643 10704
rect 0 10646 1643 10648
rect 0 10616 800 10646
rect 1577 10643 1643 10646
rect 8385 10706 8451 10709
rect 9857 10706 9923 10709
rect 8385 10704 9923 10706
rect 8385 10648 8390 10704
rect 8446 10648 9862 10704
rect 9918 10648 9923 10704
rect 8385 10646 9923 10648
rect 8385 10643 8451 10646
rect 9857 10643 9923 10646
rect 11329 10706 11395 10709
rect 12617 10706 12683 10709
rect 12801 10706 12867 10709
rect 11329 10704 12867 10706
rect 11329 10648 11334 10704
rect 11390 10648 12622 10704
rect 12678 10648 12806 10704
rect 12862 10648 12867 10704
rect 11329 10646 12867 10648
rect 11329 10643 11395 10646
rect 12617 10643 12683 10646
rect 12801 10643 12867 10646
rect 4981 10570 5047 10573
rect 9213 10570 9279 10573
rect 11053 10570 11119 10573
rect 4981 10568 9279 10570
rect 4981 10512 4986 10568
rect 5042 10512 9218 10568
rect 9274 10512 9279 10568
rect 4981 10510 9279 10512
rect 4981 10507 5047 10510
rect 9213 10507 9279 10510
rect 9492 10568 11119 10570
rect 9492 10512 11058 10568
rect 11114 10512 11119 10568
rect 9492 10510 11119 10512
rect 7189 10434 7255 10437
rect 9492 10434 9552 10510
rect 11053 10507 11119 10510
rect 11329 10570 11395 10573
rect 11697 10570 11763 10573
rect 11329 10568 11763 10570
rect 11329 10512 11334 10568
rect 11390 10512 11702 10568
rect 11758 10512 11763 10568
rect 11329 10510 11763 10512
rect 11329 10507 11395 10510
rect 11697 10507 11763 10510
rect 7189 10432 9552 10434
rect 7189 10376 7194 10432
rect 7250 10376 9552 10432
rect 7189 10374 9552 10376
rect 9673 10434 9739 10437
rect 10317 10434 10383 10437
rect 9673 10432 10383 10434
rect 9673 10376 9678 10432
rect 9734 10376 10322 10432
rect 10378 10376 10383 10432
rect 9673 10374 10383 10376
rect 7189 10371 7255 10374
rect 9673 10371 9739 10374
rect 10317 10371 10383 10374
rect 4210 10368 4526 10369
rect 4210 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4526 10368
rect 4210 10303 4526 10304
rect 12210 10368 12526 10369
rect 12210 10304 12216 10368
rect 12280 10304 12296 10368
rect 12360 10304 12376 10368
rect 12440 10304 12456 10368
rect 12520 10304 12526 10368
rect 12210 10303 12526 10304
rect 9397 10298 9463 10301
rect 9581 10298 9647 10301
rect 9397 10296 9647 10298
rect 9397 10240 9402 10296
rect 9458 10240 9586 10296
rect 9642 10240 9647 10296
rect 9397 10238 9647 10240
rect 9397 10235 9463 10238
rect 9581 10235 9647 10238
rect 2405 10162 2471 10165
rect 9857 10162 9923 10165
rect 2405 10160 9923 10162
rect 2405 10104 2410 10160
rect 2466 10104 9862 10160
rect 9918 10104 9923 10160
rect 2405 10102 9923 10104
rect 2405 10099 2471 10102
rect 9857 10099 9923 10102
rect 8477 10026 8543 10029
rect 8702 10026 8708 10028
rect 8477 10024 8708 10026
rect 8477 9968 8482 10024
rect 8538 9968 8708 10024
rect 8477 9966 8708 9968
rect 8477 9963 8543 9966
rect 8702 9964 8708 9966
rect 8772 9964 8778 10028
rect 9305 9890 9371 9893
rect 11145 9890 11211 9893
rect 9305 9888 11211 9890
rect 9305 9832 9310 9888
rect 9366 9832 11150 9888
rect 11206 9832 11211 9888
rect 9305 9830 11211 9832
rect 9305 9827 9371 9830
rect 11145 9827 11211 9830
rect 8210 9824 8526 9825
rect 0 9754 800 9784
rect 8210 9760 8216 9824
rect 8280 9760 8296 9824
rect 8360 9760 8376 9824
rect 8440 9760 8456 9824
rect 8520 9760 8526 9824
rect 8210 9759 8526 9760
rect 2129 9754 2195 9757
rect 0 9752 2195 9754
rect 0 9696 2134 9752
rect 2190 9696 2195 9752
rect 0 9694 2195 9696
rect 0 9664 800 9694
rect 2129 9691 2195 9694
rect 6637 9754 6703 9757
rect 7465 9754 7531 9757
rect 6637 9752 7531 9754
rect 6637 9696 6642 9752
rect 6698 9696 7470 9752
rect 7526 9696 7531 9752
rect 6637 9694 7531 9696
rect 6637 9691 6703 9694
rect 7465 9691 7531 9694
rect 9673 9754 9739 9757
rect 10317 9754 10383 9757
rect 9673 9752 10383 9754
rect 9673 9696 9678 9752
rect 9734 9696 10322 9752
rect 10378 9696 10383 9752
rect 9673 9694 10383 9696
rect 9673 9691 9739 9694
rect 10317 9691 10383 9694
rect 7189 9618 7255 9621
rect 11053 9618 11119 9621
rect 7189 9616 11119 9618
rect 7189 9560 7194 9616
rect 7250 9560 11058 9616
rect 11114 9560 11119 9616
rect 7189 9558 11119 9560
rect 7189 9555 7255 9558
rect 11053 9555 11119 9558
rect 5809 9482 5875 9485
rect 6821 9482 6887 9485
rect 5809 9480 6887 9482
rect 5809 9424 5814 9480
rect 5870 9424 6826 9480
rect 6882 9424 6887 9480
rect 5809 9422 6887 9424
rect 5809 9419 5875 9422
rect 6821 9419 6887 9422
rect 8702 9420 8708 9484
rect 8772 9482 8778 9484
rect 10225 9482 10291 9485
rect 8772 9480 10291 9482
rect 8772 9424 10230 9480
rect 10286 9424 10291 9480
rect 8772 9422 10291 9424
rect 8772 9420 8778 9422
rect 10225 9419 10291 9422
rect 8477 9346 8543 9349
rect 10409 9346 10475 9349
rect 8477 9344 10475 9346
rect 8477 9288 8482 9344
rect 8538 9288 10414 9344
rect 10470 9288 10475 9344
rect 8477 9286 10475 9288
rect 8477 9283 8543 9286
rect 10409 9283 10475 9286
rect 4210 9280 4526 9281
rect 4210 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4526 9280
rect 4210 9215 4526 9216
rect 12210 9280 12526 9281
rect 12210 9216 12216 9280
rect 12280 9216 12296 9280
rect 12360 9216 12376 9280
rect 12440 9216 12456 9280
rect 12520 9216 12526 9280
rect 12210 9215 12526 9216
rect 9029 9210 9095 9213
rect 9489 9210 9555 9213
rect 9029 9208 9555 9210
rect 9029 9152 9034 9208
rect 9090 9152 9494 9208
rect 9550 9152 9555 9208
rect 9029 9150 9555 9152
rect 9029 9147 9095 9150
rect 9489 9147 9555 9150
rect 8201 8938 8267 8941
rect 10225 8938 10291 8941
rect 8201 8936 10291 8938
rect 8201 8880 8206 8936
rect 8262 8880 10230 8936
rect 10286 8880 10291 8936
rect 8201 8878 10291 8880
rect 8201 8875 8267 8878
rect 10225 8875 10291 8878
rect 0 8802 800 8832
rect 2129 8802 2195 8805
rect 0 8800 2195 8802
rect 0 8744 2134 8800
rect 2190 8744 2195 8800
rect 0 8742 2195 8744
rect 0 8712 800 8742
rect 2129 8739 2195 8742
rect 12617 8802 12683 8805
rect 14200 8802 15000 8832
rect 12617 8800 15000 8802
rect 12617 8744 12622 8800
rect 12678 8744 15000 8800
rect 12617 8742 15000 8744
rect 12617 8739 12683 8742
rect 8210 8736 8526 8737
rect 8210 8672 8216 8736
rect 8280 8672 8296 8736
rect 8360 8672 8376 8736
rect 8440 8672 8456 8736
rect 8520 8672 8526 8736
rect 14200 8712 15000 8742
rect 8210 8671 8526 8672
rect 4210 8192 4526 8193
rect 4210 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4526 8192
rect 4210 8127 4526 8128
rect 12210 8192 12526 8193
rect 12210 8128 12216 8192
rect 12280 8128 12296 8192
rect 12360 8128 12376 8192
rect 12440 8128 12456 8192
rect 12520 8128 12526 8192
rect 12210 8127 12526 8128
rect 0 7986 800 8016
rect 3049 7986 3115 7989
rect 0 7984 3115 7986
rect 0 7928 3054 7984
rect 3110 7928 3115 7984
rect 0 7926 3115 7928
rect 0 7896 800 7926
rect 3049 7923 3115 7926
rect 8210 7648 8526 7649
rect 8210 7584 8216 7648
rect 8280 7584 8296 7648
rect 8360 7584 8376 7648
rect 8440 7584 8456 7648
rect 8520 7584 8526 7648
rect 8210 7583 8526 7584
rect 3785 7442 3851 7445
rect 5533 7442 5599 7445
rect 3785 7440 5599 7442
rect 3785 7384 3790 7440
rect 3846 7384 5538 7440
rect 5594 7384 5599 7440
rect 3785 7382 5599 7384
rect 3785 7379 3851 7382
rect 5533 7379 5599 7382
rect 4210 7104 4526 7105
rect 0 7034 800 7064
rect 4210 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4526 7104
rect 4210 7039 4526 7040
rect 12210 7104 12526 7105
rect 12210 7040 12216 7104
rect 12280 7040 12296 7104
rect 12360 7040 12376 7104
rect 12440 7040 12456 7104
rect 12520 7040 12526 7104
rect 12210 7039 12526 7040
rect 3877 7034 3943 7037
rect 0 7032 3943 7034
rect 0 6976 3882 7032
rect 3938 6976 3943 7032
rect 0 6974 3943 6976
rect 0 6944 800 6974
rect 3877 6971 3943 6974
rect 8210 6560 8526 6561
rect 8210 6496 8216 6560
rect 8280 6496 8296 6560
rect 8360 6496 8376 6560
rect 8440 6496 8456 6560
rect 8520 6496 8526 6560
rect 8210 6495 8526 6496
rect 2589 6354 2655 6357
rect 4061 6354 4127 6357
rect 2589 6352 4127 6354
rect 2589 6296 2594 6352
rect 2650 6296 4066 6352
rect 4122 6296 4127 6352
rect 2589 6294 4127 6296
rect 2589 6291 2655 6294
rect 4061 6291 4127 6294
rect 13537 6218 13603 6221
rect 14200 6218 15000 6248
rect 13537 6216 15000 6218
rect 13537 6160 13542 6216
rect 13598 6160 15000 6216
rect 13537 6158 15000 6160
rect 13537 6155 13603 6158
rect 14200 6128 15000 6158
rect 0 6082 800 6112
rect 1393 6082 1459 6085
rect 0 6080 1459 6082
rect 0 6024 1398 6080
rect 1454 6024 1459 6080
rect 0 6022 1459 6024
rect 0 5992 800 6022
rect 1393 6019 1459 6022
rect 4210 6016 4526 6017
rect 4210 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4526 6016
rect 4210 5951 4526 5952
rect 12210 6016 12526 6017
rect 12210 5952 12216 6016
rect 12280 5952 12296 6016
rect 12360 5952 12376 6016
rect 12440 5952 12456 6016
rect 12520 5952 12526 6016
rect 12210 5951 12526 5952
rect 8210 5472 8526 5473
rect 8210 5408 8216 5472
rect 8280 5408 8296 5472
rect 8360 5408 8376 5472
rect 8440 5408 8456 5472
rect 8520 5408 8526 5472
rect 8210 5407 8526 5408
rect 0 5130 800 5160
rect 1393 5130 1459 5133
rect 0 5128 1459 5130
rect 0 5072 1398 5128
rect 1454 5072 1459 5128
rect 0 5070 1459 5072
rect 0 5040 800 5070
rect 1393 5067 1459 5070
rect 4210 4928 4526 4929
rect 4210 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4526 4928
rect 4210 4863 4526 4864
rect 12210 4928 12526 4929
rect 12210 4864 12216 4928
rect 12280 4864 12296 4928
rect 12360 4864 12376 4928
rect 12440 4864 12456 4928
rect 12520 4864 12526 4928
rect 12210 4863 12526 4864
rect 8210 4384 8526 4385
rect 8210 4320 8216 4384
rect 8280 4320 8296 4384
rect 8360 4320 8376 4384
rect 8440 4320 8456 4384
rect 8520 4320 8526 4384
rect 8210 4319 8526 4320
rect 0 4178 800 4208
rect 3509 4178 3575 4181
rect 0 4176 3575 4178
rect 0 4120 3514 4176
rect 3570 4120 3575 4176
rect 0 4118 3575 4120
rect 0 4088 800 4118
rect 3509 4115 3575 4118
rect 3601 4042 3667 4045
rect 4889 4042 4955 4045
rect 5625 4042 5691 4045
rect 8017 4042 8083 4045
rect 3601 4040 8083 4042
rect 3601 3984 3606 4040
rect 3662 3984 4894 4040
rect 4950 3984 5630 4040
rect 5686 3984 8022 4040
rect 8078 3984 8083 4040
rect 3601 3982 8083 3984
rect 3601 3979 3667 3982
rect 4889 3979 4955 3982
rect 5625 3979 5691 3982
rect 8017 3979 8083 3982
rect 4210 3840 4526 3841
rect 4210 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4526 3840
rect 4210 3775 4526 3776
rect 12210 3840 12526 3841
rect 12210 3776 12216 3840
rect 12280 3776 12296 3840
rect 12360 3776 12376 3840
rect 12440 3776 12456 3840
rect 12520 3776 12526 3840
rect 12210 3775 12526 3776
rect 13353 3770 13419 3773
rect 14200 3770 15000 3800
rect 13353 3768 15000 3770
rect 13353 3712 13358 3768
rect 13414 3712 15000 3768
rect 13353 3710 15000 3712
rect 13353 3707 13419 3710
rect 14200 3680 15000 3710
rect 8210 3296 8526 3297
rect 0 3226 800 3256
rect 8210 3232 8216 3296
rect 8280 3232 8296 3296
rect 8360 3232 8376 3296
rect 8440 3232 8456 3296
rect 8520 3232 8526 3296
rect 8210 3231 8526 3232
rect 2129 3226 2195 3229
rect 0 3224 2195 3226
rect 0 3168 2134 3224
rect 2190 3168 2195 3224
rect 0 3166 2195 3168
rect 0 3136 800 3166
rect 2129 3163 2195 3166
rect 4210 2752 4526 2753
rect 4210 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4526 2752
rect 4210 2687 4526 2688
rect 12210 2752 12526 2753
rect 12210 2688 12216 2752
rect 12280 2688 12296 2752
rect 12360 2688 12376 2752
rect 12440 2688 12456 2752
rect 12520 2688 12526 2752
rect 12210 2687 12526 2688
rect 0 2274 800 2304
rect 1577 2274 1643 2277
rect 0 2272 1643 2274
rect 0 2216 1582 2272
rect 1638 2216 1643 2272
rect 0 2214 1643 2216
rect 0 2184 800 2214
rect 1577 2211 1643 2214
rect 8210 2208 8526 2209
rect 8210 2144 8216 2208
rect 8280 2144 8296 2208
rect 8360 2144 8376 2208
rect 8440 2144 8456 2208
rect 8520 2144 8526 2208
rect 8210 2143 8526 2144
rect 4210 1664 4526 1665
rect 4210 1600 4216 1664
rect 4280 1600 4296 1664
rect 4360 1600 4376 1664
rect 4440 1600 4456 1664
rect 4520 1600 4526 1664
rect 4210 1599 4526 1600
rect 12210 1664 12526 1665
rect 12210 1600 12216 1664
rect 12280 1600 12296 1664
rect 12360 1600 12376 1664
rect 12440 1600 12456 1664
rect 12520 1600 12526 1664
rect 12210 1599 12526 1600
rect 0 1322 800 1352
rect 2957 1322 3023 1325
rect 0 1320 3023 1322
rect 0 1264 2962 1320
rect 3018 1264 3023 1320
rect 0 1262 3023 1264
rect 0 1232 800 1262
rect 2957 1259 3023 1262
rect 11237 1322 11303 1325
rect 14200 1322 15000 1352
rect 11237 1320 15000 1322
rect 11237 1264 11242 1320
rect 11298 1264 15000 1320
rect 11237 1262 15000 1264
rect 11237 1259 11303 1262
rect 14200 1232 15000 1262
rect 8210 1120 8526 1121
rect 8210 1056 8216 1120
rect 8280 1056 8296 1120
rect 8360 1056 8376 1120
rect 8440 1056 8456 1120
rect 8520 1056 8526 1120
rect 8210 1055 8526 1056
rect 0 506 800 536
rect 1393 506 1459 509
rect 0 504 1459 506
rect 0 448 1398 504
rect 1454 448 1459 504
rect 0 446 1459 448
rect 0 416 800 446
rect 1393 443 1459 446
<< via3 >>
rect 4216 13628 4280 13632
rect 4216 13572 4220 13628
rect 4220 13572 4276 13628
rect 4276 13572 4280 13628
rect 4216 13568 4280 13572
rect 4296 13628 4360 13632
rect 4296 13572 4300 13628
rect 4300 13572 4356 13628
rect 4356 13572 4360 13628
rect 4296 13568 4360 13572
rect 4376 13628 4440 13632
rect 4376 13572 4380 13628
rect 4380 13572 4436 13628
rect 4436 13572 4440 13628
rect 4376 13568 4440 13572
rect 4456 13628 4520 13632
rect 4456 13572 4460 13628
rect 4460 13572 4516 13628
rect 4516 13572 4520 13628
rect 4456 13568 4520 13572
rect 12216 13628 12280 13632
rect 12216 13572 12220 13628
rect 12220 13572 12276 13628
rect 12276 13572 12280 13628
rect 12216 13568 12280 13572
rect 12296 13628 12360 13632
rect 12296 13572 12300 13628
rect 12300 13572 12356 13628
rect 12356 13572 12360 13628
rect 12296 13568 12360 13572
rect 12376 13628 12440 13632
rect 12376 13572 12380 13628
rect 12380 13572 12436 13628
rect 12436 13572 12440 13628
rect 12376 13568 12440 13572
rect 12456 13628 12520 13632
rect 12456 13572 12460 13628
rect 12460 13572 12516 13628
rect 12516 13572 12520 13628
rect 12456 13568 12520 13572
rect 8216 13084 8280 13088
rect 8216 13028 8220 13084
rect 8220 13028 8276 13084
rect 8276 13028 8280 13084
rect 8216 13024 8280 13028
rect 8296 13084 8360 13088
rect 8296 13028 8300 13084
rect 8300 13028 8356 13084
rect 8356 13028 8360 13084
rect 8296 13024 8360 13028
rect 8376 13084 8440 13088
rect 8376 13028 8380 13084
rect 8380 13028 8436 13084
rect 8436 13028 8440 13084
rect 8376 13024 8440 13028
rect 8456 13084 8520 13088
rect 8456 13028 8460 13084
rect 8460 13028 8516 13084
rect 8516 13028 8520 13084
rect 8456 13024 8520 13028
rect 4216 12540 4280 12544
rect 4216 12484 4220 12540
rect 4220 12484 4276 12540
rect 4276 12484 4280 12540
rect 4216 12480 4280 12484
rect 4296 12540 4360 12544
rect 4296 12484 4300 12540
rect 4300 12484 4356 12540
rect 4356 12484 4360 12540
rect 4296 12480 4360 12484
rect 4376 12540 4440 12544
rect 4376 12484 4380 12540
rect 4380 12484 4436 12540
rect 4436 12484 4440 12540
rect 4376 12480 4440 12484
rect 4456 12540 4520 12544
rect 4456 12484 4460 12540
rect 4460 12484 4516 12540
rect 4516 12484 4520 12540
rect 4456 12480 4520 12484
rect 12216 12540 12280 12544
rect 12216 12484 12220 12540
rect 12220 12484 12276 12540
rect 12276 12484 12280 12540
rect 12216 12480 12280 12484
rect 12296 12540 12360 12544
rect 12296 12484 12300 12540
rect 12300 12484 12356 12540
rect 12356 12484 12360 12540
rect 12296 12480 12360 12484
rect 12376 12540 12440 12544
rect 12376 12484 12380 12540
rect 12380 12484 12436 12540
rect 12436 12484 12440 12540
rect 12376 12480 12440 12484
rect 12456 12540 12520 12544
rect 12456 12484 12460 12540
rect 12460 12484 12516 12540
rect 12516 12484 12520 12540
rect 12456 12480 12520 12484
rect 8216 11996 8280 12000
rect 8216 11940 8220 11996
rect 8220 11940 8276 11996
rect 8276 11940 8280 11996
rect 8216 11936 8280 11940
rect 8296 11996 8360 12000
rect 8296 11940 8300 11996
rect 8300 11940 8356 11996
rect 8356 11940 8360 11996
rect 8296 11936 8360 11940
rect 8376 11996 8440 12000
rect 8376 11940 8380 11996
rect 8380 11940 8436 11996
rect 8436 11940 8440 11996
rect 8376 11936 8440 11940
rect 8456 11996 8520 12000
rect 8456 11940 8460 11996
rect 8460 11940 8516 11996
rect 8516 11940 8520 11996
rect 8456 11936 8520 11940
rect 4216 11452 4280 11456
rect 4216 11396 4220 11452
rect 4220 11396 4276 11452
rect 4276 11396 4280 11452
rect 4216 11392 4280 11396
rect 4296 11452 4360 11456
rect 4296 11396 4300 11452
rect 4300 11396 4356 11452
rect 4356 11396 4360 11452
rect 4296 11392 4360 11396
rect 4376 11452 4440 11456
rect 4376 11396 4380 11452
rect 4380 11396 4436 11452
rect 4436 11396 4440 11452
rect 4376 11392 4440 11396
rect 4456 11452 4520 11456
rect 4456 11396 4460 11452
rect 4460 11396 4516 11452
rect 4516 11396 4520 11452
rect 4456 11392 4520 11396
rect 12216 11452 12280 11456
rect 12216 11396 12220 11452
rect 12220 11396 12276 11452
rect 12276 11396 12280 11452
rect 12216 11392 12280 11396
rect 12296 11452 12360 11456
rect 12296 11396 12300 11452
rect 12300 11396 12356 11452
rect 12356 11396 12360 11452
rect 12296 11392 12360 11396
rect 12376 11452 12440 11456
rect 12376 11396 12380 11452
rect 12380 11396 12436 11452
rect 12436 11396 12440 11452
rect 12376 11392 12440 11396
rect 12456 11452 12520 11456
rect 12456 11396 12460 11452
rect 12460 11396 12516 11452
rect 12516 11396 12520 11452
rect 12456 11392 12520 11396
rect 8216 10908 8280 10912
rect 8216 10852 8220 10908
rect 8220 10852 8276 10908
rect 8276 10852 8280 10908
rect 8216 10848 8280 10852
rect 8296 10908 8360 10912
rect 8296 10852 8300 10908
rect 8300 10852 8356 10908
rect 8356 10852 8360 10908
rect 8296 10848 8360 10852
rect 8376 10908 8440 10912
rect 8376 10852 8380 10908
rect 8380 10852 8436 10908
rect 8436 10852 8440 10908
rect 8376 10848 8440 10852
rect 8456 10908 8520 10912
rect 8456 10852 8460 10908
rect 8460 10852 8516 10908
rect 8516 10852 8520 10908
rect 8456 10848 8520 10852
rect 4216 10364 4280 10368
rect 4216 10308 4220 10364
rect 4220 10308 4276 10364
rect 4276 10308 4280 10364
rect 4216 10304 4280 10308
rect 4296 10364 4360 10368
rect 4296 10308 4300 10364
rect 4300 10308 4356 10364
rect 4356 10308 4360 10364
rect 4296 10304 4360 10308
rect 4376 10364 4440 10368
rect 4376 10308 4380 10364
rect 4380 10308 4436 10364
rect 4436 10308 4440 10364
rect 4376 10304 4440 10308
rect 4456 10364 4520 10368
rect 4456 10308 4460 10364
rect 4460 10308 4516 10364
rect 4516 10308 4520 10364
rect 4456 10304 4520 10308
rect 12216 10364 12280 10368
rect 12216 10308 12220 10364
rect 12220 10308 12276 10364
rect 12276 10308 12280 10364
rect 12216 10304 12280 10308
rect 12296 10364 12360 10368
rect 12296 10308 12300 10364
rect 12300 10308 12356 10364
rect 12356 10308 12360 10364
rect 12296 10304 12360 10308
rect 12376 10364 12440 10368
rect 12376 10308 12380 10364
rect 12380 10308 12436 10364
rect 12436 10308 12440 10364
rect 12376 10304 12440 10308
rect 12456 10364 12520 10368
rect 12456 10308 12460 10364
rect 12460 10308 12516 10364
rect 12516 10308 12520 10364
rect 12456 10304 12520 10308
rect 8708 9964 8772 10028
rect 8216 9820 8280 9824
rect 8216 9764 8220 9820
rect 8220 9764 8276 9820
rect 8276 9764 8280 9820
rect 8216 9760 8280 9764
rect 8296 9820 8360 9824
rect 8296 9764 8300 9820
rect 8300 9764 8356 9820
rect 8356 9764 8360 9820
rect 8296 9760 8360 9764
rect 8376 9820 8440 9824
rect 8376 9764 8380 9820
rect 8380 9764 8436 9820
rect 8436 9764 8440 9820
rect 8376 9760 8440 9764
rect 8456 9820 8520 9824
rect 8456 9764 8460 9820
rect 8460 9764 8516 9820
rect 8516 9764 8520 9820
rect 8456 9760 8520 9764
rect 8708 9420 8772 9484
rect 4216 9276 4280 9280
rect 4216 9220 4220 9276
rect 4220 9220 4276 9276
rect 4276 9220 4280 9276
rect 4216 9216 4280 9220
rect 4296 9276 4360 9280
rect 4296 9220 4300 9276
rect 4300 9220 4356 9276
rect 4356 9220 4360 9276
rect 4296 9216 4360 9220
rect 4376 9276 4440 9280
rect 4376 9220 4380 9276
rect 4380 9220 4436 9276
rect 4436 9220 4440 9276
rect 4376 9216 4440 9220
rect 4456 9276 4520 9280
rect 4456 9220 4460 9276
rect 4460 9220 4516 9276
rect 4516 9220 4520 9276
rect 4456 9216 4520 9220
rect 12216 9276 12280 9280
rect 12216 9220 12220 9276
rect 12220 9220 12276 9276
rect 12276 9220 12280 9276
rect 12216 9216 12280 9220
rect 12296 9276 12360 9280
rect 12296 9220 12300 9276
rect 12300 9220 12356 9276
rect 12356 9220 12360 9276
rect 12296 9216 12360 9220
rect 12376 9276 12440 9280
rect 12376 9220 12380 9276
rect 12380 9220 12436 9276
rect 12436 9220 12440 9276
rect 12376 9216 12440 9220
rect 12456 9276 12520 9280
rect 12456 9220 12460 9276
rect 12460 9220 12516 9276
rect 12516 9220 12520 9276
rect 12456 9216 12520 9220
rect 8216 8732 8280 8736
rect 8216 8676 8220 8732
rect 8220 8676 8276 8732
rect 8276 8676 8280 8732
rect 8216 8672 8280 8676
rect 8296 8732 8360 8736
rect 8296 8676 8300 8732
rect 8300 8676 8356 8732
rect 8356 8676 8360 8732
rect 8296 8672 8360 8676
rect 8376 8732 8440 8736
rect 8376 8676 8380 8732
rect 8380 8676 8436 8732
rect 8436 8676 8440 8732
rect 8376 8672 8440 8676
rect 8456 8732 8520 8736
rect 8456 8676 8460 8732
rect 8460 8676 8516 8732
rect 8516 8676 8520 8732
rect 8456 8672 8520 8676
rect 4216 8188 4280 8192
rect 4216 8132 4220 8188
rect 4220 8132 4276 8188
rect 4276 8132 4280 8188
rect 4216 8128 4280 8132
rect 4296 8188 4360 8192
rect 4296 8132 4300 8188
rect 4300 8132 4356 8188
rect 4356 8132 4360 8188
rect 4296 8128 4360 8132
rect 4376 8188 4440 8192
rect 4376 8132 4380 8188
rect 4380 8132 4436 8188
rect 4436 8132 4440 8188
rect 4376 8128 4440 8132
rect 4456 8188 4520 8192
rect 4456 8132 4460 8188
rect 4460 8132 4516 8188
rect 4516 8132 4520 8188
rect 4456 8128 4520 8132
rect 12216 8188 12280 8192
rect 12216 8132 12220 8188
rect 12220 8132 12276 8188
rect 12276 8132 12280 8188
rect 12216 8128 12280 8132
rect 12296 8188 12360 8192
rect 12296 8132 12300 8188
rect 12300 8132 12356 8188
rect 12356 8132 12360 8188
rect 12296 8128 12360 8132
rect 12376 8188 12440 8192
rect 12376 8132 12380 8188
rect 12380 8132 12436 8188
rect 12436 8132 12440 8188
rect 12376 8128 12440 8132
rect 12456 8188 12520 8192
rect 12456 8132 12460 8188
rect 12460 8132 12516 8188
rect 12516 8132 12520 8188
rect 12456 8128 12520 8132
rect 8216 7644 8280 7648
rect 8216 7588 8220 7644
rect 8220 7588 8276 7644
rect 8276 7588 8280 7644
rect 8216 7584 8280 7588
rect 8296 7644 8360 7648
rect 8296 7588 8300 7644
rect 8300 7588 8356 7644
rect 8356 7588 8360 7644
rect 8296 7584 8360 7588
rect 8376 7644 8440 7648
rect 8376 7588 8380 7644
rect 8380 7588 8436 7644
rect 8436 7588 8440 7644
rect 8376 7584 8440 7588
rect 8456 7644 8520 7648
rect 8456 7588 8460 7644
rect 8460 7588 8516 7644
rect 8516 7588 8520 7644
rect 8456 7584 8520 7588
rect 4216 7100 4280 7104
rect 4216 7044 4220 7100
rect 4220 7044 4276 7100
rect 4276 7044 4280 7100
rect 4216 7040 4280 7044
rect 4296 7100 4360 7104
rect 4296 7044 4300 7100
rect 4300 7044 4356 7100
rect 4356 7044 4360 7100
rect 4296 7040 4360 7044
rect 4376 7100 4440 7104
rect 4376 7044 4380 7100
rect 4380 7044 4436 7100
rect 4436 7044 4440 7100
rect 4376 7040 4440 7044
rect 4456 7100 4520 7104
rect 4456 7044 4460 7100
rect 4460 7044 4516 7100
rect 4516 7044 4520 7100
rect 4456 7040 4520 7044
rect 12216 7100 12280 7104
rect 12216 7044 12220 7100
rect 12220 7044 12276 7100
rect 12276 7044 12280 7100
rect 12216 7040 12280 7044
rect 12296 7100 12360 7104
rect 12296 7044 12300 7100
rect 12300 7044 12356 7100
rect 12356 7044 12360 7100
rect 12296 7040 12360 7044
rect 12376 7100 12440 7104
rect 12376 7044 12380 7100
rect 12380 7044 12436 7100
rect 12436 7044 12440 7100
rect 12376 7040 12440 7044
rect 12456 7100 12520 7104
rect 12456 7044 12460 7100
rect 12460 7044 12516 7100
rect 12516 7044 12520 7100
rect 12456 7040 12520 7044
rect 8216 6556 8280 6560
rect 8216 6500 8220 6556
rect 8220 6500 8276 6556
rect 8276 6500 8280 6556
rect 8216 6496 8280 6500
rect 8296 6556 8360 6560
rect 8296 6500 8300 6556
rect 8300 6500 8356 6556
rect 8356 6500 8360 6556
rect 8296 6496 8360 6500
rect 8376 6556 8440 6560
rect 8376 6500 8380 6556
rect 8380 6500 8436 6556
rect 8436 6500 8440 6556
rect 8376 6496 8440 6500
rect 8456 6556 8520 6560
rect 8456 6500 8460 6556
rect 8460 6500 8516 6556
rect 8516 6500 8520 6556
rect 8456 6496 8520 6500
rect 4216 6012 4280 6016
rect 4216 5956 4220 6012
rect 4220 5956 4276 6012
rect 4276 5956 4280 6012
rect 4216 5952 4280 5956
rect 4296 6012 4360 6016
rect 4296 5956 4300 6012
rect 4300 5956 4356 6012
rect 4356 5956 4360 6012
rect 4296 5952 4360 5956
rect 4376 6012 4440 6016
rect 4376 5956 4380 6012
rect 4380 5956 4436 6012
rect 4436 5956 4440 6012
rect 4376 5952 4440 5956
rect 4456 6012 4520 6016
rect 4456 5956 4460 6012
rect 4460 5956 4516 6012
rect 4516 5956 4520 6012
rect 4456 5952 4520 5956
rect 12216 6012 12280 6016
rect 12216 5956 12220 6012
rect 12220 5956 12276 6012
rect 12276 5956 12280 6012
rect 12216 5952 12280 5956
rect 12296 6012 12360 6016
rect 12296 5956 12300 6012
rect 12300 5956 12356 6012
rect 12356 5956 12360 6012
rect 12296 5952 12360 5956
rect 12376 6012 12440 6016
rect 12376 5956 12380 6012
rect 12380 5956 12436 6012
rect 12436 5956 12440 6012
rect 12376 5952 12440 5956
rect 12456 6012 12520 6016
rect 12456 5956 12460 6012
rect 12460 5956 12516 6012
rect 12516 5956 12520 6012
rect 12456 5952 12520 5956
rect 8216 5468 8280 5472
rect 8216 5412 8220 5468
rect 8220 5412 8276 5468
rect 8276 5412 8280 5468
rect 8216 5408 8280 5412
rect 8296 5468 8360 5472
rect 8296 5412 8300 5468
rect 8300 5412 8356 5468
rect 8356 5412 8360 5468
rect 8296 5408 8360 5412
rect 8376 5468 8440 5472
rect 8376 5412 8380 5468
rect 8380 5412 8436 5468
rect 8436 5412 8440 5468
rect 8376 5408 8440 5412
rect 8456 5468 8520 5472
rect 8456 5412 8460 5468
rect 8460 5412 8516 5468
rect 8516 5412 8520 5468
rect 8456 5408 8520 5412
rect 4216 4924 4280 4928
rect 4216 4868 4220 4924
rect 4220 4868 4276 4924
rect 4276 4868 4280 4924
rect 4216 4864 4280 4868
rect 4296 4924 4360 4928
rect 4296 4868 4300 4924
rect 4300 4868 4356 4924
rect 4356 4868 4360 4924
rect 4296 4864 4360 4868
rect 4376 4924 4440 4928
rect 4376 4868 4380 4924
rect 4380 4868 4436 4924
rect 4436 4868 4440 4924
rect 4376 4864 4440 4868
rect 4456 4924 4520 4928
rect 4456 4868 4460 4924
rect 4460 4868 4516 4924
rect 4516 4868 4520 4924
rect 4456 4864 4520 4868
rect 12216 4924 12280 4928
rect 12216 4868 12220 4924
rect 12220 4868 12276 4924
rect 12276 4868 12280 4924
rect 12216 4864 12280 4868
rect 12296 4924 12360 4928
rect 12296 4868 12300 4924
rect 12300 4868 12356 4924
rect 12356 4868 12360 4924
rect 12296 4864 12360 4868
rect 12376 4924 12440 4928
rect 12376 4868 12380 4924
rect 12380 4868 12436 4924
rect 12436 4868 12440 4924
rect 12376 4864 12440 4868
rect 12456 4924 12520 4928
rect 12456 4868 12460 4924
rect 12460 4868 12516 4924
rect 12516 4868 12520 4924
rect 12456 4864 12520 4868
rect 8216 4380 8280 4384
rect 8216 4324 8220 4380
rect 8220 4324 8276 4380
rect 8276 4324 8280 4380
rect 8216 4320 8280 4324
rect 8296 4380 8360 4384
rect 8296 4324 8300 4380
rect 8300 4324 8356 4380
rect 8356 4324 8360 4380
rect 8296 4320 8360 4324
rect 8376 4380 8440 4384
rect 8376 4324 8380 4380
rect 8380 4324 8436 4380
rect 8436 4324 8440 4380
rect 8376 4320 8440 4324
rect 8456 4380 8520 4384
rect 8456 4324 8460 4380
rect 8460 4324 8516 4380
rect 8516 4324 8520 4380
rect 8456 4320 8520 4324
rect 4216 3836 4280 3840
rect 4216 3780 4220 3836
rect 4220 3780 4276 3836
rect 4276 3780 4280 3836
rect 4216 3776 4280 3780
rect 4296 3836 4360 3840
rect 4296 3780 4300 3836
rect 4300 3780 4356 3836
rect 4356 3780 4360 3836
rect 4296 3776 4360 3780
rect 4376 3836 4440 3840
rect 4376 3780 4380 3836
rect 4380 3780 4436 3836
rect 4436 3780 4440 3836
rect 4376 3776 4440 3780
rect 4456 3836 4520 3840
rect 4456 3780 4460 3836
rect 4460 3780 4516 3836
rect 4516 3780 4520 3836
rect 4456 3776 4520 3780
rect 12216 3836 12280 3840
rect 12216 3780 12220 3836
rect 12220 3780 12276 3836
rect 12276 3780 12280 3836
rect 12216 3776 12280 3780
rect 12296 3836 12360 3840
rect 12296 3780 12300 3836
rect 12300 3780 12356 3836
rect 12356 3780 12360 3836
rect 12296 3776 12360 3780
rect 12376 3836 12440 3840
rect 12376 3780 12380 3836
rect 12380 3780 12436 3836
rect 12436 3780 12440 3836
rect 12376 3776 12440 3780
rect 12456 3836 12520 3840
rect 12456 3780 12460 3836
rect 12460 3780 12516 3836
rect 12516 3780 12520 3836
rect 12456 3776 12520 3780
rect 8216 3292 8280 3296
rect 8216 3236 8220 3292
rect 8220 3236 8276 3292
rect 8276 3236 8280 3292
rect 8216 3232 8280 3236
rect 8296 3292 8360 3296
rect 8296 3236 8300 3292
rect 8300 3236 8356 3292
rect 8356 3236 8360 3292
rect 8296 3232 8360 3236
rect 8376 3292 8440 3296
rect 8376 3236 8380 3292
rect 8380 3236 8436 3292
rect 8436 3236 8440 3292
rect 8376 3232 8440 3236
rect 8456 3292 8520 3296
rect 8456 3236 8460 3292
rect 8460 3236 8516 3292
rect 8516 3236 8520 3292
rect 8456 3232 8520 3236
rect 4216 2748 4280 2752
rect 4216 2692 4220 2748
rect 4220 2692 4276 2748
rect 4276 2692 4280 2748
rect 4216 2688 4280 2692
rect 4296 2748 4360 2752
rect 4296 2692 4300 2748
rect 4300 2692 4356 2748
rect 4356 2692 4360 2748
rect 4296 2688 4360 2692
rect 4376 2748 4440 2752
rect 4376 2692 4380 2748
rect 4380 2692 4436 2748
rect 4436 2692 4440 2748
rect 4376 2688 4440 2692
rect 4456 2748 4520 2752
rect 4456 2692 4460 2748
rect 4460 2692 4516 2748
rect 4516 2692 4520 2748
rect 4456 2688 4520 2692
rect 12216 2748 12280 2752
rect 12216 2692 12220 2748
rect 12220 2692 12276 2748
rect 12276 2692 12280 2748
rect 12216 2688 12280 2692
rect 12296 2748 12360 2752
rect 12296 2692 12300 2748
rect 12300 2692 12356 2748
rect 12356 2692 12360 2748
rect 12296 2688 12360 2692
rect 12376 2748 12440 2752
rect 12376 2692 12380 2748
rect 12380 2692 12436 2748
rect 12436 2692 12440 2748
rect 12376 2688 12440 2692
rect 12456 2748 12520 2752
rect 12456 2692 12460 2748
rect 12460 2692 12516 2748
rect 12516 2692 12520 2748
rect 12456 2688 12520 2692
rect 8216 2204 8280 2208
rect 8216 2148 8220 2204
rect 8220 2148 8276 2204
rect 8276 2148 8280 2204
rect 8216 2144 8280 2148
rect 8296 2204 8360 2208
rect 8296 2148 8300 2204
rect 8300 2148 8356 2204
rect 8356 2148 8360 2204
rect 8296 2144 8360 2148
rect 8376 2204 8440 2208
rect 8376 2148 8380 2204
rect 8380 2148 8436 2204
rect 8436 2148 8440 2204
rect 8376 2144 8440 2148
rect 8456 2204 8520 2208
rect 8456 2148 8460 2204
rect 8460 2148 8516 2204
rect 8516 2148 8520 2204
rect 8456 2144 8520 2148
rect 4216 1660 4280 1664
rect 4216 1604 4220 1660
rect 4220 1604 4276 1660
rect 4276 1604 4280 1660
rect 4216 1600 4280 1604
rect 4296 1660 4360 1664
rect 4296 1604 4300 1660
rect 4300 1604 4356 1660
rect 4356 1604 4360 1660
rect 4296 1600 4360 1604
rect 4376 1660 4440 1664
rect 4376 1604 4380 1660
rect 4380 1604 4436 1660
rect 4436 1604 4440 1660
rect 4376 1600 4440 1604
rect 4456 1660 4520 1664
rect 4456 1604 4460 1660
rect 4460 1604 4516 1660
rect 4516 1604 4520 1660
rect 4456 1600 4520 1604
rect 12216 1660 12280 1664
rect 12216 1604 12220 1660
rect 12220 1604 12276 1660
rect 12276 1604 12280 1660
rect 12216 1600 12280 1604
rect 12296 1660 12360 1664
rect 12296 1604 12300 1660
rect 12300 1604 12356 1660
rect 12356 1604 12360 1660
rect 12296 1600 12360 1604
rect 12376 1660 12440 1664
rect 12376 1604 12380 1660
rect 12380 1604 12436 1660
rect 12436 1604 12440 1660
rect 12376 1600 12440 1604
rect 12456 1660 12520 1664
rect 12456 1604 12460 1660
rect 12460 1604 12516 1660
rect 12516 1604 12520 1660
rect 12456 1600 12520 1604
rect 8216 1116 8280 1120
rect 8216 1060 8220 1116
rect 8220 1060 8276 1116
rect 8276 1060 8280 1116
rect 8216 1056 8280 1060
rect 8296 1116 8360 1120
rect 8296 1060 8300 1116
rect 8300 1060 8356 1116
rect 8356 1060 8360 1116
rect 8296 1056 8360 1060
rect 8376 1116 8440 1120
rect 8376 1060 8380 1116
rect 8380 1060 8436 1116
rect 8436 1060 8440 1116
rect 8376 1056 8440 1060
rect 8456 1116 8520 1120
rect 8456 1060 8460 1116
rect 8460 1060 8516 1116
rect 8516 1060 8520 1116
rect 8456 1056 8520 1060
<< metal4 >>
rect 4208 13632 4528 13648
rect 4208 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4528 13632
rect 4208 12544 4528 13568
rect 4208 12480 4216 12544
rect 4280 12488 4296 12544
rect 4360 12488 4376 12544
rect 4440 12488 4456 12544
rect 4520 12480 4528 12544
rect 4208 12252 4250 12480
rect 4486 12252 4528 12480
rect 4208 11456 4528 12252
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 4208 10368 4528 11392
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 4208 9280 4528 10304
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 8192 4528 9216
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 7104 4528 8128
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 6016 4528 7040
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 4928 4528 5952
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 4488 4528 4864
rect 4208 4252 4250 4488
rect 4486 4252 4528 4488
rect 4208 3840 4528 4252
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 2752 4528 3776
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 1664 4528 2688
rect 4208 1600 4216 1664
rect 4280 1600 4296 1664
rect 4360 1600 4376 1664
rect 4440 1600 4456 1664
rect 4520 1600 4528 1664
rect 4208 1040 4528 1600
rect 8208 13088 8528 13648
rect 8208 13024 8216 13088
rect 8280 13024 8296 13088
rect 8360 13024 8376 13088
rect 8440 13024 8456 13088
rect 8520 13024 8528 13088
rect 8208 12000 8528 13024
rect 8208 11936 8216 12000
rect 8280 11936 8296 12000
rect 8360 11936 8376 12000
rect 8440 11936 8456 12000
rect 8520 11936 8528 12000
rect 8208 10912 8528 11936
rect 8208 10848 8216 10912
rect 8280 10848 8296 10912
rect 8360 10848 8376 10912
rect 8440 10848 8456 10912
rect 8520 10848 8528 10912
rect 8208 9824 8528 10848
rect 12208 13632 12528 13648
rect 12208 13568 12216 13632
rect 12280 13568 12296 13632
rect 12360 13568 12376 13632
rect 12440 13568 12456 13632
rect 12520 13568 12528 13632
rect 12208 12544 12528 13568
rect 12208 12480 12216 12544
rect 12280 12488 12296 12544
rect 12360 12488 12376 12544
rect 12440 12488 12456 12544
rect 12520 12480 12528 12544
rect 12208 12252 12250 12480
rect 12486 12252 12528 12480
rect 12208 11456 12528 12252
rect 12208 11392 12216 11456
rect 12280 11392 12296 11456
rect 12360 11392 12376 11456
rect 12440 11392 12456 11456
rect 12520 11392 12528 11456
rect 12208 10368 12528 11392
rect 12208 10304 12216 10368
rect 12280 10304 12296 10368
rect 12360 10304 12376 10368
rect 12440 10304 12456 10368
rect 12520 10304 12528 10368
rect 8707 10028 8773 10029
rect 8707 9964 8708 10028
rect 8772 9964 8773 10028
rect 8707 9963 8773 9964
rect 8208 9760 8216 9824
rect 8280 9760 8296 9824
rect 8360 9760 8376 9824
rect 8440 9760 8456 9824
rect 8520 9760 8528 9824
rect 8208 8736 8528 9760
rect 8710 9485 8770 9963
rect 8707 9484 8773 9485
rect 8707 9420 8708 9484
rect 8772 9420 8773 9484
rect 8707 9419 8773 9420
rect 8208 8672 8216 8736
rect 8280 8672 8296 8736
rect 8360 8672 8376 8736
rect 8440 8672 8456 8736
rect 8520 8672 8528 8736
rect 8208 8488 8528 8672
rect 8208 8252 8250 8488
rect 8486 8252 8528 8488
rect 8208 7648 8528 8252
rect 8208 7584 8216 7648
rect 8280 7584 8296 7648
rect 8360 7584 8376 7648
rect 8440 7584 8456 7648
rect 8520 7584 8528 7648
rect 8208 6560 8528 7584
rect 8208 6496 8216 6560
rect 8280 6496 8296 6560
rect 8360 6496 8376 6560
rect 8440 6496 8456 6560
rect 8520 6496 8528 6560
rect 8208 5472 8528 6496
rect 8208 5408 8216 5472
rect 8280 5408 8296 5472
rect 8360 5408 8376 5472
rect 8440 5408 8456 5472
rect 8520 5408 8528 5472
rect 8208 4384 8528 5408
rect 8208 4320 8216 4384
rect 8280 4320 8296 4384
rect 8360 4320 8376 4384
rect 8440 4320 8456 4384
rect 8520 4320 8528 4384
rect 8208 3296 8528 4320
rect 8208 3232 8216 3296
rect 8280 3232 8296 3296
rect 8360 3232 8376 3296
rect 8440 3232 8456 3296
rect 8520 3232 8528 3296
rect 8208 2208 8528 3232
rect 8208 2144 8216 2208
rect 8280 2144 8296 2208
rect 8360 2144 8376 2208
rect 8440 2144 8456 2208
rect 8520 2144 8528 2208
rect 8208 1120 8528 2144
rect 8208 1056 8216 1120
rect 8280 1056 8296 1120
rect 8360 1056 8376 1120
rect 8440 1056 8456 1120
rect 8520 1056 8528 1120
rect 8208 1040 8528 1056
rect 12208 9280 12528 10304
rect 12208 9216 12216 9280
rect 12280 9216 12296 9280
rect 12360 9216 12376 9280
rect 12440 9216 12456 9280
rect 12520 9216 12528 9280
rect 12208 8192 12528 9216
rect 12208 8128 12216 8192
rect 12280 8128 12296 8192
rect 12360 8128 12376 8192
rect 12440 8128 12456 8192
rect 12520 8128 12528 8192
rect 12208 7104 12528 8128
rect 12208 7040 12216 7104
rect 12280 7040 12296 7104
rect 12360 7040 12376 7104
rect 12440 7040 12456 7104
rect 12520 7040 12528 7104
rect 12208 6016 12528 7040
rect 12208 5952 12216 6016
rect 12280 5952 12296 6016
rect 12360 5952 12376 6016
rect 12440 5952 12456 6016
rect 12520 5952 12528 6016
rect 12208 4928 12528 5952
rect 12208 4864 12216 4928
rect 12280 4864 12296 4928
rect 12360 4864 12376 4928
rect 12440 4864 12456 4928
rect 12520 4864 12528 4928
rect 12208 4488 12528 4864
rect 12208 4252 12250 4488
rect 12486 4252 12528 4488
rect 12208 3840 12528 4252
rect 12208 3776 12216 3840
rect 12280 3776 12296 3840
rect 12360 3776 12376 3840
rect 12440 3776 12456 3840
rect 12520 3776 12528 3840
rect 12208 2752 12528 3776
rect 12208 2688 12216 2752
rect 12280 2688 12296 2752
rect 12360 2688 12376 2752
rect 12440 2688 12456 2752
rect 12520 2688 12528 2752
rect 12208 1664 12528 2688
rect 12208 1600 12216 1664
rect 12280 1600 12296 1664
rect 12360 1600 12376 1664
rect 12440 1600 12456 1664
rect 12520 1600 12528 1664
rect 12208 1040 12528 1600
<< via4 >>
rect 4250 12480 4280 12488
rect 4280 12480 4296 12488
rect 4296 12480 4360 12488
rect 4360 12480 4376 12488
rect 4376 12480 4440 12488
rect 4440 12480 4456 12488
rect 4456 12480 4486 12488
rect 4250 12252 4486 12480
rect 4250 4252 4486 4488
rect 12250 12480 12280 12488
rect 12280 12480 12296 12488
rect 12296 12480 12360 12488
rect 12360 12480 12376 12488
rect 12376 12480 12440 12488
rect 12440 12480 12456 12488
rect 12456 12480 12486 12488
rect 12250 12252 12486 12480
rect 8250 8252 8486 8488
rect 12250 4252 12486 4488
<< metal5 >>
rect 1056 12488 13940 12530
rect 1056 12252 4250 12488
rect 4486 12252 12250 12488
rect 12486 12252 13940 12488
rect 1056 12210 13940 12252
rect 1056 8488 13940 8530
rect 1056 8252 8250 8488
rect 8486 8252 13940 8488
rect 1056 8210 13940 8252
rect 1056 4488 13940 4530
rect 1056 4252 4250 4488
rect 4486 4252 12250 4488
rect 12486 4252 13940 4488
rect 1056 4210 13940 4252
use sky130_fd_sc_hd__diode_2  ANTENNA__207__A1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform 1 0 1564 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__213__A1
timestamp 1665323087
transform -1 0 4968 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__213__B1
timestamp 1665323087
transform -1 0 3956 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__214__B1
timestamp 1665323087
transform 1 0 1380 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__215__B1
timestamp 1665323087
transform -1 0 2668 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__216__A
timestamp 1665323087
transform -1 0 3680 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__219__A
timestamp 1665323087
transform -1 0 6624 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__222__A1
timestamp 1665323087
transform -1 0 6808 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__222__B2
timestamp 1665323087
transform -1 0 5152 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__225__B1
timestamp 1665323087
transform 1 0 1380 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__235__A
timestamp 1665323087
transform -1 0 1656 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__288__A
timestamp 1665323087
transform 1 0 7268 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__289__A1
timestamp 1665323087
transform -1 0 2300 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__289__A2
timestamp 1665323087
transform 1 0 3404 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__293__A_N
timestamp 1665323087
transform 1 0 6532 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__295__A1
timestamp 1665323087
transform 1 0 2668 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__295__A2
timestamp 1665323087
transform -1 0 2300 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__296__B
timestamp 1665323087
transform 1 0 10764 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__299__A1
timestamp 1665323087
transform 1 0 1380 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__299__A2
timestamp 1665323087
transform -1 0 1564 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__300__A1
timestamp 1665323087
transform 1 0 1380 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__300__A2
timestamp 1665323087
transform -1 0 1564 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__302__A1
timestamp 1665323087
transform 1 0 3956 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__302__A2
timestamp 1665323087
transform -1 0 3588 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__305__A1
timestamp 1665323087
transform 1 0 3128 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__305__A2
timestamp 1665323087
transform -1 0 1748 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__306__A1
timestamp 1665323087
transform 1 0 1380 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__306__A2
timestamp 1665323087
transform 1 0 1380 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__309__A1
timestamp 1665323087
transform 1 0 4416 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__309__A2
timestamp 1665323087
transform 1 0 2208 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__310__A1
timestamp 1665323087
transform 1 0 5704 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__310__A2
timestamp 1665323087
transform 1 0 4600 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__312__A1
timestamp 1665323087
transform 1 0 6532 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__312__A2
timestamp 1665323087
transform 1 0 6348 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__313__A_N
timestamp 1665323087
transform -1 0 3496 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__313__B
timestamp 1665323087
transform 1 0 3496 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__314__A1
timestamp 1665323087
transform 1 0 6348 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__316__B1
timestamp 1665323087
transform -1 0 3772 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__316__B2
timestamp 1665323087
transform 1 0 4048 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__317__A1
timestamp 1665323087
transform 1 0 4876 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__317__A2
timestamp 1665323087
transform -1 0 4876 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__319__A1
timestamp 1665323087
transform 1 0 5704 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__319__A2
timestamp 1665323087
transform -1 0 7268 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__326__A1
timestamp 1665323087
transform 1 0 7360 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__326__A2
timestamp 1665323087
transform -1 0 9568 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__334__B1
timestamp 1665323087
transform 1 0 10120 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__334__B2
timestamp 1665323087
transform 1 0 9568 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__337__A1
timestamp 1665323087
transform 1 0 13432 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__337__A2
timestamp 1665323087
transform -1 0 9016 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__341__B1
timestamp 1665323087
transform -1 0 9292 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__341__B2
timestamp 1665323087
transform 1 0 9292 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__342__A1
timestamp 1665323087
transform 1 0 11960 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__342__A2
timestamp 1665323087
transform -1 0 13616 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__343__A1
timestamp 1665323087
transform 1 0 10304 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__343__A2
timestamp 1665323087
transform 1 0 10120 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__346__B1
timestamp 1665323087
transform 1 0 8832 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__346__B2
timestamp 1665323087
transform 1 0 7820 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__348__A1
timestamp 1665323087
transform 1 0 11868 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__348__A2
timestamp 1665323087
transform 1 0 13432 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__350__B1
timestamp 1665323087
transform -1 0 9108 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__350__B2
timestamp 1665323087
transform 1 0 9108 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__351__A1
timestamp 1665323087
transform 1 0 11224 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__351__A2
timestamp 1665323087
transform 1 0 13432 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__352__A_N
timestamp 1665323087
transform 1 0 11592 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__353__A1
timestamp 1665323087
transform 1 0 13064 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__353__A2
timestamp 1665323087
transform 1 0 13248 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__354__A1
timestamp 1665323087
transform 1 0 11040 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__354__A2
timestamp 1665323087
transform -1 0 11224 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__355__A
timestamp 1665323087
transform -1 0 6532 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__355__B
timestamp 1665323087
transform -1 0 6716 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__356__A
timestamp 1665323087
transform 1 0 8648 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__357__A
timestamp 1665323087
transform 1 0 8648 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__358__A
timestamp 1665323087
transform 1 0 12880 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__359__A
timestamp 1665323087
transform 1 0 6348 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__360__A
timestamp 1665323087
transform 1 0 8372 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__361__A
timestamp 1665323087
transform 1 0 8464 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__362__A
timestamp 1665323087
transform 1 0 5612 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__363__A
timestamp 1665323087
transform 1 0 5980 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__364__A
timestamp 1665323087
transform 1 0 11040 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__365__A
timestamp 1665323087
transform 1 0 6256 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__366__A
timestamp 1665323087
transform 1 0 12696 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__367__A
timestamp 1665323087
transform 1 0 12420 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__368__A
timestamp 1665323087
transform 1 0 13340 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__369__A
timestamp 1665323087
transform 1 0 11224 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__370__A
timestamp 1665323087
transform 1 0 6900 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__371__A
timestamp 1665323087
transform 1 0 13432 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__372__A
timestamp 1665323087
transform 1 0 13064 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__373__A
timestamp 1665323087
transform 1 0 11224 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__374__A
timestamp 1665323087
transform 1 0 8188 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__375__A
timestamp 1665323087
transform 1 0 3588 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__376__A
timestamp 1665323087
transform 1 0 3680 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__377__A
timestamp 1665323087
transform 1 0 4232 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__378__A
timestamp 1665323087
transform 1 0 3772 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__394__D
timestamp 1665323087
transform -1 0 13616 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_81 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform 1 0 8556 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_90
timestamp 1665323087
transform 1 0 9384 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_3
timestamp 1665323087
transform 1 0 1380 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_50
timestamp 1665323087
transform 1 0 5704 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_59
timestamp 1665323087
transform 1 0 6532 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_3
timestamp 1665323087
transform 1 0 1380 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_35
timestamp 1665323087
transform 1 0 4324 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_2_79 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform 1 0 8372 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_2_99
timestamp 1665323087
transform 1 0 10212 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_134 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform 1 0 13432 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_3_3
timestamp 1665323087
transform 1 0 1380 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_3_49
timestamp 1665323087
transform 1 0 5612 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_76
timestamp 1665323087
transform 1 0 8096 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_3_99
timestamp 1665323087
transform 1 0 10212 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_3_109
timestamp 1665323087
transform 1 0 11132 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_3_118
timestamp 1665323087
transform 1 0 11960 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_132 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform 1 0 13248 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_31
timestamp 1665323087
transform 1 0 3956 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_55
timestamp 1665323087
transform 1 0 6164 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_62
timestamp 1665323087
transform 1 0 6808 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_90
timestamp 1665323087
transform 1 0 9384 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_132
timestamp 1665323087
transform 1 0 13248 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_78
timestamp 1665323087
transform 1 0 8280 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_5_87
timestamp 1665323087
transform 1 0 9108 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_134
timestamp 1665323087
transform 1 0 13432 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_95
timestamp 1665323087
transform 1 0 9844 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_6_120 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform 1 0 12144 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_41
timestamp 1665323087
transform 1 0 4876 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_47
timestamp 1665323087
transform 1 0 5428 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_55
timestamp 1665323087
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_89
timestamp 1665323087
transform 1 0 9292 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_7_113
timestamp 1665323087
transform 1 0 11500 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_124
timestamp 1665323087
transform 1 0 12512 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_8_24
timestamp 1665323087
transform 1 0 3312 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_8_42
timestamp 1665323087
transform 1 0 4968 0 1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_8_58 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform 1 0 6440 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_70
timestamp 1665323087
transform 1 0 7544 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_90
timestamp 1665323087
transform 1 0 9384 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_8_128
timestamp 1665323087
transform 1 0 12880 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_134
timestamp 1665323087
transform 1 0 13432 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_9_57
timestamp 1665323087
transform 1 0 6348 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_9_78
timestamp 1665323087
transform 1 0 8280 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_9_111
timestamp 1665323087
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_9_125
timestamp 1665323087
transform 1 0 12604 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_9_135
timestamp 1665323087
transform 1 0 13524 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_3
timestamp 1665323087
transform 1 0 1380 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_27
timestamp 1665323087
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_70
timestamp 1665323087
transform 1 0 7544 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_10_85
timestamp 1665323087
transform 1 0 8924 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_11_55
timestamp 1665323087
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_11_85
timestamp 1665323087
transform 1 0 8924 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_11_100
timestamp 1665323087
transform 1 0 10304 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_11_113
timestamp 1665323087
transform 1 0 11500 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_11_131
timestamp 1665323087
transform 1 0 13156 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_135
timestamp 1665323087
transform 1 0 13524 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_16
timestamp 1665323087
transform 1 0 2576 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_27
timestamp 1665323087
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_75
timestamp 1665323087
transform 1 0 8004 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_85
timestamp 1665323087
transform 1 0 8924 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_107
timestamp 1665323087
transform 1 0 10948 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_3
timestamp 1665323087
transform 1 0 1380 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_24
timestamp 1665323087
transform 1 0 3312 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_13_69
timestamp 1665323087
transform 1 0 7452 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_13_94
timestamp 1665323087
transform 1 0 9752 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_118
timestamp 1665323087
transform 1 0 11960 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_5
timestamp 1665323087
transform 1 0 1564 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_10
timestamp 1665323087
transform 1 0 2024 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_27
timestamp 1665323087
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_69
timestamp 1665323087
transform 1 0 7452 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_79
timestamp 1665323087
transform 1 0 8372 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_83
timestamp 1665323087
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_135
timestamp 1665323087
transform 1 0 13524 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_15_23
timestamp 1665323087
transform 1 0 3220 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_15_67
timestamp 1665323087
transform 1 0 7268 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_15_75
timestamp 1665323087
transform 1 0 8004 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_15_99
timestamp 1665323087
transform 1 0 10212 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_15_135
timestamp 1665323087
transform 1 0 13524 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_45
timestamp 1665323087
transform 1 0 5244 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_67
timestamp 1665323087
transform 1 0 7268 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_78
timestamp 1665323087
transform 1 0 8280 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_116
timestamp 1665323087
transform 1 0 11776 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_135
timestamp 1665323087
transform 1 0 13524 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_17_26
timestamp 1665323087
transform 1 0 3496 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_17_49
timestamp 1665323087
transform 1 0 5612 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_17_69
timestamp 1665323087
transform 1 0 7452 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_17_84
timestamp 1665323087
transform 1 0 8832 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_17_108
timestamp 1665323087
transform 1 0 11040 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_17_135
timestamp 1665323087
transform 1 0 13524 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_18_72
timestamp 1665323087
transform 1 0 7728 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_18_75
timestamp 1665323087
transform 1 0 8004 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_18_97
timestamp 1665323087
transform 1 0 10028 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_19_47
timestamp 1665323087
transform 1 0 5428 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_19_111
timestamp 1665323087
transform 1 0 11316 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_20_33
timestamp 1665323087
transform 1 0 4140 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_20_97
timestamp 1665323087
transform 1 0 10028 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_21_72
timestamp 1665323087
transform 1 0 7728 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_21_111
timestamp 1665323087
transform 1 0 11316 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_21_135
timestamp 1665323087
transform 1 0 13524 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_22_35
timestamp 1665323087
transform 1 0 4324 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_22_83
timestamp 1665323087
transform 1 0 8740 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_22_88
timestamp 1665323087
transform 1 0 9200 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_22_127
timestamp 1665323087
transform 1 0 12788 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1665323087
transform 1 0 1104 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1665323087
transform -1 0 13892 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1665323087
transform 1 0 1104 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1665323087
transform -1 0 13892 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1665323087
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1665323087
transform -1 0 13892 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1665323087
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1665323087
transform -1 0 13892 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1665323087
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1665323087
transform -1 0 13892 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1665323087
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1665323087
transform -1 0 13892 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1665323087
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1665323087
transform -1 0 13892 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1665323087
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1665323087
transform -1 0 13892 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1665323087
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1665323087
transform -1 0 13892 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1665323087
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1665323087
transform -1 0 13892 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1665323087
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1665323087
transform -1 0 13892 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1665323087
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1665323087
transform -1 0 13892 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1665323087
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1665323087
transform -1 0 13892 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1665323087
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1665323087
transform -1 0 13892 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1665323087
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1665323087
transform -1 0 13892 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1665323087
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1665323087
transform -1 0 13892 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1665323087
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1665323087
transform -1 0 13892 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1665323087
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1665323087
transform -1 0 13892 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1665323087
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1665323087
transform -1 0 13892 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1665323087
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1665323087
transform -1 0 13892 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1665323087
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1665323087
transform -1 0 13892 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1665323087
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1665323087
transform -1 0 13892 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1665323087
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1665323087
transform -1 0 13892 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_46 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform 1 0 3680 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_47
timestamp 1665323087
transform 1 0 6256 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_48
timestamp 1665323087
transform 1 0 8832 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_49
timestamp 1665323087
transform 1 0 11408 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_50
timestamp 1665323087
transform 1 0 6256 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_51
timestamp 1665323087
transform 1 0 11408 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_52
timestamp 1665323087
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_53
timestamp 1665323087
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_54
timestamp 1665323087
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_55
timestamp 1665323087
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_56
timestamp 1665323087
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_57
timestamp 1665323087
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_58
timestamp 1665323087
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_59
timestamp 1665323087
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_60
timestamp 1665323087
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_61
timestamp 1665323087
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_62
timestamp 1665323087
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_63
timestamp 1665323087
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_64
timestamp 1665323087
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_65
timestamp 1665323087
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_66
timestamp 1665323087
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_67
timestamp 1665323087
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_68
timestamp 1665323087
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_69
timestamp 1665323087
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_70
timestamp 1665323087
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_71
timestamp 1665323087
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_72
timestamp 1665323087
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_73
timestamp 1665323087
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_74
timestamp 1665323087
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_75
timestamp 1665323087
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_76
timestamp 1665323087
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_77
timestamp 1665323087
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_78
timestamp 1665323087
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_79
timestamp 1665323087
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_80
timestamp 1665323087
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_81
timestamp 1665323087
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_82
timestamp 1665323087
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_83
timestamp 1665323087
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_84
timestamp 1665323087
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_85
timestamp 1665323087
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_86
timestamp 1665323087
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_87
timestamp 1665323087
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_88
timestamp 1665323087
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_89
timestamp 1665323087
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_90
timestamp 1665323087
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_91
timestamp 1665323087
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_92
timestamp 1665323087
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_93
timestamp 1665323087
transform 1 0 6256 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_94
timestamp 1665323087
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_95
timestamp 1665323087
transform 1 0 11408 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _176_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform -1 0 11776 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _177_
timestamp 1665323087
transform 1 0 9476 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _178_
timestamp 1665323087
transform -1 0 9844 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _179_
timestamp 1665323087
transform 1 0 8096 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _180_
timestamp 1665323087
transform -1 0 11040 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_2  _181_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform -1 0 13248 0 -1 3264
box -38 -48 1234 592
use sky130_fd_sc_hd__xor2_2  _182_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform -1 0 13432 0 1 2176
box -38 -48 1234 592
use sky130_fd_sc_hd__mux2_1  _183_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform 1 0 1932 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _184_
timestamp 1665323087
transform 1 0 3496 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _185_
timestamp 1665323087
transform -1 0 5612 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _186_
timestamp 1665323087
transform 1 0 4692 0 1 1088
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _187_
timestamp 1665323087
transform 1 0 2852 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_2  _188_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform 1 0 4692 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__or2_2  _189_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform -1 0 3588 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__and2_2  _190_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform -1 0 1932 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_2  _191_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform -1 0 3496 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _192_
timestamp 1665323087
transform 1 0 3404 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__and2_2  _193_
timestamp 1665323087
transform -1 0 4968 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_2  _194_
timestamp 1665323087
transform -1 0 4784 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__or2_2  _195_
timestamp 1665323087
transform -1 0 5428 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__and2_2  _196_
timestamp 1665323087
transform 1 0 5152 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__and2_2  _197_
timestamp 1665323087
transform -1 0 5612 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__and2_2  _198_
timestamp 1665323087
transform 1 0 3772 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_2  _199_
timestamp 1665323087
transform -1 0 2852 0 1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_2  _200_
timestamp 1665323087
transform -1 0 5612 0 1 2176
box -38 -48 1234 592
use sky130_fd_sc_hd__a21o_2  _201_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform 1 0 3220 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_2  _202_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform 1 0 4048 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_2  _203_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform 1 0 3772 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_2  _204_
timestamp 1665323087
transform 1 0 1380 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__and2_2  _205_
timestamp 1665323087
transform 1 0 2484 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_2  _206_
timestamp 1665323087
transform -1 0 1840 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_2  _207_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform 1 0 1748 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_2  _208_
timestamp 1665323087
transform 1 0 5704 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_2  _209_
timestamp 1665323087
transform -1 0 3680 0 1 3264
box -38 -48 1234 592
use sky130_fd_sc_hd__or2_2  _210_
timestamp 1665323087
transform 1 0 4416 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__nand3_2  _211_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform 1 0 3680 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_2  _212_
timestamp 1665323087
transform 1 0 3036 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__a32o_2  _213_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform 1 0 2668 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__a21oi_2  _214_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform -1 0 3036 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_2  _215_
timestamp 1665323087
transform 1 0 2668 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_2  _216_
timestamp 1665323087
transform -1 0 3680 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__or3_2  _217_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform -1 0 2392 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_2  _218_
timestamp 1665323087
transform -1 0 5060 0 -1 3264
box -38 -48 1234 592
use sky130_fd_sc_hd__nand2_2  _219_
timestamp 1665323087
transform -1 0 2392 0 1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__or2_2  _220_
timestamp 1665323087
transform -1 0 3680 0 1 1088
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _221_
timestamp 1665323087
transform -1 0 3220 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__o22a_2  _222_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform 1 0 1472 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_2  _223_
timestamp 1665323087
transform 1 0 1380 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__a2111oi_2  _224_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform -1 0 2668 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__o21a_2  _225_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform 1 0 1840 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__and2_2  _226_
timestamp 1665323087
transform 1 0 2668 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__o31a_2  _227_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform -1 0 2668 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__or2_2  _228_
timestamp 1665323087
transform -1 0 10764 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__or2_2  _229_
timestamp 1665323087
transform 1 0 11500 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__or2_2  _230_
timestamp 1665323087
transform 1 0 7636 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _231_
timestamp 1665323087
transform -1 0 6348 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__or2_2  _232_
timestamp 1665323087
transform -1 0 8372 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__or4bb_2  _233_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform 1 0 8924 0 1 4352
box -38 -48 958 592
use sky130_fd_sc_hd__and3_2  _234_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform -1 0 10028 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__and2_2  _235_
timestamp 1665323087
transform -1 0 2760 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__or3b_2  _236_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform 1 0 1840 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__or3_2  _237_
timestamp 1665323087
transform -1 0 1932 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__and4_2  _238_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform -1 0 9936 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_2  _239_
timestamp 1665323087
transform -1 0 9108 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _240_
timestamp 1665323087
transform 1 0 9752 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _241_
timestamp 1665323087
transform -1 0 10304 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__or4_2  _242_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform 1 0 8924 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__o31a_2  _243_
timestamp 1665323087
transform -1 0 11316 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_2  _244_
timestamp 1665323087
transform -1 0 8280 0 -1 6528
box -38 -48 1234 592
use sky130_fd_sc_hd__nor2_2  _245_
timestamp 1665323087
transform -1 0 9384 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__and2_2  _246_
timestamp 1665323087
transform -1 0 8188 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_2  _247_
timestamp 1665323087
transform -1 0 8832 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _248_
timestamp 1665323087
transform -1 0 6808 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _249_
timestamp 1665323087
transform -1 0 10304 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_2  _250_
timestamp 1665323087
transform 1 0 7728 0 -1 8704
box -38 -48 1234 592
use sky130_fd_sc_hd__a21bo_2  _251_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform -1 0 8832 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__a32o_2  _252_
timestamp 1665323087
transform 1 0 8924 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__a32o_2  _253_
timestamp 1665323087
transform 1 0 6900 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__xnor2_2  _254_
timestamp 1665323087
transform -1 0 7268 0 1 7616
box -38 -48 1234 592
use sky130_fd_sc_hd__and2_2  _255_
timestamp 1665323087
transform -1 0 6900 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_2  _256_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform 1 0 6808 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_2  _257_
timestamp 1665323087
transform 1 0 7268 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_2  _258_
timestamp 1665323087
transform 1 0 8188 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_2  _259_
timestamp 1665323087
transform 1 0 8556 0 -1 6528
box -38 -48 1234 592
use sky130_fd_sc_hd__mux2_1  _260_
timestamp 1665323087
transform 1 0 9752 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__xor2_2  _261_
timestamp 1665323087
transform 1 0 7728 0 -1 7616
box -38 -48 1234 592
use sky130_fd_sc_hd__mux2_1  _262_
timestamp 1665323087
transform -1 0 10028 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__a21oi_2  _263_
timestamp 1665323087
transform 1 0 9200 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_2  _264_
timestamp 1665323087
transform -1 0 10948 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_2  _265_
timestamp 1665323087
transform 1 0 9844 0 -1 8704
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_2  _266_
timestamp 1665323087
transform 1 0 9016 0 1 7616
box -38 -48 1234 592
use sky130_fd_sc_hd__o2bb2a_2  _267_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform 1 0 9476 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_2  _268_
timestamp 1665323087
transform -1 0 9292 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_2  _269_
timestamp 1665323087
transform 1 0 6808 0 -1 5440
box -38 -48 1234 592
use sky130_fd_sc_hd__mux2_1  _270_
timestamp 1665323087
transform 1 0 8004 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_2  _271_
timestamp 1665323087
transform -1 0 11040 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_2  _272_
timestamp 1665323087
transform -1 0 10580 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__and3_2  _273_
timestamp 1665323087
transform 1 0 5704 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__and2_2  _274_
timestamp 1665323087
transform -1 0 6440 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_2  _275_
timestamp 1665323087
transform 1 0 5244 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__nand2b_2  _276_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform 1 0 5520 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_2  _277_
timestamp 1665323087
transform 1 0 5704 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_2  _278_
timestamp 1665323087
transform 1 0 6348 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_2  _279_
timestamp 1665323087
transform 1 0 6348 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__or2_2  _280_
timestamp 1665323087
transform 1 0 7636 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_2  _281_
timestamp 1665323087
transform 1 0 6992 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_2  _282_
timestamp 1665323087
transform 1 0 6716 0 1 1088
box -38 -48 1234 592
use sky130_fd_sc_hd__a21oi_2  _283_
timestamp 1665323087
transform 1 0 7544 0 1 2176
box -38 -48 682 592
use sky130_fd_sc_hd__nand3_2  _284_
timestamp 1665323087
transform 1 0 5520 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _285_
timestamp 1665323087
transform 1 0 10304 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _286_
timestamp 1665323087
transform 1 0 8924 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__or2_2  _287_
timestamp 1665323087
transform -1 0 9384 0 1 1088
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _288_
timestamp 1665323087
transform -1 0 7268 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_2  _289_
timestamp 1665323087
transform -1 0 4416 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__or3_2  _290_
timestamp 1665323087
transform -1 0 9476 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_2  _291_
timestamp 1665323087
transform -1 0 9384 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _292_
timestamp 1665323087
transform -1 0 8832 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__and2b_2  _293_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform -1 0 6992 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__and3_2  _294_
timestamp 1665323087
transform -1 0 6256 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_2  _295_
timestamp 1665323087
transform -1 0 3680 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_2  _296_
timestamp 1665323087
transform 1 0 10580 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__or2_2  _297_
timestamp 1665323087
transform 1 0 5336 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__or3_2  _298_
timestamp 1665323087
transform 1 0 8280 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_2  _299_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform -1 0 2116 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_2  _300_
timestamp 1665323087
transform -1 0 3128 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_2  _301_
timestamp 1665323087
transform -1 0 6256 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_2  _302_
timestamp 1665323087
transform -1 0 2208 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__or2_2  _303_
timestamp 1665323087
transform -1 0 7912 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_2  _304_
timestamp 1665323087
transform -1 0 6992 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_2  _305_
timestamp 1665323087
transform -1 0 3496 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_2  _306_
timestamp 1665323087
transform -1 0 4600 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__or3_2  _307_
timestamp 1665323087
transform -1 0 9568 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__or2_2  _308_
timestamp 1665323087
transform -1 0 7728 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_2  _309_
timestamp 1665323087
transform -1 0 7360 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _310_
timestamp 1665323087
transform 1 0 6532 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__o22a_2  _311_
timestamp 1665323087
transform 1 0 6716 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _312_
timestamp 1665323087
transform 1 0 6716 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__nand2b_2  _313_
timestamp 1665323087
transform 1 0 4232 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__o31a_2  _314_
timestamp 1665323087
transform -1 0 7268 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__or2_2  _315_
timestamp 1665323087
transform -1 0 7452 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_2  _316_
timestamp 1665323087
transform 1 0 5428 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_2  _317_
timestamp 1665323087
transform 1 0 5796 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__or2_2  _318_
timestamp 1665323087
transform -1 0 6808 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_2  _319_
timestamp 1665323087
transform -1 0 7084 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_2  _320_
timestamp 1665323087
transform 1 0 8096 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_2  _321_
timestamp 1665323087
transform 1 0 7360 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_2  _322_
timestamp 1665323087
transform 1 0 7544 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_2  _323_
timestamp 1665323087
transform 1 0 11040 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__or2_2  _324_
timestamp 1665323087
transform 1 0 9568 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__or2_2  _325_
timestamp 1665323087
transform -1 0 11316 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_2  _326_
timestamp 1665323087
transform -1 0 8280 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__or2_2  _327_
timestamp 1665323087
transform 1 0 10304 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__or2_2  _328_
timestamp 1665323087
transform -1 0 9384 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_2  _329_
timestamp 1665323087
transform 1 0 7912 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_2  _330_
timestamp 1665323087
transform 1 0 6992 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__o22a_2  _331_
timestamp 1665323087
transform -1 0 8832 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__and3_2  _332_
timestamp 1665323087
transform 1 0 7452 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__and3_2  _333_
timestamp 1665323087
transform 1 0 8556 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__a32o_2  _334_
timestamp 1665323087
transform 1 0 9752 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__o22a_2  _335_
timestamp 1665323087
transform -1 0 10028 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__and3_2  _336_
timestamp 1665323087
transform 1 0 9292 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_2  _337_
timestamp 1665323087
transform -1 0 11316 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_2  _338_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform 1 0 9476 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__or2_2  _339_
timestamp 1665323087
transform 1 0 10580 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__and3_2  _340_
timestamp 1665323087
transform 1 0 10304 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__a32o_2  _341_
timestamp 1665323087
transform 1 0 10120 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_2  _342_
timestamp 1665323087
transform -1 0 12236 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _343_
timestamp 1665323087
transform -1 0 8740 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_2  _344_
timestamp 1665323087
transform -1 0 12144 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_2  _345_
timestamp 1665323087
transform -1 0 11408 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_2  _346_
timestamp 1665323087
transform 1 0 8004 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__or3_2  _347_
timestamp 1665323087
transform 1 0 10028 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_2  _348_
timestamp 1665323087
transform 1 0 10304 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__or2_2  _349_
timestamp 1665323087
transform 1 0 11500 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_2  _350_
timestamp 1665323087
transform -1 0 11868 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_2  _351_
timestamp 1665323087
transform 1 0 11960 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_2  _352_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform 1 0 11776 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_2  _353_
timestamp 1665323087
transform 1 0 12420 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_2  _354_
timestamp 1665323087
transform 1 0 11224 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_2  _355_
timestamp 1665323087
transform -1 0 4232 0 1 1088
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _356_
timestamp 1665323087
transform -1 0 10948 0 -1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _357_
timestamp 1665323087
transform -1 0 10212 0 1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _358_
timestamp 1665323087
transform -1 0 12420 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _359_
timestamp 1665323087
transform 1 0 5796 0 -1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _360_
timestamp 1665323087
transform -1 0 8372 0 1 1088
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _361_
timestamp 1665323087
transform -1 0 9384 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _362_
timestamp 1665323087
transform 1 0 5796 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _363_
timestamp 1665323087
transform -1 0 5980 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _364_
timestamp 1665323087
transform -1 0 12420 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _365_
timestamp 1665323087
transform 1 0 6440 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _366_
timestamp 1665323087
transform -1 0 12696 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _367_
timestamp 1665323087
transform -1 0 11960 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _368_
timestamp 1665323087
transform -1 0 12420 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _369_
timestamp 1665323087
transform -1 0 11960 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _370_
timestamp 1665323087
transform 1 0 6440 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _371_
timestamp 1665323087
transform -1 0 11408 0 -1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _372_
timestamp 1665323087
transform 1 0 12420 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _373_
timestamp 1665323087
transform 1 0 11500 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _374_
timestamp 1665323087
transform 1 0 1472 0 1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _375_
timestamp 1665323087
transform 1 0 4232 0 1 1088
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _376_
timestamp 1665323087
transform 1 0 3864 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _377_
timestamp 1665323087
transform -1 0 4232 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _378_
timestamp 1665323087
transform -1 0 3128 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__dfrtp_2  _379_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform 1 0 8556 0 -1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _380_
timestamp 1665323087
transform 1 0 8280 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _381_
timestamp 1665323087
transform 1 0 10304 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _382_
timestamp 1665323087
transform 1 0 5612 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _383_
timestamp 1665323087
transform -1 0 8556 0 -1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _384_
timestamp 1665323087
transform -1 0 8832 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _385_
timestamp 1665323087
transform -1 0 8280 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _386_
timestamp 1665323087
transform 1 0 4324 0 -1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _387_
timestamp 1665323087
transform 1 0 10028 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _388_
timestamp 1665323087
transform 1 0 6900 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _389_
timestamp 1665323087
transform 1 0 10212 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _390_
timestamp 1665323087
transform 1 0 10304 0 1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _391_
timestamp 1665323087
transform 1 0 10028 0 1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _392_
timestamp 1665323087
transform 1 0 9476 0 -1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _393_
timestamp 1665323087
transform 1 0 5612 0 1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _394_
timestamp 1665323087
transform 1 0 9476 0 1 1088
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _395_
timestamp 1665323087
transform 1 0 11500 0 1 1088
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _396_
timestamp 1665323087
transform 1 0 11500 0 -1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _397_
timestamp 1665323087
transform -1 0 3588 0 -1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _398_
timestamp 1665323087
transform 1 0 3772 0 -1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _399_
timestamp 1665323087
transform -1 0 5704 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _400_
timestamp 1665323087
transform 1 0 2760 0 -1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _401_
timestamp 1665323087
transform 1 0 1472 0 1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__clkbuf_16  clockp_buffer_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform -1 0 3220 0 1 1088
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clockp_buffer_1
timestamp 1665323087
transform 1 0 1472 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[0\].id.delaybuf0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform 1 0 5704 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[0\].id.delaybuf1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform -1 0 5060 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[0\].id.delayen0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform 1 0 4140 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[0\].id.delayen1
timestamp 1665323087
transform -1 0 5704 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__einvn_8  ringosc.dstage\[0\].id.delayenb0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform 1 0 3588 0 -1 8704
box -38 -48 1694 592
use sky130_fd_sc_hd__einvn_4  ringosc.dstage\[0\].id.delayenb1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform -1 0 6256 0 -1 8704
box -38 -48 1050 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[0\].id.delayint0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform -1 0 4692 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[1\].id.delaybuf0
timestamp 1665323087
transform 1 0 4876 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[1\].id.delaybuf1
timestamp 1665323087
transform 1 0 5980 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[1\].id.delayen0
timestamp 1665323087
transform 1 0 4048 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[1\].id.delayen1
timestamp 1665323087
transform -1 0 5980 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__einvn_8  ringosc.dstage\[1\].id.delayenb0
timestamp 1665323087
transform 1 0 3680 0 -1 9792
box -38 -48 1694 592
use sky130_fd_sc_hd__einvn_4  ringosc.dstage\[1\].id.delayenb1
timestamp 1665323087
transform -1 0 5704 0 1 8704
box -38 -48 1050 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[1\].id.delayint0
timestamp 1665323087
transform -1 0 5336 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[2\].id.delaybuf0
timestamp 1665323087
transform -1 0 3680 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[2\].id.delaybuf1
timestamp 1665323087
transform 1 0 3312 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[2\].id.delayen0
timestamp 1665323087
transform 1 0 1748 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[2\].id.delayen1
timestamp 1665323087
transform 1 0 2392 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__einvn_8  ringosc.dstage\[2\].id.delayenb0
timestamp 1665323087
transform 1 0 1564 0 -1 9792
box -38 -48 1694 592
use sky130_fd_sc_hd__einvn_4  ringosc.dstage\[2\].id.delayenb1
timestamp 1665323087
transform 1 0 2300 0 1 8704
box -38 -48 1050 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[2\].id.delayint0
timestamp 1665323087
transform 1 0 3772 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[3\].id.delaybuf0
timestamp 1665323087
transform -1 0 2668 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[3\].id.delaybuf1
timestamp 1665323087
transform 1 0 2392 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[3\].id.delayen0
timestamp 1665323087
transform -1 0 2484 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[3\].id.delayen1
timestamp 1665323087
transform 1 0 1564 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__einvn_8  ringosc.dstage\[3\].id.delayenb0
timestamp 1665323087
transform 1 0 1380 0 1 10880
box -38 -48 1694 592
use sky130_fd_sc_hd__einvn_4  ringosc.dstage\[3\].id.delayenb1
timestamp 1665323087
transform 1 0 1380 0 1 11968
box -38 -48 1050 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[3\].id.delayint0
timestamp 1665323087
transform -1 0 1840 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[4\].id.delaybuf0
timestamp 1665323087
transform 1 0 3772 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[4\].id.delaybuf1
timestamp 1665323087
transform 1 0 3772 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[4\].id.delayen0
timestamp 1665323087
transform 1 0 2392 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[4\].id.delayen1
timestamp 1665323087
transform 1 0 3036 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__einvn_8  ringosc.dstage\[4\].id.delayenb0
timestamp 1665323087
transform 1 0 2208 0 -1 13056
box -38 -48 1694 592
use sky130_fd_sc_hd__einvn_4  ringosc.dstage\[4\].id.delayenb1
timestamp 1665323087
transform 1 0 2668 0 1 11968
box -38 -48 1050 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[4\].id.delayint0
timestamp 1665323087
transform 1 0 4048 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[5\].id.delaybuf0
timestamp 1665323087
transform 1 0 3680 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[5\].id.delaybuf1
timestamp 1665323087
transform 1 0 5336 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[5\].id.delayen0
timestamp 1665323087
transform 1 0 3036 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[5\].id.delayen1
timestamp 1665323087
transform -1 0 4876 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__einvn_8  ringosc.dstage\[5\].id.delayenb0
timestamp 1665323087
transform 1 0 3772 0 1 10880
box -38 -48 1694 592
use sky130_fd_sc_hd__einvn_4  ringosc.dstage\[5\].id.delayenb1
timestamp 1665323087
transform -1 0 5060 0 -1 10880
box -38 -48 1050 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[5\].id.delayint0
timestamp 1665323087
transform -1 0 4048 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[6\].id.delaybuf0
timestamp 1665323087
transform 1 0 5060 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[6\].id.delaybuf1
timestamp 1665323087
transform 1 0 6348 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[6\].id.delayen0
timestamp 1665323087
transform -1 0 6532 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[6\].id.delayen1
timestamp 1665323087
transform 1 0 5060 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__einvn_8  ringosc.dstage\[6\].id.delayenb0
timestamp 1665323087
transform 1 0 4600 0 -1 13056
box -38 -48 1694 592
use sky130_fd_sc_hd__einvn_4  ringosc.dstage\[6\].id.delayenb1
timestamp 1665323087
transform 1 0 4876 0 1 11968
box -38 -48 1050 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[6\].id.delayint0
timestamp 1665323087
transform -1 0 5060 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[7\].id.delaybuf0
timestamp 1665323087
transform 1 0 5888 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[7\].id.delaybuf1
timestamp 1665323087
transform 1 0 8924 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[7\].id.delayen0
timestamp 1665323087
transform 1 0 9384 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[7\].id.delayen1
timestamp 1665323087
transform 1 0 7360 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__einvn_8  ringosc.dstage\[7\].id.delayenb0
timestamp 1665323087
transform 1 0 9016 0 -1 13056
box -38 -48 1694 592
use sky130_fd_sc_hd__einvn_4  ringosc.dstage\[7\].id.delayenb1
timestamp 1665323087
transform 1 0 7820 0 -1 13056
box -38 -48 1050 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[7\].id.delayint0
timestamp 1665323087
transform 1 0 9844 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[8\].id.delaybuf0
timestamp 1665323087
transform 1 0 10764 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[8\].id.delaybuf1
timestamp 1665323087
transform -1 0 11408 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[8\].id.delayen0
timestamp 1665323087
transform 1 0 12144 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[8\].id.delayen1
timestamp 1665323087
transform -1 0 12144 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__einvn_8  ringosc.dstage\[8\].id.delayenb0
timestamp 1665323087
transform 1 0 11500 0 -1 13056
box -38 -48 1694 592
use sky130_fd_sc_hd__einvn_4  ringosc.dstage\[8\].id.delayenb1
timestamp 1665323087
transform 1 0 10948 0 1 11968
box -38 -48 1050 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[8\].id.delayint0
timestamp 1665323087
transform -1 0 10764 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[9\].id.delaybuf0
timestamp 1665323087
transform -1 0 13524 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[9\].id.delaybuf1
timestamp 1665323087
transform 1 0 12880 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[9\].id.delayen0
timestamp 1665323087
transform 1 0 12788 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[9\].id.delayen1
timestamp 1665323087
transform 1 0 12144 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__einvn_8  ringosc.dstage\[9\].id.delayenb0
timestamp 1665323087
transform 1 0 11960 0 1 11968
box -38 -48 1694 592
use sky130_fd_sc_hd__einvn_4  ringosc.dstage\[9\].id.delayenb1
timestamp 1665323087
transform 1 0 12052 0 1 10880
box -38 -48 1050 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[9\].id.delayint0
timestamp 1665323087
transform 1 0 13156 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[10\].id.delaybuf0
timestamp 1665323087
transform -1 0 13432 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[10\].id.delaybuf1
timestamp 1665323087
transform -1 0 12328 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[10\].id.delayen0
timestamp 1665323087
transform 1 0 12880 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[10\].id.delayen1
timestamp 1665323087
transform 1 0 12236 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__einvn_8  ringosc.dstage\[10\].id.delayenb0
timestamp 1665323087
transform 1 0 11868 0 1 9792
box -38 -48 1694 592
use sky130_fd_sc_hd__einvn_4  ringosc.dstage\[10\].id.delayenb1
timestamp 1665323087
transform 1 0 12144 0 -1 9792
box -38 -48 1050 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[10\].id.delayint0
timestamp 1665323087
transform -1 0 11408 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[11\].id.delaybuf0
timestamp 1665323087
transform 1 0 13156 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[11\].id.delaybuf1
timestamp 1665323087
transform 1 0 13340 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[11\].id.delayen0
timestamp 1665323087
transform 1 0 12696 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[11\].id.delayen1
timestamp 1665323087
transform 1 0 12696 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__einvn_8  ringosc.dstage\[11\].id.delayenb0
timestamp 1665323087
transform 1 0 11960 0 1 6528
box -38 -48 1694 592
use sky130_fd_sc_hd__einvn_4  ringosc.dstage\[11\].id.delayenb1
timestamp 1665323087
transform 1 0 12604 0 -1 5440
box -38 -48 1050 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[11\].id.delayint0
timestamp 1665323087
transform 1 0 13156 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  ringosc.ibufp00 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform -1 0 5520 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_8  ringosc.ibufp01 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform -1 0 5612 0 1 6528
box -38 -48 1234 592
use sky130_fd_sc_hd__clkinv_2  ringosc.ibufp10
timestamp 1665323087
transform -1 0 2024 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_8  ringosc.ibufp11
timestamp 1665323087
transform 1 0 1380 0 1 7616
box -38 -48 1234 592
use sky130_fd_sc_hd__conb_1  ringosc.iss.const1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform 1 0 12880 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__or2_2  ringosc.iss.ctrlen0
timestamp 1665323087
transform 1 0 11316 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.iss.delaybuf0
timestamp 1665323087
transform 1 0 13248 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_2  ringosc.iss.delayen0
timestamp 1665323087
transform 1 0 11776 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__einvp_2  ringosc.iss.delayen1
timestamp 1665323087
transform 1 0 12604 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__einvn_8  ringosc.iss.delayenb0
timestamp 1665323087
transform 1 0 11776 0 1 7616
box -38 -48 1694 592
use sky130_fd_sc_hd__einvn_4  ringosc.iss.delayenb1
timestamp 1665323087
transform 1 0 12328 0 -1 8704
box -38 -48 1050 592
use sky130_fd_sc_hd__clkinv_1  ringosc.iss.delayint0
timestamp 1665323087
transform 1 0 13340 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_1  ringosc.iss.reseten0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform 1 0 12420 0 -1 7616
box -38 -48 498 592
<< labels >>
flabel metal4 s 8208 1040 8528 13648 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal5 s 1056 8210 13940 8530 0 FreeSans 2560 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 4208 1040 4528 13648 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 12208 1040 12528 13648 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal5 s 1056 4210 13940 4530 0 FreeSans 2560 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal5 s 1056 12210 13940 12530 0 FreeSans 2560 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal3 s 0 416 800 536 0 FreeSans 480 0 0 0 clockp[0]
port 2 nsew signal tristate
flabel metal3 s 0 1232 800 1352 0 FreeSans 480 0 0 0 clockp[1]
port 3 nsew signal tristate
flabel metal3 s 0 7896 800 8016 0 FreeSans 480 0 0 0 dco
port 4 nsew signal input
flabel metal3 s 0 2184 800 2304 0 FreeSans 480 0 0 0 div[0]
port 5 nsew signal input
flabel metal3 s 0 3136 800 3256 0 FreeSans 480 0 0 0 div[1]
port 6 nsew signal input
flabel metal3 s 0 4088 800 4208 0 FreeSans 480 0 0 0 div[2]
port 7 nsew signal input
flabel metal3 s 0 5040 800 5160 0 FreeSans 480 0 0 0 div[3]
port 8 nsew signal input
flabel metal3 s 0 5992 800 6112 0 FreeSans 480 0 0 0 div[4]
port 9 nsew signal input
flabel metal3 s 0 6944 800 7064 0 FreeSans 480 0 0 0 enable
port 10 nsew signal input
flabel metal3 s 0 8712 800 8832 0 FreeSans 480 0 0 0 ext_trim[0]
port 11 nsew signal input
flabel metal2 s 3974 14200 4030 15000 0 FreeSans 224 90 0 0 ext_trim[10]
port 12 nsew signal input
flabel metal2 s 5170 14200 5226 15000 0 FreeSans 224 90 0 0 ext_trim[11]
port 13 nsew signal input
flabel metal2 s 6274 14200 6330 15000 0 FreeSans 224 90 0 0 ext_trim[12]
port 14 nsew signal input
flabel metal2 s 7470 14200 7526 15000 0 FreeSans 224 90 0 0 ext_trim[13]
port 15 nsew signal input
flabel metal2 s 8574 14200 8630 15000 0 FreeSans 224 90 0 0 ext_trim[14]
port 16 nsew signal input
flabel metal2 s 9770 14200 9826 15000 0 FreeSans 224 90 0 0 ext_trim[15]
port 17 nsew signal input
flabel metal2 s 10874 14200 10930 15000 0 FreeSans 224 90 0 0 ext_trim[16]
port 18 nsew signal input
flabel metal2 s 12070 14200 12126 15000 0 FreeSans 224 90 0 0 ext_trim[17]
port 19 nsew signal input
flabel metal2 s 13174 14200 13230 15000 0 FreeSans 224 90 0 0 ext_trim[18]
port 20 nsew signal input
flabel metal2 s 14370 14200 14426 15000 0 FreeSans 224 90 0 0 ext_trim[19]
port 21 nsew signal input
flabel metal3 s 0 9664 800 9784 0 FreeSans 480 0 0 0 ext_trim[1]
port 22 nsew signal input
flabel metal3 s 14200 13608 15000 13728 0 FreeSans 480 0 0 0 ext_trim[20]
port 23 nsew signal input
flabel metal3 s 14200 11160 15000 11280 0 FreeSans 480 0 0 0 ext_trim[21]
port 24 nsew signal input
flabel metal3 s 14200 8712 15000 8832 0 FreeSans 480 0 0 0 ext_trim[22]
port 25 nsew signal input
flabel metal3 s 14200 6128 15000 6248 0 FreeSans 480 0 0 0 ext_trim[23]
port 26 nsew signal input
flabel metal3 s 14200 3680 15000 3800 0 FreeSans 480 0 0 0 ext_trim[24]
port 27 nsew signal input
flabel metal3 s 14200 1232 15000 1352 0 FreeSans 480 0 0 0 ext_trim[25]
port 28 nsew signal input
flabel metal3 s 0 10616 800 10736 0 FreeSans 480 0 0 0 ext_trim[2]
port 29 nsew signal input
flabel metal3 s 0 11568 800 11688 0 FreeSans 480 0 0 0 ext_trim[3]
port 30 nsew signal input
flabel metal3 s 0 12520 800 12640 0 FreeSans 480 0 0 0 ext_trim[4]
port 31 nsew signal input
flabel metal3 s 0 13472 800 13592 0 FreeSans 480 0 0 0 ext_trim[5]
port 32 nsew signal input
flabel metal3 s 0 14424 800 14544 0 FreeSans 480 0 0 0 ext_trim[6]
port 33 nsew signal input
flabel metal2 s 570 14200 626 15000 0 FreeSans 224 90 0 0 ext_trim[7]
port 34 nsew signal input
flabel metal2 s 1674 14200 1730 15000 0 FreeSans 224 90 0 0 ext_trim[8]
port 35 nsew signal input
flabel metal2 s 2870 14200 2926 15000 0 FreeSans 224 90 0 0 ext_trim[9]
port 36 nsew signal input
flabel metal2 s 11150 0 11206 800 0 FreeSans 224 90 0 0 osc
port 37 nsew signal input
flabel metal2 s 3698 0 3754 800 0 FreeSans 224 90 0 0 resetb
port 38 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 15000 15000
<< end >>
