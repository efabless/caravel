magic
tech sky130A
magscale 1 2
timestamp 1651019111
<< metal1 >>
rect 195330 1007088 195336 1007140
rect 195388 1007128 195394 1007140
rect 203886 1007128 203892 1007140
rect 195388 1007100 203892 1007128
rect 195388 1007088 195394 1007100
rect 203886 1007088 203892 1007100
rect 203944 1007088 203950 1007140
rect 92606 1006544 92612 1006596
rect 92664 1006584 92670 1006596
rect 99926 1006584 99932 1006596
rect 92664 1006556 99932 1006584
rect 92664 1006544 92670 1006556
rect 99926 1006544 99932 1006556
rect 99984 1006544 99990 1006596
rect 95970 1006476 95976 1006528
rect 96028 1006516 96034 1006528
rect 104802 1006516 104808 1006528
rect 96028 1006488 104808 1006516
rect 96028 1006476 96034 1006488
rect 104802 1006476 104808 1006488
rect 104860 1006476 104866 1006528
rect 249058 1006476 249064 1006528
rect 249116 1006516 249122 1006528
rect 258166 1006516 258172 1006528
rect 249116 1006488 258172 1006516
rect 249116 1006476 249122 1006488
rect 258166 1006476 258172 1006488
rect 258224 1006476 258230 1006528
rect 302878 1006476 302884 1006528
rect 302936 1006516 302942 1006528
rect 308122 1006516 308128 1006528
rect 302936 1006488 308128 1006516
rect 302936 1006476 302942 1006488
rect 308122 1006476 308128 1006488
rect 308180 1006476 308186 1006528
rect 428366 1006476 428372 1006528
rect 428424 1006516 428430 1006528
rect 428424 1006488 437474 1006516
rect 428424 1006476 428430 1006488
rect 93210 1006408 93216 1006460
rect 93268 1006448 93274 1006460
rect 104342 1006448 104348 1006460
rect 93268 1006420 104348 1006448
rect 93268 1006408 93274 1006420
rect 104342 1006408 104348 1006420
rect 104400 1006408 104406 1006460
rect 253290 1006408 253296 1006460
rect 253348 1006448 253354 1006460
rect 253348 1006420 258074 1006448
rect 253348 1006408 253354 1006420
rect 99098 1006340 99104 1006392
rect 99156 1006380 99162 1006392
rect 126238 1006380 126244 1006392
rect 99156 1006352 126244 1006380
rect 99156 1006340 99162 1006352
rect 126238 1006340 126244 1006352
rect 126296 1006340 126302 1006392
rect 149698 1006340 149704 1006392
rect 149756 1006380 149762 1006392
rect 150894 1006380 150900 1006392
rect 149756 1006352 150900 1006380
rect 149756 1006340 149762 1006352
rect 150894 1006340 150900 1006352
rect 150952 1006380 150958 1006392
rect 150952 1006352 157334 1006380
rect 150952 1006340 150958 1006352
rect 93118 1006272 93124 1006324
rect 93176 1006312 93182 1006324
rect 100662 1006312 100668 1006324
rect 93176 1006284 100668 1006312
rect 93176 1006272 93182 1006284
rect 100662 1006272 100668 1006284
rect 100720 1006272 100726 1006324
rect 146938 1006272 146944 1006324
rect 146996 1006312 147002 1006324
rect 154114 1006312 154120 1006324
rect 146996 1006284 154120 1006312
rect 146996 1006272 147002 1006284
rect 154114 1006272 154120 1006284
rect 154172 1006272 154178 1006324
rect 145558 1006204 145564 1006256
rect 145616 1006244 145622 1006256
rect 151722 1006244 151728 1006256
rect 145616 1006216 151728 1006244
rect 145616 1006204 145622 1006216
rect 151722 1006204 151728 1006216
rect 151780 1006204 151786 1006256
rect 157306 1006244 157334 1006352
rect 201862 1006340 201868 1006392
rect 201920 1006380 201926 1006392
rect 228358 1006380 228364 1006392
rect 201920 1006352 228364 1006380
rect 201920 1006340 201926 1006352
rect 228358 1006340 228364 1006352
rect 228416 1006340 228422 1006392
rect 248322 1006340 248328 1006392
rect 248380 1006380 248386 1006392
rect 254854 1006380 254860 1006392
rect 248380 1006352 254860 1006380
rect 248380 1006340 248386 1006352
rect 254854 1006340 254860 1006352
rect 254912 1006340 254918 1006392
rect 177298 1006312 177304 1006324
rect 161446 1006284 177304 1006312
rect 161446 1006244 161474 1006284
rect 177298 1006272 177304 1006284
rect 177356 1006272 177362 1006324
rect 195146 1006272 195152 1006324
rect 195204 1006312 195210 1006324
rect 202690 1006312 202696 1006324
rect 195204 1006284 202696 1006312
rect 195204 1006272 195210 1006284
rect 202690 1006272 202696 1006284
rect 202748 1006272 202754 1006324
rect 207658 1006272 207664 1006324
rect 207716 1006312 207722 1006324
rect 210050 1006312 210056 1006324
rect 207716 1006284 210056 1006312
rect 207716 1006272 207722 1006284
rect 210050 1006272 210056 1006284
rect 210108 1006272 210114 1006324
rect 258046 1006312 258074 1006420
rect 301498 1006408 301504 1006460
rect 301556 1006448 301562 1006460
rect 307294 1006448 307300 1006460
rect 301556 1006420 307300 1006448
rect 301556 1006408 301562 1006420
rect 307294 1006408 307300 1006420
rect 307352 1006408 307358 1006460
rect 358170 1006408 358176 1006460
rect 358228 1006448 358234 1006460
rect 369118 1006448 369124 1006460
rect 358228 1006420 369124 1006448
rect 358228 1006408 358234 1006420
rect 369118 1006408 369124 1006420
rect 369176 1006408 369182 1006460
rect 427538 1006408 427544 1006460
rect 427596 1006448 427602 1006460
rect 427596 1006420 432644 1006448
rect 427596 1006408 427602 1006420
rect 356054 1006340 356060 1006392
rect 356112 1006380 356118 1006392
rect 380158 1006380 380164 1006392
rect 356112 1006352 380164 1006380
rect 356112 1006340 356118 1006352
rect 380158 1006340 380164 1006352
rect 380216 1006340 380222 1006392
rect 280798 1006312 280804 1006324
rect 258046 1006284 280804 1006312
rect 280798 1006272 280804 1006284
rect 280856 1006272 280862 1006324
rect 298738 1006272 298744 1006324
rect 298796 1006312 298802 1006324
rect 310606 1006312 310612 1006324
rect 298796 1006284 310612 1006312
rect 298796 1006272 298802 1006284
rect 310606 1006272 310612 1006284
rect 310664 1006272 310670 1006324
rect 357710 1006272 357716 1006324
rect 357768 1006312 357774 1006324
rect 374638 1006312 374644 1006324
rect 357768 1006284 374644 1006312
rect 357768 1006272 357774 1006284
rect 374638 1006272 374644 1006284
rect 374696 1006272 374702 1006324
rect 432616 1006312 432644 1006420
rect 437446 1006380 437474 1006488
rect 437446 1006352 441614 1006380
rect 441586 1006312 441614 1006352
rect 504542 1006340 504548 1006392
rect 504600 1006380 504606 1006392
rect 514202 1006380 514208 1006392
rect 504600 1006352 514208 1006380
rect 504600 1006340 504606 1006352
rect 514202 1006340 514208 1006352
rect 514260 1006340 514266 1006392
rect 445754 1006312 445760 1006324
rect 432616 1006284 437474 1006312
rect 441586 1006284 445760 1006312
rect 157306 1006216 161474 1006244
rect 196618 1006204 196624 1006256
rect 196676 1006244 196682 1006256
rect 204346 1006244 204352 1006256
rect 196676 1006216 204352 1006244
rect 196676 1006204 196682 1006216
rect 204346 1006204 204352 1006216
rect 204404 1006204 204410 1006256
rect 249150 1006204 249156 1006256
rect 249208 1006244 249214 1006256
rect 257338 1006244 257344 1006256
rect 249208 1006216 257344 1006244
rect 249208 1006204 249214 1006216
rect 257338 1006204 257344 1006216
rect 257396 1006204 257402 1006256
rect 300302 1006204 300308 1006256
rect 300360 1006244 300366 1006256
rect 306466 1006244 306472 1006256
rect 300360 1006216 306472 1006244
rect 300360 1006204 300366 1006216
rect 306466 1006204 306472 1006216
rect 306524 1006204 306530 1006256
rect 358906 1006204 358912 1006256
rect 358964 1006244 358970 1006256
rect 376018 1006244 376024 1006256
rect 358964 1006216 376024 1006244
rect 358964 1006204 358970 1006216
rect 376018 1006204 376024 1006216
rect 376076 1006204 376082 1006256
rect 437446 1006244 437474 1006284
rect 445754 1006272 445760 1006284
rect 445812 1006272 445818 1006324
rect 555970 1006272 555976 1006324
rect 556028 1006312 556034 1006324
rect 556028 1006284 572714 1006312
rect 556028 1006272 556034 1006284
rect 456058 1006244 456064 1006256
rect 437446 1006216 456064 1006244
rect 456058 1006204 456064 1006216
rect 456116 1006204 456122 1006256
rect 505370 1006204 505376 1006256
rect 505428 1006244 505434 1006256
rect 514110 1006244 514116 1006256
rect 505428 1006216 514116 1006244
rect 505428 1006204 505434 1006216
rect 514110 1006204 514116 1006216
rect 514168 1006204 514174 1006256
rect 94682 1006136 94688 1006188
rect 94740 1006176 94746 1006188
rect 103606 1006176 103612 1006188
rect 94740 1006148 103612 1006176
rect 94740 1006136 94746 1006148
rect 103606 1006136 103612 1006148
rect 103664 1006136 103670 1006188
rect 147030 1006136 147036 1006188
rect 147088 1006176 147094 1006188
rect 152090 1006176 152096 1006188
rect 147088 1006148 152096 1006176
rect 147088 1006136 147094 1006148
rect 152090 1006136 152096 1006148
rect 152148 1006136 152154 1006188
rect 197354 1006136 197360 1006188
rect 197412 1006176 197418 1006188
rect 197412 1006148 203748 1006176
rect 197412 1006136 197418 1006148
rect 98270 1006068 98276 1006120
rect 98328 1006108 98334 1006120
rect 99098 1006108 99104 1006120
rect 98328 1006080 99104 1006108
rect 98328 1006068 98334 1006080
rect 99098 1006068 99104 1006080
rect 99156 1006068 99162 1006120
rect 102778 1006068 102784 1006120
rect 102836 1006108 102842 1006120
rect 108850 1006108 108856 1006120
rect 102836 1006080 108856 1006108
rect 102836 1006068 102842 1006080
rect 108850 1006068 108856 1006080
rect 108908 1006068 108914 1006120
rect 154482 1006068 154488 1006120
rect 154540 1006108 154546 1006120
rect 160646 1006108 160652 1006120
rect 154540 1006080 160652 1006108
rect 154540 1006068 154546 1006080
rect 160646 1006068 160652 1006080
rect 160704 1006068 160710 1006120
rect 197998 1006068 198004 1006120
rect 198056 1006108 198062 1006120
rect 198056 1006080 200114 1006108
rect 198056 1006068 198062 1006080
rect 94498 1006000 94504 1006052
rect 94556 1006040 94562 1006052
rect 103146 1006040 103152 1006052
rect 94556 1006012 103152 1006040
rect 94556 1006000 94562 1006012
rect 103146 1006000 103152 1006012
rect 103204 1006000 103210 1006052
rect 144178 1006000 144184 1006052
rect 144236 1006040 144242 1006052
rect 150894 1006040 150900 1006052
rect 144236 1006012 150900 1006040
rect 144236 1006000 144242 1006012
rect 150894 1006000 150900 1006012
rect 150952 1006000 150958 1006052
rect 159082 1006000 159088 1006052
rect 159140 1006040 159146 1006052
rect 162118 1006040 162124 1006052
rect 159140 1006012 162124 1006040
rect 159140 1006000 159146 1006012
rect 162118 1006000 162124 1006012
rect 162176 1006000 162182 1006052
rect 200086 1006040 200114 1006080
rect 201034 1006068 201040 1006120
rect 201092 1006108 201098 1006120
rect 201862 1006108 201868 1006120
rect 201092 1006080 201868 1006108
rect 201092 1006068 201098 1006080
rect 201862 1006068 201868 1006080
rect 201920 1006068 201926 1006120
rect 203720 1006108 203748 1006148
rect 204990 1006136 204996 1006188
rect 205048 1006176 205054 1006188
rect 210418 1006176 210424 1006188
rect 205048 1006148 210424 1006176
rect 205048 1006136 205054 1006148
rect 210418 1006136 210424 1006148
rect 210476 1006136 210482 1006188
rect 247678 1006136 247684 1006188
rect 247736 1006176 247742 1006188
rect 255314 1006176 255320 1006188
rect 247736 1006148 255320 1006176
rect 247736 1006136 247742 1006148
rect 255314 1006136 255320 1006148
rect 255372 1006136 255378 1006188
rect 425146 1006136 425152 1006188
rect 425204 1006176 425210 1006188
rect 449250 1006176 449256 1006188
rect 425204 1006148 449256 1006176
rect 425204 1006136 425210 1006148
rect 449250 1006136 449256 1006148
rect 449308 1006136 449314 1006188
rect 505002 1006136 505008 1006188
rect 505060 1006176 505066 1006188
rect 516778 1006176 516784 1006188
rect 505060 1006148 516784 1006176
rect 505060 1006136 505066 1006148
rect 516778 1006136 516784 1006148
rect 516836 1006136 516842 1006188
rect 557166 1006136 557172 1006188
rect 557224 1006176 557230 1006188
rect 565170 1006176 565176 1006188
rect 557224 1006148 565176 1006176
rect 557224 1006136 557230 1006148
rect 565170 1006136 565176 1006148
rect 565228 1006136 565234 1006188
rect 207198 1006108 207204 1006120
rect 203720 1006080 207204 1006108
rect 207198 1006068 207204 1006080
rect 207256 1006068 207262 1006120
rect 209590 1006068 209596 1006120
rect 209648 1006108 209654 1006120
rect 228450 1006108 228456 1006120
rect 209648 1006080 228456 1006108
rect 209648 1006068 209654 1006080
rect 228450 1006068 228456 1006080
rect 228508 1006068 228514 1006120
rect 248414 1006068 248420 1006120
rect 248472 1006108 248478 1006120
rect 248472 1006080 253934 1006108
rect 248472 1006068 248478 1006080
rect 207566 1006040 207572 1006052
rect 200086 1006012 207572 1006040
rect 207566 1006000 207572 1006012
rect 207624 1006000 207630 1006052
rect 252462 1006000 252468 1006052
rect 252520 1006040 252526 1006052
rect 253290 1006040 253296 1006052
rect 252520 1006012 253296 1006040
rect 252520 1006000 252526 1006012
rect 253290 1006000 253296 1006012
rect 253348 1006000 253354 1006052
rect 253906 1006040 253934 1006080
rect 254670 1006068 254676 1006120
rect 254728 1006108 254734 1006120
rect 258534 1006108 258540 1006120
rect 254728 1006080 258540 1006108
rect 254728 1006068 254734 1006080
rect 258534 1006068 258540 1006080
rect 258592 1006068 258598 1006120
rect 303522 1006068 303528 1006120
rect 303580 1006108 303586 1006120
rect 304074 1006108 304080 1006120
rect 303580 1006080 304080 1006108
rect 303580 1006068 303586 1006080
rect 304074 1006068 304080 1006080
rect 304132 1006108 304138 1006120
rect 304902 1006108 304908 1006120
rect 304132 1006080 304908 1006108
rect 304132 1006068 304138 1006080
rect 304902 1006068 304908 1006080
rect 304960 1006068 304966 1006120
rect 356882 1006068 356888 1006120
rect 356940 1006108 356946 1006120
rect 360838 1006108 360844 1006120
rect 356940 1006080 360844 1006108
rect 356940 1006068 356946 1006080
rect 360838 1006068 360844 1006080
rect 360896 1006068 360902 1006120
rect 361390 1006068 361396 1006120
rect 361448 1006108 361454 1006120
rect 368474 1006108 368480 1006120
rect 361448 1006080 368480 1006108
rect 361448 1006068 361454 1006080
rect 368474 1006068 368480 1006080
rect 368532 1006068 368538 1006120
rect 369118 1006068 369124 1006120
rect 369176 1006108 369182 1006120
rect 380894 1006108 380900 1006120
rect 369176 1006080 380900 1006108
rect 369176 1006068 369182 1006080
rect 380894 1006068 380900 1006080
rect 380952 1006068 380958 1006120
rect 420822 1006068 420828 1006120
rect 420880 1006108 420886 1006120
rect 422662 1006108 422668 1006120
rect 420880 1006080 422668 1006108
rect 420880 1006068 420886 1006080
rect 422662 1006068 422668 1006080
rect 422720 1006068 422726 1006120
rect 427998 1006068 428004 1006120
rect 428056 1006108 428062 1006120
rect 465718 1006108 465724 1006120
rect 428056 1006080 465724 1006108
rect 428056 1006068 428062 1006080
rect 465718 1006068 465724 1006080
rect 465776 1006068 465782 1006120
rect 502518 1006068 502524 1006120
rect 502576 1006108 502582 1006120
rect 502576 1006080 509234 1006108
rect 502576 1006068 502582 1006080
rect 256970 1006040 256976 1006052
rect 253906 1006012 256976 1006040
rect 256970 1006000 256976 1006012
rect 257028 1006000 257034 1006052
rect 257338 1006000 257344 1006052
rect 257396 1006040 257402 1006052
rect 258994 1006040 259000 1006052
rect 257396 1006012 259000 1006040
rect 257396 1006000 257402 1006012
rect 258994 1006000 259000 1006012
rect 259052 1006000 259058 1006052
rect 261018 1006000 261024 1006052
rect 261076 1006040 261082 1006052
rect 269758 1006040 269764 1006052
rect 261076 1006012 269764 1006040
rect 261076 1006000 261082 1006012
rect 269758 1006000 269764 1006012
rect 269816 1006000 269822 1006052
rect 298830 1006000 298836 1006052
rect 298888 1006040 298894 1006052
rect 305270 1006040 305276 1006052
rect 298888 1006012 305276 1006040
rect 298888 1006000 298894 1006012
rect 305270 1006000 305276 1006012
rect 305328 1006000 305334 1006052
rect 315114 1006000 315120 1006052
rect 315172 1006040 315178 1006052
rect 319438 1006040 319444 1006052
rect 315172 1006012 319444 1006040
rect 315172 1006000 315178 1006012
rect 319438 1006000 319444 1006012
rect 319496 1006000 319502 1006052
rect 353110 1006000 353116 1006052
rect 353168 1006040 353174 1006052
rect 354490 1006040 354496 1006052
rect 353168 1006012 354496 1006040
rect 353168 1006000 353174 1006012
rect 354490 1006000 354496 1006012
rect 354548 1006000 354554 1006052
rect 358538 1006000 358544 1006052
rect 358596 1006040 358602 1006052
rect 362218 1006040 362224 1006052
rect 358596 1006012 362224 1006040
rect 358596 1006000 358602 1006012
rect 362218 1006000 362224 1006012
rect 362276 1006000 362282 1006052
rect 423490 1006000 423496 1006052
rect 423548 1006040 423554 1006052
rect 426342 1006040 426348 1006052
rect 423548 1006012 426348 1006040
rect 423548 1006000 423554 1006012
rect 426342 1006000 426348 1006012
rect 426400 1006000 426406 1006052
rect 430022 1006000 430028 1006052
rect 430080 1006040 430086 1006052
rect 468478 1006040 468484 1006052
rect 430080 1006012 468484 1006040
rect 430080 1006000 430086 1006012
rect 468478 1006000 468484 1006012
rect 468536 1006000 468542 1006052
rect 498102 1006000 498108 1006052
rect 498160 1006040 498166 1006052
rect 499666 1006040 499672 1006052
rect 498160 1006012 499672 1006040
rect 498160 1006000 498166 1006012
rect 499666 1006000 499672 1006012
rect 499724 1006000 499730 1006052
rect 500494 1006000 500500 1006052
rect 500552 1006040 500558 1006052
rect 504358 1006040 504364 1006052
rect 500552 1006012 504364 1006040
rect 500552 1006000 500558 1006012
rect 504358 1006000 504364 1006012
rect 504416 1006000 504422 1006052
rect 509206 1006040 509234 1006080
rect 518894 1006040 518900 1006052
rect 509206 1006012 518900 1006040
rect 518894 1006000 518900 1006012
rect 518952 1006000 518958 1006052
rect 549162 1006000 549168 1006052
rect 549220 1006040 549226 1006052
rect 550266 1006040 550272 1006052
rect 549220 1006012 550272 1006040
rect 549220 1006000 549226 1006012
rect 550266 1006000 550272 1006012
rect 550324 1006040 550330 1006052
rect 551094 1006040 551100 1006052
rect 550324 1006012 551100 1006040
rect 550324 1006000 550330 1006012
rect 551094 1006000 551100 1006012
rect 551152 1006000 551158 1006052
rect 552290 1006000 552296 1006052
rect 552348 1006040 552354 1006052
rect 556706 1006040 556712 1006052
rect 552348 1006012 556712 1006040
rect 552348 1006000 552354 1006012
rect 556706 1006000 556712 1006012
rect 556764 1006000 556770 1006052
rect 556798 1006000 556804 1006052
rect 556856 1006040 556862 1006052
rect 570598 1006040 570604 1006052
rect 556856 1006012 570604 1006040
rect 556856 1006000 556862 1006012
rect 570598 1006000 570604 1006012
rect 570656 1006000 570662 1006052
rect 572686 1006040 572714 1006284
rect 573358 1006040 573364 1006052
rect 572686 1006012 573364 1006040
rect 573358 1006000 573364 1006012
rect 573416 1006000 573422 1006052
rect 143718 1005388 143724 1005440
rect 143776 1005428 143782 1005440
rect 169018 1005428 169024 1005440
rect 143776 1005400 169024 1005428
rect 143776 1005388 143782 1005400
rect 169018 1005388 169024 1005400
rect 169076 1005388 169082 1005440
rect 361022 1005388 361028 1005440
rect 361080 1005428 361086 1005440
rect 371878 1005428 371884 1005440
rect 361080 1005400 371884 1005428
rect 361080 1005388 361086 1005400
rect 371878 1005388 371884 1005400
rect 371936 1005388 371942 1005440
rect 360562 1005320 360568 1005372
rect 360620 1005360 360626 1005372
rect 378778 1005360 378784 1005372
rect 360620 1005332 378784 1005360
rect 360620 1005320 360626 1005332
rect 378778 1005320 378784 1005332
rect 378836 1005320 378842 1005372
rect 360194 1005252 360200 1005304
rect 360252 1005292 360258 1005304
rect 381538 1005292 381544 1005304
rect 360252 1005264 381544 1005292
rect 360252 1005252 360258 1005264
rect 381538 1005252 381544 1005264
rect 381596 1005252 381602 1005304
rect 426342 1005252 426348 1005304
rect 426400 1005292 426406 1005304
rect 462958 1005292 462964 1005304
rect 426400 1005264 462964 1005292
rect 426400 1005252 426406 1005264
rect 462958 1005252 462964 1005264
rect 463016 1005252 463022 1005304
rect 503346 1005252 503352 1005304
rect 503404 1005292 503410 1005304
rect 518986 1005292 518992 1005304
rect 503404 1005264 518992 1005292
rect 503404 1005252 503410 1005264
rect 518986 1005252 518992 1005264
rect 519044 1005252 519050 1005304
rect 508682 1005048 508688 1005100
rect 508740 1005088 508746 1005100
rect 511258 1005088 511264 1005100
rect 508740 1005060 511264 1005088
rect 508740 1005048 508746 1005060
rect 511258 1005048 511264 1005060
rect 511316 1005048 511322 1005100
rect 507026 1004980 507032 1005032
rect 507084 1005020 507090 1005032
rect 509786 1005020 509792 1005032
rect 507084 1004992 509792 1005020
rect 507084 1004980 507090 1004992
rect 509786 1004980 509792 1004992
rect 509844 1004980 509850 1005032
rect 508222 1004912 508228 1004964
rect 508280 1004952 508286 1004964
rect 510614 1004952 510620 1004964
rect 508280 1004924 510620 1004952
rect 508280 1004912 508286 1004924
rect 510614 1004912 510620 1004924
rect 510672 1004912 510678 1004964
rect 159818 1004844 159824 1004896
rect 159876 1004884 159882 1004896
rect 162302 1004884 162308 1004896
rect 159876 1004856 162308 1004884
rect 159876 1004844 159882 1004856
rect 162302 1004844 162308 1004856
rect 162360 1004844 162366 1004896
rect 363414 1004844 363420 1004896
rect 363472 1004884 363478 1004896
rect 366358 1004884 366364 1004896
rect 363472 1004856 366364 1004884
rect 363472 1004844 363478 1004856
rect 366358 1004844 366364 1004856
rect 366416 1004844 366422 1004896
rect 159450 1004776 159456 1004828
rect 159508 1004816 159514 1004828
rect 161474 1004816 161480 1004828
rect 159508 1004788 161480 1004816
rect 159508 1004776 159514 1004788
rect 161474 1004776 161480 1004788
rect 161532 1004776 161538 1004828
rect 208762 1004776 208768 1004828
rect 208820 1004816 208826 1004828
rect 211798 1004816 211804 1004828
rect 208820 1004788 211804 1004816
rect 208820 1004776 208826 1004788
rect 211798 1004776 211804 1004788
rect 211856 1004776 211862 1004828
rect 304258 1004776 304264 1004828
rect 304316 1004816 304322 1004828
rect 306926 1004816 306932 1004828
rect 304316 1004788 306932 1004816
rect 304316 1004776 304322 1004788
rect 306926 1004776 306932 1004788
rect 306984 1004776 306990 1004828
rect 313826 1004776 313832 1004828
rect 313884 1004816 313890 1004828
rect 316034 1004816 316040 1004828
rect 313884 1004788 316040 1004816
rect 313884 1004776 313890 1004788
rect 316034 1004776 316040 1004788
rect 316092 1004776 316098 1004828
rect 364242 1004776 364248 1004828
rect 364300 1004816 364306 1004828
rect 366542 1004816 366548 1004828
rect 364300 1004788 366548 1004816
rect 364300 1004776 364306 1004788
rect 366542 1004776 366548 1004788
rect 366600 1004776 366606 1004828
rect 499482 1004776 499488 1004828
rect 499540 1004816 499546 1004828
rect 501322 1004816 501328 1004828
rect 499540 1004788 501328 1004816
rect 499540 1004776 499546 1004788
rect 501322 1004776 501328 1004788
rect 501380 1004776 501386 1004828
rect 507854 1004776 507860 1004828
rect 507912 1004816 507918 1004828
rect 510062 1004816 510068 1004828
rect 507912 1004788 510068 1004816
rect 507912 1004776 507918 1004788
rect 510062 1004776 510068 1004788
rect 510120 1004776 510126 1004828
rect 160278 1004708 160284 1004760
rect 160336 1004748 160342 1004760
rect 163498 1004748 163504 1004760
rect 160336 1004720 163504 1004748
rect 160336 1004708 160342 1004720
rect 163498 1004708 163504 1004720
rect 163556 1004708 163562 1004760
rect 209222 1004708 209228 1004760
rect 209280 1004748 209286 1004760
rect 211154 1004748 211160 1004760
rect 209280 1004720 211160 1004748
rect 209280 1004708 209286 1004720
rect 211154 1004708 211160 1004720
rect 211212 1004708 211218 1004760
rect 305822 1004708 305828 1004760
rect 305880 1004748 305886 1004760
rect 308582 1004748 308588 1004760
rect 305880 1004720 308588 1004748
rect 305880 1004708 305886 1004720
rect 308582 1004708 308588 1004720
rect 308640 1004708 308646 1004760
rect 314654 1004708 314660 1004760
rect 314712 1004748 314718 1004760
rect 316678 1004748 316684 1004760
rect 314712 1004720 316684 1004748
rect 314712 1004708 314718 1004720
rect 316678 1004708 316684 1004720
rect 316736 1004708 316742 1004760
rect 354306 1004708 354312 1004760
rect 354364 1004748 354370 1004760
rect 356882 1004748 356888 1004760
rect 354364 1004720 356888 1004748
rect 354364 1004708 354370 1004720
rect 356882 1004708 356888 1004720
rect 356940 1004708 356946 1004760
rect 361850 1004708 361856 1004760
rect 361908 1004748 361914 1004760
rect 364978 1004748 364984 1004760
rect 361908 1004720 364984 1004748
rect 361908 1004708 361914 1004720
rect 364978 1004708 364984 1004720
rect 365036 1004708 365042 1004760
rect 499022 1004708 499028 1004760
rect 499080 1004748 499086 1004760
rect 500862 1004748 500868 1004760
rect 499080 1004720 500868 1004748
rect 499080 1004708 499086 1004720
rect 500862 1004708 500868 1004720
rect 500920 1004708 500926 1004760
rect 509050 1004708 509056 1004760
rect 509108 1004748 509114 1004760
rect 510706 1004748 510712 1004760
rect 509108 1004720 510712 1004748
rect 509108 1004708 509114 1004720
rect 510706 1004708 510712 1004720
rect 510764 1004708 510770 1004760
rect 556338 1004708 556344 1004760
rect 556396 1004748 556402 1004760
rect 559742 1004748 559748 1004760
rect 556396 1004720 559748 1004748
rect 556396 1004708 556402 1004720
rect 559742 1004708 559748 1004720
rect 559800 1004708 559806 1004760
rect 94590 1004640 94596 1004692
rect 94648 1004680 94654 1004692
rect 103146 1004680 103152 1004692
rect 94648 1004652 103152 1004680
rect 94648 1004640 94654 1004652
rect 103146 1004640 103152 1004652
rect 103204 1004640 103210 1004692
rect 160646 1004640 160652 1004692
rect 160704 1004680 160710 1004692
rect 162946 1004680 162952 1004692
rect 160704 1004652 162952 1004680
rect 160704 1004640 160710 1004652
rect 162946 1004640 162952 1004652
rect 163004 1004640 163010 1004692
rect 199378 1004640 199384 1004692
rect 199436 1004680 199442 1004692
rect 202230 1004680 202236 1004692
rect 199436 1004652 202236 1004680
rect 199436 1004640 199442 1004652
rect 202230 1004640 202236 1004652
rect 202288 1004640 202294 1004692
rect 208394 1004640 208400 1004692
rect 208452 1004680 208458 1004692
rect 209774 1004680 209780 1004692
rect 208452 1004652 209780 1004680
rect 208452 1004640 208458 1004652
rect 209774 1004640 209780 1004652
rect 209832 1004640 209838 1004692
rect 305638 1004640 305644 1004692
rect 305696 1004680 305702 1004692
rect 307754 1004680 307760 1004692
rect 305696 1004652 307760 1004680
rect 305696 1004640 305702 1004652
rect 307754 1004640 307760 1004652
rect 307812 1004640 307818 1004692
rect 315482 1004640 315488 1004692
rect 315540 1004680 315546 1004692
rect 318058 1004680 318064 1004692
rect 315540 1004652 318064 1004680
rect 315540 1004640 315546 1004652
rect 318058 1004640 318064 1004652
rect 318116 1004640 318122 1004692
rect 354582 1004640 354588 1004692
rect 354640 1004680 354646 1004692
rect 356054 1004680 356060 1004692
rect 354640 1004652 356060 1004680
rect 354640 1004640 354646 1004652
rect 356054 1004640 356060 1004652
rect 356112 1004640 356118 1004692
rect 362586 1004640 362592 1004692
rect 362644 1004680 362650 1004692
rect 365162 1004680 365168 1004692
rect 362644 1004652 365168 1004680
rect 362644 1004640 362650 1004652
rect 365162 1004640 365168 1004652
rect 365220 1004640 365226 1004692
rect 499206 1004640 499212 1004692
rect 499264 1004680 499270 1004692
rect 500494 1004680 500500 1004692
rect 499264 1004652 500500 1004680
rect 499264 1004640 499270 1004652
rect 500494 1004640 500500 1004652
rect 500552 1004640 500558 1004692
rect 507394 1004640 507400 1004692
rect 507452 1004680 507458 1004692
rect 509234 1004680 509240 1004692
rect 507452 1004652 509240 1004680
rect 507452 1004640 507458 1004652
rect 509234 1004640 509240 1004652
rect 509292 1004640 509298 1004692
rect 557626 1004640 557632 1004692
rect 557684 1004680 557690 1004692
rect 559558 1004680 559564 1004692
rect 557684 1004652 559564 1004680
rect 557684 1004640 557690 1004652
rect 559558 1004640 559564 1004652
rect 559616 1004640 559622 1004692
rect 298922 1004572 298928 1004624
rect 298980 1004612 298986 1004624
rect 308950 1004612 308956 1004624
rect 298980 1004584 308956 1004612
rect 298980 1004572 298986 1004584
rect 308950 1004572 308956 1004584
rect 309008 1004572 309014 1004624
rect 422018 1004572 422024 1004624
rect 422076 1004612 422082 1004624
rect 423858 1004612 423864 1004624
rect 422076 1004584 423864 1004612
rect 422076 1004572 422082 1004584
rect 423858 1004572 423864 1004584
rect 423916 1004572 423922 1004624
rect 424686 1004028 424692 1004080
rect 424744 1004068 424750 1004080
rect 451274 1004068 451280 1004080
rect 424744 1004040 451280 1004068
rect 424744 1004028 424750 1004040
rect 451274 1004028 451280 1004040
rect 451332 1004028 451338 1004080
rect 423490 1003892 423496 1003944
rect 423548 1003932 423554 1003944
rect 454310 1003932 454316 1003944
rect 423548 1003904 454316 1003932
rect 423548 1003892 423554 1003904
rect 454310 1003892 454316 1003904
rect 454368 1003892 454374 1003944
rect 503714 1003892 503720 1003944
rect 503772 1003932 503778 1003944
rect 519262 1003932 519268 1003944
rect 503772 1003904 519268 1003932
rect 503772 1003892 503778 1003904
rect 519262 1003892 519268 1003904
rect 519320 1003892 519326 1003944
rect 92514 1003280 92520 1003332
rect 92572 1003320 92578 1003332
rect 99466 1003320 99472 1003332
rect 92572 1003292 99472 1003320
rect 92572 1003280 92578 1003292
rect 99466 1003280 99472 1003292
rect 99524 1003280 99530 1003332
rect 380894 1003280 380900 1003332
rect 380952 1003320 380958 1003332
rect 383562 1003320 383568 1003332
rect 380952 1003292 383568 1003320
rect 380952 1003280 380958 1003292
rect 383562 1003280 383568 1003292
rect 383620 1003280 383626 1003332
rect 553394 1003280 553400 1003332
rect 553452 1003320 553458 1003332
rect 554682 1003320 554688 1003332
rect 553452 1003292 554688 1003320
rect 553452 1003280 553458 1003292
rect 554682 1003280 554688 1003292
rect 554740 1003280 554746 1003332
rect 445754 1003212 445760 1003264
rect 445812 1003252 445818 1003264
rect 449802 1003252 449808 1003264
rect 445812 1003224 449808 1003252
rect 445812 1003212 445818 1003224
rect 449802 1003212 449808 1003224
rect 449860 1003212 449866 1003264
rect 553946 1002600 553952 1002652
rect 554004 1002640 554010 1002652
rect 564986 1002640 564992 1002652
rect 554004 1002612 564992 1002640
rect 554004 1002600 554010 1002612
rect 564986 1002600 564992 1002612
rect 565044 1002600 565050 1002652
rect 144086 1002532 144092 1002584
rect 144144 1002572 144150 1002584
rect 154574 1002572 154580 1002584
rect 144144 1002544 154580 1002572
rect 144144 1002532 144150 1002544
rect 154574 1002532 154580 1002544
rect 154632 1002532 154638 1002584
rect 354582 1002532 354588 1002584
rect 354640 1002572 354646 1002584
rect 359182 1002572 359188 1002584
rect 354640 1002544 359188 1002572
rect 354640 1002532 354646 1002544
rect 359182 1002532 359188 1002544
rect 359240 1002532 359246 1002584
rect 425974 1002532 425980 1002584
rect 426032 1002572 426038 1002584
rect 469306 1002572 469312 1002584
rect 426032 1002544 469312 1002572
rect 426032 1002532 426038 1002544
rect 469306 1002532 469312 1002544
rect 469364 1002532 469370 1002584
rect 554314 1002532 554320 1002584
rect 554372 1002572 554378 1002584
rect 567286 1002572 567292 1002584
rect 554372 1002544 567292 1002572
rect 554372 1002532 554378 1002544
rect 567286 1002532 567292 1002544
rect 567344 1002532 567350 1002584
rect 559190 1002396 559196 1002448
rect 559248 1002436 559254 1002448
rect 562502 1002436 562508 1002448
rect 559248 1002408 562508 1002436
rect 559248 1002396 559254 1002408
rect 562502 1002396 562508 1002408
rect 562560 1002396 562566 1002448
rect 106826 1002328 106832 1002380
rect 106884 1002368 106890 1002380
rect 109862 1002368 109868 1002380
rect 106884 1002340 109868 1002368
rect 106884 1002328 106890 1002340
rect 109862 1002328 109868 1002340
rect 109920 1002328 109926 1002380
rect 560846 1002328 560852 1002380
rect 560904 1002368 560910 1002380
rect 565078 1002368 565084 1002380
rect 560904 1002340 565084 1002368
rect 560904 1002328 560910 1002340
rect 565078 1002328 565084 1002340
rect 565136 1002328 565142 1002380
rect 106182 1002260 106188 1002312
rect 106240 1002300 106246 1002312
rect 108482 1002300 108488 1002312
rect 106240 1002272 108488 1002300
rect 106240 1002260 106246 1002272
rect 108482 1002260 108488 1002272
rect 108540 1002260 108546 1002312
rect 261846 1002260 261852 1002312
rect 261904 1002300 261910 1002312
rect 264238 1002300 264244 1002312
rect 261904 1002272 264244 1002300
rect 261904 1002260 261910 1002272
rect 264238 1002260 264244 1002272
rect 264296 1002260 264302 1002312
rect 558454 1002260 558460 1002312
rect 558512 1002300 558518 1002312
rect 560938 1002300 560944 1002312
rect 558512 1002272 560944 1002300
rect 558512 1002260 558518 1002272
rect 560938 1002260 560944 1002272
rect 560996 1002260 561002 1002312
rect 95878 1002192 95884 1002244
rect 95936 1002232 95942 1002244
rect 101490 1002232 101496 1002244
rect 95936 1002204 101496 1002232
rect 95936 1002192 95942 1002204
rect 101490 1002192 101496 1002204
rect 101548 1002192 101554 1002244
rect 105998 1002192 106004 1002244
rect 106056 1002232 106062 1002244
rect 108298 1002232 108304 1002244
rect 106056 1002204 108304 1002232
rect 106056 1002192 106062 1002204
rect 108298 1002192 108304 1002204
rect 108356 1002192 108362 1002244
rect 158254 1002192 158260 1002244
rect 158312 1002232 158318 1002244
rect 160738 1002232 160744 1002244
rect 158312 1002204 160744 1002232
rect 158312 1002192 158318 1002204
rect 160738 1002192 160744 1002204
rect 160796 1002192 160802 1002244
rect 202138 1002192 202144 1002244
rect 202196 1002232 202202 1002244
rect 205174 1002232 205180 1002244
rect 202196 1002204 205180 1002232
rect 202196 1002192 202202 1002204
rect 205174 1002192 205180 1002204
rect 205232 1002192 205238 1002244
rect 211614 1002192 211620 1002244
rect 211672 1002232 211678 1002244
rect 215938 1002232 215944 1002244
rect 211672 1002204 215944 1002232
rect 211672 1002192 211678 1002204
rect 215938 1002192 215944 1002204
rect 215996 1002192 216002 1002244
rect 252462 1002192 252468 1002244
rect 252520 1002232 252526 1002244
rect 254486 1002232 254492 1002244
rect 252520 1002204 254492 1002232
rect 252520 1002192 252526 1002204
rect 254486 1002192 254492 1002204
rect 254544 1002192 254550 1002244
rect 261478 1002192 261484 1002244
rect 261536 1002232 261542 1002244
rect 263594 1002232 263600 1002244
rect 261536 1002204 263600 1002232
rect 261536 1002192 261542 1002204
rect 263594 1002192 263600 1002204
rect 263652 1002192 263658 1002244
rect 559650 1002192 559656 1002244
rect 559708 1002232 559714 1002244
rect 561766 1002232 561772 1002244
rect 559708 1002204 561772 1002232
rect 559708 1002192 559714 1002204
rect 561766 1002192 561772 1002204
rect 561824 1002192 561830 1002244
rect 97350 1002124 97356 1002176
rect 97408 1002164 97414 1002176
rect 102318 1002164 102324 1002176
rect 97408 1002136 102324 1002164
rect 97408 1002124 97414 1002136
rect 102318 1002124 102324 1002136
rect 102376 1002124 102382 1002176
rect 105630 1002124 105636 1002176
rect 105688 1002164 105694 1002176
rect 107930 1002164 107936 1002176
rect 105688 1002136 107936 1002164
rect 105688 1002124 105694 1002136
rect 107930 1002124 107936 1002136
rect 107988 1002124 107994 1002176
rect 108022 1002124 108028 1002176
rect 108080 1002164 108086 1002176
rect 110506 1002164 110512 1002176
rect 108080 1002136 110512 1002164
rect 108080 1002124 108086 1002136
rect 110506 1002124 110512 1002136
rect 110564 1002124 110570 1002176
rect 157794 1002124 157800 1002176
rect 157852 1002164 157858 1002176
rect 160186 1002164 160192 1002176
rect 157852 1002136 160192 1002164
rect 157852 1002124 157858 1002136
rect 160186 1002124 160192 1002136
rect 160244 1002124 160250 1002176
rect 200942 1002124 200948 1002176
rect 201000 1002164 201006 1002176
rect 203518 1002164 203524 1002176
rect 201000 1002136 203524 1002164
rect 201000 1002124 201006 1002136
rect 203518 1002124 203524 1002136
rect 203576 1002124 203582 1002176
rect 210418 1002124 210424 1002176
rect 210476 1002164 210482 1002176
rect 213178 1002164 213184 1002176
rect 210476 1002136 213184 1002164
rect 210476 1002124 210482 1002136
rect 213178 1002124 213184 1002136
rect 213236 1002124 213242 1002176
rect 253750 1002124 253756 1002176
rect 253808 1002164 253814 1002176
rect 256142 1002164 256148 1002176
rect 253808 1002136 256148 1002164
rect 253808 1002124 253814 1002136
rect 256142 1002124 256148 1002136
rect 256200 1002124 256206 1002176
rect 260834 1002124 260840 1002176
rect 260892 1002164 260898 1002176
rect 261846 1002164 261852 1002176
rect 260892 1002136 261852 1002164
rect 260892 1002124 260898 1002136
rect 261846 1002124 261852 1002136
rect 261904 1002124 261910 1002176
rect 262674 1002124 262680 1002176
rect 262732 1002164 262738 1002176
rect 265802 1002164 265808 1002176
rect 262732 1002136 265808 1002164
rect 262732 1002124 262738 1002136
rect 265802 1002124 265808 1002136
rect 265860 1002124 265866 1002176
rect 550266 1002124 550272 1002176
rect 550324 1002164 550330 1002176
rect 553118 1002164 553124 1002176
rect 550324 1002136 553124 1002164
rect 550324 1002124 550330 1002136
rect 553118 1002124 553124 1002136
rect 553176 1002124 553182 1002176
rect 560478 1002124 560484 1002176
rect 560536 1002164 560542 1002176
rect 563054 1002164 563060 1002176
rect 560536 1002136 563060 1002164
rect 560536 1002124 560542 1002136
rect 563054 1002124 563060 1002136
rect 563112 1002124 563118 1002176
rect 97258 1002056 97264 1002108
rect 97316 1002096 97322 1002108
rect 100294 1002096 100300 1002108
rect 97316 1002068 100300 1002096
rect 97316 1002056 97322 1002068
rect 100294 1002056 100300 1002068
rect 100352 1002056 100358 1002108
rect 107654 1002056 107660 1002108
rect 107712 1002096 107718 1002108
rect 109586 1002096 109592 1002108
rect 107712 1002068 109592 1002096
rect 107712 1002056 107718 1002068
rect 109586 1002056 109592 1002068
rect 109644 1002056 109650 1002108
rect 157426 1002056 157432 1002108
rect 157484 1002096 157490 1002108
rect 159358 1002096 159364 1002108
rect 157484 1002068 159364 1002096
rect 157484 1002056 157490 1002068
rect 159358 1002056 159364 1002068
rect 159416 1002056 159422 1002108
rect 203702 1002056 203708 1002108
rect 203760 1002096 203766 1002108
rect 205910 1002096 205916 1002108
rect 203760 1002068 205916 1002096
rect 203760 1002056 203766 1002068
rect 205910 1002056 205916 1002068
rect 205968 1002056 205974 1002108
rect 211246 1002056 211252 1002108
rect 211304 1002096 211310 1002108
rect 213362 1002096 213368 1002108
rect 211304 1002068 213368 1002096
rect 211304 1002056 211310 1002068
rect 213362 1002056 213368 1002068
rect 213420 1002056 213426 1002108
rect 253842 1002056 253848 1002108
rect 253900 1002096 253906 1002108
rect 255682 1002096 255688 1002108
rect 253900 1002068 255688 1002096
rect 253900 1002056 253906 1002068
rect 255682 1002056 255688 1002068
rect 255740 1002056 255746 1002108
rect 259822 1002056 259828 1002108
rect 259880 1002096 259886 1002108
rect 261478 1002096 261484 1002108
rect 259880 1002068 261484 1002096
rect 259880 1002056 259886 1002068
rect 261478 1002056 261484 1002068
rect 261536 1002056 261542 1002108
rect 263502 1002056 263508 1002108
rect 263560 1002096 263566 1002108
rect 266998 1002096 267004 1002108
rect 263560 1002068 267004 1002096
rect 263560 1002056 263566 1002068
rect 266998 1002056 267004 1002068
rect 267056 1002056 267062 1002108
rect 310146 1002056 310152 1002108
rect 310204 1002096 310210 1002108
rect 311894 1002096 311900 1002108
rect 310204 1002068 311900 1002096
rect 310204 1002056 310210 1002068
rect 311894 1002056 311900 1002068
rect 311952 1002056 311958 1002108
rect 365070 1002056 365076 1002108
rect 365128 1002096 365134 1002108
rect 367922 1002096 367928 1002108
rect 365128 1002068 367928 1002096
rect 365128 1002056 365134 1002068
rect 367922 1002056 367928 1002068
rect 367980 1002056 367986 1002108
rect 423306 1002056 423312 1002108
rect 423364 1002096 423370 1002108
rect 425974 1002096 425980 1002108
rect 423364 1002068 425980 1002096
rect 423364 1002056 423370 1002068
rect 425974 1002056 425980 1002068
rect 426032 1002056 426038 1002108
rect 502150 1002056 502156 1002108
rect 502208 1002096 502214 1002108
rect 503714 1002096 503720 1002108
rect 502208 1002068 503720 1002096
rect 502208 1002056 502214 1002068
rect 503714 1002056 503720 1002068
rect 503772 1002056 503778 1002108
rect 509510 1002056 509516 1002108
rect 509568 1002096 509574 1002108
rect 514018 1002096 514024 1002108
rect 509568 1002068 514024 1002096
rect 509568 1002056 509574 1002068
rect 514018 1002056 514024 1002068
rect 514076 1002056 514082 1002108
rect 550358 1002056 550364 1002108
rect 550416 1002096 550422 1002108
rect 552290 1002096 552296 1002108
rect 550416 1002068 552296 1002096
rect 550416 1002056 550422 1002068
rect 552290 1002056 552296 1002068
rect 552348 1002056 552354 1002108
rect 560018 1002056 560024 1002108
rect 560076 1002096 560082 1002108
rect 562318 1002096 562324 1002108
rect 560076 1002068 562324 1002096
rect 560076 1002056 560082 1002068
rect 562318 1002056 562324 1002068
rect 562376 1002056 562382 1002108
rect 92330 1001988 92336 1002040
rect 92388 1002028 92394 1002040
rect 92606 1002028 92612 1002040
rect 92388 1002000 92612 1002028
rect 92388 1001988 92394 1002000
rect 92606 1001988 92612 1002000
rect 92664 1001988 92670 1002040
rect 98638 1001988 98644 1002040
rect 98696 1002028 98702 1002040
rect 101122 1002028 101128 1002040
rect 98696 1002000 101128 1002028
rect 98696 1001988 98702 1002000
rect 101122 1001988 101128 1002000
rect 101180 1001988 101186 1002040
rect 104342 1001988 104348 1002040
rect 104400 1002028 104406 1002040
rect 106642 1002028 106648 1002040
rect 104400 1002000 106648 1002028
rect 104400 1001988 104406 1002000
rect 106642 1001988 106648 1002000
rect 106700 1001988 106706 1002040
rect 107194 1001988 107200 1002040
rect 107252 1002028 107258 1002040
rect 109034 1002028 109040 1002040
rect 107252 1002000 109040 1002028
rect 107252 1001988 107258 1002000
rect 109034 1001988 109040 1002000
rect 109092 1001988 109098 1002040
rect 109678 1001988 109684 1002040
rect 109736 1002028 109742 1002040
rect 111794 1002028 111800 1002040
rect 109736 1002000 111800 1002028
rect 109736 1001988 109742 1002000
rect 111794 1001988 111800 1002000
rect 111852 1001988 111858 1002040
rect 158622 1001988 158628 1002040
rect 158680 1002028 158686 1002040
rect 160094 1002028 160100 1002040
rect 158680 1002000 160100 1002028
rect 158680 1001988 158686 1002000
rect 160094 1001988 160100 1002000
rect 160152 1001988 160158 1002040
rect 200298 1001988 200304 1002040
rect 200356 1002028 200362 1002040
rect 203058 1002028 203064 1002040
rect 200356 1002000 203064 1002028
rect 200356 1001988 200362 1002000
rect 203058 1001988 203064 1002000
rect 203116 1001988 203122 1002040
rect 203518 1001988 203524 1002040
rect 203576 1002028 203582 1002040
rect 205542 1002028 205548 1002040
rect 203576 1002000 205548 1002028
rect 203576 1001988 203582 1002000
rect 205542 1001988 205548 1002000
rect 205600 1001988 205606 1002040
rect 212534 1001988 212540 1002040
rect 212592 1002028 212598 1002040
rect 214558 1002028 214564 1002040
rect 212592 1002000 214564 1002028
rect 212592 1001988 212598 1002000
rect 214558 1001988 214564 1002000
rect 214616 1001988 214622 1002040
rect 260190 1001988 260196 1002040
rect 260248 1002028 260254 1002040
rect 262858 1002028 262864 1002040
rect 260248 1002000 262864 1002028
rect 260248 1001988 260254 1002000
rect 262858 1001988 262864 1002000
rect 262916 1001988 262922 1002040
rect 263042 1001988 263048 1002040
rect 263100 1002028 263106 1002040
rect 265618 1002028 265624 1002040
rect 263100 1002000 265624 1002028
rect 263100 1001988 263106 1002000
rect 265618 1001988 265624 1002000
rect 265676 1001988 265682 1002040
rect 300118 1001988 300124 1002040
rect 300176 1002028 300182 1002040
rect 306098 1002028 306104 1002040
rect 300176 1002000 306104 1002028
rect 300176 1001988 300182 1002000
rect 306098 1001988 306104 1002000
rect 306156 1001988 306162 1002040
rect 307018 1001988 307024 1002040
rect 307076 1002028 307082 1002040
rect 309318 1002028 309324 1002040
rect 307076 1002000 309324 1002028
rect 307076 1001988 307082 1002000
rect 309318 1001988 309324 1002000
rect 309376 1001988 309382 1002040
rect 312262 1001988 312268 1002040
rect 312320 1002028 312326 1002040
rect 314654 1002028 314660 1002040
rect 312320 1002000 314660 1002028
rect 312320 1001988 312326 1002000
rect 314654 1001988 314660 1002000
rect 314712 1001988 314718 1002040
rect 357158 1001988 357164 1002040
rect 357216 1002028 357222 1002040
rect 359366 1002028 359372 1002040
rect 357216 1002000 359372 1002028
rect 357216 1001988 357222 1002000
rect 359366 1001988 359372 1002000
rect 359424 1001988 359430 1002040
rect 365898 1001988 365904 1002040
rect 365956 1002028 365962 1002040
rect 369118 1002028 369124 1002040
rect 365956 1002000 369124 1002028
rect 365956 1001988 365962 1002000
rect 369118 1001988 369124 1002000
rect 369176 1001988 369182 1002040
rect 424962 1001988 424968 1002040
rect 425020 1002028 425026 1002040
rect 426342 1002028 426348 1002040
rect 425020 1002000 426348 1002028
rect 425020 1001988 425026 1002000
rect 426342 1001988 426348 1002000
rect 426400 1001988 426406 1002040
rect 505830 1001988 505836 1002040
rect 505888 1002028 505894 1002040
rect 508682 1002028 508688 1002040
rect 505888 1002000 508688 1002028
rect 505888 1001988 505894 1002000
rect 508682 1001988 508688 1002000
rect 508740 1001988 508746 1002040
rect 509878 1001988 509884 1002040
rect 509936 1002028 509942 1002040
rect 512822 1002028 512828 1002040
rect 509936 1002000 512828 1002028
rect 509936 1001988 509942 1002000
rect 512822 1001988 512828 1002000
rect 512880 1001988 512886 1002040
rect 550450 1001988 550456 1002040
rect 550508 1002028 550514 1002040
rect 552658 1002028 552664 1002040
rect 550508 1002000 552664 1002028
rect 550508 1001988 550514 1002000
rect 552658 1001988 552664 1002000
rect 552716 1001988 552722 1002040
rect 553118 1001988 553124 1002040
rect 553176 1002028 553182 1002040
rect 555142 1002028 555148 1002040
rect 553176 1002000 555148 1002028
rect 553176 1001988 553182 1002000
rect 555142 1001988 555148 1002000
rect 555200 1001988 555206 1002040
rect 557994 1001988 558000 1002040
rect 558052 1002028 558058 1002040
rect 560570 1002028 560576 1002040
rect 558052 1002000 560576 1002028
rect 558052 1001988 558058 1002000
rect 560570 1001988 560576 1002000
rect 560628 1001988 560634 1002040
rect 561674 1001988 561680 1002040
rect 561732 1002028 561738 1002040
rect 563698 1002028 563704 1002040
rect 561732 1002000 563704 1002028
rect 561732 1001988 561738 1002000
rect 563698 1001988 563704 1002000
rect 563756 1001988 563762 1002040
rect 100018 1001920 100024 1001972
rect 100076 1001960 100082 1001972
rect 101950 1001960 101956 1001972
rect 100076 1001932 101956 1001960
rect 100076 1001920 100082 1001932
rect 101950 1001920 101956 1001932
rect 102008 1001920 102014 1001972
rect 106458 1001920 106464 1001972
rect 106516 1001960 106522 1001972
rect 107746 1001960 107752 1001972
rect 106516 1001932 107752 1001960
rect 106516 1001920 106522 1001932
rect 107746 1001920 107752 1001932
rect 107804 1001920 107810 1001972
rect 108482 1001920 108488 1001972
rect 108540 1001960 108546 1001972
rect 111058 1001960 111064 1001972
rect 108540 1001932 111064 1001960
rect 108540 1001920 108546 1001932
rect 111058 1001920 111064 1001932
rect 111116 1001920 111122 1001972
rect 156966 1001920 156972 1001972
rect 157024 1001960 157030 1001972
rect 158714 1001960 158720 1001972
rect 157024 1001932 158720 1001960
rect 157024 1001920 157030 1001932
rect 158714 1001920 158720 1001932
rect 158772 1001920 158778 1001972
rect 195146 1001920 195152 1001972
rect 195204 1001960 195210 1001972
rect 197354 1001960 197360 1001972
rect 195204 1001932 197360 1001960
rect 195204 1001920 195210 1001932
rect 197354 1001920 197360 1001932
rect 197412 1001920 197418 1001972
rect 202322 1001920 202328 1001972
rect 202380 1001960 202386 1001972
rect 204714 1001960 204720 1001972
rect 202380 1001932 204720 1001960
rect 202380 1001920 202386 1001932
rect 204714 1001920 204720 1001932
rect 204772 1001920 204778 1001972
rect 204898 1001920 204904 1001972
rect 204956 1001960 204962 1001972
rect 206738 1001960 206744 1001972
rect 204956 1001932 206744 1001960
rect 204956 1001920 204962 1001932
rect 206738 1001920 206744 1001932
rect 206796 1001920 206802 1001972
rect 212074 1001920 212080 1001972
rect 212132 1001960 212138 1001972
rect 213914 1001960 213920 1001972
rect 212132 1001932 213920 1001960
rect 212132 1001920 212138 1001932
rect 213914 1001920 213920 1001932
rect 213972 1001920 213978 1001972
rect 251818 1001920 251824 1001972
rect 251876 1001960 251882 1001972
rect 254118 1001960 254124 1001972
rect 251876 1001932 254124 1001960
rect 251876 1001920 251882 1001932
rect 254118 1001920 254124 1001932
rect 254176 1001920 254182 1001972
rect 254578 1001920 254584 1001972
rect 254636 1001960 254642 1001972
rect 256510 1001960 256516 1001972
rect 254636 1001932 256516 1001960
rect 254636 1001920 254642 1001932
rect 256510 1001920 256516 1001932
rect 256568 1001920 256574 1001972
rect 260650 1001920 260656 1001972
rect 260708 1001960 260714 1001972
rect 262214 1001960 262220 1001972
rect 260708 1001932 262220 1001960
rect 260708 1001920 260714 1001932
rect 262214 1001920 262220 1001932
rect 262272 1001920 262278 1001972
rect 263870 1001920 263876 1001972
rect 263928 1001960 263934 1001972
rect 267090 1001960 267096 1001972
rect 263928 1001932 267096 1001960
rect 263928 1001920 263934 1001932
rect 267090 1001920 267096 1001932
rect 267148 1001920 267154 1001972
rect 300210 1001920 300216 1001972
rect 300268 1001960 300274 1001972
rect 305730 1001960 305736 1001972
rect 300268 1001932 305736 1001960
rect 300268 1001920 300274 1001932
rect 305730 1001920 305736 1001932
rect 305788 1001920 305794 1001972
rect 311434 1001920 311440 1001972
rect 311492 1001960 311498 1001972
rect 313550 1001960 313556 1001972
rect 311492 1001932 313556 1001960
rect 311492 1001920 311498 1001932
rect 313550 1001920 313556 1001932
rect 313608 1001920 313614 1001972
rect 357342 1001920 357348 1001972
rect 357400 1001960 357406 1001972
rect 358906 1001960 358912 1001972
rect 357400 1001932 358912 1001960
rect 357400 1001920 357406 1001932
rect 358906 1001920 358912 1001932
rect 358964 1001920 358970 1001972
rect 365438 1001920 365444 1001972
rect 365496 1001960 365502 1001972
rect 367738 1001960 367744 1001972
rect 365496 1001932 367744 1001960
rect 365496 1001920 365502 1001932
rect 367738 1001920 367744 1001932
rect 367796 1001920 367802 1001972
rect 420822 1001920 420828 1001972
rect 420880 1001960 420886 1001972
rect 421466 1001960 421472 1001972
rect 420880 1001932 421472 1001960
rect 420880 1001920 420886 1001932
rect 421466 1001920 421472 1001932
rect 421524 1001920 421530 1001972
rect 423398 1001920 423404 1001972
rect 423456 1001960 423462 1001972
rect 425146 1001960 425152 1001972
rect 423456 1001932 425152 1001960
rect 423456 1001920 423462 1001932
rect 425146 1001920 425152 1001932
rect 425204 1001920 425210 1001972
rect 425698 1001920 425704 1001972
rect 425756 1001960 425762 1001972
rect 426802 1001960 426808 1001972
rect 425756 1001932 426808 1001960
rect 425756 1001920 425762 1001932
rect 426802 1001920 426808 1001932
rect 426860 1001920 426866 1001972
rect 506198 1001920 506204 1001972
rect 506256 1001960 506262 1001972
rect 508498 1001960 508504 1001972
rect 506256 1001932 508504 1001960
rect 506256 1001920 506262 1001932
rect 508498 1001920 508504 1001932
rect 508556 1001920 508562 1001972
rect 510338 1001920 510344 1001972
rect 510396 1001960 510402 1001972
rect 512638 1001960 512644 1001972
rect 510396 1001932 512644 1001960
rect 510396 1001920 510402 1001932
rect 512638 1001920 512644 1001932
rect 512696 1001920 512702 1001972
rect 549070 1001920 549076 1001972
rect 549128 1001960 549134 1001972
rect 551462 1001960 551468 1001972
rect 549128 1001932 551468 1001960
rect 549128 1001920 549134 1001932
rect 551462 1001920 551468 1001932
rect 551520 1001920 551526 1001972
rect 551922 1001920 551928 1001972
rect 551980 1001960 551986 1001972
rect 553486 1001960 553492 1001972
rect 551980 1001932 553492 1001960
rect 551980 1001920 551986 1001932
rect 553486 1001920 553492 1001932
rect 553544 1001920 553550 1001972
rect 558822 1001920 558828 1001972
rect 558880 1001960 558886 1001972
rect 560294 1001960 560300 1001972
rect 558880 1001932 560300 1001960
rect 558880 1001920 558886 1001932
rect 560294 1001920 560300 1001932
rect 560352 1001920 560358 1001972
rect 561306 1001920 561312 1001972
rect 561364 1001960 561370 1001972
rect 563882 1001960 563888 1001972
rect 561364 1001932 563888 1001960
rect 561364 1001920 561370 1001932
rect 563882 1001920 563888 1001932
rect 563940 1001920 563946 1001972
rect 298370 1001852 298376 1001904
rect 298428 1001892 298434 1001904
rect 310146 1001892 310152 1001904
rect 298428 1001864 310152 1001892
rect 298428 1001852 298434 1001864
rect 310146 1001852 310152 1001864
rect 310204 1001852 310210 1001904
rect 518894 1001852 518900 1001904
rect 518952 1001892 518958 1001904
rect 523862 1001892 523868 1001904
rect 518952 1001864 523868 1001892
rect 518952 1001852 518958 1001864
rect 523862 1001852 523868 1001864
rect 523920 1001852 523926 1001904
rect 449250 1001784 449256 1001836
rect 449308 1001824 449314 1001836
rect 452562 1001824 452568 1001836
rect 449308 1001796 452568 1001824
rect 449308 1001784 449314 1001796
rect 452562 1001784 452568 1001796
rect 452620 1001784 452626 1001836
rect 424962 1001240 424968 1001292
rect 425020 1001280 425026 1001292
rect 447134 1001280 447140 1001292
rect 425020 1001252 447140 1001280
rect 425020 1001240 425026 1001252
rect 447134 1001240 447140 1001252
rect 447192 1001240 447198 1001292
rect 92422 1001172 92428 1001224
rect 92480 1001212 92486 1001224
rect 98638 1001212 98644 1001224
rect 92480 1001184 98644 1001212
rect 92480 1001172 92486 1001184
rect 98638 1001172 98644 1001184
rect 98696 1001172 98702 1001224
rect 195422 1001172 195428 1001224
rect 195480 1001212 195486 1001224
rect 200942 1001212 200948 1001224
rect 195480 1001184 200948 1001212
rect 195480 1001172 195486 1001184
rect 200942 1001172 200948 1001184
rect 201000 1001172 201006 1001224
rect 423306 1001172 423312 1001224
rect 423364 1001212 423370 1001224
rect 469214 1001212 469220 1001224
rect 423364 1001184 469220 1001212
rect 423364 1001172 423370 1001184
rect 469214 1001172 469220 1001184
rect 469272 1001172 469278 1001224
rect 299382 1000560 299388 1000612
rect 299440 1000600 299446 1000612
rect 302878 1000600 302884 1000612
rect 299440 1000572 302884 1000600
rect 299440 1000560 299446 1000572
rect 302878 1000560 302884 1000572
rect 302936 1000560 302942 1000612
rect 92698 1000492 92704 1000544
rect 92756 1000532 92762 1000544
rect 94682 1000532 94688 1000544
rect 92756 1000504 94688 1000532
rect 92756 1000492 92762 1000504
rect 94682 1000492 94688 1000504
rect 94740 1000492 94746 1000544
rect 152734 1000492 152740 1000544
rect 152792 1000532 152798 1000544
rect 154942 1000532 154948 1000544
rect 152792 1000504 154948 1000532
rect 152792 1000492 152798 1000504
rect 154942 1000492 154948 1000504
rect 155000 1000492 155006 1000544
rect 298554 1000492 298560 1000544
rect 298612 1000532 298618 1000544
rect 300302 1000532 300308 1000544
rect 298612 1000504 300308 1000532
rect 298612 1000492 298618 1000504
rect 300302 1000492 300308 1000504
rect 300360 1000492 300366 1000544
rect 611354 1000492 611360 1000544
rect 611412 1000532 611418 1000544
rect 625706 1000532 625712 1000544
rect 611412 1000504 625712 1000532
rect 611412 1000492 611418 1000504
rect 625706 1000492 625712 1000504
rect 625764 1000492 625770 1000544
rect 514202 1000424 514208 1000476
rect 514260 1000464 514266 1000476
rect 520182 1000464 520188 1000476
rect 514260 1000436 520188 1000464
rect 514260 1000424 514266 1000436
rect 520182 1000424 520188 1000436
rect 520240 1000424 520246 1000476
rect 451274 1000220 451280 1000272
rect 451332 1000260 451338 1000272
rect 459554 1000260 459560 1000272
rect 451332 1000232 459560 1000260
rect 451332 1000220 451338 1000232
rect 459554 1000220 459560 1000232
rect 459612 1000220 459618 1000272
rect 247034 999948 247040 1000000
rect 247092 999988 247098 1000000
rect 252462 999988 252468 1000000
rect 247092 999960 252468 999988
rect 247092 999948 247098 999960
rect 252462 999948 252468 999960
rect 252520 999948 252526 1000000
rect 551922 999812 551928 999864
rect 551980 999852 551986 999864
rect 568206 999852 568212 999864
rect 551980 999824 568212 999852
rect 551980 999812 551986 999824
rect 568206 999812 568212 999824
rect 568264 999812 568270 999864
rect 143810 999744 143816 999796
rect 143868 999784 143874 999796
rect 155770 999784 155776 999796
rect 143868 999756 155776 999784
rect 143868 999744 143874 999756
rect 155770 999744 155776 999756
rect 155828 999744 155834 999796
rect 428826 999744 428832 999796
rect 428884 999784 428890 999796
rect 469398 999784 469404 999796
rect 428884 999756 469404 999784
rect 428884 999744 428890 999756
rect 469398 999744 469404 999756
rect 469456 999744 469462 999796
rect 499482 999744 499488 999796
rect 499540 999784 499546 999796
rect 504266 999784 504272 999796
rect 499540 999756 504272 999784
rect 499540 999744 499546 999756
rect 504266 999744 504272 999756
rect 504324 999744 504330 999796
rect 508682 999744 508688 999796
rect 508740 999784 508746 999796
rect 513926 999784 513932 999796
rect 508740 999756 513932 999784
rect 508740 999744 508746 999756
rect 513926 999744 513932 999756
rect 513984 999744 513990 999796
rect 550266 999744 550272 999796
rect 550324 999784 550330 999796
rect 567930 999784 567936 999796
rect 550324 999756 567936 999784
rect 550324 999744 550330 999756
rect 567930 999744 567936 999756
rect 567988 999744 567994 999796
rect 247126 999472 247132 999524
rect 247184 999512 247190 999524
rect 253750 999512 253756 999524
rect 247184 999484 253756 999512
rect 247184 999472 247190 999484
rect 253750 999472 253756 999484
rect 253808 999472 253814 999524
rect 249702 999132 249708 999184
rect 249760 999172 249766 999184
rect 254670 999172 254676 999184
rect 249760 999144 254676 999172
rect 249760 999132 249766 999144
rect 254670 999132 254676 999144
rect 254728 999132 254734 999184
rect 469306 999132 469312 999184
rect 469364 999172 469370 999184
rect 472066 999172 472072 999184
rect 469364 999144 472072 999172
rect 469364 999132 469370 999144
rect 472066 999132 472072 999144
rect 472124 999132 472130 999184
rect 92330 999064 92336 999116
rect 92388 999104 92394 999116
rect 94590 999104 94596 999116
rect 92388 999076 94596 999104
rect 92388 999064 92394 999076
rect 94590 999064 94596 999076
rect 94648 999064 94654 999116
rect 250714 999064 250720 999116
rect 250772 999104 250778 999116
rect 253842 999104 253848 999116
rect 250772 999076 253848 999104
rect 250772 999064 250778 999076
rect 253842 999064 253848 999076
rect 253900 999064 253906 999116
rect 514110 999064 514116 999116
rect 514168 999104 514174 999116
rect 520090 999104 520096 999116
rect 514168 999076 520096 999104
rect 514168 999064 514174 999076
rect 520090 999064 520096 999076
rect 520148 999064 520154 999116
rect 357158 998996 357164 999048
rect 357216 999036 357222 999048
rect 361574 999036 361580 999048
rect 357216 999008 361580 999036
rect 357216 998996 357222 999008
rect 361574 998996 361580 999008
rect 361632 998996 361638 999048
rect 469214 998860 469220 998912
rect 469272 998900 469278 998912
rect 472250 998900 472256 998912
rect 469272 998872 472256 998900
rect 469272 998860 469278 998872
rect 472250 998860 472256 998872
rect 472308 998860 472314 998912
rect 516778 998656 516784 998708
rect 516836 998696 516842 998708
rect 524046 998696 524052 998708
rect 516836 998668 524052 998696
rect 516836 998656 516842 998668
rect 524046 998656 524052 998668
rect 524104 998656 524110 998708
rect 452562 998588 452568 998640
rect 452620 998628 452626 998640
rect 459646 998628 459652 998640
rect 452620 998600 459652 998628
rect 452620 998588 452626 998600
rect 459646 998588 459652 998600
rect 459704 998588 459710 998640
rect 499022 998588 499028 998640
rect 499080 998628 499086 998640
rect 516870 998628 516876 998640
rect 499080 998600 516876 998628
rect 499080 998588 499086 998600
rect 516870 998588 516876 998600
rect 516928 998588 516934 998640
rect 423398 998520 423404 998572
rect 423456 998560 423462 998572
rect 472158 998560 472164 998572
rect 423456 998532 472164 998560
rect 423456 998520 423462 998532
rect 472158 998520 472164 998532
rect 472216 998520 472222 998572
rect 499206 998520 499212 998572
rect 499264 998560 499270 998572
rect 516962 998560 516968 998572
rect 499264 998532 516968 998560
rect 499264 998520 499270 998532
rect 516962 998520 516968 998532
rect 517020 998520 517026 998572
rect 368474 998452 368480 998504
rect 368532 998492 368538 998504
rect 383378 998492 383384 998504
rect 368532 998464 383384 998492
rect 368532 998452 368538 998464
rect 383378 998452 383384 998464
rect 383436 998452 383442 998504
rect 425698 998452 425704 998504
rect 425756 998492 425762 998504
rect 472618 998492 472624 998504
rect 425756 998464 472624 998492
rect 425756 998452 425762 998464
rect 472618 998452 472624 998464
rect 472676 998452 472682 998504
rect 504358 998452 504364 998504
rect 504416 998492 504422 998504
rect 522390 998492 522396 998504
rect 504416 998464 522396 998492
rect 504416 998452 504422 998464
rect 522390 998452 522396 998464
rect 522448 998452 522454 998504
rect 360838 998384 360844 998436
rect 360896 998424 360902 998436
rect 380894 998424 380900 998436
rect 360896 998396 380900 998424
rect 360896 998384 360902 998396
rect 380894 998384 380900 998396
rect 380952 998384 380958 998436
rect 422018 998384 422024 998436
rect 422076 998424 422082 998436
rect 422076 998396 451274 998424
rect 422076 998384 422082 998396
rect 451246 998220 451274 998396
rect 465718 998384 465724 998436
rect 465776 998424 465782 998436
rect 472526 998424 472532 998436
rect 465776 998396 472532 998424
rect 465776 998384 465782 998396
rect 472526 998384 472532 998396
rect 472584 998384 472590 998436
rect 502150 998384 502156 998436
rect 502208 998424 502214 998436
rect 524046 998424 524052 998436
rect 502208 998396 524052 998424
rect 502208 998384 502214 998396
rect 524046 998384 524052 998396
rect 524104 998384 524110 998436
rect 549070 998384 549076 998436
rect 549128 998424 549134 998436
rect 572714 998424 572720 998436
rect 549128 998396 572720 998424
rect 549128 998384 549134 998396
rect 572714 998384 572720 998396
rect 572772 998384 572778 998436
rect 472342 998220 472348 998232
rect 451246 998192 472348 998220
rect 472342 998180 472348 998192
rect 472400 998180 472406 998232
rect 430850 998112 430856 998164
rect 430908 998152 430914 998164
rect 433978 998152 433984 998164
rect 430908 998124 433984 998152
rect 430908 998112 430914 998124
rect 433978 998112 433984 998124
rect 434036 998112 434042 998164
rect 149054 998044 149060 998096
rect 149112 998084 149118 998096
rect 152918 998084 152924 998096
rect 149112 998056 152924 998084
rect 149112 998044 149118 998056
rect 152918 998044 152924 998056
rect 152976 998044 152982 998096
rect 431678 998044 431684 998096
rect 431736 998084 431742 998096
rect 434162 998084 434168 998096
rect 431736 998056 434168 998084
rect 431736 998044 431742 998056
rect 434162 998044 434168 998056
rect 434220 998044 434226 998096
rect 148318 997976 148324 998028
rect 148376 998016 148382 998028
rect 151262 998016 151268 998028
rect 148376 997988 151268 998016
rect 148376 997976 148382 997988
rect 151262 997976 151268 997988
rect 151320 997976 151326 998028
rect 429654 997976 429660 998028
rect 429712 998016 429718 998028
rect 431954 998016 431960 998028
rect 429712 997988 431960 998016
rect 429712 997976 429718 997988
rect 431954 997976 431960 997988
rect 432012 997976 432018 998028
rect 151078 997908 151084 997960
rect 151136 997948 151142 997960
rect 153746 997948 153752 997960
rect 151136 997920 153752 997948
rect 151136 997908 151142 997920
rect 153746 997908 153752 997920
rect 153804 997908 153810 997960
rect 246666 997908 246672 997960
rect 246724 997948 246730 997960
rect 248414 997948 248420 997960
rect 246724 997920 248420 997948
rect 246724 997908 246730 997920
rect 248414 997908 248420 997920
rect 248472 997908 248478 997960
rect 428458 997908 428464 997960
rect 428516 997948 428522 997960
rect 430850 997948 430856 997960
rect 428516 997920 430856 997948
rect 428516 997908 428522 997920
rect 430850 997908 430856 997920
rect 430908 997908 430914 997960
rect 432874 997908 432880 997960
rect 432932 997948 432938 997960
rect 436738 997948 436744 997960
rect 432932 997920 436744 997948
rect 432932 997908 432938 997920
rect 436738 997908 436744 997920
rect 436796 997908 436802 997960
rect 518986 997908 518992 997960
rect 519044 997948 519050 997960
rect 523954 997948 523960 997960
rect 519044 997920 523960 997948
rect 519044 997908 519050 997920
rect 523954 997908 523960 997920
rect 524012 997908 524018 997960
rect 92606 997840 92612 997892
rect 92664 997880 92670 997892
rect 94498 997880 94504 997892
rect 92664 997852 94504 997880
rect 92664 997840 92670 997852
rect 94498 997840 94504 997852
rect 94556 997840 94562 997892
rect 150342 997840 150348 997892
rect 150400 997880 150406 997892
rect 152550 997880 152556 997892
rect 150400 997852 152556 997880
rect 150400 997840 150406 997852
rect 152550 997840 152556 997852
rect 152608 997840 152614 997892
rect 298278 997840 298284 997892
rect 298336 997880 298342 997892
rect 298336 997852 306374 997880
rect 298336 997840 298342 997852
rect 151262 997772 151268 997824
rect 151320 997812 151326 997824
rect 153378 997812 153384 997824
rect 151320 997784 153384 997812
rect 151320 997772 151326 997784
rect 153378 997772 153384 997784
rect 153436 997772 153442 997824
rect 246758 997772 246764 997824
rect 246816 997812 246822 997824
rect 253658 997812 253664 997824
rect 246816 997784 253664 997812
rect 246816 997772 246822 997784
rect 253658 997772 253664 997784
rect 253716 997772 253722 997824
rect 303246 997772 303252 997824
rect 303304 997812 303310 997824
rect 305822 997812 305828 997824
rect 303304 997784 305828 997812
rect 303304 997772 303310 997784
rect 305822 997772 305828 997784
rect 305880 997772 305886 997824
rect 306346 997812 306374 997852
rect 430390 997840 430396 997892
rect 430448 997880 430454 997892
rect 432138 997880 432144 997892
rect 430448 997852 432144 997880
rect 430448 997840 430454 997852
rect 432138 997840 432144 997852
rect 432196 997840 432202 997892
rect 432414 997840 432420 997892
rect 432472 997880 432478 997892
rect 435542 997880 435548 997892
rect 432472 997852 435548 997880
rect 432472 997840 432478 997852
rect 435542 997840 435548 997852
rect 435600 997840 435606 997892
rect 328362 997812 328368 997824
rect 306346 997784 328368 997812
rect 328362 997772 328368 997784
rect 328420 997772 328426 997824
rect 378778 997772 378784 997824
rect 378836 997812 378842 997824
rect 383470 997812 383476 997824
rect 378836 997784 383476 997812
rect 378836 997772 378842 997784
rect 383470 997772 383476 997784
rect 383528 997772 383534 997824
rect 429194 997772 429200 997824
rect 429252 997812 429258 997824
rect 431218 997812 431224 997824
rect 429252 997784 431224 997812
rect 429252 997772 429258 997784
rect 431218 997772 431224 997784
rect 431276 997772 431282 997824
rect 432046 997772 432052 997824
rect 432104 997812 432110 997824
rect 433334 997812 433340 997824
rect 432104 997784 433340 997812
rect 432104 997772 432110 997784
rect 433334 997772 433340 997784
rect 433392 997772 433398 997824
rect 625798 997812 625804 997824
rect 612752 997784 625804 997812
rect 109862 997704 109868 997756
rect 109920 997744 109926 997756
rect 117222 997744 117228 997756
rect 109920 997716 117228 997744
rect 109920 997704 109926 997716
rect 117222 997704 117228 997716
rect 117280 997704 117286 997756
rect 160738 997704 160744 997756
rect 160796 997744 160802 997756
rect 167546 997744 167552 997756
rect 160796 997716 167552 997744
rect 160796 997704 160802 997716
rect 167546 997704 167552 997716
rect 167604 997704 167610 997756
rect 195238 997704 195244 997756
rect 195296 997744 195302 997756
rect 211154 997744 211160 997756
rect 195296 997716 211160 997744
rect 195296 997704 195302 997716
rect 211154 997704 211160 997716
rect 211212 997704 211218 997756
rect 213362 997704 213368 997756
rect 213420 997744 213426 997756
rect 218882 997744 218888 997756
rect 213420 997716 218888 997744
rect 213420 997704 213426 997716
rect 218882 997704 218888 997716
rect 218940 997704 218946 997756
rect 246574 997704 246580 997756
rect 246632 997744 246638 997756
rect 260834 997744 260840 997756
rect 246632 997716 260840 997744
rect 246632 997704 246638 997716
rect 260834 997704 260840 997716
rect 260892 997704 260898 997756
rect 265802 997704 265808 997756
rect 265860 997744 265866 997756
rect 270402 997744 270408 997756
rect 265860 997716 270408 997744
rect 265860 997704 265866 997716
rect 270402 997704 270408 997716
rect 270460 997704 270466 997756
rect 298738 997704 298744 997756
rect 298796 997744 298802 997756
rect 316034 997744 316040 997756
rect 298796 997716 316040 997744
rect 298796 997704 298802 997716
rect 316034 997704 316040 997716
rect 316092 997704 316098 997756
rect 362218 997704 362224 997756
rect 362276 997744 362282 997756
rect 372338 997744 372344 997756
rect 362276 997716 372344 997744
rect 362276 997704 362282 997716
rect 372338 997704 372344 997716
rect 372396 997704 372402 997756
rect 399938 997704 399944 997756
rect 399996 997744 400002 997756
rect 433426 997744 433432 997756
rect 399996 997716 433432 997744
rect 399996 997704 400002 997716
rect 433426 997704 433432 997716
rect 433484 997704 433490 997756
rect 434162 997704 434168 997756
rect 434220 997744 434226 997756
rect 439682 997744 439688 997756
rect 434220 997716 439688 997744
rect 434220 997704 434226 997716
rect 439682 997704 439688 997716
rect 439740 997704 439746 997756
rect 488902 997704 488908 997756
rect 488960 997744 488966 997756
rect 510706 997744 510712 997756
rect 488960 997716 510712 997744
rect 488960 997704 488966 997716
rect 510706 997704 510712 997716
rect 510764 997704 510770 997756
rect 513926 997704 513932 997756
rect 513984 997744 513990 997756
rect 516686 997744 516692 997756
rect 513984 997716 516692 997744
rect 513984 997704 513990 997716
rect 516686 997704 516692 997716
rect 516744 997704 516750 997756
rect 540882 997704 540888 997756
rect 540940 997744 540946 997756
rect 563054 997744 563060 997756
rect 540940 997716 563060 997744
rect 540940 997704 540946 997716
rect 563054 997704 563060 997716
rect 563112 997704 563118 997756
rect 567286 997704 567292 997756
rect 567344 997744 567350 997756
rect 612752 997744 612780 997784
rect 625798 997772 625804 997784
rect 625856 997772 625862 997824
rect 567344 997716 612780 997744
rect 567344 997704 567350 997716
rect 111058 997636 111064 997688
rect 111116 997676 111122 997688
rect 116302 997676 116308 997688
rect 111116 997648 116308 997676
rect 111116 997636 111122 997648
rect 116302 997636 116308 997648
rect 116360 997636 116366 997688
rect 144822 997636 144828 997688
rect 144880 997676 144886 997688
rect 160186 997676 160192 997688
rect 144880 997648 160192 997676
rect 144880 997636 144886 997648
rect 160186 997636 160192 997648
rect 160244 997636 160250 997688
rect 162302 997636 162308 997688
rect 162360 997676 162366 997688
rect 167638 997676 167644 997688
rect 162360 997648 167644 997676
rect 162360 997636 162366 997648
rect 167638 997636 167644 997648
rect 167696 997636 167702 997688
rect 201402 997636 201408 997688
rect 201460 997676 201466 997688
rect 203702 997676 203708 997688
rect 201460 997648 203708 997676
rect 201460 997636 201466 997648
rect 203702 997636 203708 997648
rect 203760 997636 203766 997688
rect 366542 997636 366548 997688
rect 366600 997676 366606 997688
rect 372430 997676 372436 997688
rect 366600 997648 372436 997676
rect 366600 997636 366606 997648
rect 372430 997636 372436 997648
rect 372488 997636 372494 997688
rect 400030 997636 400036 997688
rect 400088 997676 400094 997688
rect 432138 997676 432144 997688
rect 400088 997648 432144 997676
rect 400088 997636 400094 997648
rect 432138 997636 432144 997648
rect 432196 997636 432202 997688
rect 511258 997636 511264 997688
rect 511316 997676 511322 997688
rect 516778 997676 516784 997688
rect 511316 997648 516784 997676
rect 511316 997636 511322 997648
rect 516778 997636 516784 997648
rect 516836 997636 516842 997688
rect 568206 997636 568212 997688
rect 568264 997676 568270 997688
rect 611354 997676 611360 997688
rect 568264 997648 611360 997676
rect 568264 997636 568270 997648
rect 611354 997636 611360 997648
rect 611412 997636 611418 997688
rect 144730 997568 144736 997620
rect 144788 997608 144794 997620
rect 161474 997608 161480 997620
rect 144788 997580 161480 997608
rect 144788 997568 144794 997580
rect 161474 997568 161480 997580
rect 161532 997568 161538 997620
rect 365162 997568 365168 997620
rect 365220 997608 365226 997620
rect 372522 997608 372528 997620
rect 365220 997580 372528 997608
rect 365220 997568 365226 997580
rect 372522 997568 372528 997580
rect 372580 997568 372586 997620
rect 550358 997568 550364 997620
rect 550416 997608 550422 997620
rect 550416 997580 590700 997608
rect 550416 997568 550422 997580
rect 564986 997500 564992 997552
rect 565044 997540 565050 997552
rect 565044 997532 590534 997540
rect 565044 997512 590476 997532
rect 565044 997500 565050 997512
rect 565170 997432 565176 997484
rect 565228 997472 565234 997484
rect 590470 997480 590476 997512
rect 590528 997480 590534 997532
rect 565228 997444 590376 997472
rect 565228 997432 565234 997444
rect 590348 997432 590376 997444
rect 590562 997432 590568 997444
rect 590348 997404 590568 997432
rect 590562 997392 590568 997404
rect 590620 997392 590626 997444
rect 143994 997296 144000 997348
rect 144052 997336 144058 997348
rect 147030 997336 147036 997348
rect 144052 997308 147036 997336
rect 144052 997296 144058 997308
rect 147030 997296 147036 997308
rect 147088 997296 147094 997348
rect 202046 997296 202052 997348
rect 202104 997336 202110 997348
rect 204898 997336 204904 997348
rect 202104 997308 204904 997336
rect 202104 997296 202110 997308
rect 204898 997296 204904 997308
rect 204956 997296 204962 997348
rect 590378 997284 590384 997336
rect 590436 997324 590442 997336
rect 590672 997324 590700 997580
rect 590436 997296 590700 997324
rect 590436 997284 590442 997296
rect 200206 997228 200212 997280
rect 200264 997268 200270 997280
rect 204990 997268 204996 997280
rect 200264 997240 204996 997268
rect 200264 997228 200270 997240
rect 204990 997228 204996 997240
rect 205048 997228 205054 997280
rect 573358 997160 573364 997212
rect 573416 997200 573422 997212
rect 620278 997200 620284 997212
rect 573416 997172 620284 997200
rect 573416 997160 573422 997172
rect 620278 997160 620284 997172
rect 620336 997160 620342 997212
rect 559742 997092 559748 997144
rect 559800 997132 559806 997144
rect 618162 997132 618168 997144
rect 559800 997104 618168 997132
rect 559800 997092 559806 997104
rect 618162 997092 618168 997104
rect 618220 997092 618226 997144
rect 328362 997024 328368 997076
rect 328420 997064 328426 997076
rect 381170 997064 381176 997076
rect 328420 997036 381176 997064
rect 328420 997024 328426 997036
rect 381170 997024 381176 997036
rect 381228 997024 381234 997076
rect 550450 997024 550456 997076
rect 550508 997064 550514 997076
rect 622394 997064 622400 997076
rect 550508 997036 622400 997064
rect 550508 997024 550514 997036
rect 622394 997024 622400 997036
rect 622452 997024 622458 997076
rect 195238 996820 195244 996872
rect 195296 996860 195302 996872
rect 199378 996860 199384 996872
rect 195296 996832 199384 996860
rect 195296 996820 195302 996832
rect 199378 996820 199384 996832
rect 199436 996820 199442 996872
rect 195974 996752 195980 996804
rect 196032 996792 196038 996804
rect 202322 996792 202328 996804
rect 196032 996764 202328 996792
rect 196032 996752 196038 996764
rect 202322 996752 202328 996764
rect 202380 996752 202386 996804
rect 303246 996412 303252 996464
rect 303304 996452 303310 996464
rect 304258 996452 304264 996464
rect 303304 996424 304264 996452
rect 303304 996412 303310 996424
rect 304258 996412 304264 996424
rect 304316 996412 304322 996464
rect 299290 996344 299296 996396
rect 299348 996384 299354 996396
rect 305638 996384 305644 996396
rect 299348 996356 305644 996384
rect 299348 996344 299354 996356
rect 305638 996344 305644 996356
rect 305696 996344 305702 996396
rect 159358 996140 159364 996192
rect 159416 996180 159422 996192
rect 209774 996180 209780 996192
rect 159416 996172 178862 996180
rect 195126 996172 209780 996180
rect 159416 996152 209780 996172
rect 159416 996140 159422 996152
rect 178832 996144 195160 996152
rect 209774 996140 209780 996152
rect 209832 996140 209838 996192
rect 262858 996140 262864 996192
rect 262916 996180 262922 996192
rect 313550 996180 313556 996192
rect 262916 996172 281886 996180
rect 298146 996172 313556 996180
rect 262916 996152 313556 996172
rect 262916 996140 262922 996152
rect 281856 996144 298172 996152
rect 313550 996140 313556 996152
rect 313608 996140 313614 996192
rect 364978 996140 364984 996192
rect 365036 996180 365042 996192
rect 431954 996180 431960 996192
rect 365036 996172 383692 996180
rect 399908 996172 431960 996180
rect 365036 996152 431960 996172
rect 365036 996140 365042 996152
rect 383662 996144 399940 996152
rect 431954 996140 431960 996152
rect 432012 996140 432018 996192
rect 433978 996140 433984 996192
rect 434036 996180 434042 996192
rect 510614 996180 510620 996192
rect 434036 996172 472732 996180
rect 488908 996172 510620 996180
rect 434036 996152 510620 996172
rect 434036 996140 434042 996152
rect 472700 996144 488940 996152
rect 510614 996140 510620 996152
rect 510672 996140 510678 996192
rect 556706 996140 556712 996192
rect 556764 996180 556770 996192
rect 556764 996152 625154 996180
rect 556764 996140 556770 996152
rect 108298 996072 108304 996124
rect 108356 996112 108362 996124
rect 158714 996112 158720 996124
rect 108356 996084 158720 996112
rect 108356 996072 108362 996084
rect 158714 996072 158720 996084
rect 158772 996072 158778 996124
rect 162118 996072 162124 996124
rect 162176 996112 162182 996124
rect 207658 996112 207664 996124
rect 162176 996084 207664 996112
rect 162176 996072 162182 996084
rect 207658 996072 207664 996084
rect 207716 996072 207722 996124
rect 211798 996072 211804 996124
rect 211856 996112 211862 996124
rect 261478 996112 261484 996124
rect 211856 996084 261484 996112
rect 211856 996072 211862 996084
rect 261478 996072 261484 996084
rect 261536 996072 261542 996124
rect 264238 996072 264244 996124
rect 264296 996112 264302 996124
rect 313366 996112 313372 996124
rect 264296 996084 313372 996112
rect 264296 996072 264302 996084
rect 313366 996072 313372 996084
rect 313424 996072 313430 996124
rect 366358 996072 366364 996124
rect 366416 996112 366422 996124
rect 428458 996112 428464 996124
rect 366416 996084 428464 996112
rect 366416 996072 366422 996084
rect 428458 996072 428464 996084
rect 428516 996072 428522 996124
rect 431218 996072 431224 996124
rect 431276 996112 431282 996124
rect 506566 996112 506572 996124
rect 431276 996084 506572 996112
rect 431276 996072 431282 996084
rect 506566 996072 506572 996084
rect 506624 996072 506630 996124
rect 508498 996072 508504 996124
rect 508556 996112 508562 996124
rect 560570 996112 560576 996124
rect 508556 996084 560576 996112
rect 508556 996072 508562 996084
rect 560570 996072 560576 996084
rect 560628 996072 560634 996124
rect 109586 996004 109592 996056
rect 109644 996044 109650 996056
rect 160094 996044 160100 996056
rect 109644 996016 160100 996044
rect 109644 996004 109650 996016
rect 160094 996004 160100 996016
rect 160152 996004 160158 996056
rect 228450 996004 228456 996056
rect 228508 996044 228514 996056
rect 262214 996044 262220 996056
rect 228508 996016 262220 996044
rect 228508 996004 228514 996016
rect 262214 996004 262220 996016
rect 262272 996004 262278 996056
rect 269758 996004 269764 996056
rect 269816 996044 269822 996056
rect 314654 996044 314660 996056
rect 269816 996016 314660 996044
rect 269816 996004 269822 996016
rect 314654 996004 314660 996016
rect 314712 996004 314718 996056
rect 361574 996004 361580 996056
rect 361632 996044 361638 996056
rect 361632 996016 373994 996044
rect 361632 996004 361638 996016
rect 298922 995976 298928 995988
rect 290660 995948 298928 995976
rect 150342 995908 150348 995920
rect 139228 995880 150348 995908
rect 139228 995852 139256 995880
rect 150342 995868 150348 995880
rect 150400 995868 150406 995920
rect 213178 995868 213184 995920
rect 213236 995908 213242 995920
rect 263594 995908 263600 995920
rect 213236 995880 263600 995908
rect 213236 995868 213242 995880
rect 263594 995868 263600 995880
rect 263652 995868 263658 995920
rect 290660 995852 290688 995948
rect 298922 995936 298928 995948
rect 298980 995936 298986 995988
rect 298462 995908 298468 995920
rect 291120 995880 298468 995908
rect 291120 995852 291148 995880
rect 298462 995868 298468 995880
rect 298520 995868 298526 995920
rect 373966 995908 373994 996016
rect 468478 996004 468484 996056
rect 468536 996044 468542 996056
rect 509234 996044 509240 996056
rect 468536 996016 509240 996044
rect 468536 996004 468542 996016
rect 509234 996004 509240 996016
rect 509292 996004 509298 996056
rect 510062 996004 510068 996056
rect 510120 996044 510126 996056
rect 561766 996044 561772 996056
rect 510120 996016 561772 996044
rect 510120 996004 510126 996016
rect 561766 996004 561772 996016
rect 561824 996004 561830 996056
rect 504266 995936 504272 995988
rect 504324 995976 504330 995988
rect 504324 995948 532372 995976
rect 504324 995936 504330 995948
rect 373966 995880 391796 995908
rect 391768 995852 391796 995880
rect 472342 995868 472348 995920
rect 472400 995908 472406 995920
rect 472400 995880 478276 995908
rect 472400 995868 472406 995880
rect 478248 995852 478276 995880
rect 509786 995868 509792 995920
rect 509844 995908 509850 995920
rect 509844 995880 528554 995908
rect 509844 995868 509850 995880
rect 85298 995800 85304 995852
rect 85356 995840 85362 995852
rect 92238 995840 92244 995852
rect 85356 995812 92244 995840
rect 85356 995800 85362 995812
rect 92238 995800 92244 995812
rect 92296 995800 92302 995852
rect 139210 995800 139216 995852
rect 139268 995800 139274 995852
rect 140498 995800 140504 995852
rect 140556 995840 140562 995852
rect 143718 995840 143724 995852
rect 140556 995812 143724 995840
rect 140556 995800 140562 995812
rect 143718 995800 143724 995812
rect 143776 995800 143782 995852
rect 192478 995800 192484 995852
rect 192536 995840 192542 995852
rect 195146 995840 195152 995852
rect 192536 995812 195152 995840
rect 192536 995800 192542 995812
rect 195146 995800 195152 995812
rect 195204 995800 195210 995852
rect 242066 995800 242072 995852
rect 242124 995840 242130 995852
rect 247678 995840 247684 995852
rect 242124 995812 247684 995840
rect 242124 995800 242130 995812
rect 247678 995800 247684 995812
rect 247736 995800 247742 995852
rect 290642 995800 290648 995852
rect 290700 995800 290706 995852
rect 291102 995800 291108 995852
rect 291160 995800 291166 995852
rect 292482 995800 292488 995852
rect 292540 995840 292546 995852
rect 298830 995840 298836 995852
rect 292540 995812 298836 995840
rect 292540 995800 292546 995812
rect 298830 995800 298836 995812
rect 298888 995800 298894 995852
rect 383378 995800 383384 995852
rect 383436 995840 383442 995852
rect 385678 995840 385684 995852
rect 383436 995812 385684 995840
rect 383436 995800 383442 995812
rect 385678 995800 385684 995812
rect 385736 995800 385742 995852
rect 391750 995800 391756 995852
rect 391808 995800 391814 995852
rect 472526 995800 472532 995852
rect 472584 995840 472590 995852
rect 473354 995840 473360 995852
rect 472584 995812 473360 995840
rect 472584 995800 472590 995812
rect 473354 995800 473360 995812
rect 473412 995800 473418 995852
rect 478230 995800 478236 995852
rect 478288 995800 478294 995852
rect 523954 995800 523960 995852
rect 524012 995840 524018 995852
rect 525334 995840 525340 995852
rect 524012 995812 525340 995840
rect 524012 995800 524018 995812
rect 525334 995800 525340 995812
rect 525392 995800 525398 995852
rect 91554 995732 91560 995784
rect 91612 995772 91618 995784
rect 92330 995772 92336 995784
rect 91612 995744 92336 995772
rect 91612 995732 91618 995744
rect 92330 995732 92336 995744
rect 92388 995732 92394 995784
rect 141050 995732 141056 995784
rect 141108 995772 141114 995784
rect 143810 995772 143816 995784
rect 141108 995744 143816 995772
rect 141108 995732 141114 995744
rect 143810 995732 143816 995744
rect 143868 995732 143874 995784
rect 190454 995732 190460 995784
rect 190512 995772 190518 995784
rect 195330 995772 195336 995784
rect 190512 995744 195336 995772
rect 190512 995732 190518 995744
rect 195330 995732 195336 995744
rect 195388 995732 195394 995784
rect 245562 995732 245568 995784
rect 245620 995772 245626 995784
rect 246666 995772 246672 995784
rect 245620 995744 246672 995772
rect 245620 995732 245626 995744
rect 246666 995732 246672 995744
rect 246724 995732 246730 995784
rect 297266 995732 297272 995784
rect 297324 995772 297330 995784
rect 298042 995772 298048 995784
rect 297324 995744 298048 995772
rect 297324 995732 297330 995744
rect 298042 995732 298048 995744
rect 298100 995732 298106 995784
rect 383634 995732 383640 995784
rect 383692 995772 383698 995784
rect 384390 995772 384396 995784
rect 383692 995744 384396 995772
rect 383692 995732 383698 995744
rect 384390 995732 384396 995744
rect 384448 995732 384454 995784
rect 432046 995732 432052 995784
rect 432104 995772 432110 995784
rect 439774 995772 439780 995784
rect 432104 995744 439780 995772
rect 432104 995732 432110 995744
rect 439774 995732 439780 995744
rect 439832 995732 439838 995784
rect 472434 995732 472440 995784
rect 472492 995772 472498 995784
rect 474734 995772 474740 995784
rect 472492 995744 474740 995772
rect 472492 995732 472498 995744
rect 474734 995732 474740 995744
rect 474792 995732 474798 995784
rect 524138 995732 524144 995784
rect 524196 995772 524202 995784
rect 524782 995772 524788 995784
rect 524196 995744 524788 995772
rect 524196 995732 524202 995744
rect 524782 995732 524788 995744
rect 524840 995732 524846 995784
rect 528526 995772 528554 995880
rect 532344 995840 532372 995948
rect 560294 995908 560300 995920
rect 538186 995880 560300 995908
rect 533430 995840 533436 995852
rect 532344 995812 533436 995840
rect 533430 995800 533436 995812
rect 533488 995800 533494 995852
rect 538186 995772 538214 995880
rect 560294 995868 560300 995880
rect 560352 995868 560358 995920
rect 557534 995800 557540 995852
rect 557592 995840 557598 995852
rect 568206 995840 568212 995852
rect 557592 995812 568212 995840
rect 557592 995800 557598 995812
rect 568206 995800 568212 995812
rect 568264 995800 568270 995852
rect 625126 995840 625154 996152
rect 634722 995840 634728 995852
rect 625126 995812 634728 995840
rect 634722 995800 634728 995812
rect 634780 995800 634786 995852
rect 528526 995744 538214 995772
rect 625798 995732 625804 995784
rect 625856 995772 625862 995784
rect 627178 995772 627184 995784
rect 625856 995744 627184 995772
rect 625856 995732 625862 995744
rect 627178 995732 627184 995744
rect 627236 995732 627242 995784
rect 87874 995664 87880 995716
rect 87932 995704 87938 995716
rect 92422 995704 92428 995716
rect 87932 995676 92428 995704
rect 87932 995664 87938 995676
rect 92422 995664 92428 995676
rect 92480 995664 92486 995716
rect 136266 995664 136272 995716
rect 136324 995704 136330 995716
rect 144086 995704 144092 995716
rect 136324 995676 144092 995704
rect 136324 995664 136330 995676
rect 144086 995664 144092 995676
rect 144144 995664 144150 995716
rect 235258 995664 235264 995716
rect 235316 995704 235322 995716
rect 247126 995704 247132 995716
rect 235316 995676 247132 995704
rect 235316 995664 235322 995676
rect 247126 995664 247132 995676
rect 247184 995664 247190 995716
rect 294874 995664 294880 995716
rect 294932 995704 294938 995716
rect 298278 995704 298284 995716
rect 294932 995676 298284 995704
rect 294932 995664 294938 995676
rect 298278 995664 298284 995676
rect 298336 995664 298342 995716
rect 383726 995664 383732 995716
rect 383784 995704 383790 995716
rect 388622 995704 388628 995716
rect 383784 995676 388628 995704
rect 383784 995664 383790 995676
rect 388622 995664 388628 995676
rect 388680 995664 388686 995716
rect 472250 995664 472256 995716
rect 472308 995704 472314 995716
rect 473998 995704 474004 995716
rect 472308 995676 474004 995704
rect 472308 995664 472314 995676
rect 473998 995664 474004 995676
rect 474056 995664 474062 995716
rect 523862 995664 523868 995716
rect 523920 995704 523926 995716
rect 529014 995704 529020 995716
rect 523920 995676 529020 995704
rect 523920 995664 523926 995676
rect 529014 995664 529020 995676
rect 529072 995664 529078 995716
rect 625706 995664 625712 995716
rect 625764 995704 625770 995716
rect 630858 995704 630864 995716
rect 625764 995676 630864 995704
rect 625764 995664 625770 995676
rect 630858 995664 630864 995676
rect 630916 995664 630922 995716
rect 169018 995596 169024 995648
rect 169076 995636 169082 995648
rect 184290 995636 184296 995648
rect 169076 995608 184296 995636
rect 169076 995596 169082 995608
rect 184290 995596 184296 995608
rect 184348 995596 184354 995648
rect 240870 995596 240876 995648
rect 240928 995636 240934 995648
rect 246758 995636 246764 995648
rect 240928 995608 246764 995636
rect 240928 995596 240934 995608
rect 246758 995596 246764 995608
rect 246816 995596 246822 995648
rect 295426 995596 295432 995648
rect 295484 995636 295490 995648
rect 298370 995636 298376 995648
rect 295484 995608 298376 995636
rect 295484 995596 295490 995608
rect 298370 995596 298376 995608
rect 298428 995596 298434 995648
rect 472158 995596 472164 995648
rect 472216 995636 472222 995648
rect 477678 995636 477684 995648
rect 472216 995608 477684 995636
rect 472216 995596 472222 995608
rect 477678 995596 477684 995608
rect 477736 995596 477742 995648
rect 472066 995528 472072 995580
rect 472124 995568 472130 995580
rect 476942 995568 476948 995580
rect 472124 995540 476948 995568
rect 472124 995528 472130 995540
rect 476942 995528 476948 995540
rect 477000 995528 477006 995580
rect 288066 995460 288072 995512
rect 288124 995500 288130 995512
rect 300118 995500 300124 995512
rect 288124 995472 300124 995500
rect 288124 995460 288130 995472
rect 300118 995460 300124 995472
rect 300176 995460 300182 995512
rect 286778 995392 286784 995444
rect 286836 995432 286842 995444
rect 299290 995432 299296 995444
rect 286836 995404 299296 995432
rect 286836 995392 286842 995404
rect 299290 995392 299296 995404
rect 299348 995392 299354 995444
rect 81250 995324 81256 995376
rect 81308 995364 81314 995376
rect 95878 995364 95884 995376
rect 81308 995336 95884 995364
rect 81308 995324 81314 995336
rect 95878 995324 95884 995336
rect 95936 995324 95942 995376
rect 287514 995324 287520 995376
rect 287572 995364 287578 995376
rect 301498 995364 301504 995376
rect 287572 995336 301504 995364
rect 287572 995324 287578 995336
rect 301498 995324 301504 995336
rect 301556 995324 301562 995376
rect 78306 995256 78312 995308
rect 78364 995296 78370 995308
rect 95970 995296 95976 995308
rect 78364 995268 95976 995296
rect 78364 995256 78370 995268
rect 95970 995256 95976 995268
rect 96028 995256 96034 995308
rect 133414 995256 133420 995308
rect 133472 995296 133478 995308
rect 145558 995296 145564 995308
rect 133472 995268 145564 995296
rect 133472 995256 133478 995268
rect 145558 995256 145564 995268
rect 145616 995256 145622 995308
rect 239260 995256 239266 995308
rect 239318 995296 239324 995308
rect 251818 995296 251824 995308
rect 239318 995268 251824 995296
rect 239318 995256 239324 995268
rect 251818 995256 251824 995268
rect 251876 995256 251882 995308
rect 359182 995256 359188 995308
rect 359240 995296 359246 995308
rect 392670 995296 392676 995308
rect 359240 995268 392676 995296
rect 359240 995256 359246 995268
rect 392670 995256 392676 995268
rect 392728 995256 392734 995308
rect 572714 995256 572720 995308
rect 572772 995296 572778 995308
rect 636148 995296 636154 995308
rect 572772 995268 636154 995296
rect 572772 995256 572778 995268
rect 636148 995256 636154 995268
rect 636206 995256 636212 995308
rect 80698 995188 80704 995240
rect 80756 995228 80762 995240
rect 100018 995228 100024 995240
rect 80756 995200 100024 995228
rect 80756 995188 80762 995200
rect 100018 995188 100024 995200
rect 100076 995188 100082 995240
rect 184152 995188 184158 995240
rect 184210 995228 184216 995240
rect 196618 995228 196624 995240
rect 184210 995200 196624 995228
rect 184210 995188 184216 995200
rect 196618 995188 196624 995200
rect 196676 995188 196682 995240
rect 235580 995188 235586 995240
rect 235638 995228 235644 995240
rect 250714 995228 250720 995240
rect 235638 995200 250720 995228
rect 235638 995188 235644 995200
rect 250714 995188 250720 995200
rect 250772 995188 250778 995240
rect 284110 995188 284116 995240
rect 284168 995228 284174 995240
rect 298646 995228 298652 995240
rect 284168 995200 298652 995228
rect 284168 995188 284174 995200
rect 298646 995188 298652 995200
rect 298704 995188 298710 995240
rect 567930 995188 567936 995240
rect 567988 995228 567994 995240
rect 637344 995228 637350 995240
rect 567988 995200 637350 995228
rect 567988 995188 567994 995200
rect 637344 995188 637350 995200
rect 637402 995188 637408 995240
rect 77662 995120 77668 995172
rect 77720 995160 77726 995172
rect 97350 995160 97356 995172
rect 77720 995132 97356 995160
rect 77720 995120 77726 995132
rect 97350 995120 97356 995132
rect 97408 995120 97414 995172
rect 129090 995120 129096 995172
rect 129148 995160 129154 995172
rect 151078 995160 151084 995172
rect 129148 995132 151084 995160
rect 129148 995120 129154 995132
rect 151078 995120 151084 995132
rect 151136 995120 151142 995172
rect 187602 995120 187608 995172
rect 187660 995160 187666 995172
rect 201402 995160 201408 995172
rect 187660 995132 201408 995160
rect 187660 995120 187666 995132
rect 201402 995120 201408 995132
rect 201460 995120 201466 995172
rect 231578 995120 231584 995172
rect 231636 995160 231642 995172
rect 249058 995160 249064 995172
rect 231636 995132 249064 995160
rect 231636 995120 231642 995132
rect 249058 995120 249064 995132
rect 249116 995120 249122 995172
rect 283466 995120 283472 995172
rect 283524 995160 283530 995172
rect 299382 995160 299388 995172
rect 283524 995132 299388 995160
rect 283524 995120 283530 995132
rect 299382 995120 299388 995132
rect 299440 995120 299446 995172
rect 354306 995120 354312 995172
rect 354364 995160 354370 995172
rect 393222 995160 393228 995172
rect 354364 995132 393228 995160
rect 354364 995120 354370 995132
rect 393222 995120 393228 995132
rect 393280 995120 393286 995172
rect 520090 995120 520096 995172
rect 520148 995160 520154 995172
rect 537386 995160 537392 995172
rect 520148 995132 537392 995160
rect 520148 995120 520154 995132
rect 537386 995120 537392 995132
rect 537444 995120 537450 995172
rect 570598 995120 570604 995172
rect 570656 995160 570662 995172
rect 638954 995160 638960 995172
rect 570656 995132 638960 995160
rect 570656 995120 570662 995132
rect 638954 995120 638960 995132
rect 639012 995120 639018 995172
rect 77018 995052 77024 995104
rect 77076 995092 77082 995104
rect 106642 995092 106648 995104
rect 77076 995064 106648 995092
rect 77076 995052 77082 995064
rect 106642 995052 106648 995064
rect 106700 995052 106706 995104
rect 129734 995052 129740 995104
rect 129792 995092 129798 995104
rect 155218 995092 155224 995104
rect 129792 995064 155224 995092
rect 129792 995052 129798 995064
rect 155218 995052 155224 995064
rect 155276 995052 155282 995104
rect 181438 995052 181444 995104
rect 181496 995092 181502 995104
rect 197998 995092 198004 995104
rect 181496 995064 198004 995092
rect 181496 995052 181502 995064
rect 197998 995052 198004 995064
rect 198056 995052 198062 995104
rect 232222 995052 232228 995104
rect 232280 995092 232286 995104
rect 254578 995092 254584 995104
rect 232280 995064 254584 995092
rect 232280 995052 232286 995064
rect 254578 995052 254584 995064
rect 254636 995052 254642 995104
rect 282822 995052 282828 995104
rect 282880 995092 282886 995104
rect 311894 995092 311900 995104
rect 282880 995064 311900 995092
rect 282880 995052 282886 995064
rect 311894 995052 311900 995064
rect 311952 995052 311958 995104
rect 371878 995052 371884 995104
rect 371936 995092 371942 995104
rect 396994 995092 397000 995104
rect 371936 995064 397000 995092
rect 371936 995052 371942 995064
rect 396994 995052 397000 995064
rect 397052 995052 397058 995104
rect 501966 995052 501972 995104
rect 502024 995092 502030 995104
rect 528738 995092 528744 995104
rect 502024 995064 528744 995092
rect 502024 995052 502030 995064
rect 528738 995052 528744 995064
rect 528796 995052 528802 995104
rect 553118 995052 553124 995104
rect 553176 995092 553182 995104
rect 633986 995092 633992 995104
rect 553176 995064 633992 995092
rect 553176 995052 553182 995064
rect 633986 995052 633992 995064
rect 634044 995052 634050 995104
rect 640702 995092 640708 995104
rect 634786 995064 640708 995092
rect 88702 994984 88708 995036
rect 88760 995024 88766 995036
rect 121730 995024 121736 995036
rect 88760 994996 121736 995024
rect 88760 994984 88766 994996
rect 121730 994984 121736 994996
rect 121788 994984 121794 995036
rect 180702 994984 180708 995036
rect 180760 995024 180766 995036
rect 202138 995024 202144 995036
rect 180760 994996 202144 995024
rect 180760 994984 180766 994996
rect 202138 994984 202144 994996
rect 202196 994984 202202 995036
rect 243262 994984 243268 995036
rect 243320 995024 243326 995036
rect 316402 995024 316408 995036
rect 243320 994996 316408 995024
rect 243320 994984 243326 994996
rect 316402 994984 316408 994996
rect 316460 994984 316466 995036
rect 357342 994984 357348 995036
rect 357400 995024 357406 995036
rect 398834 995024 398840 995036
rect 357400 994996 398840 995024
rect 357400 994984 357406 994996
rect 398834 994984 398840 994996
rect 398892 994984 398898 995036
rect 447134 994984 447140 995036
rect 447192 995024 447198 995036
rect 487798 995024 487804 995036
rect 447192 994996 487804 995024
rect 447192 994984 447198 994996
rect 487798 994984 487804 994996
rect 487856 994984 487862 995036
rect 501690 994984 501696 995036
rect 501748 995024 501754 995036
rect 535546 995024 535552 995036
rect 501748 994996 535552 995024
rect 501748 994984 501754 994996
rect 535546 994984 535552 994996
rect 535604 994984 535610 995036
rect 553394 994984 553400 995036
rect 553452 995024 553458 995036
rect 634786 995024 634814 995064
rect 640702 995052 640708 995064
rect 640760 995052 640766 995104
rect 553452 994996 634814 995024
rect 553452 994984 553458 994996
rect 638862 994984 638868 995036
rect 638920 995024 638926 995036
rect 640794 995024 640800 995036
rect 638920 994996 640800 995024
rect 638920 994984 638926 994996
rect 640794 994984 640800 994996
rect 640852 994984 640858 995036
rect 319438 992944 319444 992996
rect 319496 992984 319502 992996
rect 332594 992984 332600 992996
rect 319496 992956 332600 992984
rect 319496 992944 319502 992956
rect 332594 992944 332600 992956
rect 332652 992944 332658 992996
rect 367922 992944 367928 992996
rect 367980 992984 367986 992996
rect 429930 992984 429936 992996
rect 367980 992956 429936 992984
rect 367980 992944 367986 992956
rect 429930 992944 429936 992956
rect 429988 992944 429994 992996
rect 562502 992944 562508 992996
rect 562560 992984 562566 992996
rect 661678 992984 661684 992996
rect 562560 992956 661684 992984
rect 562560 992944 562566 992956
rect 661678 992944 661684 992956
rect 661736 992944 661742 992996
rect 48958 992876 48964 992928
rect 49016 992916 49022 992928
rect 110506 992916 110512 992928
rect 49016 992888 110512 992916
rect 49016 992876 49022 992888
rect 110506 992876 110512 992888
rect 110564 992876 110570 992928
rect 215294 992876 215300 992928
rect 215352 992916 215358 992928
rect 251450 992916 251456 992928
rect 215352 992888 251456 992916
rect 215352 992876 215358 992888
rect 251450 992876 251456 992888
rect 251508 992876 251514 992928
rect 265618 992876 265624 992928
rect 265676 992916 265682 992928
rect 300026 992916 300032 992928
rect 265676 992888 300032 992916
rect 265676 992876 265682 992888
rect 300026 992876 300032 992888
rect 300084 992876 300090 992928
rect 316678 992876 316684 992928
rect 316736 992916 316742 992928
rect 364978 992916 364984 992928
rect 316736 992888 364984 992916
rect 316736 992876 316742 992888
rect 364978 992876 364984 992888
rect 365036 992876 365042 992928
rect 420822 992876 420828 992928
rect 420880 992916 420886 992928
rect 666738 992916 666744 992928
rect 420880 992888 666744 992916
rect 420880 992876 420886 992888
rect 666738 992876 666744 992888
rect 666796 992876 666802 992928
rect 47578 991516 47584 991568
rect 47636 991556 47642 991568
rect 107746 991556 107752 991568
rect 47636 991528 107752 991556
rect 47636 991516 47642 991528
rect 107746 991516 107752 991528
rect 107804 991516 107810 991568
rect 512822 991516 512828 991568
rect 512880 991556 512886 991568
rect 527634 991556 527640 991568
rect 512880 991528 527640 991556
rect 512880 991516 512886 991528
rect 527634 991516 527640 991528
rect 527692 991516 527698 991568
rect 559558 991516 559564 991568
rect 559616 991556 559622 991568
rect 660298 991556 660304 991568
rect 559616 991528 660304 991556
rect 559616 991516 559622 991528
rect 660298 991516 660304 991528
rect 660356 991516 660362 991568
rect 44818 991448 44824 991500
rect 44876 991488 44882 991500
rect 109034 991488 109040 991500
rect 44876 991460 109040 991488
rect 44876 991448 44882 991460
rect 109034 991448 109040 991460
rect 109092 991448 109098 991500
rect 138290 991448 138296 991500
rect 138348 991488 138354 991500
rect 162946 991488 162952 991500
rect 138348 991460 162952 991488
rect 138348 991448 138354 991460
rect 162946 991448 162952 991460
rect 163004 991448 163010 991500
rect 203150 991448 203156 991500
rect 203208 991488 203214 991500
rect 213914 991488 213920 991500
rect 203208 991460 213920 991488
rect 203208 991448 203214 991460
rect 213914 991448 213920 991460
rect 213972 991448 213978 991500
rect 367738 991448 367744 991500
rect 367796 991488 367802 991500
rect 397822 991488 397828 991500
rect 367796 991460 397828 991488
rect 367796 991448 367802 991460
rect 397822 991448 397828 991460
rect 397880 991448 397886 991500
rect 435542 991448 435548 991500
rect 435600 991488 435606 991500
rect 495158 991488 495164 991500
rect 435600 991460 495164 991488
rect 435600 991448 435606 991460
rect 495158 991448 495164 991460
rect 495216 991448 495222 991500
rect 498102 991448 498108 991500
rect 498160 991488 498166 991500
rect 666554 991488 666560 991500
rect 498160 991460 666560 991488
rect 498160 991448 498166 991460
rect 666554 991448 666560 991460
rect 666612 991448 666618 991500
rect 214558 991176 214564 991228
rect 214616 991216 214622 991228
rect 219434 991216 219440 991228
rect 214616 991188 219440 991216
rect 214616 991176 214622 991188
rect 219434 991176 219440 991188
rect 219492 991176 219498 991228
rect 184290 990836 184296 990888
rect 184348 990876 184354 990888
rect 186958 990876 186964 990888
rect 184348 990848 186964 990876
rect 184348 990836 184354 990848
rect 186958 990836 186964 990848
rect 187016 990836 187022 990888
rect 267090 990836 267096 990888
rect 267148 990876 267154 990888
rect 268746 990876 268752 990888
rect 267148 990848 268752 990876
rect 267148 990836 267154 990848
rect 268746 990836 268752 990848
rect 268804 990836 268810 990888
rect 560938 990224 560944 990276
rect 560996 990264 561002 990276
rect 658918 990264 658924 990276
rect 560996 990236 658924 990264
rect 560996 990224 561002 990236
rect 658918 990224 658924 990236
rect 658976 990224 658982 990276
rect 562318 990156 562324 990208
rect 562376 990196 562382 990208
rect 669958 990196 669964 990208
rect 562376 990168 669964 990196
rect 562376 990156 562382 990168
rect 669958 990156 669964 990168
rect 670016 990156 670022 990208
rect 50338 990088 50344 990140
rect 50396 990128 50402 990140
rect 107930 990128 107936 990140
rect 50396 990100 107936 990128
rect 50396 990088 50402 990100
rect 107930 990088 107936 990100
rect 107988 990088 107994 990140
rect 353110 990088 353116 990140
rect 353168 990128 353174 990140
rect 666830 990128 666836 990140
rect 353168 990100 666836 990128
rect 353168 990088 353174 990100
rect 666830 990088 666836 990100
rect 666888 990088 666894 990140
rect 512638 988728 512644 988780
rect 512696 988768 512702 988780
rect 543826 988768 543832 988780
rect 512696 988740 543832 988768
rect 512696 988728 512702 988740
rect 543826 988728 543832 988740
rect 543884 988728 543890 988780
rect 563882 988728 563888 988780
rect 563940 988768 563946 988780
rect 592494 988768 592500 988780
rect 563940 988740 592500 988768
rect 563940 988728 563946 988740
rect 592494 988728 592500 988740
rect 592552 988728 592558 988780
rect 435358 987368 435364 987420
rect 435416 987408 435422 987420
rect 478966 987408 478972 987420
rect 435416 987380 478972 987408
rect 435416 987368 435422 987380
rect 478966 987368 478972 987380
rect 479024 987368 479030 987420
rect 563698 987368 563704 987420
rect 563756 987408 563762 987420
rect 608778 987408 608784 987420
rect 563756 987380 608784 987408
rect 563756 987368 563762 987380
rect 608778 987368 608784 987380
rect 608836 987368 608842 987420
rect 266998 986620 267004 986672
rect 267056 986660 267062 986672
rect 268102 986660 268108 986672
rect 267056 986632 268108 986660
rect 267056 986620 267062 986632
rect 268102 986620 268108 986632
rect 268160 986620 268166 986672
rect 89622 986008 89628 986060
rect 89680 986048 89686 986060
rect 111794 986048 111800 986060
rect 89680 986020 111800 986048
rect 89680 986008 89686 986020
rect 111794 986008 111800 986020
rect 111852 986008 111858 986060
rect 73430 985940 73436 985992
rect 73488 985980 73494 985992
rect 102778 985980 102784 985992
rect 73488 985952 102784 985980
rect 73488 985940 73494 985952
rect 102778 985940 102784 985952
rect 102836 985940 102842 985992
rect 215938 985940 215944 985992
rect 215996 985980 216002 985992
rect 235626 985980 235632 985992
rect 215996 985952 235632 985980
rect 215996 985940 216002 985952
rect 235626 985940 235632 985952
rect 235684 985940 235690 985992
rect 268746 985940 268752 985992
rect 268804 985980 268810 985992
rect 284294 985980 284300 985992
rect 268804 985952 284300 985980
rect 268804 985940 268810 985952
rect 284294 985940 284300 985952
rect 284352 985940 284358 985992
rect 318058 985940 318064 985992
rect 318116 985980 318122 985992
rect 349154 985980 349160 985992
rect 318116 985952 349160 985980
rect 318116 985940 318122 985952
rect 349154 985940 349160 985952
rect 349212 985940 349218 985992
rect 369118 985940 369124 985992
rect 369176 985980 369182 985992
rect 414106 985980 414112 985992
rect 369176 985952 414112 985980
rect 369176 985940 369182 985952
rect 414106 985940 414112 985952
rect 414164 985940 414170 985992
rect 436738 985940 436744 985992
rect 436796 985980 436802 985992
rect 462774 985980 462780 985992
rect 436796 985952 462780 985980
rect 436796 985940 436802 985952
rect 462774 985940 462780 985952
rect 462832 985940 462838 985992
rect 514018 985940 514024 985992
rect 514076 985980 514082 985992
rect 560110 985980 560116 985992
rect 514076 985952 560116 985980
rect 514076 985940 514082 985952
rect 560110 985940 560116 985952
rect 560168 985940 560174 985992
rect 565078 985940 565084 985992
rect 565136 985980 565142 985992
rect 624970 985980 624976 985992
rect 565136 985952 624976 985980
rect 565136 985940 565142 985952
rect 624970 985940 624976 985952
rect 625028 985940 625034 985992
rect 163498 985872 163504 985924
rect 163556 985912 163562 985924
rect 170766 985912 170772 985924
rect 163556 985884 170772 985912
rect 163556 985872 163562 985884
rect 170766 985872 170772 985884
rect 170824 985872 170830 985924
rect 549162 984920 549168 984972
rect 549220 984960 549226 984972
rect 666646 984960 666652 984972
rect 549220 984932 666652 984960
rect 549220 984920 549226 984932
rect 666646 984920 666652 984932
rect 666704 984920 666710 984972
rect 303522 984852 303528 984904
rect 303580 984892 303586 984904
rect 665450 984892 665456 984904
rect 303580 984864 665456 984892
rect 303580 984852 303586 984864
rect 665450 984852 665456 984864
rect 665508 984852 665514 984904
rect 280798 984784 280804 984836
rect 280856 984824 280862 984836
rect 650086 984824 650092 984836
rect 280856 984796 650092 984824
rect 280856 984784 280862 984796
rect 650086 984784 650092 984796
rect 650144 984784 650150 984836
rect 228358 984716 228364 984768
rect 228416 984756 228422 984768
rect 651466 984756 651472 984768
rect 228416 984728 651472 984756
rect 228416 984716 228422 984728
rect 651466 984716 651472 984728
rect 651524 984716 651530 984768
rect 177298 984648 177304 984700
rect 177356 984688 177362 984700
rect 649994 984688 650000 984700
rect 177356 984660 650000 984688
rect 177356 984648 177362 984660
rect 649994 984648 650000 984660
rect 650052 984648 650058 984700
rect 126238 984580 126244 984632
rect 126296 984620 126302 984632
rect 651374 984620 651380 984632
rect 126296 984592 651380 984620
rect 126296 984580 126302 984592
rect 651374 984580 651380 984592
rect 651432 984580 651438 984632
rect 42702 975672 42708 975724
rect 42760 975712 42766 975724
rect 62114 975712 62120 975724
rect 42760 975684 62120 975712
rect 42760 975672 42766 975684
rect 62114 975672 62120 975684
rect 62172 975672 62178 975724
rect 651650 975672 651656 975724
rect 651708 975712 651714 975724
rect 671338 975712 671344 975724
rect 651708 975684 671344 975712
rect 651708 975672 651714 975684
rect 671338 975672 671344 975684
rect 671396 975672 671402 975724
rect 42150 967240 42156 967292
rect 42208 967280 42214 967292
rect 42702 967280 42708 967292
rect 42208 967252 42708 967280
rect 42208 967240 42214 967252
rect 42702 967240 42708 967252
rect 42760 967240 42766 967292
rect 42150 963976 42156 964028
rect 42208 964016 42214 964028
rect 42794 964016 42800 964028
rect 42208 963988 42800 964016
rect 42208 963976 42214 963988
rect 42794 963976 42800 963988
rect 42852 963976 42858 964028
rect 42150 962820 42156 962872
rect 42208 962860 42214 962872
rect 42886 962860 42892 962872
rect 42208 962832 42892 962860
rect 42208 962820 42214 962832
rect 42886 962820 42892 962832
rect 42944 962820 42950 962872
rect 674834 962684 674840 962736
rect 674892 962724 674898 962736
rect 675478 962724 675484 962736
rect 674892 962696 675484 962724
rect 674892 962684 674898 962696
rect 675478 962684 675484 962696
rect 675536 962684 675542 962736
rect 675018 962004 675024 962056
rect 675076 962044 675082 962056
rect 675386 962044 675392 962056
rect 675076 962016 675392 962044
rect 675076 962004 675082 962016
rect 675386 962004 675392 962016
rect 675444 962004 675450 962056
rect 47670 961868 47676 961920
rect 47728 961908 47734 961920
rect 62114 961908 62120 961920
rect 47728 961880 62120 961908
rect 47728 961868 47734 961880
rect 62114 961868 62120 961880
rect 62172 961868 62178 961920
rect 42058 959692 42064 959744
rect 42116 959732 42122 959744
rect 44174 959732 44180 959744
rect 42116 959704 44180 959732
rect 42116 959692 42122 959704
rect 44174 959692 44180 959704
rect 44232 959692 44238 959744
rect 42150 959080 42156 959132
rect 42208 959120 42214 959132
rect 42978 959120 42984 959132
rect 42208 959092 42984 959120
rect 42208 959080 42214 959092
rect 42978 959080 42984 959092
rect 43036 959080 43042 959132
rect 673270 958332 673276 958384
rect 673328 958372 673334 958384
rect 675386 958372 675392 958384
rect 673328 958344 675392 958372
rect 673328 958332 673334 958344
rect 675386 958332 675392 958344
rect 675444 958332 675450 958384
rect 659010 957788 659016 957840
rect 659068 957828 659074 957840
rect 674834 957828 674840 957840
rect 659068 957800 674840 957828
rect 659068 957788 659074 957800
rect 674834 957788 674840 957800
rect 674892 957788 674898 957840
rect 674742 956972 674748 957024
rect 674800 957012 674806 957024
rect 675386 957012 675392 957024
rect 674800 956984 675392 957012
rect 674800 956972 674806 956984
rect 675386 956972 675392 956984
rect 675444 956972 675450 957024
rect 672350 956496 672356 956548
rect 672408 956536 672414 956548
rect 675018 956536 675024 956548
rect 672408 956508 675024 956536
rect 672408 956496 672414 956508
rect 675018 956496 675024 956508
rect 675076 956496 675082 956548
rect 674558 955680 674564 955732
rect 674616 955720 674622 955732
rect 675478 955720 675484 955732
rect 674616 955692 675484 955720
rect 674616 955680 674622 955692
rect 675478 955680 675484 955692
rect 675536 955680 675542 955732
rect 42334 955544 42340 955596
rect 42392 955584 42398 955596
rect 42702 955584 42708 955596
rect 42392 955556 42708 955584
rect 42392 955544 42398 955556
rect 42702 955544 42708 955556
rect 42760 955544 42766 955596
rect 674834 955476 674840 955528
rect 674892 955516 674898 955528
rect 675478 955516 675484 955528
rect 674892 955488 675484 955516
rect 674892 955476 674898 955488
rect 675478 955476 675484 955488
rect 675536 955476 675542 955528
rect 42242 954252 42248 954304
rect 42300 954292 42306 954304
rect 42702 954292 42708 954304
rect 42300 954264 42708 954292
rect 42300 954252 42306 954264
rect 42702 954252 42708 954264
rect 42760 954252 42766 954304
rect 36538 952212 36544 952264
rect 36596 952252 36602 952264
rect 42334 952252 42340 952264
rect 36596 952224 42340 952252
rect 36596 952212 36602 952224
rect 42334 952212 42340 952224
rect 42392 952212 42398 952264
rect 675754 952008 675760 952060
rect 675812 952008 675818 952060
rect 675772 951788 675800 952008
rect 675754 951736 675760 951788
rect 675812 951736 675818 951788
rect 31018 951464 31024 951516
rect 31076 951504 31082 951516
rect 41874 951504 41880 951516
rect 31076 951476 41880 951504
rect 31076 951464 31082 951476
rect 41874 951464 41880 951476
rect 41932 951464 41938 951516
rect 675754 949424 675760 949476
rect 675812 949464 675818 949476
rect 678238 949464 678244 949476
rect 675812 949436 678244 949464
rect 675812 949424 675818 949436
rect 678238 949424 678244 949436
rect 678296 949424 678302 949476
rect 651558 948064 651564 948116
rect 651616 948104 651622 948116
rect 674190 948104 674196 948116
rect 651616 948076 674196 948104
rect 651616 948064 651622 948076
rect 674190 948064 674196 948076
rect 674248 948064 674254 948116
rect 34514 945956 34520 946008
rect 34572 945996 34578 946008
rect 62114 945996 62120 946008
rect 34572 945968 62120 945996
rect 34572 945956 34578 945968
rect 62114 945956 62120 945968
rect 62172 945956 62178 946008
rect 35802 943236 35808 943288
rect 35860 943276 35866 943288
rect 48406 943276 48412 943288
rect 35860 943248 48412 943276
rect 35860 943236 35866 943248
rect 48406 943236 48412 943248
rect 48464 943236 48470 943288
rect 35710 943168 35716 943220
rect 35768 943208 35774 943220
rect 47670 943208 47676 943220
rect 35768 943180 47676 943208
rect 35768 943168 35774 943180
rect 47670 943168 47676 943180
rect 47728 943168 47734 943220
rect 41782 941808 41788 941860
rect 41840 941848 41846 941860
rect 42058 941848 42064 941860
rect 41840 941820 42064 941848
rect 41840 941808 41846 941820
rect 42058 941808 42064 941820
rect 42116 941808 42122 941860
rect 652018 939768 652024 939820
rect 652076 939808 652082 939820
rect 676030 939808 676036 939820
rect 652076 939780 676036 939808
rect 652076 939768 652082 939780
rect 676030 939768 676036 939780
rect 676088 939768 676094 939820
rect 674190 939156 674196 939208
rect 674248 939196 674254 939208
rect 676030 939196 676036 939208
rect 674248 939168 676036 939196
rect 674248 939156 674254 939168
rect 676030 939156 676036 939168
rect 676088 939156 676094 939208
rect 671338 938680 671344 938732
rect 671396 938720 671402 938732
rect 676214 938720 676220 938732
rect 671396 938692 676220 938720
rect 671396 938680 671402 938692
rect 676214 938680 676220 938692
rect 676272 938680 676278 938732
rect 669958 938544 669964 938596
rect 670016 938584 670022 938596
rect 676030 938584 676036 938596
rect 670016 938556 676036 938584
rect 670016 938544 670022 938556
rect 676030 938544 676036 938556
rect 676088 938544 676094 938596
rect 661678 937320 661684 937372
rect 661736 937360 661742 937372
rect 676214 937360 676220 937372
rect 661736 937332 676220 937360
rect 661736 937320 661742 937332
rect 676214 937320 676220 937332
rect 676272 937320 676278 937372
rect 658918 937184 658924 937236
rect 658976 937224 658982 937236
rect 676214 937224 676220 937236
rect 658976 937196 676220 937224
rect 658976 937184 658982 937196
rect 676214 937184 676220 937196
rect 676272 937184 676278 937236
rect 672626 937116 672632 937168
rect 672684 937156 672690 937168
rect 676122 937156 676128 937168
rect 672684 937128 676128 937156
rect 672684 937116 672690 937128
rect 676122 937116 676128 937128
rect 676180 937116 676186 937168
rect 673178 937048 673184 937100
rect 673236 937088 673242 937100
rect 676030 937088 676036 937100
rect 673236 937060 676036 937088
rect 673236 937048 673242 937060
rect 676030 937048 676036 937060
rect 676088 937048 676094 937100
rect 48406 936980 48412 937032
rect 48464 937020 48470 937032
rect 62114 937020 62120 937032
rect 48464 936992 62120 937020
rect 48464 936980 48470 936992
rect 62114 936980 62120 936992
rect 62172 936980 62178 937032
rect 651558 936980 651564 937032
rect 651616 937020 651622 937032
rect 659010 937020 659016 937032
rect 651616 936992 659016 937020
rect 651616 936980 651622 936992
rect 659010 936980 659016 936992
rect 659068 936980 659074 937032
rect 673638 936640 673644 936692
rect 673696 936680 673702 936692
rect 676030 936680 676036 936692
rect 673696 936652 676036 936680
rect 673696 936640 673702 936652
rect 676030 936640 676036 936652
rect 676088 936640 676094 936692
rect 674650 935824 674656 935876
rect 674708 935864 674714 935876
rect 676030 935864 676036 935876
rect 674708 935836 676036 935864
rect 674708 935824 674714 935836
rect 676030 935824 676036 935836
rect 676088 935824 676094 935876
rect 660298 935620 660304 935672
rect 660356 935660 660362 935672
rect 676214 935660 676220 935672
rect 660356 935632 676220 935660
rect 660356 935620 660362 935632
rect 676214 935620 676220 935632
rect 676272 935620 676278 935672
rect 39942 932084 39948 932136
rect 40000 932124 40006 932136
rect 41874 932124 41880 932136
rect 40000 932096 41880 932124
rect 40000 932084 40006 932096
rect 41874 932084 41880 932096
rect 41932 932084 41938 932136
rect 674558 931948 674564 932000
rect 674616 931988 674622 932000
rect 676214 931988 676220 932000
rect 674616 931960 676220 931988
rect 674616 931948 674622 931960
rect 676214 931948 676220 931960
rect 676272 931948 676278 932000
rect 673270 930248 673276 930300
rect 673328 930288 673334 930300
rect 676214 930288 676220 930300
rect 673328 930260 676220 930288
rect 673328 930248 673334 930260
rect 676214 930248 676220 930260
rect 676272 930248 676278 930300
rect 669958 927392 669964 927444
rect 670016 927432 670022 927444
rect 683114 927432 683120 927444
rect 670016 927404 683120 927432
rect 670016 927392 670022 927404
rect 683114 927392 683120 927404
rect 683172 927392 683178 927444
rect 51718 923244 51724 923296
rect 51776 923284 51782 923296
rect 62114 923284 62120 923296
rect 51776 923256 62120 923284
rect 51776 923244 51782 923256
rect 62114 923244 62120 923256
rect 62172 923244 62178 923296
rect 651558 921816 651564 921868
rect 651616 921856 651622 921868
rect 664438 921856 664444 921868
rect 651616 921828 664444 921856
rect 651616 921816 651622 921828
rect 664438 921816 664444 921828
rect 664496 921816 664502 921868
rect 40678 909440 40684 909492
rect 40736 909480 40742 909492
rect 62114 909480 62120 909492
rect 40736 909452 62120 909480
rect 40736 909440 40742 909452
rect 62114 909440 62120 909452
rect 62172 909440 62178 909492
rect 651558 909440 651564 909492
rect 651616 909480 651622 909492
rect 661678 909480 661684 909492
rect 651616 909452 661684 909480
rect 651616 909440 651622 909452
rect 661678 909440 661684 909452
rect 661736 909440 661742 909492
rect 53098 896996 53104 897048
rect 53156 897036 53162 897048
rect 62114 897036 62120 897048
rect 53156 897008 62120 897036
rect 53156 896996 53162 897008
rect 62114 896996 62120 897008
rect 62172 896996 62178 897048
rect 651558 895636 651564 895688
rect 651616 895676 651622 895688
rect 660298 895676 660304 895688
rect 651616 895648 660304 895676
rect 651616 895636 651622 895648
rect 660298 895636 660304 895648
rect 660356 895636 660362 895688
rect 44818 884620 44824 884672
rect 44876 884660 44882 884672
rect 62114 884660 62120 884672
rect 44876 884632 62120 884660
rect 44876 884620 44882 884632
rect 62114 884620 62120 884632
rect 62172 884620 62178 884672
rect 671982 879044 671988 879096
rect 672040 879084 672046 879096
rect 675294 879084 675300 879096
rect 672040 879056 675300 879084
rect 672040 879044 672046 879056
rect 675294 879044 675300 879056
rect 675352 879044 675358 879096
rect 673086 873536 673092 873588
rect 673144 873576 673150 873588
rect 675386 873576 675392 873588
rect 673144 873548 675392 873576
rect 673144 873536 673150 873548
rect 675386 873536 675392 873548
rect 675444 873536 675450 873588
rect 55950 870816 55956 870868
rect 56008 870856 56014 870868
rect 62114 870856 62120 870868
rect 56008 870828 62120 870856
rect 56008 870816 56014 870828
rect 62114 870816 62120 870828
rect 62172 870816 62178 870868
rect 674374 869796 674380 869848
rect 674432 869836 674438 869848
rect 675386 869836 675392 869848
rect 674432 869808 675392 869836
rect 674432 869796 674438 869808
rect 675386 869796 675392 869808
rect 675444 869796 675450 869848
rect 672994 869592 673000 869644
rect 673052 869632 673058 869644
rect 675386 869632 675392 869644
rect 673052 869604 675392 869632
rect 673052 869592 673058 869604
rect 675386 869592 675392 869604
rect 675444 869592 675450 869644
rect 651558 869388 651564 869440
rect 651616 869428 651622 869440
rect 671338 869428 671344 869440
rect 651616 869400 671344 869428
rect 651616 869388 651622 869400
rect 671338 869388 671344 869400
rect 671396 869388 671402 869440
rect 672902 868980 672908 869032
rect 672960 869020 672966 869032
rect 675386 869020 675392 869032
rect 672960 868992 675392 869020
rect 672960 868980 672966 868992
rect 675386 868980 675392 868992
rect 675444 868980 675450 869032
rect 652018 868640 652024 868692
rect 652076 868680 652082 868692
rect 674926 868680 674932 868692
rect 652076 868652 674932 868680
rect 652076 868640 652082 868652
rect 674926 868640 674932 868652
rect 674984 868640 674990 868692
rect 674558 868028 674564 868080
rect 674616 868068 674622 868080
rect 675386 868068 675392 868080
rect 674616 868040 675392 868068
rect 674616 868028 674622 868040
rect 675386 868028 675392 868040
rect 675444 868028 675450 868080
rect 674466 866804 674472 866856
rect 674524 866844 674530 866856
rect 675386 866844 675392 866856
rect 674524 866816 675392 866844
rect 674524 866804 674530 866816
rect 675386 866804 675392 866816
rect 675444 866804 675450 866856
rect 674926 866192 674932 866244
rect 674984 866232 674990 866244
rect 675386 866232 675392 866244
rect 674984 866204 675392 866232
rect 674984 866192 674990 866204
rect 675386 866192 675392 866204
rect 675444 866192 675450 866244
rect 672810 862792 672816 862844
rect 672868 862832 672874 862844
rect 675478 862832 675484 862844
rect 672868 862804 675484 862832
rect 672868 862792 672874 862804
rect 675478 862792 675484 862804
rect 675536 862792 675542 862844
rect 43622 858372 43628 858424
rect 43680 858412 43686 858424
rect 62114 858412 62120 858424
rect 43680 858384 62120 858412
rect 43680 858372 43686 858384
rect 62114 858372 62120 858384
rect 62172 858372 62178 858424
rect 652570 855584 652576 855636
rect 652628 855624 652634 855636
rect 672718 855624 672724 855636
rect 652628 855596 672724 855624
rect 652628 855584 652634 855596
rect 672718 855584 672724 855596
rect 672776 855584 672782 855636
rect 54478 844568 54484 844620
rect 54536 844608 54542 844620
rect 62114 844608 62120 844620
rect 54536 844580 62120 844608
rect 54536 844568 54542 844580
rect 62114 844568 62120 844580
rect 62172 844568 62178 844620
rect 651558 841780 651564 841832
rect 651616 841820 651622 841832
rect 663058 841820 663064 841832
rect 651616 841792 663064 841820
rect 651616 841780 651622 841792
rect 663058 841780 663064 841792
rect 663116 841780 663122 841832
rect 50430 832124 50436 832176
rect 50488 832164 50494 832176
rect 62114 832164 62120 832176
rect 50488 832136 62120 832164
rect 50488 832124 50494 832136
rect 62114 832124 62120 832136
rect 62172 832124 62178 832176
rect 651558 829404 651564 829456
rect 651616 829444 651622 829456
rect 659010 829444 659016 829456
rect 651616 829416 659016 829444
rect 651616 829404 651622 829416
rect 659010 829404 659016 829416
rect 659068 829404 659074 829456
rect 47578 818320 47584 818372
rect 47636 818360 47642 818372
rect 62114 818360 62120 818372
rect 47636 818332 62120 818360
rect 47636 818320 47642 818332
rect 62114 818320 62120 818332
rect 62172 818320 62178 818372
rect 41322 817504 41328 817556
rect 41380 817544 41386 817556
rect 44818 817544 44824 817556
rect 41380 817516 44824 817544
rect 41380 817504 41386 817516
rect 44818 817504 44824 817516
rect 44876 817504 44882 817556
rect 41230 817368 41236 817420
rect 41288 817408 41294 817420
rect 53098 817408 53104 817420
rect 41288 817380 53104 817408
rect 41288 817368 41294 817380
rect 53098 817368 53104 817380
rect 53156 817368 53162 817420
rect 651558 815600 651564 815652
rect 651616 815640 651622 815652
rect 665818 815640 665824 815652
rect 651616 815612 665824 815640
rect 651616 815600 651622 815612
rect 665818 815600 665824 815612
rect 665876 815600 665882 815652
rect 41506 814852 41512 814904
rect 41564 814892 41570 814904
rect 41782 814892 41788 814904
rect 41564 814864 41788 814892
rect 41564 814852 41570 814864
rect 41782 814852 41788 814864
rect 41840 814852 41846 814904
rect 35802 806420 35808 806472
rect 35860 806460 35866 806472
rect 41874 806460 41880 806472
rect 35860 806432 41880 806460
rect 35860 806420 35866 806432
rect 41874 806420 41880 806432
rect 41932 806420 41938 806472
rect 50338 805944 50344 805996
rect 50396 805984 50402 805996
rect 62114 805984 62120 805996
rect 50396 805956 62120 805984
rect 50396 805944 50402 805956
rect 62114 805944 62120 805956
rect 62172 805944 62178 805996
rect 42150 803836 42156 803888
rect 42208 803876 42214 803888
rect 42610 803876 42616 803888
rect 42208 803848 42616 803876
rect 42208 803836 42214 803848
rect 42610 803836 42616 803848
rect 42668 803836 42674 803888
rect 42058 803768 42064 803820
rect 42116 803808 42122 803820
rect 42702 803808 42708 803820
rect 42116 803780 42708 803808
rect 42116 803768 42122 803780
rect 42702 803768 42708 803780
rect 42760 803768 42766 803820
rect 651558 803156 651564 803208
rect 651616 803196 651622 803208
rect 658918 803196 658924 803208
rect 651616 803168 658924 803196
rect 651616 803156 651622 803168
rect 658918 803156 658924 803168
rect 658976 803156 658982 803208
rect 35250 801116 35256 801168
rect 35308 801156 35314 801168
rect 43070 801156 43076 801168
rect 35308 801128 43076 801156
rect 35308 801116 35314 801128
rect 43070 801116 43076 801128
rect 43128 801116 43134 801168
rect 32398 801048 32404 801100
rect 32456 801088 32462 801100
rect 42886 801088 42892 801100
rect 32456 801060 42892 801088
rect 32456 801048 32462 801060
rect 42886 801048 42892 801060
rect 42944 801048 42950 801100
rect 40678 800504 40684 800556
rect 40736 800544 40742 800556
rect 42978 800544 42984 800556
rect 40736 800516 42984 800544
rect 40736 800504 40742 800516
rect 42978 800504 42984 800516
rect 43036 800504 43042 800556
rect 42150 799960 42156 800012
rect 42208 800000 42214 800012
rect 42334 800000 42340 800012
rect 42208 799972 42340 800000
rect 42208 799960 42214 799972
rect 42334 799960 42340 799972
rect 42392 799960 42398 800012
rect 51718 799728 51724 799740
rect 42720 799700 51724 799728
rect 42720 799128 42748 799700
rect 51718 799688 51724 799700
rect 51776 799688 51782 799740
rect 42702 799076 42708 799128
rect 42760 799076 42766 799128
rect 42150 798124 42156 798176
rect 42208 798164 42214 798176
rect 42610 798164 42616 798176
rect 42208 798136 42616 798164
rect 42208 798124 42214 798136
rect 42610 798124 42616 798136
rect 42668 798124 42674 798176
rect 42150 797240 42156 797292
rect 42208 797280 42214 797292
rect 42702 797280 42708 797292
rect 42208 797252 42708 797280
rect 42208 797240 42214 797252
rect 42702 797240 42708 797252
rect 42760 797240 42766 797292
rect 42150 796288 42156 796340
rect 42208 796328 42214 796340
rect 42702 796328 42708 796340
rect 42208 796300 42708 796328
rect 42208 796288 42214 796300
rect 42702 796288 42708 796300
rect 42760 796288 42766 796340
rect 42150 794996 42156 795048
rect 42208 795036 42214 795048
rect 42426 795036 42432 795048
rect 42208 795008 42432 795036
rect 42208 794996 42214 795008
rect 42426 794996 42432 795008
rect 42484 794996 42490 795048
rect 42426 794860 42432 794912
rect 42484 794900 42490 794912
rect 42978 794900 42984 794912
rect 42484 794872 42984 794900
rect 42484 794860 42490 794872
rect 42978 794860 42984 794872
rect 43036 794860 43042 794912
rect 43162 794860 43168 794912
rect 43220 794900 43226 794912
rect 44450 794900 44456 794912
rect 43220 794872 44456 794900
rect 43220 794860 43226 794872
rect 44450 794860 44456 794872
rect 44508 794860 44514 794912
rect 42150 794248 42156 794300
rect 42208 794288 42214 794300
rect 42702 794288 42708 794300
rect 42208 794260 42708 794288
rect 42208 794248 42214 794260
rect 42702 794248 42708 794260
rect 42760 794248 42766 794300
rect 42150 793772 42156 793824
rect 42208 793812 42214 793824
rect 43162 793812 43168 793824
rect 42208 793784 43168 793812
rect 42208 793772 42214 793784
rect 43162 793772 43168 793784
rect 43220 793772 43226 793824
rect 44818 793500 44824 793552
rect 44876 793540 44882 793552
rect 62114 793540 62120 793552
rect 44876 793512 62120 793540
rect 44876 793500 44882 793512
rect 62114 793500 62120 793512
rect 62172 793500 62178 793552
rect 42150 793160 42156 793212
rect 42208 793200 42214 793212
rect 42426 793200 42432 793212
rect 42208 793172 42432 793200
rect 42208 793160 42214 793172
rect 42426 793160 42432 793172
rect 42484 793160 42490 793212
rect 42426 793024 42432 793076
rect 42484 793064 42490 793076
rect 44358 793064 44364 793076
rect 42484 793036 44364 793064
rect 42484 793024 42490 793036
rect 44358 793024 44364 793036
rect 44416 793024 44422 793076
rect 42150 790644 42156 790696
rect 42208 790684 42214 790696
rect 42702 790684 42708 790696
rect 42208 790656 42708 790684
rect 42208 790644 42214 790656
rect 42702 790644 42708 790656
rect 42760 790644 42766 790696
rect 42150 790100 42156 790152
rect 42208 790140 42214 790152
rect 42426 790140 42432 790152
rect 42208 790112 42432 790140
rect 42208 790100 42214 790112
rect 42426 790100 42432 790112
rect 42484 790100 42490 790152
rect 42150 789420 42156 789472
rect 42208 789460 42214 789472
rect 42334 789460 42340 789472
rect 42208 789432 42340 789460
rect 42208 789420 42214 789432
rect 42334 789420 42340 789432
rect 42392 789420 42398 789472
rect 651650 789352 651656 789404
rect 651708 789392 651714 789404
rect 661770 789392 661776 789404
rect 651708 789364 661776 789392
rect 651708 789352 651714 789364
rect 661770 789352 661776 789364
rect 661828 789352 661834 789404
rect 674282 787312 674288 787364
rect 674340 787352 674346 787364
rect 675386 787352 675392 787364
rect 674340 787324 675392 787352
rect 674340 787312 674346 787324
rect 675386 787312 675392 787324
rect 675444 787312 675450 787364
rect 42058 786428 42064 786480
rect 42116 786468 42122 786480
rect 42426 786468 42432 786480
rect 42116 786440 42432 786468
rect 42116 786428 42122 786440
rect 42426 786428 42432 786440
rect 42484 786428 42490 786480
rect 42150 785612 42156 785664
rect 42208 785652 42214 785664
rect 42702 785652 42708 785664
rect 42208 785624 42708 785652
rect 42208 785612 42214 785624
rect 42702 785612 42708 785624
rect 42760 785612 42766 785664
rect 674190 784252 674196 784304
rect 674248 784292 674254 784304
rect 675386 784292 675392 784304
rect 674248 784264 675392 784292
rect 674248 784252 674254 784264
rect 675386 784252 675392 784264
rect 675444 784252 675450 784304
rect 674006 782892 674012 782944
rect 674064 782932 674070 782944
rect 675478 782932 675484 782944
rect 674064 782904 675484 782932
rect 674064 782892 674070 782904
rect 675478 782892 675484 782904
rect 675536 782892 675542 782944
rect 671890 780716 671896 780768
rect 671948 780756 671954 780768
rect 675478 780756 675484 780768
rect 671948 780728 675484 780756
rect 671948 780716 671954 780728
rect 675478 780716 675484 780728
rect 675536 780716 675542 780768
rect 673270 779968 673276 780020
rect 673328 780008 673334 780020
rect 675478 780008 675484 780020
rect 673328 779980 675484 780008
rect 673328 779968 673334 779980
rect 675478 779968 675484 779980
rect 675536 779968 675542 780020
rect 51718 779696 51724 779748
rect 51776 779736 51782 779748
rect 62114 779736 62120 779748
rect 51776 779708 62120 779736
rect 51776 779696 51782 779708
rect 62114 779696 62120 779708
rect 62172 779696 62178 779748
rect 672534 779288 672540 779340
rect 672592 779328 672598 779340
rect 675386 779328 675392 779340
rect 672592 779300 675392 779328
rect 672592 779288 672598 779300
rect 675386 779288 675392 779300
rect 675444 779288 675450 779340
rect 659010 778948 659016 779000
rect 659068 778988 659074 779000
rect 674742 778988 674748 779000
rect 659068 778960 674748 778988
rect 659068 778948 659074 778960
rect 674742 778948 674748 778960
rect 674800 778948 674806 779000
rect 673730 778608 673736 778660
rect 673788 778648 673794 778660
rect 675478 778648 675484 778660
rect 673788 778620 675484 778648
rect 673788 778608 673794 778620
rect 675478 778608 675484 778620
rect 675536 778608 675542 778660
rect 673914 777316 673920 777368
rect 673972 777356 673978 777368
rect 675386 777356 675392 777368
rect 673972 777328 675392 777356
rect 673972 777316 673978 777328
rect 675386 777316 675392 777328
rect 675444 777316 675450 777368
rect 674742 777044 674748 777096
rect 674800 777084 674806 777096
rect 675386 777084 675392 777096
rect 674800 777056 675392 777084
rect 674800 777044 674806 777056
rect 675386 777044 675392 777056
rect 675444 777044 675450 777096
rect 651558 775548 651564 775600
rect 651616 775588 651622 775600
rect 659010 775588 659016 775600
rect 651616 775560 659016 775588
rect 651616 775548 651622 775560
rect 659010 775548 659016 775560
rect 659068 775548 659074 775600
rect 670510 775548 670516 775600
rect 670568 775588 670574 775600
rect 675386 775588 675392 775600
rect 670568 775560 675392 775588
rect 670568 775548 670574 775560
rect 675386 775548 675392 775560
rect 675444 775548 675450 775600
rect 35802 774188 35808 774240
rect 35860 774228 35866 774240
rect 54478 774228 54484 774240
rect 35860 774200 54484 774228
rect 35860 774188 35866 774200
rect 54478 774188 54484 774200
rect 54536 774188 54542 774240
rect 672442 773576 672448 773628
rect 672500 773616 672506 773628
rect 675478 773616 675484 773628
rect 672500 773588 675484 773616
rect 672500 773576 672506 773588
rect 675478 773576 675484 773588
rect 675536 773576 675542 773628
rect 48958 767320 48964 767372
rect 49016 767360 49022 767372
rect 62114 767360 62120 767372
rect 49016 767332 62120 767360
rect 49016 767320 49022 767332
rect 62114 767320 62120 767332
rect 62172 767320 62178 767372
rect 675202 766572 675208 766624
rect 675260 766612 675266 766624
rect 675662 766612 675668 766624
rect 675260 766584 675668 766612
rect 675260 766572 675266 766584
rect 675662 766572 675668 766584
rect 675720 766572 675726 766624
rect 651558 763172 651564 763224
rect 651616 763212 651622 763224
rect 664530 763212 664536 763224
rect 651616 763184 664536 763212
rect 651616 763172 651622 763184
rect 664530 763172 664536 763184
rect 664588 763172 664594 763224
rect 41506 761744 41512 761796
rect 41564 761784 41570 761796
rect 55858 761784 55864 761796
rect 41564 761756 55864 761784
rect 41564 761744 41570 761756
rect 55858 761744 55864 761756
rect 55916 761744 55922 761796
rect 664438 760792 664444 760844
rect 664496 760832 664502 760844
rect 676214 760832 676220 760844
rect 664496 760804 676220 760832
rect 664496 760792 664502 760804
rect 676214 760792 676220 760804
rect 676272 760792 676278 760844
rect 661678 760656 661684 760708
rect 661736 760696 661742 760708
rect 676122 760696 676128 760708
rect 661736 760668 676128 760696
rect 661736 760656 661742 760668
rect 676122 760656 676128 760668
rect 676180 760656 676186 760708
rect 660298 760520 660304 760572
rect 660356 760560 660362 760572
rect 676030 760560 676036 760572
rect 660356 760532 676036 760560
rect 660356 760520 660362 760532
rect 676030 760520 676036 760532
rect 676088 760520 676094 760572
rect 31018 759636 31024 759688
rect 31076 759676 31082 759688
rect 41874 759676 41880 759688
rect 31076 759648 41880 759676
rect 31076 759636 31082 759648
rect 41874 759636 41880 759648
rect 41932 759636 41938 759688
rect 672626 759296 672632 759348
rect 672684 759336 672690 759348
rect 676214 759336 676220 759348
rect 672684 759308 676220 759336
rect 672684 759296 672690 759308
rect 676214 759296 676220 759308
rect 676272 759296 676278 759348
rect 673178 759160 673184 759212
rect 673236 759200 673242 759212
rect 676214 759200 676220 759212
rect 673236 759172 676220 759200
rect 673236 759160 673242 759172
rect 676214 759160 676220 759172
rect 676272 759160 676278 759212
rect 673822 759024 673828 759076
rect 673880 759064 673886 759076
rect 676030 759064 676036 759076
rect 673880 759036 676036 759064
rect 673880 759024 673886 759036
rect 676030 759024 676036 759036
rect 676088 759024 676094 759076
rect 673638 758820 673644 758872
rect 673696 758860 673702 758872
rect 676214 758860 676220 758872
rect 673696 758832 676220 758860
rect 673696 758820 673702 758832
rect 676214 758820 676220 758832
rect 676272 758820 676278 758872
rect 33778 758480 33784 758532
rect 33836 758520 33842 758532
rect 41782 758520 41788 758532
rect 33836 758492 41788 758520
rect 33836 758480 33842 758492
rect 41782 758480 41788 758492
rect 41840 758480 41846 758532
rect 32490 758344 32496 758396
rect 32548 758384 32554 758396
rect 42702 758384 42708 758396
rect 32548 758356 42708 758384
rect 32548 758344 32554 758356
rect 42702 758344 42708 758356
rect 42760 758344 42766 758396
rect 32398 758276 32404 758328
rect 32456 758316 32462 758328
rect 42426 758316 42432 758328
rect 32456 758288 42432 758316
rect 32456 758276 32462 758288
rect 42426 758276 42432 758288
rect 42484 758276 42490 758328
rect 673546 758208 673552 758260
rect 673604 758248 673610 758260
rect 676030 758248 676036 758260
rect 673604 758220 676036 758248
rect 673604 758208 673610 758220
rect 676030 758208 676036 758220
rect 676088 758208 676094 758260
rect 41874 756984 41880 757036
rect 41932 756984 41938 757036
rect 41892 756764 41920 756984
rect 42426 756848 42432 756900
rect 42484 756888 42490 756900
rect 55950 756888 55956 756900
rect 42484 756860 55956 756888
rect 42484 756848 42490 756860
rect 55950 756848 55956 756860
rect 56008 756848 56014 756900
rect 41874 756712 41880 756764
rect 41932 756712 41938 756764
rect 42702 756508 42708 756560
rect 42760 756548 42766 756560
rect 42978 756548 42984 756560
rect 42760 756520 42984 756548
rect 42760 756508 42766 756520
rect 42978 756508 42984 756520
rect 43036 756508 43042 756560
rect 673362 756236 673368 756288
rect 673420 756276 673426 756288
rect 676214 756276 676220 756288
rect 673420 756248 676220 756276
rect 673420 756236 673426 756248
rect 676214 756236 676220 756248
rect 676272 756236 676278 756288
rect 674374 755556 674380 755608
rect 674432 755596 674438 755608
rect 676214 755596 676220 755608
rect 674432 755568 676220 755596
rect 674432 755556 674438 755568
rect 676214 755556 676220 755568
rect 676272 755556 676278 755608
rect 42426 755488 42432 755540
rect 42484 755528 42490 755540
rect 42484 755500 42748 755528
rect 42484 755488 42490 755500
rect 42610 755216 42616 755268
rect 42668 755256 42674 755268
rect 42720 755256 42748 755500
rect 42668 755228 42748 755256
rect 42668 755216 42674 755228
rect 672810 755080 672816 755132
rect 672868 755120 672874 755132
rect 676214 755120 676220 755132
rect 672868 755092 676220 755120
rect 672868 755080 672874 755092
rect 676214 755080 676220 755092
rect 676272 755080 676278 755132
rect 671982 754944 671988 754996
rect 672040 754984 672046 754996
rect 676122 754984 676128 754996
rect 672040 754956 676128 754984
rect 672040 754944 672046 754956
rect 676122 754944 676128 754956
rect 676180 754944 676186 754996
rect 42058 754264 42064 754316
rect 42116 754304 42122 754316
rect 42610 754304 42616 754316
rect 42116 754276 42616 754304
rect 42116 754264 42122 754276
rect 42610 754264 42616 754276
rect 42668 754264 42674 754316
rect 673086 753584 673092 753636
rect 673144 753624 673150 753636
rect 676214 753624 676220 753636
rect 673144 753596 676220 753624
rect 673144 753584 673150 753596
rect 676214 753584 676220 753596
rect 676272 753584 676278 753636
rect 43622 753516 43628 753568
rect 43680 753556 43686 753568
rect 62114 753556 62120 753568
rect 43680 753528 62120 753556
rect 43680 753516 43686 753528
rect 62114 753516 62120 753528
rect 62172 753516 62178 753568
rect 674466 753380 674472 753432
rect 674524 753420 674530 753432
rect 676030 753420 676036 753432
rect 674524 753392 676036 753420
rect 674524 753380 674530 753392
rect 676030 753380 676036 753392
rect 676088 753380 676094 753432
rect 672994 752360 673000 752412
rect 673052 752400 673058 752412
rect 676214 752400 676220 752412
rect 673052 752372 676220 752400
rect 673052 752360 673058 752372
rect 676214 752360 676220 752372
rect 676272 752360 676278 752412
rect 672902 752224 672908 752276
rect 672960 752264 672966 752276
rect 676122 752264 676128 752276
rect 672960 752236 676128 752264
rect 672960 752224 672966 752236
rect 676122 752224 676128 752236
rect 676180 752224 676186 752276
rect 674558 751884 674564 751936
rect 674616 751924 674622 751936
rect 676214 751924 676220 751936
rect 674616 751896 676220 751924
rect 674616 751884 674622 751896
rect 676214 751884 676220 751896
rect 676272 751884 676278 751936
rect 42150 751748 42156 751800
rect 42208 751788 42214 751800
rect 42610 751788 42616 751800
rect 42208 751760 42616 751788
rect 42208 751748 42214 751760
rect 42610 751748 42616 751760
rect 42668 751748 42674 751800
rect 42610 751612 42616 751664
rect 42668 751652 42674 751664
rect 42978 751652 42984 751664
rect 42668 751624 42984 751652
rect 42668 751612 42674 751624
rect 42978 751612 42984 751624
rect 43036 751612 43042 751664
rect 42150 751068 42156 751120
rect 42208 751108 42214 751120
rect 43254 751108 43260 751120
rect 42208 751080 43260 751108
rect 42208 751068 42214 751080
rect 43254 751068 43260 751080
rect 43312 751068 43318 751120
rect 42150 749776 42156 749828
rect 42208 749816 42214 749828
rect 43162 749816 43168 749828
rect 42208 749788 43168 749816
rect 42208 749776 42214 749788
rect 43162 749776 43168 749788
rect 43220 749776 43226 749828
rect 42978 749368 42984 749420
rect 43036 749408 43042 749420
rect 44450 749408 44456 749420
rect 43036 749380 44456 749408
rect 43036 749368 43042 749380
rect 44450 749368 44456 749380
rect 44508 749368 44514 749420
rect 651558 749368 651564 749420
rect 651616 749408 651622 749420
rect 668578 749408 668584 749420
rect 651616 749380 668584 749408
rect 651616 749368 651622 749380
rect 668578 749368 668584 749380
rect 668636 749368 668642 749420
rect 670050 749368 670056 749420
rect 670108 749408 670114 749420
rect 683114 749408 683120 749420
rect 670108 749380 683120 749408
rect 670108 749368 670114 749380
rect 683114 749368 683120 749380
rect 683172 749368 683178 749420
rect 43070 747940 43076 747992
rect 43128 747980 43134 747992
rect 44358 747980 44364 747992
rect 43128 747952 44364 747980
rect 43128 747940 43134 747952
rect 44358 747940 44364 747952
rect 44416 747940 44422 747992
rect 42978 747028 42984 747040
rect 42076 747000 42984 747028
rect 42076 746972 42104 747000
rect 42978 746988 42984 747000
rect 43036 746988 43042 747040
rect 42058 746920 42064 746972
rect 42116 746920 42122 746972
rect 42150 746920 42156 746972
rect 42208 746960 42214 746972
rect 42610 746960 42616 746972
rect 42208 746932 42616 746960
rect 42208 746920 42214 746932
rect 42610 746920 42616 746932
rect 42668 746920 42674 746972
rect 42150 746036 42156 746088
rect 42208 746076 42214 746088
rect 43070 746076 43076 746088
rect 42208 746048 43076 746076
rect 42208 746036 42214 746048
rect 43070 746036 43076 746048
rect 43128 746036 43134 746088
rect 42150 745628 42156 745680
rect 42208 745668 42214 745680
rect 42702 745668 42708 745680
rect 42208 745640 42708 745668
rect 42208 745628 42214 745640
rect 42702 745628 42708 745640
rect 42760 745628 42766 745680
rect 42702 745492 42708 745544
rect 42760 745532 42766 745544
rect 42886 745532 42892 745544
rect 42760 745504 42892 745532
rect 42760 745492 42766 745504
rect 42886 745492 42892 745504
rect 42944 745492 42950 745544
rect 670602 743792 670608 743844
rect 670660 743832 670666 743844
rect 670660 743804 675432 743832
rect 670660 743792 670666 743804
rect 675404 743776 675432 743804
rect 42150 743724 42156 743776
rect 42208 743764 42214 743776
rect 42702 743764 42708 743776
rect 42208 743736 42708 743764
rect 42208 743724 42214 743736
rect 42702 743724 42708 743736
rect 42760 743724 42766 743776
rect 675386 743724 675392 743776
rect 675444 743724 675450 743776
rect 42150 743248 42156 743300
rect 42208 743288 42214 743300
rect 42610 743288 42616 743300
rect 42208 743260 42616 743288
rect 42208 743248 42214 743260
rect 42610 743248 42616 743260
rect 42668 743248 42674 743300
rect 673178 742500 673184 742552
rect 673236 742540 673242 742552
rect 675386 742540 675392 742552
rect 673236 742512 675392 742540
rect 673236 742500 673242 742512
rect 675386 742500 675392 742512
rect 675444 742500 675450 742552
rect 54478 741072 54484 741124
rect 54536 741112 54542 741124
rect 62114 741112 62120 741124
rect 54536 741084 62120 741112
rect 54536 741072 54542 741084
rect 62114 741072 62120 741084
rect 62172 741072 62178 741124
rect 674834 739916 674840 739968
rect 674892 739956 674898 739968
rect 675386 739956 675392 739968
rect 674892 739928 675392 739956
rect 674892 739916 674898 739928
rect 675386 739916 675392 739928
rect 675444 739916 675450 739968
rect 672994 739100 673000 739152
rect 673052 739140 673058 739152
rect 675386 739140 675392 739152
rect 673052 739112 675392 739140
rect 673052 739100 673058 739112
rect 675386 739100 675392 739112
rect 675444 739100 675450 739152
rect 673086 738624 673092 738676
rect 673144 738664 673150 738676
rect 675386 738664 675392 738676
rect 673144 738636 675392 738664
rect 673144 738624 673150 738636
rect 675386 738624 675392 738636
rect 675444 738624 675450 738676
rect 673638 738216 673644 738268
rect 673696 738256 673702 738268
rect 675386 738256 675392 738268
rect 673696 738228 675392 738256
rect 673696 738216 673702 738228
rect 675386 738216 675392 738228
rect 675444 738216 675450 738268
rect 674374 735632 674380 735684
rect 674432 735672 674438 735684
rect 675386 735672 675392 735684
rect 674432 735644 675392 735672
rect 674432 735632 674438 735644
rect 675386 735632 675392 735644
rect 675444 735632 675450 735684
rect 651558 735564 651564 735616
rect 651616 735604 651622 735616
rect 660298 735604 660304 735616
rect 651616 735576 660304 735604
rect 651616 735564 651622 735576
rect 660298 735564 660304 735576
rect 660356 735564 660362 735616
rect 672902 734952 672908 735004
rect 672960 734992 672966 735004
rect 675386 734992 675392 735004
rect 672960 734964 675392 734992
rect 672960 734952 672966 734964
rect 675386 734952 675392 734964
rect 675444 734952 675450 735004
rect 659010 734816 659016 734868
rect 659068 734856 659074 734868
rect 674650 734856 674656 734868
rect 659068 734828 674656 734856
rect 659068 734816 659074 734828
rect 674650 734816 674656 734828
rect 674708 734816 674714 734868
rect 672626 733864 672632 733916
rect 672684 733904 672690 733916
rect 675386 733904 675392 733916
rect 672684 733876 675392 733904
rect 672684 733864 672690 733876
rect 675386 733864 675392 733876
rect 675444 733864 675450 733916
rect 674650 732028 674656 732080
rect 674708 732068 674714 732080
rect 675386 732068 675392 732080
rect 674708 732040 675392 732068
rect 674708 732028 674714 732040
rect 675386 732028 675392 732040
rect 675444 732028 675450 732080
rect 31386 731348 31392 731400
rect 31444 731388 31450 731400
rect 44542 731388 44548 731400
rect 31444 731360 44548 731388
rect 31444 731348 31450 731360
rect 44542 731348 44548 731360
rect 44600 731348 44606 731400
rect 31478 731212 31484 731264
rect 31536 731252 31542 731264
rect 44818 731252 44824 731264
rect 31536 731224 44824 731252
rect 31536 731212 31542 731224
rect 44818 731212 44824 731224
rect 44876 731212 44882 731264
rect 31570 731076 31576 731128
rect 31628 731116 31634 731128
rect 50338 731116 50344 731128
rect 31628 731088 50344 731116
rect 31628 731076 31634 731088
rect 50338 731076 50344 731088
rect 50396 731076 50402 731128
rect 31662 730940 31668 730992
rect 31720 730980 31726 730992
rect 51718 730980 51724 730992
rect 31720 730952 51724 730980
rect 31720 730940 31726 730952
rect 51718 730940 51724 730952
rect 51776 730940 51782 730992
rect 671798 730464 671804 730516
rect 671856 730504 671862 730516
rect 675386 730504 675392 730516
rect 671856 730476 675392 730504
rect 671856 730464 671862 730476
rect 675386 730464 675392 730476
rect 675444 730464 675450 730516
rect 674650 728628 674656 728680
rect 674708 728668 674714 728680
rect 675478 728668 675484 728680
rect 674708 728640 675484 728668
rect 674708 728628 674714 728640
rect 675478 728628 675484 728640
rect 675536 728628 675542 728680
rect 51718 727268 51724 727320
rect 51776 727308 51782 727320
rect 62114 727308 62120 727320
rect 51776 727280 62120 727308
rect 51776 727268 51782 727280
rect 62114 727268 62120 727280
rect 62172 727268 62178 727320
rect 652018 723120 652024 723172
rect 652076 723160 652082 723172
rect 668670 723160 668676 723172
rect 652076 723132 668676 723160
rect 652076 723120 652082 723132
rect 668670 723120 668676 723132
rect 668728 723120 668734 723172
rect 41506 719652 41512 719704
rect 41564 719692 41570 719704
rect 50338 719692 50344 719704
rect 41564 719664 50344 719692
rect 41564 719652 41570 719664
rect 50338 719652 50344 719664
rect 50396 719652 50402 719704
rect 35802 716864 35808 716916
rect 35860 716904 35866 716916
rect 42426 716904 42432 716916
rect 35860 716876 42432 716904
rect 35860 716864 35866 716876
rect 42426 716864 42432 716876
rect 42484 716864 42490 716916
rect 672718 716524 672724 716576
rect 672776 716564 672782 716576
rect 676030 716564 676036 716576
rect 672776 716536 676036 716564
rect 672776 716524 672782 716536
rect 676030 716524 676036 716536
rect 676088 716524 676094 716576
rect 40770 716184 40776 716236
rect 40828 716224 40834 716236
rect 41874 716224 41880 716236
rect 40828 716196 41880 716224
rect 40828 716184 40834 716196
rect 41874 716184 41880 716196
rect 41932 716184 41938 716236
rect 671338 716116 671344 716168
rect 671396 716156 671402 716168
rect 676030 716156 676036 716168
rect 671396 716128 676036 716156
rect 671396 716116 671402 716128
rect 676030 716116 676036 716128
rect 676088 716116 676094 716168
rect 35710 715504 35716 715556
rect 35768 715544 35774 715556
rect 42518 715544 42524 715556
rect 35768 715516 42524 715544
rect 35768 715504 35774 715516
rect 42518 715504 42524 715516
rect 42576 715504 42582 715556
rect 663058 714960 663064 715012
rect 663116 715000 663122 715012
rect 676030 715000 676036 715012
rect 663116 714972 676036 715000
rect 663116 714960 663122 714972
rect 676030 714960 676036 714972
rect 676088 714960 676094 715012
rect 50430 714824 50436 714876
rect 50488 714864 50494 714876
rect 62114 714864 62120 714876
rect 50488 714836 62120 714864
rect 50488 714824 50494 714836
rect 62114 714824 62120 714836
rect 62172 714824 62178 714876
rect 673822 714484 673828 714536
rect 673880 714524 673886 714536
rect 676030 714524 676036 714536
rect 673880 714496 676036 714524
rect 673880 714484 673886 714496
rect 676030 714484 676036 714496
rect 676088 714484 676094 714536
rect 40678 714212 40684 714264
rect 40736 714252 40742 714264
rect 42794 714252 42800 714264
rect 40736 714224 42800 714252
rect 40736 714212 40742 714224
rect 42794 714212 42800 714224
rect 42852 714212 42858 714264
rect 40862 714144 40868 714196
rect 40920 714184 40926 714196
rect 42886 714184 42892 714196
rect 40920 714156 42892 714184
rect 40920 714144 40926 714156
rect 42886 714144 42892 714156
rect 42944 714144 42950 714196
rect 673822 714008 673828 714060
rect 673880 714048 673886 714060
rect 676030 714048 676036 714060
rect 673880 714020 676036 714048
rect 673880 714008 673886 714020
rect 676030 714008 676036 714020
rect 676088 714008 676094 714060
rect 41874 713804 41880 713856
rect 41932 713804 41938 713856
rect 41892 713584 41920 713804
rect 673546 713668 673552 713720
rect 673604 713708 673610 713720
rect 676030 713708 676036 713720
rect 673604 713680 676036 713708
rect 673604 713668 673610 713680
rect 676030 713668 676036 713680
rect 676088 713668 676094 713720
rect 41874 713532 41880 713584
rect 41932 713532 41938 713584
rect 674558 713192 674564 713244
rect 674616 713232 674622 713244
rect 676030 713232 676036 713244
rect 674616 713204 676036 713232
rect 674616 713192 674622 713204
rect 676030 713192 676036 713204
rect 676088 713192 676094 713244
rect 673362 712852 673368 712904
rect 673420 712892 673426 712904
rect 676030 712892 676036 712904
rect 673420 712864 676036 712892
rect 673420 712852 673426 712864
rect 676030 712852 676036 712864
rect 676088 712852 676094 712904
rect 672166 712376 672172 712428
rect 672224 712416 672230 712428
rect 676030 712416 676036 712428
rect 672224 712388 676036 712416
rect 672224 712376 672230 712388
rect 676030 712376 676036 712388
rect 676088 712376 676094 712428
rect 43070 712104 43076 712156
rect 43128 712144 43134 712156
rect 47578 712144 47584 712156
rect 43128 712116 47584 712144
rect 43128 712104 43134 712116
rect 47578 712104 47584 712116
rect 47636 712104 47642 712156
rect 42150 711628 42156 711680
rect 42208 711668 42214 711680
rect 42794 711668 42800 711680
rect 42208 711640 42800 711668
rect 42208 711628 42214 711640
rect 42794 711628 42800 711640
rect 42852 711628 42858 711680
rect 670510 711628 670516 711680
rect 670568 711668 670574 711680
rect 676030 711668 676036 711680
rect 670568 711640 676036 711668
rect 670568 711628 670574 711640
rect 676030 711628 676036 711640
rect 676088 711628 676094 711680
rect 42518 710948 42524 711000
rect 42576 710988 42582 711000
rect 42794 710988 42800 711000
rect 42576 710960 42800 710988
rect 42576 710948 42582 710960
rect 42794 710948 42800 710960
rect 42852 710948 42858 711000
rect 42150 710880 42156 710932
rect 42208 710920 42214 710932
rect 43070 710920 43076 710932
rect 42208 710892 43076 710920
rect 42208 710880 42214 710892
rect 43070 710880 43076 710892
rect 43128 710880 43134 710932
rect 671890 710404 671896 710456
rect 671948 710444 671954 710456
rect 676030 710444 676036 710456
rect 671948 710416 676036 710444
rect 671948 710404 671954 710416
rect 676030 710404 676036 710416
rect 676088 710404 676094 710456
rect 672442 709996 672448 710048
rect 672500 710036 672506 710048
rect 676030 710036 676036 710048
rect 672500 710008 676036 710036
rect 672500 709996 672506 710008
rect 676030 709996 676036 710008
rect 676088 709996 676094 710048
rect 42150 709860 42156 709912
rect 42208 709900 42214 709912
rect 42886 709900 42892 709912
rect 42208 709872 42892 709900
rect 42208 709860 42214 709872
rect 42886 709860 42892 709872
rect 42944 709860 42950 709912
rect 674282 709588 674288 709640
rect 674340 709628 674346 709640
rect 676030 709628 676036 709640
rect 674340 709600 676036 709628
rect 674340 709588 674346 709600
rect 676030 709588 676036 709600
rect 676088 709588 676094 709640
rect 42886 709316 42892 709368
rect 42944 709356 42950 709368
rect 44174 709356 44180 709368
rect 42944 709328 44180 709356
rect 42944 709316 42950 709328
rect 44174 709316 44180 709328
rect 44232 709316 44238 709368
rect 651558 709316 651564 709368
rect 651616 709356 651622 709368
rect 671430 709356 671436 709368
rect 651616 709328 671436 709356
rect 651616 709316 651622 709328
rect 671430 709316 671436 709328
rect 671488 709316 671494 709368
rect 674190 709180 674196 709232
rect 674248 709220 674254 709232
rect 676030 709220 676036 709232
rect 674248 709192 676036 709220
rect 674248 709180 674254 709192
rect 676030 709180 676036 709192
rect 676088 709180 676094 709232
rect 676030 709044 676036 709096
rect 676088 709084 676094 709096
rect 676950 709084 676956 709096
rect 676088 709056 676956 709084
rect 676088 709044 676094 709056
rect 676950 709044 676956 709056
rect 677008 709044 677014 709096
rect 42150 708568 42156 708620
rect 42208 708608 42214 708620
rect 42518 708608 42524 708620
rect 42208 708580 42524 708608
rect 42208 708568 42214 708580
rect 42518 708568 42524 708580
rect 42576 708568 42582 708620
rect 673914 708364 673920 708416
rect 673972 708404 673978 708416
rect 676030 708404 676036 708416
rect 673972 708376 676036 708404
rect 673972 708364 673978 708376
rect 676030 708364 676036 708376
rect 676088 708364 676094 708416
rect 42150 708024 42156 708076
rect 42208 708064 42214 708076
rect 42978 708064 42984 708076
rect 42208 708036 42984 708064
rect 42208 708024 42214 708036
rect 42978 708024 42984 708036
rect 43036 708024 43042 708076
rect 672534 707956 672540 708008
rect 672592 707996 672598 708008
rect 676030 707996 676036 708008
rect 672592 707968 676036 707996
rect 672592 707956 672598 707968
rect 676030 707956 676036 707968
rect 676088 707956 676094 708008
rect 674006 707548 674012 707600
rect 674064 707588 674070 707600
rect 676030 707588 676036 707600
rect 674064 707560 676036 707588
rect 674064 707548 674070 707560
rect 676030 707548 676036 707560
rect 676088 707548 676094 707600
rect 42150 707208 42156 707260
rect 42208 707248 42214 707260
rect 42886 707248 42892 707260
rect 42208 707220 42892 707248
rect 42208 707208 42214 707220
rect 42886 707208 42892 707220
rect 42944 707208 42950 707260
rect 673730 706732 673736 706784
rect 673788 706772 673794 706784
rect 675938 706772 675944 706784
rect 673788 706744 675944 706772
rect 673788 706732 673794 706744
rect 675938 706732 675944 706744
rect 675996 706732 676002 706784
rect 673270 706664 673276 706716
rect 673328 706704 673334 706716
rect 676030 706704 676036 706716
rect 673328 706676 676036 706704
rect 673328 706664 673334 706676
rect 676030 706664 676036 706676
rect 676088 706664 676094 706716
rect 44450 706636 44456 706648
rect 42536 706608 44456 706636
rect 42426 706052 42432 706104
rect 42484 706092 42490 706104
rect 42536 706092 42564 706608
rect 44450 706596 44456 706608
rect 44508 706596 44514 706648
rect 42484 706064 42564 706092
rect 42484 706052 42490 706064
rect 42058 704216 42064 704268
rect 42116 704256 42122 704268
rect 42426 704256 42432 704268
rect 42116 704228 42432 704256
rect 42116 704216 42122 704228
rect 42426 704216 42432 704228
rect 42484 704216 42490 704268
rect 672718 703808 672724 703860
rect 672776 703848 672782 703860
rect 676030 703848 676036 703860
rect 672776 703820 676036 703848
rect 672776 703808 672782 703820
rect 676030 703808 676036 703820
rect 676088 703808 676094 703860
rect 42150 703672 42156 703724
rect 42208 703712 42214 703724
rect 42794 703712 42800 703724
rect 42208 703684 42800 703712
rect 42208 703672 42214 703684
rect 42794 703672 42800 703684
rect 42852 703672 42858 703724
rect 42794 701020 42800 701072
rect 42852 701060 42858 701072
rect 44358 701060 44364 701072
rect 42852 701032 44364 701060
rect 42852 701020 42858 701032
rect 44358 701020 44364 701032
rect 44416 701020 44422 701072
rect 42150 700408 42156 700460
rect 42208 700448 42214 700460
rect 42426 700448 42432 700460
rect 42208 700420 42432 700448
rect 42208 700408 42214 700420
rect 42426 700408 42432 700420
rect 42484 700408 42490 700460
rect 42150 699864 42156 699916
rect 42208 699904 42214 699916
rect 42702 699904 42708 699916
rect 42208 699876 42708 699904
rect 42208 699864 42214 699876
rect 42702 699864 42708 699876
rect 42760 699864 42766 699916
rect 671982 698164 671988 698216
rect 672040 698204 672046 698216
rect 675386 698204 675392 698216
rect 672040 698176 675392 698204
rect 672040 698164 672046 698176
rect 675386 698164 675392 698176
rect 675444 698164 675450 698216
rect 672258 697348 672264 697400
rect 672316 697388 672322 697400
rect 675386 697388 675392 697400
rect 672316 697360 675392 697388
rect 672316 697348 672322 697360
rect 675386 697348 675392 697360
rect 675444 697348 675450 697400
rect 30282 696192 30288 696244
rect 30340 696232 30346 696244
rect 43622 696232 43628 696244
rect 30340 696204 43628 696232
rect 30340 696192 30346 696204
rect 43622 696192 43628 696204
rect 43680 696192 43686 696244
rect 674466 694288 674472 694340
rect 674524 694328 674530 694340
rect 675478 694328 675484 694340
rect 674524 694300 675484 694328
rect 674524 694288 674530 694300
rect 675478 694288 675484 694300
rect 675536 694288 675542 694340
rect 673546 692996 673552 693048
rect 673604 693036 673610 693048
rect 675478 693036 675484 693048
rect 673604 693008 675484 693036
rect 673604 692996 673610 693008
rect 675478 692996 675484 693008
rect 675536 692996 675542 693048
rect 673362 690412 673368 690464
rect 673420 690452 673426 690464
rect 675386 690452 675392 690464
rect 673420 690424 675392 690452
rect 673420 690412 673426 690424
rect 675386 690412 675392 690424
rect 675444 690412 675450 690464
rect 674006 690004 674012 690056
rect 674064 690044 674070 690056
rect 675386 690044 675392 690056
rect 674064 690016 675392 690044
rect 674064 690004 674070 690016
rect 675386 690004 675392 690016
rect 675444 690004 675450 690056
rect 672810 689324 672816 689376
rect 672868 689364 672874 689376
rect 675478 689364 675484 689376
rect 672868 689336 675484 689364
rect 672868 689324 672874 689336
rect 675478 689324 675484 689336
rect 675536 689324 675542 689376
rect 674190 688712 674196 688764
rect 674248 688752 674254 688764
rect 675386 688752 675392 688764
rect 674248 688724 675392 688752
rect 674248 688712 674254 688724
rect 675386 688712 675392 688724
rect 675444 688712 675450 688764
rect 43714 688644 43720 688696
rect 43772 688684 43778 688696
rect 62114 688684 62120 688696
rect 43772 688656 62120 688684
rect 43772 688644 43778 688656
rect 62114 688644 62120 688656
rect 62172 688644 62178 688696
rect 668670 688644 668676 688696
rect 668728 688684 668734 688696
rect 674282 688684 674288 688696
rect 668728 688656 674288 688684
rect 668728 688644 668734 688656
rect 674282 688644 674288 688656
rect 674340 688644 674346 688696
rect 35802 687896 35808 687948
rect 35860 687936 35866 687948
rect 51718 687936 51724 687948
rect 35860 687908 51724 687936
rect 35860 687896 35866 687908
rect 51718 687896 51724 687908
rect 51776 687896 51782 687948
rect 35618 687760 35624 687812
rect 35676 687800 35682 687812
rect 54478 687800 54484 687812
rect 35676 687772 54484 687800
rect 35676 687760 35682 687772
rect 54478 687760 54484 687772
rect 54536 687760 54542 687812
rect 674282 687012 674288 687064
rect 674340 687052 674346 687064
rect 675478 687052 675484 687064
rect 674340 687024 675484 687052
rect 674340 687012 674346 687024
rect 675478 687012 675484 687024
rect 675536 687012 675542 687064
rect 673914 684224 673920 684276
rect 673972 684264 673978 684276
rect 675386 684264 675392 684276
rect 673972 684236 675392 684264
rect 673972 684224 673978 684236
rect 675386 684224 675392 684236
rect 675444 684224 675450 684276
rect 651834 683136 651840 683188
rect 651892 683176 651898 683188
rect 659010 683176 659016 683188
rect 651892 683148 659016 683176
rect 651892 683136 651898 683148
rect 659010 683136 659016 683148
rect 659068 683136 659074 683188
rect 40678 683000 40684 683052
rect 40736 683040 40742 683052
rect 41690 683040 41696 683052
rect 40736 683012 41696 683040
rect 40736 683000 40742 683012
rect 41690 683000 41696 683012
rect 41748 683000 41754 683052
rect 40770 681776 40776 681828
rect 40828 681816 40834 681828
rect 41690 681816 41696 681828
rect 40828 681788 41696 681816
rect 40828 681776 40834 681788
rect 41690 681776 41696 681788
rect 41748 681776 41754 681828
rect 30466 676812 30472 676864
rect 30524 676852 30530 676864
rect 51718 676852 51724 676864
rect 30524 676824 51724 676852
rect 30524 676812 30530 676824
rect 51718 676812 51724 676824
rect 51776 676812 51782 676864
rect 55950 674840 55956 674892
rect 56008 674880 56014 674892
rect 62114 674880 62120 674892
rect 56008 674852 62120 674880
rect 56008 674840 56014 674852
rect 62114 674840 62120 674852
rect 62172 674840 62178 674892
rect 35158 672800 35164 672852
rect 35216 672840 35222 672852
rect 42426 672840 42432 672852
rect 35216 672812 42432 672840
rect 35216 672800 35222 672812
rect 42426 672800 42432 672812
rect 42484 672800 42490 672852
rect 31018 672732 31024 672784
rect 31076 672772 31082 672784
rect 41874 672772 41880 672784
rect 31076 672744 41880 672772
rect 31076 672732 31082 672744
rect 41874 672732 41880 672744
rect 41932 672732 41938 672784
rect 40770 670964 40776 671016
rect 40828 671004 40834 671016
rect 42058 671004 42064 671016
rect 40828 670976 42064 671004
rect 40828 670964 40834 670976
rect 42058 670964 42064 670976
rect 42116 670964 42122 671016
rect 40678 670896 40684 670948
rect 40736 670936 40742 670948
rect 41782 670936 41788 670948
rect 40736 670908 41788 670936
rect 40736 670896 40742 670908
rect 41782 670896 41788 670908
rect 41840 670896 41846 670948
rect 665818 670896 665824 670948
rect 665876 670936 665882 670948
rect 676030 670936 676036 670948
rect 665876 670908 676036 670936
rect 665876 670896 665882 670908
rect 676030 670896 676036 670908
rect 676088 670896 676094 670948
rect 658918 670760 658924 670812
rect 658976 670800 658982 670812
rect 676214 670800 676220 670812
rect 658976 670772 676220 670800
rect 658976 670760 658982 670772
rect 676214 670760 676220 670772
rect 676272 670760 676278 670812
rect 41874 670556 41880 670608
rect 41932 670556 41938 670608
rect 41966 670556 41972 670608
rect 42024 670596 42030 670608
rect 42886 670596 42892 670608
rect 42024 670568 42892 670596
rect 42024 670556 42030 670568
rect 42886 670556 42892 670568
rect 42944 670556 42950 670608
rect 41892 670404 41920 670556
rect 41874 670352 41880 670404
rect 41932 670352 41938 670404
rect 42702 670012 42708 670064
rect 42760 670052 42766 670064
rect 48958 670052 48964 670064
rect 42760 670024 48964 670052
rect 42760 670012 42766 670024
rect 48958 670012 48964 670024
rect 49016 670012 49022 670064
rect 673822 669468 673828 669520
rect 673880 669508 673886 669520
rect 676030 669508 676036 669520
rect 673880 669480 676036 669508
rect 673880 669468 673886 669480
rect 676030 669468 676036 669480
rect 676088 669468 676094 669520
rect 661770 669400 661776 669452
rect 661828 669440 661834 669452
rect 676122 669440 676128 669452
rect 661828 669412 676128 669440
rect 661828 669400 661834 669412
rect 676122 669400 676128 669412
rect 676180 669400 676186 669452
rect 651558 669332 651564 669384
rect 651616 669372 651622 669384
rect 658918 669372 658924 669384
rect 651616 669344 658924 669372
rect 651616 669332 651622 669344
rect 658918 669332 658924 669344
rect 658976 669332 658982 669384
rect 672442 669332 672448 669384
rect 672500 669372 672506 669384
rect 676214 669372 676220 669384
rect 672500 669344 676220 669372
rect 672500 669332 672506 669344
rect 676214 669332 676220 669344
rect 676272 669332 676278 669384
rect 674558 668516 674564 668568
rect 674616 668556 674622 668568
rect 676030 668556 676036 668568
rect 674616 668528 676036 668556
rect 674616 668516 674622 668528
rect 676030 668516 676036 668528
rect 676088 668516 676094 668568
rect 672534 667904 672540 667956
rect 672592 667944 672598 667956
rect 676214 667944 676220 667956
rect 672592 667916 676220 667944
rect 672592 667904 672598 667916
rect 676214 667904 676220 667916
rect 676272 667904 676278 667956
rect 42150 667836 42156 667888
rect 42208 667876 42214 667888
rect 42702 667876 42708 667888
rect 42208 667848 42708 667876
rect 42208 667836 42214 667848
rect 42702 667836 42708 667848
rect 42760 667836 42766 667888
rect 42794 667768 42800 667820
rect 42852 667768 42858 667820
rect 42812 667616 42840 667768
rect 42794 667564 42800 667616
rect 42852 667564 42858 667616
rect 673822 667224 673828 667276
rect 673880 667264 673886 667276
rect 676030 667264 676036 667276
rect 673880 667236 676036 667264
rect 673880 667224 673886 667236
rect 676030 667224 676036 667236
rect 676088 667224 676094 667276
rect 42150 666680 42156 666732
rect 42208 666720 42214 666732
rect 44174 666720 44180 666732
rect 42208 666692 44180 666720
rect 42208 666680 42214 666692
rect 44174 666680 44180 666692
rect 44232 666680 44238 666732
rect 672166 666680 672172 666732
rect 672224 666720 672230 666732
rect 676214 666720 676220 666732
rect 672224 666692 676220 666720
rect 672224 666680 672230 666692
rect 676214 666680 676220 666692
rect 676272 666680 676278 666732
rect 671798 665456 671804 665508
rect 671856 665496 671862 665508
rect 676122 665496 676128 665508
rect 671856 665468 676128 665496
rect 671856 665456 671862 665468
rect 676122 665456 676128 665468
rect 676180 665456 676186 665508
rect 670602 665320 670608 665372
rect 670660 665360 670666 665372
rect 676214 665360 676220 665372
rect 670660 665332 676220 665360
rect 670660 665320 670666 665332
rect 676214 665320 676220 665332
rect 676272 665320 676278 665372
rect 674374 665252 674380 665304
rect 674432 665292 674438 665304
rect 676030 665292 676036 665304
rect 674432 665264 676036 665292
rect 674432 665252 674438 665264
rect 676030 665252 676036 665264
rect 676088 665252 676094 665304
rect 42886 665184 42892 665236
rect 42944 665224 42950 665236
rect 44450 665224 44456 665236
rect 42944 665196 44456 665224
rect 42944 665184 42950 665196
rect 44450 665184 44456 665196
rect 44508 665184 44514 665236
rect 674650 664980 674656 665032
rect 674708 665020 674714 665032
rect 676214 665020 676220 665032
rect 674708 664992 676220 665020
rect 674708 664980 674714 664992
rect 676214 664980 676220 664992
rect 676272 664980 676278 665032
rect 42150 663960 42156 664012
rect 42208 664000 42214 664012
rect 42886 664000 42892 664012
rect 42208 663972 42892 664000
rect 42208 663960 42214 663972
rect 42886 663960 42892 663972
rect 42944 663960 42950 664012
rect 673178 663960 673184 664012
rect 673236 664000 673242 664012
rect 676214 664000 676220 664012
rect 673236 663972 676220 664000
rect 673236 663960 673242 663972
rect 676214 663960 676220 663972
rect 676272 663960 676278 664012
rect 42702 663756 42708 663808
rect 42760 663796 42766 663808
rect 42886 663796 42892 663808
rect 42760 663768 42892 663796
rect 42760 663756 42766 663768
rect 42886 663756 42892 663768
rect 42944 663756 42950 663808
rect 672994 663756 673000 663808
rect 673052 663796 673058 663808
rect 676214 663796 676220 663808
rect 673052 663768 676220 663796
rect 673052 663756 673058 663768
rect 676214 663756 676220 663768
rect 676272 663756 676278 663808
rect 42794 662600 42800 662652
rect 42852 662640 42858 662652
rect 43070 662640 43076 662652
rect 42852 662612 43076 662640
rect 42852 662600 42858 662612
rect 43070 662600 43076 662612
rect 43128 662600 43134 662652
rect 42702 662396 42708 662448
rect 42760 662436 42766 662448
rect 42978 662436 42984 662448
rect 42760 662408 42984 662436
rect 42760 662396 42766 662408
rect 42978 662396 42984 662408
rect 43036 662396 43042 662448
rect 47578 662396 47584 662448
rect 47636 662436 47642 662448
rect 62114 662436 62120 662448
rect 47636 662408 62120 662436
rect 47636 662396 47642 662408
rect 62114 662396 62120 662408
rect 62172 662396 62178 662448
rect 673086 662396 673092 662448
rect 673144 662436 673150 662448
rect 676214 662436 676220 662448
rect 673144 662408 676220 662436
rect 673144 662396 673150 662408
rect 676214 662396 676220 662408
rect 676272 662396 676278 662448
rect 673638 662328 673644 662380
rect 673696 662368 673702 662380
rect 676030 662368 676036 662380
rect 673696 662340 676036 662368
rect 673696 662328 673702 662340
rect 676030 662328 676036 662340
rect 676088 662328 676094 662380
rect 672902 661240 672908 661292
rect 672960 661280 672966 661292
rect 676214 661280 676220 661292
rect 672960 661252 676220 661280
rect 672960 661240 672966 661252
rect 676214 661240 676220 661252
rect 676272 661240 676278 661292
rect 672626 661104 672632 661156
rect 672684 661144 672690 661156
rect 676122 661144 676128 661156
rect 672684 661116 676128 661144
rect 672684 661104 672690 661116
rect 676122 661104 676128 661116
rect 676180 661104 676186 661156
rect 42150 661036 42156 661088
rect 42208 661076 42214 661088
rect 42794 661076 42800 661088
rect 42208 661048 42800 661076
rect 42208 661036 42214 661048
rect 42794 661036 42800 661048
rect 42852 661036 42858 661088
rect 42150 659676 42156 659728
rect 42208 659716 42214 659728
rect 42886 659716 42892 659728
rect 42208 659688 42892 659716
rect 42208 659676 42214 659688
rect 42886 659676 42892 659688
rect 42944 659676 42950 659728
rect 674190 659676 674196 659728
rect 674248 659716 674254 659728
rect 683114 659716 683120 659728
rect 674248 659688 683120 659716
rect 674248 659676 674254 659688
rect 683114 659676 683120 659688
rect 683172 659676 683178 659728
rect 42150 658996 42156 659048
rect 42208 659036 42214 659048
rect 42702 659036 42708 659048
rect 42208 659008 42708 659036
rect 42208 658996 42214 659008
rect 42702 658996 42708 659008
rect 42760 658996 42766 659048
rect 42150 657228 42156 657280
rect 42208 657268 42214 657280
rect 42518 657268 42524 657280
rect 42208 657240 42524 657268
rect 42208 657228 42214 657240
rect 42518 657228 42524 657240
rect 42576 657228 42582 657280
rect 651558 656888 651564 656940
rect 651616 656928 651622 656940
rect 663058 656928 663064 656940
rect 651616 656900 663064 656928
rect 651616 656888 651622 656900
rect 663058 656888 663064 656900
rect 663116 656888 663122 656940
rect 42150 656820 42156 656872
rect 42208 656860 42214 656872
rect 43070 656860 43076 656872
rect 42208 656832 43076 656860
rect 42208 656820 42214 656832
rect 43070 656820 43076 656832
rect 43128 656820 43134 656872
rect 42150 656140 42156 656192
rect 42208 656180 42214 656192
rect 42334 656180 42340 656192
rect 42208 656152 42340 656180
rect 42208 656140 42214 656152
rect 42334 656140 42340 656152
rect 42392 656140 42398 656192
rect 675202 653760 675208 653812
rect 675260 653800 675266 653812
rect 675478 653800 675484 653812
rect 675260 653772 675484 653800
rect 675260 653760 675266 653772
rect 675478 653760 675484 653772
rect 675536 653760 675542 653812
rect 671890 652740 671896 652792
rect 671948 652780 671954 652792
rect 675386 652780 675392 652792
rect 671948 652752 675392 652780
rect 671948 652740 671954 652752
rect 675386 652740 675392 652752
rect 675444 652740 675450 652792
rect 674650 652128 674656 652180
rect 674708 652168 674714 652180
rect 675478 652168 675484 652180
rect 674708 652140 675484 652168
rect 674708 652128 674714 652140
rect 675478 652128 675484 652140
rect 675536 652128 675542 652180
rect 671798 651516 671804 651568
rect 671856 651556 671862 651568
rect 675386 651556 675392 651568
rect 671856 651528 675392 651556
rect 671856 651516 671862 651528
rect 675386 651516 675392 651528
rect 675444 651516 675450 651568
rect 674374 649068 674380 649120
rect 674432 649108 674438 649120
rect 675386 649108 675392 649120
rect 674432 649080 675392 649108
rect 674432 649068 674438 649080
rect 675386 649068 675392 649080
rect 675444 649068 675450 649120
rect 43622 647844 43628 647896
rect 43680 647884 43686 647896
rect 62114 647884 62120 647896
rect 43680 647856 62120 647884
rect 43680 647844 43686 647856
rect 62114 647844 62120 647856
rect 62172 647844 62178 647896
rect 673178 647708 673184 647760
rect 673236 647748 673242 647760
rect 675478 647748 675484 647760
rect 673236 647720 675484 647748
rect 673236 647708 673242 647720
rect 675478 647708 675484 647720
rect 675536 647708 675542 647760
rect 673730 645396 673736 645448
rect 673788 645436 673794 645448
rect 675386 645436 675392 645448
rect 673788 645408 675392 645436
rect 673788 645396 673794 645408
rect 675386 645396 675392 645408
rect 675444 645396 675450 645448
rect 672994 644988 673000 645040
rect 673052 645028 673058 645040
rect 675386 645028 675392 645040
rect 673052 645000 675392 645028
rect 673052 644988 673058 645000
rect 675386 644988 675392 645000
rect 675444 644988 675450 645040
rect 35618 644580 35624 644632
rect 35676 644620 35682 644632
rect 43714 644620 43720 644632
rect 35676 644592 43720 644620
rect 35676 644580 35682 644592
rect 43714 644580 43720 644592
rect 43772 644580 43778 644632
rect 35802 644512 35808 644564
rect 35860 644552 35866 644564
rect 55950 644552 55956 644564
rect 35860 644524 55956 644552
rect 35860 644512 35866 644524
rect 55950 644512 55956 644524
rect 56008 644512 56014 644564
rect 658918 643696 658924 643748
rect 658976 643736 658982 643748
rect 674558 643736 674564 643748
rect 658976 643708 674564 643736
rect 658976 643696 658982 643708
rect 674558 643696 674564 643708
rect 674616 643696 674622 643748
rect 673086 643356 673092 643408
rect 673144 643396 673150 643408
rect 675386 643396 675392 643408
rect 673144 643368 675392 643396
rect 673144 643356 673150 643368
rect 675386 643356 675392 643368
rect 675444 643356 675450 643408
rect 651558 643084 651564 643136
rect 651616 643124 651622 643136
rect 668670 643124 668676 643136
rect 651616 643096 668676 643124
rect 651616 643084 651622 643096
rect 668670 643084 668676 643096
rect 668728 643084 668734 643136
rect 674558 641860 674564 641912
rect 674616 641900 674622 641912
rect 675386 641900 675392 641912
rect 674616 641872 675392 641900
rect 674616 641860 674622 641872
rect 675386 641860 675392 641872
rect 675444 641860 675450 641912
rect 670510 640296 670516 640348
rect 670568 640336 670574 640348
rect 675386 640336 675392 640348
rect 670568 640308 675392 640336
rect 670568 640296 670574 640308
rect 675386 640296 675392 640308
rect 675444 640296 675450 640348
rect 673270 639072 673276 639124
rect 673328 639112 673334 639124
rect 675386 639112 675392 639124
rect 673328 639084 675392 639112
rect 673328 639072 673334 639084
rect 675386 639072 675392 639084
rect 675444 639072 675450 639124
rect 55950 636216 55956 636268
rect 56008 636256 56014 636268
rect 62114 636256 62120 636268
rect 56008 636228 62120 636256
rect 56008 636216 56014 636228
rect 62114 636216 62120 636228
rect 62172 636216 62178 636268
rect 675478 633768 675484 633820
rect 675536 633808 675542 633820
rect 681090 633808 681096 633820
rect 675536 633780 681096 633808
rect 675536 633768 675542 633780
rect 681090 633768 681096 633780
rect 681148 633768 681154 633820
rect 32398 629892 32404 629944
rect 32456 629932 32462 629944
rect 41782 629932 41788 629944
rect 32456 629904 41788 629932
rect 32456 629892 32462 629904
rect 41782 629892 41788 629904
rect 41840 629892 41846 629944
rect 651558 629280 651564 629332
rect 651616 629320 651622 629332
rect 661678 629320 661684 629332
rect 651616 629292 661684 629320
rect 651616 629280 651622 629292
rect 661678 629280 661684 629292
rect 661736 629280 661742 629332
rect 39298 629212 39304 629264
rect 39356 629252 39362 629264
rect 42518 629252 42524 629264
rect 39356 629224 42524 629252
rect 39356 629212 39362 629224
rect 42518 629212 42524 629224
rect 42576 629212 42582 629264
rect 41782 627376 41788 627428
rect 41840 627376 41846 627428
rect 41800 627088 41828 627376
rect 42886 627172 42892 627224
rect 42944 627212 42950 627224
rect 50430 627212 50436 627224
rect 42944 627184 50436 627212
rect 42944 627172 42950 627184
rect 50430 627172 50436 627184
rect 50488 627172 50494 627224
rect 41782 627036 41788 627088
rect 41840 627036 41846 627088
rect 668578 625472 668584 625524
rect 668636 625512 668642 625524
rect 676122 625512 676128 625524
rect 668636 625484 676128 625512
rect 668636 625472 668642 625484
rect 676122 625472 676128 625484
rect 676180 625472 676186 625524
rect 664530 625336 664536 625388
rect 664588 625376 664594 625388
rect 676214 625376 676220 625388
rect 664588 625348 676220 625376
rect 664588 625336 664594 625348
rect 676214 625336 676220 625348
rect 676272 625336 676278 625388
rect 42150 625268 42156 625320
rect 42208 625308 42214 625320
rect 42518 625308 42524 625320
rect 42208 625280 42524 625308
rect 42208 625268 42214 625280
rect 42518 625268 42524 625280
rect 42576 625268 42582 625320
rect 660298 625132 660304 625184
rect 660356 625172 660362 625184
rect 676214 625172 676220 625184
rect 660356 625144 676220 625172
rect 660356 625132 660362 625144
rect 676214 625132 676220 625144
rect 676272 625132 676278 625184
rect 42150 624656 42156 624708
rect 42208 624696 42214 624708
rect 42886 624696 42892 624708
rect 42208 624668 42892 624696
rect 42208 624656 42214 624668
rect 42886 624656 42892 624668
rect 42944 624656 42950 624708
rect 672442 624112 672448 624164
rect 672500 624152 672506 624164
rect 676214 624152 676220 624164
rect 672500 624124 676220 624152
rect 672500 624112 672506 624124
rect 676214 624112 676220 624124
rect 676272 624112 676278 624164
rect 672534 623908 672540 623960
rect 672592 623948 672598 623960
rect 676214 623948 676220 623960
rect 672592 623920 676220 623948
rect 672592 623908 672598 623920
rect 676214 623908 676220 623920
rect 676272 623908 676278 623960
rect 42518 623840 42524 623892
rect 42576 623840 42582 623892
rect 672442 623840 672448 623892
rect 672500 623880 672506 623892
rect 676122 623880 676128 623892
rect 672500 623852 676128 623880
rect 672500 623840 672506 623852
rect 676122 623840 676128 623852
rect 676180 623840 676186 623892
rect 42150 623432 42156 623484
rect 42208 623472 42214 623484
rect 42536 623472 42564 623840
rect 51810 623772 51816 623824
rect 51868 623812 51874 623824
rect 62114 623812 62120 623824
rect 51868 623784 62120 623812
rect 51868 623772 51874 623784
rect 62114 623772 62120 623784
rect 62172 623772 62178 623824
rect 672534 623772 672540 623824
rect 672592 623812 672598 623824
rect 676030 623812 676036 623824
rect 672592 623784 676036 623812
rect 672592 623772 672598 623784
rect 676030 623772 676036 623784
rect 676088 623772 676094 623824
rect 674742 623636 674748 623688
rect 674800 623676 674806 623688
rect 676214 623676 676220 623688
rect 674800 623648 676220 623676
rect 674800 623636 674806 623648
rect 676214 623636 676220 623648
rect 676272 623636 676278 623688
rect 42208 623444 42564 623472
rect 42208 623432 42214 623444
rect 673454 623024 673460 623076
rect 673512 623064 673518 623076
rect 676030 623064 676036 623076
rect 673512 623036 676036 623064
rect 673512 623024 673518 623036
rect 676030 623024 676036 623036
rect 676088 623024 676094 623076
rect 673822 622820 673828 622872
rect 673880 622860 673886 622872
rect 676214 622860 676220 622872
rect 673880 622832 676220 622860
rect 673880 622820 673886 622832
rect 676214 622820 676220 622832
rect 676272 622820 676278 622872
rect 44542 622452 44548 622464
rect 42628 622424 44548 622452
rect 42058 622140 42064 622192
rect 42116 622180 42122 622192
rect 42518 622180 42524 622192
rect 42116 622152 42524 622180
rect 42116 622140 42122 622152
rect 42518 622140 42524 622152
rect 42576 622140 42582 622192
rect 42518 622004 42524 622056
rect 42576 622044 42582 622056
rect 42628 622044 42656 622424
rect 44542 622412 44548 622424
rect 44600 622412 44606 622464
rect 673822 622208 673828 622260
rect 673880 622248 673886 622260
rect 676030 622248 676036 622260
rect 673880 622220 676036 622248
rect 673880 622208 673886 622220
rect 676030 622208 676036 622220
rect 676088 622208 676094 622260
rect 42576 622016 42656 622044
rect 42576 622004 42582 622016
rect 671982 621120 671988 621172
rect 672040 621160 672046 621172
rect 676214 621160 676220 621172
rect 672040 621132 676220 621160
rect 672040 621120 672046 621132
rect 676214 621120 676220 621132
rect 676272 621120 676278 621172
rect 42518 621052 42524 621104
rect 42576 621052 42582 621104
rect 42536 621024 42564 621052
rect 42076 620996 42564 621024
rect 42076 620832 42104 620996
rect 42518 620916 42524 620968
rect 42576 620956 42582 620968
rect 42794 620956 42800 620968
rect 42576 620928 42800 620956
rect 42576 620916 42582 620928
rect 42794 620916 42800 620928
rect 42852 620916 42858 620968
rect 42058 620780 42064 620832
rect 42116 620780 42122 620832
rect 42058 620304 42064 620356
rect 42116 620344 42122 620356
rect 42978 620344 42984 620356
rect 42116 620316 42984 620344
rect 42116 620304 42122 620316
rect 42978 620304 42984 620316
rect 43036 620304 43042 620356
rect 673914 619828 673920 619880
rect 673972 619868 673978 619880
rect 676030 619868 676036 619880
rect 673972 619840 676036 619868
rect 673972 619828 673978 619840
rect 676030 619828 676036 619840
rect 676088 619828 676094 619880
rect 673362 619760 673368 619812
rect 673420 619800 673426 619812
rect 676214 619800 676220 619812
rect 673420 619772 676220 619800
rect 673420 619760 673426 619772
rect 676214 619760 676220 619772
rect 676272 619760 676278 619812
rect 674466 619012 674472 619064
rect 674524 619052 674530 619064
rect 676030 619052 676036 619064
rect 674524 619024 676036 619052
rect 674524 619012 674530 619024
rect 676030 619012 676036 619024
rect 676088 619012 676094 619064
rect 672258 618400 672264 618452
rect 672316 618440 672322 618452
rect 676214 618440 676220 618452
rect 672316 618412 676220 618440
rect 672316 618400 672322 618412
rect 676214 618400 676220 618412
rect 676272 618400 676278 618452
rect 44450 618304 44456 618316
rect 42628 618276 44456 618304
rect 42150 617856 42156 617908
rect 42208 617896 42214 617908
rect 42518 617896 42524 617908
rect 42208 617868 42524 617896
rect 42208 617856 42214 617868
rect 42518 617856 42524 617868
rect 42576 617856 42582 617908
rect 42518 617720 42524 617772
rect 42576 617760 42582 617772
rect 42628 617760 42656 618276
rect 44450 618264 44456 618276
rect 44508 618264 44514 618316
rect 42576 617732 42656 617760
rect 42576 617720 42582 617732
rect 673546 617380 673552 617432
rect 673604 617420 673610 617432
rect 676030 617420 676036 617432
rect 673604 617392 676036 617420
rect 673604 617380 673610 617392
rect 676030 617380 676036 617392
rect 676088 617380 676094 617432
rect 42058 617108 42064 617160
rect 42116 617148 42122 617160
rect 42518 617148 42524 617160
rect 42116 617120 42524 617148
rect 42116 617108 42122 617120
rect 42518 617108 42524 617120
rect 42576 617108 42582 617160
rect 674006 616972 674012 617024
rect 674064 617012 674070 617024
rect 676030 617012 676036 617024
rect 674064 616984 676036 617012
rect 674064 616972 674070 616984
rect 676030 616972 676036 616984
rect 676088 616972 676094 617024
rect 652386 616836 652392 616888
rect 652444 616876 652450 616888
rect 658918 616876 658924 616888
rect 652444 616848 658924 616876
rect 652444 616836 652450 616848
rect 658918 616836 658924 616848
rect 658976 616836 658982 616888
rect 672810 616836 672816 616888
rect 672868 616876 672874 616888
rect 676214 616876 676220 616888
rect 672868 616848 676220 616876
rect 672868 616836 672874 616848
rect 676214 616836 676220 616848
rect 676272 616836 676278 616888
rect 674282 616700 674288 616752
rect 674340 616740 674346 616752
rect 676214 616740 676220 616752
rect 674340 616712 676220 616740
rect 674340 616700 674346 616712
rect 676214 616700 676220 616712
rect 676272 616700 676278 616752
rect 42150 614184 42156 614236
rect 42208 614224 42214 614236
rect 42518 614224 42524 614236
rect 42208 614196 42524 614224
rect 42208 614184 42214 614196
rect 42518 614184 42524 614196
rect 42576 614184 42582 614236
rect 671338 614116 671344 614168
rect 671396 614156 671402 614168
rect 683114 614156 683120 614168
rect 671396 614128 683120 614156
rect 671396 614116 671402 614128
rect 683114 614116 683120 614128
rect 683172 614116 683178 614168
rect 42150 612756 42156 612808
rect 42208 612796 42214 612808
rect 42518 612796 42524 612808
rect 42208 612768 42524 612796
rect 42208 612756 42214 612768
rect 42518 612756 42524 612768
rect 42576 612756 42582 612808
rect 48958 609968 48964 610020
rect 49016 610008 49022 610020
rect 62114 610008 62120 610020
rect 49016 609980 62120 610008
rect 49016 609968 49022 609980
rect 62114 609968 62120 609980
rect 62172 609968 62178 610020
rect 670602 607996 670608 608048
rect 670660 608036 670666 608048
rect 675386 608036 675392 608048
rect 670660 608008 675392 608036
rect 670660 607996 670666 608008
rect 675386 607996 675392 608008
rect 675444 607996 675450 608048
rect 673362 607588 673368 607640
rect 673420 607628 673426 607640
rect 675386 607628 675392 607640
rect 673420 607600 675392 607628
rect 673420 607588 673426 607600
rect 675386 607588 675392 607600
rect 675444 607588 675450 607640
rect 675202 604528 675208 604580
rect 675260 604568 675266 604580
rect 675386 604568 675392 604580
rect 675260 604540 675392 604568
rect 675260 604528 675266 604540
rect 675386 604528 675392 604540
rect 675444 604528 675450 604580
rect 674466 604324 674472 604376
rect 674524 604364 674530 604376
rect 675386 604364 675392 604376
rect 674524 604336 675392 604364
rect 674524 604324 674530 604336
rect 675386 604324 675392 604336
rect 675444 604324 675450 604376
rect 674558 603236 674564 603288
rect 674616 603276 674622 603288
rect 675478 603276 675484 603288
rect 674616 603248 675484 603276
rect 674616 603236 674622 603248
rect 675478 603236 675484 603248
rect 675536 603236 675542 603288
rect 651558 603100 651564 603152
rect 651616 603140 651622 603152
rect 660298 603140 660304 603152
rect 651616 603112 660304 603140
rect 651616 603100 651622 603112
rect 660298 603100 660304 603112
rect 660356 603100 660362 603152
rect 673546 603032 673552 603084
rect 673604 603072 673610 603084
rect 675386 603072 675392 603084
rect 673604 603044 675392 603072
rect 673604 603032 673610 603044
rect 675386 603032 675392 603044
rect 675444 603032 675450 603084
rect 35802 601672 35808 601724
rect 35860 601712 35866 601724
rect 55950 601712 55956 601724
rect 35860 601684 55956 601712
rect 35860 601672 35866 601684
rect 55950 601672 55956 601684
rect 56008 601672 56014 601724
rect 35710 601604 35716 601656
rect 35768 601644 35774 601656
rect 43622 601644 43628 601656
rect 35768 601616 43628 601644
rect 35768 601604 35774 601616
rect 43622 601604 43628 601616
rect 43680 601604 43686 601656
rect 35618 601468 35624 601520
rect 35676 601508 35682 601520
rect 44174 601508 44180 601520
rect 35676 601480 44180 601508
rect 35676 601468 35682 601480
rect 44174 601468 44180 601480
rect 44232 601468 44238 601520
rect 35802 601332 35808 601384
rect 35860 601372 35866 601384
rect 51810 601372 51816 601384
rect 35860 601344 51816 601372
rect 35860 601332 35866 601344
rect 51810 601332 51816 601344
rect 51868 601332 51874 601384
rect 672810 600380 672816 600432
rect 672868 600420 672874 600432
rect 675478 600420 675484 600432
rect 672868 600392 675484 600420
rect 672868 600380 672874 600392
rect 675478 600380 675484 600392
rect 675536 600380 675542 600432
rect 674282 599768 674288 599820
rect 674340 599808 674346 599820
rect 675478 599808 675484 599820
rect 674340 599780 675484 599808
rect 674340 599768 674346 599780
rect 675478 599768 675484 599780
rect 675536 599768 675542 599820
rect 658918 599564 658924 599616
rect 658976 599604 658982 599616
rect 674742 599604 674748 599616
rect 658976 599576 674748 599604
rect 658976 599564 658982 599576
rect 674742 599564 674748 599576
rect 674800 599564 674806 599616
rect 674006 598408 674012 598460
rect 674064 598448 674070 598460
rect 675478 598448 675484 598460
rect 674064 598420 675484 598448
rect 674064 598408 674070 598420
rect 675478 598408 675484 598420
rect 675536 598408 675542 598460
rect 672902 597728 672908 597780
rect 672960 597768 672966 597780
rect 675478 597768 675484 597780
rect 672960 597740 675484 597768
rect 672960 597728 672966 597740
rect 675478 597728 675484 597740
rect 675536 597728 675542 597780
rect 50430 597524 50436 597576
rect 50488 597564 50494 597576
rect 62114 597564 62120 597576
rect 50488 597536 62120 597564
rect 50488 597524 50494 597536
rect 62114 597524 62120 597536
rect 62172 597524 62178 597576
rect 674742 596844 674748 596896
rect 674800 596884 674806 596896
rect 675386 596884 675392 596896
rect 674800 596856 675392 596884
rect 674800 596844 674806 596856
rect 675386 596844 675392 596856
rect 675444 596844 675450 596896
rect 672626 593376 672632 593428
rect 672684 593416 672690 593428
rect 675478 593416 675484 593428
rect 672684 593388 675484 593416
rect 672684 593376 672690 593388
rect 675478 593376 675484 593388
rect 675536 593376 675542 593428
rect 651558 590656 651564 590708
rect 651616 590696 651622 590708
rect 664438 590696 664444 590708
rect 651616 590668 664444 590696
rect 651616 590656 651622 590668
rect 664438 590656 664444 590668
rect 664496 590656 664502 590708
rect 41506 589908 41512 589960
rect 41564 589948 41570 589960
rect 53098 589948 53104 589960
rect 41564 589920 53104 589948
rect 41564 589908 41570 589920
rect 53098 589908 53104 589920
rect 53156 589908 53162 589960
rect 33778 585896 33784 585948
rect 33836 585936 33842 585948
rect 41874 585936 41880 585948
rect 33836 585908 41880 585936
rect 33836 585896 33842 585908
rect 41874 585896 41880 585908
rect 41932 585896 41938 585948
rect 32398 585760 32404 585812
rect 32456 585800 32462 585812
rect 41598 585800 41604 585812
rect 32456 585772 41604 585800
rect 32456 585760 32462 585772
rect 41598 585760 41604 585772
rect 41656 585760 41662 585812
rect 41874 584196 41880 584248
rect 41932 584196 41938 584248
rect 42058 584196 42064 584248
rect 42116 584236 42122 584248
rect 42702 584236 42708 584248
rect 42116 584208 42708 584236
rect 42116 584196 42122 584208
rect 42702 584196 42708 584208
rect 42760 584196 42766 584248
rect 41892 583976 41920 584196
rect 41874 583924 41880 583976
rect 41932 583924 41938 583976
rect 51810 583720 51816 583772
rect 51868 583760 51874 583772
rect 62114 583760 62120 583772
rect 51868 583732 62120 583760
rect 51868 583720 51874 583732
rect 62114 583720 62120 583732
rect 62172 583720 62178 583772
rect 42150 581272 42156 581324
rect 42208 581312 42214 581324
rect 47578 581312 47584 581324
rect 42208 581284 47584 581312
rect 42208 581272 42214 581284
rect 47578 581272 47584 581284
rect 47636 581272 47642 581324
rect 652018 581000 652024 581052
rect 652076 581040 652082 581052
rect 676030 581040 676036 581052
rect 652076 581012 676036 581040
rect 652076 581000 652082 581012
rect 676030 581000 676036 581012
rect 676088 581000 676094 581052
rect 672442 580048 672448 580100
rect 672500 580088 672506 580100
rect 676214 580088 676220 580100
rect 672500 580060 676220 580088
rect 672500 580048 672506 580060
rect 676214 580048 676220 580060
rect 676272 580048 676278 580100
rect 671430 579912 671436 579964
rect 671488 579952 671494 579964
rect 676122 579952 676128 579964
rect 671488 579924 676128 579952
rect 671488 579912 671494 579924
rect 676122 579912 676128 579924
rect 676180 579912 676186 579964
rect 659010 579776 659016 579828
rect 659068 579816 659074 579828
rect 676030 579816 676036 579828
rect 659068 579788 676036 579816
rect 659068 579776 659074 579788
rect 676030 579776 676036 579788
rect 676088 579776 676094 579828
rect 42978 579640 42984 579692
rect 43036 579680 43042 579692
rect 44634 579680 44640 579692
rect 43036 579652 44640 579680
rect 43036 579640 43042 579652
rect 44634 579640 44640 579652
rect 44692 579640 44698 579692
rect 42150 578416 42156 578468
rect 42208 578456 42214 578468
rect 42978 578456 42984 578468
rect 42208 578428 42984 578456
rect 42208 578416 42214 578428
rect 42978 578416 42984 578428
rect 43036 578416 43042 578468
rect 672534 578416 672540 578468
rect 672592 578456 672598 578468
rect 676214 578456 676220 578468
rect 672592 578428 676220 578456
rect 672592 578416 672598 578428
rect 676214 578416 676220 578428
rect 676272 578416 676278 578468
rect 672442 578280 672448 578332
rect 672500 578320 672506 578332
rect 676306 578320 676312 578332
rect 672500 578292 676312 578320
rect 672500 578280 672506 578292
rect 676306 578280 676312 578292
rect 676364 578280 676370 578332
rect 42978 578212 42984 578264
rect 43036 578252 43042 578264
rect 44358 578252 44364 578264
rect 43036 578224 44364 578252
rect 43036 578212 43042 578224
rect 44358 578212 44364 578224
rect 44416 578212 44422 578264
rect 672534 578212 672540 578264
rect 672592 578252 672598 578264
rect 676122 578252 676128 578264
rect 672592 578224 676128 578252
rect 672592 578212 672598 578224
rect 676122 578212 676128 578224
rect 676180 578212 676186 578264
rect 673454 578144 673460 578196
rect 673512 578184 673518 578196
rect 676030 578184 676036 578196
rect 673512 578156 676036 578184
rect 673512 578144 673518 578156
rect 676030 578144 676036 578156
rect 676088 578144 676094 578196
rect 673914 577600 673920 577652
rect 673972 577640 673978 577652
rect 676214 577640 676220 577652
rect 673972 577612 676220 577640
rect 673972 577600 673978 577612
rect 676214 577600 676220 577612
rect 676272 577600 676278 577652
rect 673822 577396 673828 577448
rect 673880 577436 673886 577448
rect 676030 577436 676036 577448
rect 673880 577408 676036 577436
rect 673880 577396 673886 577408
rect 676030 577396 676036 577408
rect 676088 577396 676094 577448
rect 42150 576920 42156 576972
rect 42208 576960 42214 576972
rect 42978 576960 42984 576972
rect 42208 576932 42984 576960
rect 42208 576920 42214 576932
rect 42978 576920 42984 576932
rect 43036 576920 43042 576972
rect 673638 576920 673644 576972
rect 673696 576960 673702 576972
rect 676030 576960 676036 576972
rect 673696 576932 676036 576960
rect 673696 576920 673702 576932
rect 676030 576920 676036 576932
rect 676088 576920 676094 576972
rect 44450 576892 44456 576904
rect 42168 576864 44456 576892
rect 42168 576632 42196 576864
rect 44450 576852 44456 576864
rect 44508 576852 44514 576904
rect 651558 576852 651564 576904
rect 651616 576892 651622 576904
rect 659010 576892 659016 576904
rect 651616 576864 659016 576892
rect 651616 576852 651622 576864
rect 659010 576852 659016 576864
rect 659068 576852 659074 576904
rect 42150 576580 42156 576632
rect 42208 576580 42214 576632
rect 42702 576376 42708 576428
rect 42760 576376 42766 576428
rect 42426 576308 42432 576360
rect 42484 576348 42490 576360
rect 42720 576348 42748 576376
rect 42484 576320 42748 576348
rect 42484 576308 42490 576320
rect 42150 576172 42156 576224
rect 42208 576212 42214 576224
rect 42208 576184 42380 576212
rect 42208 576172 42214 576184
rect 42352 576020 42380 576184
rect 42334 575968 42340 576020
rect 42392 575968 42398 576020
rect 671890 575832 671896 575884
rect 671948 575872 671954 575884
rect 676030 575872 676036 575884
rect 671948 575844 676036 575872
rect 671948 575832 671954 575844
rect 676030 575832 676036 575844
rect 676088 575832 676094 575884
rect 671798 575696 671804 575748
rect 671856 575736 671862 575748
rect 676122 575736 676128 575748
rect 671856 575708 676128 575736
rect 671856 575696 671862 575708
rect 676122 575696 676128 575708
rect 676180 575696 676186 575748
rect 670510 575560 670516 575612
rect 670568 575600 670574 575612
rect 676214 575600 676220 575612
rect 670568 575572 676220 575600
rect 670568 575560 670574 575572
rect 676214 575560 676220 575572
rect 676272 575560 676278 575612
rect 673730 574948 673736 575000
rect 673788 574988 673794 575000
rect 676030 574988 676036 575000
rect 673788 574960 676036 574988
rect 673788 574948 673794 574960
rect 676030 574948 676036 574960
rect 676088 574948 676094 575000
rect 42150 574676 42156 574728
rect 42208 574716 42214 574728
rect 42334 574716 42340 574728
rect 42208 574688 42340 574716
rect 42208 574676 42214 574688
rect 42334 574676 42340 574688
rect 42392 574676 42398 574728
rect 673270 574200 673276 574252
rect 673328 574240 673334 574252
rect 676214 574240 676220 574252
rect 673328 574212 676220 574240
rect 673328 574200 673334 574212
rect 676214 574200 676220 574212
rect 676272 574200 676278 574252
rect 42334 574132 42340 574184
rect 42392 574172 42398 574184
rect 42702 574172 42708 574184
rect 42392 574144 42708 574172
rect 42392 574132 42398 574144
rect 42702 574132 42708 574144
rect 42760 574132 42766 574184
rect 674650 574132 674656 574184
rect 674708 574172 674714 574184
rect 676030 574172 676036 574184
rect 674708 574144 676036 574172
rect 674708 574132 674714 574144
rect 676030 574132 676036 574144
rect 676088 574132 676094 574184
rect 674374 573724 674380 573776
rect 674432 573764 674438 573776
rect 676030 573764 676036 573776
rect 674432 573736 676036 573764
rect 674432 573724 674438 573736
rect 676030 573724 676036 573736
rect 676088 573724 676094 573776
rect 42150 573452 42156 573504
rect 42208 573492 42214 573504
rect 42886 573492 42892 573504
rect 42208 573464 42892 573492
rect 42208 573452 42214 573464
rect 42886 573452 42892 573464
rect 42944 573452 42950 573504
rect 41966 572704 41972 572756
rect 42024 572744 42030 572756
rect 42702 572744 42708 572756
rect 42024 572716 42708 572744
rect 42024 572704 42030 572716
rect 42702 572704 42708 572716
rect 42760 572704 42766 572756
rect 673178 571616 673184 571668
rect 673236 571656 673242 571668
rect 676214 571656 676220 571668
rect 673236 571628 676220 571656
rect 673236 571616 673242 571628
rect 676214 571616 676220 571628
rect 676272 571616 676278 571668
rect 42334 571480 42340 571532
rect 42392 571480 42398 571532
rect 672994 571480 673000 571532
rect 673052 571520 673058 571532
rect 676214 571520 676220 571532
rect 673052 571492 676220 571520
rect 673052 571480 673058 571492
rect 676214 571480 676220 571492
rect 676272 571480 676278 571532
rect 42058 570868 42064 570920
rect 42116 570908 42122 570920
rect 42352 570908 42380 571480
rect 43714 571344 43720 571396
rect 43772 571384 43778 571396
rect 62114 571384 62120 571396
rect 43772 571356 62120 571384
rect 43772 571344 43778 571356
rect 62114 571344 62120 571356
rect 62172 571344 62178 571396
rect 42116 570880 42380 570908
rect 42116 570868 42122 570880
rect 673086 569916 673092 569968
rect 673144 569956 673150 569968
rect 676214 569956 676220 569968
rect 673144 569928 676220 569956
rect 673144 569916 673150 569928
rect 676214 569916 676220 569928
rect 676272 569916 676278 569968
rect 42058 569576 42064 569628
rect 42116 569616 42122 569628
rect 42702 569616 42708 569628
rect 42116 569588 42708 569616
rect 42116 569576 42122 569588
rect 42702 569576 42708 569588
rect 42760 569576 42766 569628
rect 671430 568556 671436 568608
rect 671488 568596 671494 568608
rect 683114 568596 683120 568608
rect 671488 568568 683120 568596
rect 671488 568556 671494 568568
rect 683114 568556 683120 568568
rect 683172 568556 683178 568608
rect 35618 566448 35624 566500
rect 35676 566488 35682 566500
rect 43714 566488 43720 566500
rect 35676 566460 43720 566488
rect 35676 566448 35682 566460
rect 43714 566448 43720 566460
rect 43772 566448 43778 566500
rect 652110 563048 652116 563100
rect 652168 563088 652174 563100
rect 658918 563088 658924 563100
rect 652168 563060 658924 563088
rect 652168 563048 652174 563060
rect 658918 563048 658924 563060
rect 658976 563048 658982 563100
rect 671982 561892 671988 561944
rect 672040 561932 672046 561944
rect 675386 561932 675392 561944
rect 672040 561904 675392 561932
rect 672040 561892 672046 561904
rect 675386 561892 675392 561904
rect 675444 561892 675450 561944
rect 673270 559104 673276 559156
rect 673328 559144 673334 559156
rect 675386 559144 675392 559156
rect 673328 559116 675392 559144
rect 673328 559104 673334 559116
rect 675386 559104 675392 559116
rect 675444 559104 675450 559156
rect 35710 558288 35716 558340
rect 35768 558328 35774 558340
rect 50430 558328 50436 558340
rect 35768 558300 50436 558328
rect 35768 558288 35774 558300
rect 50430 558288 50436 558300
rect 50488 558288 50494 558340
rect 35802 558152 35808 558204
rect 35860 558192 35866 558204
rect 51810 558192 51816 558204
rect 35860 558164 51816 558192
rect 35860 558152 35866 558164
rect 51810 558152 51816 558164
rect 51868 558152 51874 558204
rect 47578 557540 47584 557592
rect 47636 557580 47642 557592
rect 62114 557580 62120 557592
rect 47636 557552 62120 557580
rect 47636 557540 47642 557552
rect 62114 557540 62120 557552
rect 62172 557540 62178 557592
rect 673178 557540 673184 557592
rect 673236 557580 673242 557592
rect 675478 557580 675484 557592
rect 673236 557552 675484 557580
rect 673236 557540 673242 557552
rect 675478 557540 675484 557552
rect 675536 557540 675542 557592
rect 674742 555228 674748 555280
rect 674800 555268 674806 555280
rect 675386 555268 675392 555280
rect 674800 555240 675392 555268
rect 674800 555228 674806 555240
rect 675386 555228 675392 555240
rect 675444 555228 675450 555280
rect 673086 554752 673092 554804
rect 673144 554792 673150 554804
rect 675294 554792 675300 554804
rect 673144 554764 675300 554792
rect 673144 554752 673150 554764
rect 675294 554752 675300 554764
rect 675352 554752 675358 554804
rect 658918 554004 658924 554056
rect 658976 554044 658982 554056
rect 675294 554044 675300 554056
rect 658976 554016 675300 554044
rect 658976 554004 658982 554016
rect 675294 554004 675300 554016
rect 675352 554004 675358 554056
rect 674374 553392 674380 553444
rect 674432 553432 674438 553444
rect 675386 553432 675392 553444
rect 674432 553404 675392 553432
rect 674432 553392 674438 553404
rect 675386 553392 675392 553404
rect 675444 553392 675450 553444
rect 651558 550604 651564 550656
rect 651616 550644 651622 550656
rect 661770 550644 661776 550656
rect 651616 550616 661776 550644
rect 651616 550604 651622 550616
rect 661770 550604 661776 550616
rect 661828 550604 661834 550656
rect 674650 549312 674656 549364
rect 674708 549352 674714 549364
rect 674926 549352 674932 549364
rect 674708 549324 674932 549352
rect 674708 549312 674714 549324
rect 674926 549312 674932 549324
rect 674984 549312 674990 549364
rect 674926 549176 674932 549228
rect 674984 549216 674990 549228
rect 675294 549216 675300 549228
rect 674984 549188 675300 549216
rect 674984 549176 674990 549188
rect 675294 549176 675300 549188
rect 675352 549176 675358 549228
rect 674742 548468 674748 548480
rect 674392 548440 674748 548468
rect 674392 547936 674420 548440
rect 674742 548428 674748 548440
rect 674800 548428 674806 548480
rect 674742 548292 674748 548344
rect 674800 548332 674806 548344
rect 675294 548332 675300 548344
rect 674800 548304 675300 548332
rect 674800 548292 674806 548304
rect 675294 548292 675300 548304
rect 675352 548292 675358 548344
rect 674650 547952 674656 548004
rect 674708 547992 674714 548004
rect 675754 547992 675760 548004
rect 674708 547964 675760 547992
rect 674708 547952 674714 547964
rect 675754 547952 675760 547964
rect 675812 547952 675818 548004
rect 674374 547884 674380 547936
rect 674432 547884 674438 547936
rect 31662 547136 31668 547188
rect 31720 547176 31726 547188
rect 35802 547176 35808 547188
rect 31720 547148 35808 547176
rect 31720 547136 31726 547148
rect 35802 547136 35808 547148
rect 35860 547176 35866 547188
rect 53190 547176 53196 547188
rect 35860 547148 53196 547176
rect 35860 547136 35866 547148
rect 53190 547136 53196 547148
rect 53248 547136 53254 547188
rect 43622 545096 43628 545148
rect 43680 545136 43686 545148
rect 62114 545136 62120 545148
rect 43680 545108 62120 545136
rect 43680 545096 43686 545108
rect 62114 545096 62120 545108
rect 62172 545096 62178 545148
rect 31018 542988 31024 543040
rect 31076 543028 31082 543040
rect 41782 543028 41788 543040
rect 31076 543000 41788 543028
rect 31076 542988 31082 543000
rect 41782 542988 41788 543000
rect 41840 542988 41846 543040
rect 40678 542308 40684 542360
rect 40736 542348 40742 542360
rect 42702 542348 42708 542360
rect 40736 542320 42708 542348
rect 40736 542308 40742 542320
rect 42702 542308 42708 542320
rect 42760 542308 42766 542360
rect 41782 541016 41788 541068
rect 41840 541016 41846 541068
rect 41800 540796 41828 541016
rect 41782 540744 41788 540796
rect 41840 540744 41846 540796
rect 42978 540200 42984 540252
rect 43036 540240 43042 540252
rect 48958 540240 48964 540252
rect 43036 540212 48964 540240
rect 43036 540200 43042 540212
rect 48958 540200 48964 540212
rect 49016 540200 49022 540252
rect 42058 538908 42064 538960
rect 42116 538948 42122 538960
rect 42702 538948 42708 538960
rect 42116 538920 42708 538948
rect 42116 538908 42122 538920
rect 42702 538908 42708 538920
rect 42760 538908 42766 538960
rect 42978 538404 42984 538416
rect 42168 538376 42984 538404
rect 42168 538280 42196 538376
rect 42978 538364 42984 538376
rect 43036 538364 43042 538416
rect 42150 538228 42156 538280
rect 42208 538228 42214 538280
rect 42978 538228 42984 538280
rect 43036 538268 43042 538280
rect 44174 538268 44180 538280
rect 43036 538240 44180 538268
rect 43036 538228 43042 538240
rect 44174 538228 44180 538240
rect 44232 538228 44238 538280
rect 42058 537072 42064 537124
rect 42116 537112 42122 537124
rect 42978 537112 42984 537124
rect 42116 537084 42984 537112
rect 42116 537072 42122 537084
rect 42978 537072 42984 537084
rect 43036 537072 43042 537124
rect 42610 536800 42616 536852
rect 42668 536840 42674 536852
rect 44542 536840 44548 536852
rect 42668 536812 44548 536840
rect 42668 536800 42674 536812
rect 44542 536800 44548 536812
rect 44600 536800 44606 536852
rect 651558 536800 651564 536852
rect 651616 536840 651622 536852
rect 660390 536840 660396 536852
rect 651616 536812 660396 536840
rect 651616 536800 651622 536812
rect 660390 536800 660396 536812
rect 660448 536800 660454 536852
rect 42610 535984 42616 536036
rect 42668 535984 42674 536036
rect 42150 535780 42156 535832
rect 42208 535820 42214 535832
rect 42628 535820 42656 535984
rect 42208 535792 42656 535820
rect 42208 535780 42214 535792
rect 668670 535712 668676 535764
rect 668728 535752 668734 535764
rect 676214 535752 676220 535764
rect 668728 535724 676220 535752
rect 668728 535712 668734 535724
rect 676214 535712 676220 535724
rect 676272 535712 676278 535764
rect 663058 535576 663064 535628
rect 663116 535616 663122 535628
rect 676030 535616 676036 535628
rect 663116 535588 676036 535616
rect 663116 535576 663122 535588
rect 676030 535576 676036 535588
rect 676088 535576 676094 535628
rect 42058 535236 42064 535288
rect 42116 535276 42122 535288
rect 43070 535276 43076 535288
rect 42116 535248 43076 535276
rect 42116 535236 42122 535248
rect 43070 535236 43076 535248
rect 43128 535236 43134 535288
rect 672442 534488 672448 534540
rect 672500 534528 672506 534540
rect 676214 534528 676220 534540
rect 672500 534500 676220 534528
rect 672500 534488 672506 534500
rect 676214 534488 676220 534500
rect 676272 534488 676278 534540
rect 672534 534352 672540 534404
rect 672592 534392 672598 534404
rect 676214 534392 676220 534404
rect 672592 534364 676220 534392
rect 672592 534352 672598 534364
rect 676214 534352 676220 534364
rect 676272 534352 676278 534404
rect 661678 534216 661684 534268
rect 661736 534256 661742 534268
rect 676122 534256 676128 534268
rect 661736 534228 676128 534256
rect 661736 534216 661742 534228
rect 676122 534216 676128 534228
rect 676180 534216 676186 534268
rect 42150 533944 42156 533996
rect 42208 533984 42214 533996
rect 42610 533984 42616 533996
rect 42208 533956 42616 533984
rect 42208 533944 42214 533956
rect 42610 533944 42616 533956
rect 42668 533944 42674 533996
rect 673914 533264 673920 533316
rect 673972 533304 673978 533316
rect 676030 533304 676036 533316
rect 673972 533276 676036 533304
rect 673972 533264 673978 533276
rect 676030 533264 676036 533276
rect 676088 533264 676094 533316
rect 55950 532720 55956 532772
rect 56008 532760 56014 532772
rect 62114 532760 62120 532772
rect 56008 532732 62120 532760
rect 56008 532720 56014 532732
rect 62114 532720 62120 532732
rect 62172 532720 62178 532772
rect 673638 532652 673644 532704
rect 673696 532692 673702 532704
rect 676214 532692 676220 532704
rect 673696 532664 676220 532692
rect 673696 532652 673702 532664
rect 676214 532652 676220 532664
rect 676272 532652 676278 532704
rect 44450 531332 44456 531344
rect 42720 531304 44456 531332
rect 42150 530884 42156 530936
rect 42208 530924 42214 530936
rect 42610 530924 42616 530936
rect 42208 530896 42616 530924
rect 42208 530884 42214 530896
rect 42610 530884 42616 530896
rect 42668 530884 42674 530936
rect 42610 530748 42616 530800
rect 42668 530788 42674 530800
rect 42720 530788 42748 531304
rect 44450 531292 44456 531304
rect 44508 531292 44514 531344
rect 42668 530760 42748 530788
rect 42668 530748 42674 530760
rect 672810 530136 672816 530188
rect 672868 530176 672874 530188
rect 676214 530176 676220 530188
rect 672868 530148 676220 530176
rect 672868 530136 672874 530148
rect 676214 530136 676220 530148
rect 676272 530136 676278 530188
rect 42150 530068 42156 530120
rect 42208 530108 42214 530120
rect 42610 530108 42616 530120
rect 42208 530080 42616 530108
rect 42208 530068 42214 530080
rect 42610 530068 42616 530080
rect 42668 530068 42674 530120
rect 670602 530000 670608 530052
rect 670660 530040 670666 530052
rect 676122 530040 676128 530052
rect 670660 530012 676128 530040
rect 670660 530000 670666 530012
rect 676122 530000 676128 530012
rect 676180 530000 676186 530052
rect 42334 529632 42340 529644
rect 42260 529604 42340 529632
rect 42150 529456 42156 529508
rect 42208 529496 42214 529508
rect 42260 529496 42288 529604
rect 42334 529592 42340 529604
rect 42392 529592 42398 529644
rect 42208 529468 42288 529496
rect 42208 529456 42214 529468
rect 674466 528980 674472 529032
rect 674524 529020 674530 529032
rect 676398 529020 676404 529032
rect 674524 528992 676404 529020
rect 674524 528980 674530 528992
rect 676398 528980 676404 528992
rect 676456 528980 676462 529032
rect 673362 528776 673368 528828
rect 673420 528816 673426 528828
rect 676214 528816 676220 528828
rect 673420 528788 676220 528816
rect 673420 528776 673426 528788
rect 676214 528776 676220 528788
rect 676272 528776 676278 528828
rect 672626 528640 672632 528692
rect 672684 528680 672690 528692
rect 676122 528680 676128 528692
rect 672684 528652 676128 528680
rect 672684 528640 672690 528652
rect 676122 528640 676128 528652
rect 676180 528640 676186 528692
rect 674558 528368 674564 528420
rect 674616 528408 674622 528420
rect 675846 528408 675852 528420
rect 674616 528380 675852 528408
rect 674616 528368 674622 528380
rect 675846 528368 675852 528380
rect 675904 528368 675910 528420
rect 672902 527416 672908 527468
rect 672960 527456 672966 527468
rect 676214 527456 676220 527468
rect 672960 527428 676220 527456
rect 672960 527416 672966 527428
rect 676214 527416 676220 527428
rect 676272 527416 676278 527468
rect 42058 527212 42064 527264
rect 42116 527252 42122 527264
rect 42334 527252 42340 527264
rect 42116 527224 42340 527252
rect 42116 527212 42122 527224
rect 42334 527212 42340 527224
rect 42392 527212 42398 527264
rect 42150 527144 42156 527196
rect 42208 527184 42214 527196
rect 42886 527184 42892 527196
rect 42208 527156 42892 527184
rect 42208 527144 42214 527156
rect 42886 527144 42892 527156
rect 42944 527144 42950 527196
rect 673546 527076 673552 527128
rect 673604 527116 673610 527128
rect 675846 527116 675852 527128
rect 673604 527088 675852 527116
rect 673604 527076 673610 527088
rect 675846 527076 675852 527088
rect 675904 527076 675910 527128
rect 674282 526940 674288 526992
rect 674340 526980 674346 526992
rect 676214 526980 676220 526992
rect 674340 526952 676220 526980
rect 674340 526940 674346 526952
rect 676214 526940 676220 526952
rect 676272 526940 676278 526992
rect 42150 526600 42156 526652
rect 42208 526640 42214 526652
rect 42610 526640 42616 526652
rect 42208 526612 42616 526640
rect 42208 526600 42214 526612
rect 42610 526600 42616 526612
rect 42668 526600 42674 526652
rect 674006 526532 674012 526584
rect 674064 526572 674070 526584
rect 676214 526572 676220 526584
rect 674064 526544 676220 526572
rect 674064 526532 674070 526544
rect 676214 526532 676220 526544
rect 676272 526532 676278 526584
rect 674466 524424 674472 524476
rect 674524 524464 674530 524476
rect 683114 524464 683120 524476
rect 674524 524436 683120 524464
rect 674524 524424 674530 524436
rect 683114 524424 683120 524436
rect 683172 524424 683178 524476
rect 651558 522996 651564 523048
rect 651616 523036 651622 523048
rect 663242 523036 663248 523048
rect 651616 523008 663248 523036
rect 651616 522996 651622 523008
rect 663242 522996 663248 523008
rect 663300 522996 663306 523048
rect 677318 520276 677324 520328
rect 677376 520316 677382 520328
rect 683850 520316 683856 520328
rect 677376 520288 683856 520316
rect 677376 520276 677382 520288
rect 683850 520276 683856 520288
rect 683908 520276 683914 520328
rect 40678 518916 40684 518968
rect 40736 518956 40742 518968
rect 62114 518956 62120 518968
rect 40736 518928 62120 518956
rect 40736 518916 40742 518928
rect 62114 518916 62120 518928
rect 62172 518916 62178 518968
rect 651558 510620 651564 510672
rect 651616 510660 651622 510672
rect 661678 510660 661684 510672
rect 651616 510632 661684 510660
rect 651616 510620 651622 510632
rect 661678 510620 661684 510632
rect 661736 510620 661742 510672
rect 48958 506472 48964 506524
rect 49016 506512 49022 506524
rect 62114 506512 62120 506524
rect 49016 506484 62120 506512
rect 49016 506472 49022 506484
rect 62114 506472 62120 506484
rect 62172 506472 62178 506524
rect 675018 500896 675024 500948
rect 675076 500936 675082 500948
rect 680998 500936 681004 500948
rect 675076 500908 681004 500936
rect 675076 500896 675082 500908
rect 680998 500896 681004 500908
rect 681056 500896 681062 500948
rect 674926 498244 674932 498296
rect 674984 498284 674990 498296
rect 679710 498284 679716 498296
rect 674984 498256 679716 498284
rect 674984 498244 674990 498256
rect 679710 498244 679716 498256
rect 679768 498244 679774 498296
rect 675754 498176 675760 498228
rect 675812 498216 675818 498228
rect 679618 498216 679624 498228
rect 675812 498188 679624 498216
rect 675812 498176 675818 498188
rect 679618 498176 679624 498188
rect 679676 498176 679682 498228
rect 651558 496816 651564 496868
rect 651616 496856 651622 496868
rect 658918 496856 658924 496868
rect 651616 496828 658924 496856
rect 651616 496816 651622 496828
rect 658918 496816 658924 496828
rect 658976 496816 658982 496868
rect 46198 491920 46204 491972
rect 46256 491960 46262 491972
rect 62114 491960 62120 491972
rect 46256 491932 62120 491960
rect 46256 491920 46262 491932
rect 62114 491920 62120 491932
rect 62172 491920 62178 491972
rect 664438 491648 664444 491700
rect 664496 491688 664502 491700
rect 675846 491688 675852 491700
rect 664496 491660 675852 491688
rect 664496 491648 664502 491660
rect 675846 491648 675852 491660
rect 675904 491648 675910 491700
rect 660298 491512 660304 491564
rect 660356 491552 660362 491564
rect 675938 491552 675944 491564
rect 660356 491524 675944 491552
rect 660356 491512 660362 491524
rect 675938 491512 675944 491524
rect 675996 491512 676002 491564
rect 659010 491376 659016 491428
rect 659068 491416 659074 491428
rect 675938 491416 675944 491428
rect 659068 491388 675944 491416
rect 659068 491376 659074 491388
rect 675938 491376 675944 491388
rect 675996 491376 676002 491428
rect 675938 490152 675944 490204
rect 675996 490192 676002 490204
rect 676122 490192 676128 490204
rect 675996 490164 676128 490192
rect 675996 490152 676002 490164
rect 676122 490152 676128 490164
rect 676180 490152 676186 490204
rect 676030 488792 676036 488844
rect 676088 488832 676094 488844
rect 677318 488832 677324 488844
rect 676088 488804 677324 488832
rect 676088 488792 676094 488804
rect 677318 488792 677324 488804
rect 677376 488792 677382 488844
rect 676030 488452 676036 488504
rect 676088 488492 676094 488504
rect 677226 488492 677232 488504
rect 676088 488464 677232 488492
rect 676088 488452 676094 488464
rect 677226 488452 677232 488464
rect 677284 488452 677290 488504
rect 676030 487976 676036 488028
rect 676088 488016 676094 488028
rect 677226 488016 677232 488028
rect 676088 487988 677232 488016
rect 676088 487976 676094 487988
rect 677226 487976 677232 487988
rect 677284 487976 677290 488028
rect 676030 486820 676036 486872
rect 676088 486860 676094 486872
rect 677502 486860 677508 486872
rect 676088 486832 677508 486860
rect 676088 486820 676094 486832
rect 677502 486820 677508 486832
rect 677560 486820 677566 486872
rect 674374 486004 674380 486056
rect 674432 486044 674438 486056
rect 676030 486044 676036 486056
rect 674432 486016 676036 486044
rect 674432 486004 674438 486016
rect 676030 486004 676036 486016
rect 676088 486004 676094 486056
rect 671982 485188 671988 485240
rect 672040 485228 672046 485240
rect 675938 485228 675944 485240
rect 672040 485200 675944 485228
rect 672040 485188 672046 485200
rect 675938 485188 675944 485200
rect 675996 485188 676002 485240
rect 673270 484780 673276 484832
rect 673328 484820 673334 484832
rect 675938 484820 675944 484832
rect 673328 484792 675944 484820
rect 673328 484780 673334 484792
rect 675938 484780 675944 484792
rect 675996 484780 676002 484832
rect 651558 484372 651564 484424
rect 651616 484412 651622 484424
rect 660482 484412 660488 484424
rect 651616 484384 660488 484412
rect 651616 484372 651622 484384
rect 660482 484372 660488 484384
rect 660540 484372 660546 484424
rect 673178 483148 673184 483200
rect 673236 483188 673242 483200
rect 675938 483188 675944 483200
rect 673236 483160 675944 483188
rect 673236 483148 673242 483160
rect 675938 483148 675944 483160
rect 675996 483148 676002 483200
rect 673086 482740 673092 482792
rect 673144 482780 673150 482792
rect 675938 482780 675944 482792
rect 673144 482752 675944 482780
rect 673144 482740 673150 482752
rect 675938 482740 675944 482752
rect 675996 482740 676002 482792
rect 44818 480224 44824 480276
rect 44876 480264 44882 480276
rect 62114 480264 62120 480276
rect 44876 480236 62120 480264
rect 44876 480224 44882 480236
rect 62114 480224 62120 480236
rect 62172 480224 62178 480276
rect 674282 480224 674288 480276
rect 674340 480264 674346 480276
rect 678974 480264 678980 480276
rect 674340 480236 678980 480264
rect 674340 480224 674346 480236
rect 678974 480224 678980 480236
rect 679032 480224 679038 480276
rect 668578 475804 668584 475856
rect 668636 475844 668642 475856
rect 674466 475844 674472 475856
rect 668636 475816 674472 475844
rect 668636 475804 668642 475816
rect 674466 475804 674472 475816
rect 674524 475804 674530 475856
rect 668670 474512 668676 474564
rect 668728 474552 668734 474564
rect 671430 474552 671436 474564
rect 668728 474524 671436 474552
rect 668728 474512 668734 474524
rect 671430 474512 671436 474524
rect 671488 474512 671494 474564
rect 651650 470568 651656 470620
rect 651708 470608 651714 470620
rect 664530 470608 664536 470620
rect 651708 470580 664536 470608
rect 651708 470568 651714 470580
rect 664530 470568 664536 470580
rect 664588 470568 664594 470620
rect 51810 466420 51816 466472
rect 51868 466460 51874 466472
rect 62114 466460 62120 466472
rect 51868 466432 62120 466460
rect 51868 466420 51874 466432
rect 62114 466420 62120 466432
rect 62172 466420 62178 466472
rect 651558 456764 651564 456816
rect 651616 456804 651622 456816
rect 663150 456804 663156 456816
rect 651616 456776 663156 456804
rect 651616 456764 651622 456776
rect 663150 456764 663156 456776
rect 663208 456764 663214 456816
rect 50430 454044 50436 454096
rect 50488 454084 50494 454096
rect 62114 454084 62120 454096
rect 50488 454056 62120 454084
rect 50488 454044 50494 454056
rect 62114 454044 62120 454056
rect 62172 454044 62178 454096
rect 651558 444388 651564 444440
rect 651616 444428 651622 444440
rect 659010 444428 659016 444440
rect 651616 444400 659016 444428
rect 651616 444388 651622 444400
rect 659010 444388 659016 444400
rect 659068 444388 659074 444440
rect 43714 440240 43720 440292
rect 43772 440280 43778 440292
rect 62114 440280 62120 440292
rect 43772 440252 62120 440280
rect 43772 440240 43778 440252
rect 62114 440240 62120 440252
rect 62172 440240 62178 440292
rect 40678 432556 40684 432608
rect 40736 432596 40742 432608
rect 41782 432596 41788 432608
rect 40736 432568 41788 432596
rect 40736 432556 40742 432568
rect 41782 432556 41788 432568
rect 41840 432556 41846 432608
rect 43162 430584 43168 430636
rect 43220 430624 43226 430636
rect 55950 430624 55956 430636
rect 43220 430596 55956 430624
rect 43220 430584 43226 430596
rect 55950 430584 55956 430596
rect 56008 430584 56014 430636
rect 651558 430584 651564 430636
rect 651616 430624 651622 430636
rect 660298 430624 660304 430636
rect 651616 430596 660304 430624
rect 651616 430584 651622 430596
rect 660298 430584 660304 430596
rect 660356 430584 660362 430636
rect 46290 427796 46296 427848
rect 46348 427836 46354 427848
rect 62114 427836 62120 427848
rect 46348 427808 62120 427836
rect 46348 427796 46354 427808
rect 62114 427796 62120 427808
rect 62172 427796 62178 427848
rect 41782 419432 41788 419484
rect 41840 419472 41846 419484
rect 43622 419472 43628 419484
rect 41840 419444 43628 419472
rect 41840 419432 41846 419444
rect 43622 419432 43628 419444
rect 43680 419432 43686 419484
rect 651558 416780 651564 416832
rect 651616 416820 651622 416832
rect 663058 416820 663064 416832
rect 651616 416792 663064 416820
rect 651616 416780 651622 416792
rect 663058 416780 663064 416792
rect 663116 416780 663122 416832
rect 55950 415420 55956 415472
rect 56008 415460 56014 415472
rect 62114 415460 62120 415472
rect 56008 415432 62120 415460
rect 56008 415420 56014 415432
rect 62114 415420 62120 415432
rect 62172 415420 62178 415472
rect 32490 414808 32496 414860
rect 32548 414848 32554 414860
rect 41874 414848 41880 414860
rect 32548 414820 41880 414848
rect 32548 414808 32554 414820
rect 41874 414808 41880 414820
rect 41932 414808 41938 414860
rect 31018 414672 31024 414724
rect 31076 414712 31082 414724
rect 42518 414712 42524 414724
rect 31076 414684 42524 414712
rect 31076 414672 31082 414684
rect 42518 414672 42524 414684
rect 42576 414672 42582 414724
rect 41874 413380 41880 413432
rect 41932 413380 41938 413432
rect 41892 413160 41920 413380
rect 41874 413108 41880 413160
rect 41932 413108 41938 413160
rect 42150 410660 42156 410712
rect 42208 410700 42214 410712
rect 47578 410700 47584 410712
rect 42208 410672 47584 410700
rect 42208 410660 42214 410672
rect 47578 410660 47584 410672
rect 47636 410660 47642 410712
rect 42058 408144 42064 408196
rect 42116 408184 42122 408196
rect 44634 408184 44640 408196
rect 42116 408156 44640 408184
rect 42116 408144 42122 408156
rect 44634 408144 44640 408156
rect 44692 408144 44698 408196
rect 42150 407600 42156 407652
rect 42208 407640 42214 407652
rect 42518 407640 42524 407652
rect 42208 407612 42524 407640
rect 42208 407600 42214 407612
rect 42518 407600 42524 407612
rect 42576 407600 42582 407652
rect 42058 406784 42064 406836
rect 42116 406824 42122 406836
rect 42978 406824 42984 406836
rect 42116 406796 42984 406824
rect 42116 406784 42122 406796
rect 42978 406784 42984 406796
rect 43036 406784 43042 406836
rect 652018 404336 652024 404388
rect 652076 404376 652082 404388
rect 661862 404376 661868 404388
rect 652076 404348 661868 404376
rect 652076 404336 652082 404348
rect 661862 404336 661868 404348
rect 661920 404336 661926 404388
rect 42150 403860 42156 403912
rect 42208 403900 42214 403912
rect 44450 403900 44456 403912
rect 42208 403872 44456 403900
rect 42208 403860 42214 403872
rect 44450 403860 44456 403872
rect 44508 403860 44514 403912
rect 663242 403384 663248 403436
rect 663300 403424 663306 403436
rect 676398 403424 676404 403436
rect 663300 403396 676404 403424
rect 663300 403384 663306 403396
rect 676398 403384 676404 403396
rect 676456 403384 676462 403436
rect 661770 403248 661776 403300
rect 661828 403288 661834 403300
rect 676214 403288 676220 403300
rect 661828 403260 676220 403288
rect 661828 403248 661834 403260
rect 676214 403248 676220 403260
rect 676272 403248 676278 403300
rect 660390 403112 660396 403164
rect 660448 403152 660454 403164
rect 676306 403152 676312 403164
rect 660448 403124 676312 403152
rect 660448 403112 660454 403124
rect 676306 403112 676312 403124
rect 676364 403112 676370 403164
rect 42150 402908 42156 402960
rect 42208 402948 42214 402960
rect 42886 402948 42892 402960
rect 42208 402920 42892 402948
rect 42208 402908 42214 402920
rect 42886 402908 42892 402920
rect 42944 402908 42950 402960
rect 47578 401616 47584 401668
rect 47636 401656 47642 401668
rect 62114 401656 62120 401668
rect 47636 401628 62120 401656
rect 47636 401616 47642 401628
rect 62114 401616 62120 401628
rect 62172 401616 62178 401668
rect 673270 401616 673276 401668
rect 673328 401656 673334 401668
rect 676214 401656 676220 401668
rect 673328 401628 676220 401656
rect 673328 401616 673334 401628
rect 676214 401616 676220 401628
rect 676272 401616 676278 401668
rect 673362 400188 673368 400240
rect 673420 400228 673426 400240
rect 676214 400228 676220 400240
rect 673420 400200 676220 400228
rect 673420 400188 673426 400200
rect 676214 400188 676220 400200
rect 676272 400188 676278 400240
rect 674650 399576 674656 399628
rect 674708 399616 674714 399628
rect 676214 399616 676220 399628
rect 674708 399588 676220 399616
rect 674708 399576 674714 399588
rect 676214 399576 676220 399588
rect 676272 399576 676278 399628
rect 675018 398216 675024 398268
rect 675076 398256 675082 398268
rect 676030 398256 676036 398268
rect 675076 398228 676036 398256
rect 675076 398216 675082 398228
rect 676030 398216 676036 398228
rect 676088 398216 676094 398268
rect 674926 397468 674932 397520
rect 674984 397508 674990 397520
rect 676030 397508 676036 397520
rect 674984 397480 676036 397508
rect 674984 397468 674990 397480
rect 676030 397468 676036 397480
rect 676088 397468 676094 397520
rect 674558 394272 674564 394324
rect 674616 394312 674622 394324
rect 676214 394312 676220 394324
rect 674616 394284 676220 394312
rect 674616 394272 674622 394284
rect 676214 394272 676220 394284
rect 676272 394272 676278 394324
rect 673178 393320 673184 393372
rect 673236 393360 673242 393372
rect 676214 393360 676220 393372
rect 673236 393332 676220 393360
rect 673236 393320 673242 393332
rect 676214 393320 676220 393332
rect 676272 393320 676278 393372
rect 670142 391960 670148 392012
rect 670200 392000 670206 392012
rect 683114 392000 683120 392012
rect 670200 391972 683120 392000
rect 670200 391960 670206 391972
rect 683114 391960 683120 391972
rect 683172 391960 683178 392012
rect 651558 390532 651564 390584
rect 651616 390572 651622 390584
rect 664438 390572 664444 390584
rect 651616 390544 664444 390572
rect 651616 390532 651622 390544
rect 664438 390532 664444 390544
rect 664496 390532 664502 390584
rect 45002 389172 45008 389224
rect 45060 389212 45066 389224
rect 62114 389212 62120 389224
rect 45060 389184 62120 389212
rect 45060 389172 45066 389184
rect 62114 389172 62120 389184
rect 62172 389172 62178 389224
rect 675202 389104 675208 389156
rect 675260 389144 675266 389156
rect 676950 389144 676956 389156
rect 675260 389116 676956 389144
rect 675260 389104 675266 389116
rect 676950 389104 676956 389116
rect 677008 389104 677014 389156
rect 35710 387744 35716 387796
rect 35768 387784 35774 387796
rect 44174 387784 44180 387796
rect 35768 387756 44180 387784
rect 35768 387744 35774 387756
rect 44174 387744 44180 387756
rect 44232 387744 44238 387796
rect 35802 387608 35808 387660
rect 35860 387648 35866 387660
rect 44818 387648 44824 387660
rect 35860 387620 44824 387648
rect 35860 387608 35866 387620
rect 44818 387608 44824 387620
rect 44876 387608 44882 387660
rect 675110 387540 675116 387592
rect 675168 387580 675174 387592
rect 676490 387580 676496 387592
rect 675168 387552 676496 387580
rect 675168 387540 675174 387552
rect 676490 387540 676496 387552
rect 676548 387540 676554 387592
rect 35618 387472 35624 387524
rect 35676 387512 35682 387524
rect 46198 387512 46204 387524
rect 35676 387484 46204 387512
rect 35676 387472 35682 387484
rect 46198 387472 46204 387484
rect 46256 387472 46262 387524
rect 35802 387336 35808 387388
rect 35860 387376 35866 387388
rect 51810 387376 51816 387388
rect 35860 387348 51816 387376
rect 35860 387336 35866 387348
rect 51810 387336 51816 387348
rect 51868 387336 51874 387388
rect 675294 387064 675300 387116
rect 675352 387104 675358 387116
rect 678238 387104 678244 387116
rect 675352 387076 678244 387104
rect 675352 387064 675358 387076
rect 678238 387064 678244 387076
rect 678296 387064 678302 387116
rect 675018 386112 675024 386164
rect 675076 386152 675082 386164
rect 675386 386152 675392 386164
rect 675076 386124 675392 386152
rect 675076 386112 675082 386124
rect 675386 386112 675392 386124
rect 675444 386112 675450 386164
rect 675018 385976 675024 386028
rect 675076 386016 675082 386028
rect 675294 386016 675300 386028
rect 675076 385988 675300 386016
rect 675076 385976 675082 385988
rect 675294 385976 675300 385988
rect 675352 385976 675358 386028
rect 675018 383868 675024 383920
rect 675076 383908 675082 383920
rect 675294 383908 675300 383920
rect 675076 383880 675300 383908
rect 675076 383868 675082 383880
rect 675294 383868 675300 383880
rect 675352 383868 675358 383920
rect 674926 383052 674932 383104
rect 674984 383092 674990 383104
rect 675386 383092 675392 383104
rect 674984 383064 675392 383092
rect 674984 383052 674990 383064
rect 675386 383052 675392 383064
rect 675444 383052 675450 383104
rect 675110 381080 675116 381132
rect 675168 381120 675174 381132
rect 675386 381120 675392 381132
rect 675168 381092 675392 381120
rect 675168 381080 675174 381092
rect 675386 381080 675392 381092
rect 675444 381080 675450 381132
rect 651558 378156 651564 378208
rect 651616 378196 651622 378208
rect 665818 378196 665824 378208
rect 651616 378168 665824 378196
rect 651616 378156 651622 378168
rect 665818 378156 665824 378168
rect 665876 378156 665882 378208
rect 674558 377952 674564 378004
rect 674616 377992 674622 378004
rect 675478 377992 675484 378004
rect 674616 377964 675484 377992
rect 674616 377952 674622 377964
rect 675478 377952 675484 377964
rect 675536 377952 675542 378004
rect 673178 376592 673184 376644
rect 673236 376632 673242 376644
rect 675478 376632 675484 376644
rect 673236 376604 675484 376632
rect 673236 376592 673242 376604
rect 675478 376592 675484 376604
rect 675536 376592 675542 376644
rect 35802 376048 35808 376100
rect 35860 376088 35866 376100
rect 41506 376088 41512 376100
rect 35860 376060 41512 376088
rect 35860 376048 35866 376060
rect 41506 376048 41512 376060
rect 41564 376088 41570 376100
rect 44818 376088 44824 376100
rect 41564 376060 44824 376088
rect 41564 376048 41570 376060
rect 44818 376048 44824 376060
rect 44876 376048 44882 376100
rect 49050 375368 49056 375420
rect 49108 375408 49114 375420
rect 62114 375408 62120 375420
rect 49108 375380 62120 375408
rect 49108 375368 49114 375380
rect 62114 375368 62120 375380
rect 62172 375368 62178 375420
rect 31018 371832 31024 371884
rect 31076 371872 31082 371884
rect 42334 371872 42340 371884
rect 31076 371844 42340 371872
rect 31076 371832 31082 371844
rect 42334 371832 42340 371844
rect 42392 371832 42398 371884
rect 40862 371220 40868 371272
rect 40920 371260 40926 371272
rect 42702 371260 42708 371272
rect 40920 371232 42708 371260
rect 40920 371220 40926 371232
rect 42702 371220 42708 371232
rect 42760 371220 42766 371272
rect 40678 370540 40684 370592
rect 40736 370580 40742 370592
rect 41782 370580 41788 370592
rect 40736 370552 41788 370580
rect 40736 370540 40742 370552
rect 41782 370540 41788 370552
rect 41840 370540 41846 370592
rect 42150 369656 42156 369708
rect 42208 369696 42214 369708
rect 42334 369696 42340 369708
rect 42208 369668 42340 369696
rect 42208 369656 42214 369668
rect 42334 369656 42340 369668
rect 42392 369656 42398 369708
rect 42150 368092 42156 368144
rect 42208 368132 42214 368144
rect 42702 368132 42708 368144
rect 42208 368104 42708 368132
rect 42208 368092 42214 368104
rect 42702 368092 42708 368104
rect 42760 368092 42766 368144
rect 42150 366800 42156 366852
rect 42208 366840 42214 366852
rect 42702 366840 42708 366852
rect 42208 366812 42708 366840
rect 42208 366800 42214 366812
rect 42702 366800 42708 366812
rect 42760 366800 42766 366852
rect 42150 364964 42156 365016
rect 42208 365004 42214 365016
rect 44542 365004 44548 365016
rect 42208 364976 44548 365004
rect 42208 364964 42214 364976
rect 44542 364964 44548 364976
rect 44600 364964 44606 365016
rect 652018 364352 652024 364404
rect 652076 364392 652082 364404
rect 660390 364392 660396 364404
rect 652076 364364 660396 364392
rect 652076 364352 652082 364364
rect 660390 364352 660396 364364
rect 660448 364352 660454 364404
rect 42150 364284 42156 364336
rect 42208 364324 42214 364336
rect 44450 364324 44456 364336
rect 42208 364296 44456 364324
rect 42208 364284 42214 364296
rect 44450 364284 44456 364296
rect 44508 364284 44514 364336
rect 42702 364216 42708 364268
rect 42760 364256 42766 364268
rect 48958 364256 48964 364268
rect 42760 364228 48964 364256
rect 42760 364216 42766 364228
rect 48958 364216 48964 364228
rect 49016 364216 49022 364268
rect 56042 362924 56048 362976
rect 56100 362964 56106 362976
rect 62114 362964 62120 362976
rect 56100 362936 62120 362964
rect 56100 362924 56106 362936
rect 62114 362924 62120 362936
rect 62172 362924 62178 362976
rect 42058 360680 42064 360732
rect 42116 360720 42122 360732
rect 43070 360720 43076 360732
rect 42116 360692 43076 360720
rect 42116 360680 42122 360692
rect 43070 360680 43076 360692
rect 43128 360680 43134 360732
rect 42150 359456 42156 359508
rect 42208 359496 42214 359508
rect 42978 359496 42984 359508
rect 42208 359468 42984 359496
rect 42208 359456 42214 359468
rect 42978 359456 42984 359468
rect 43036 359456 43042 359508
rect 661678 357824 661684 357876
rect 661736 357864 661742 357876
rect 675938 357864 675944 357876
rect 661736 357836 675944 357864
rect 661736 357824 661742 357836
rect 675938 357824 675944 357836
rect 675996 357824 676002 357876
rect 660482 357688 660488 357740
rect 660540 357728 660546 357740
rect 676030 357728 676036 357740
rect 660540 357700 676036 357728
rect 660540 357688 660546 357700
rect 676030 357688 676036 357700
rect 676088 357688 676094 357740
rect 658918 357552 658924 357604
rect 658976 357592 658982 357604
rect 675846 357592 675852 357604
rect 658976 357564 675852 357592
rect 658976 357552 658982 357564
rect 675846 357552 675852 357564
rect 675904 357552 675910 357604
rect 673270 357484 673276 357536
rect 673328 357524 673334 357536
rect 676030 357524 676036 357536
rect 673328 357496 676036 357524
rect 673328 357484 673334 357496
rect 676030 357484 676036 357496
rect 676088 357484 676094 357536
rect 673270 357008 673276 357060
rect 673328 357048 673334 357060
rect 676030 357048 676036 357060
rect 673328 357020 676036 357048
rect 673328 357008 673334 357020
rect 676030 357008 676036 357020
rect 676088 357008 676094 357060
rect 673362 356668 673368 356720
rect 673420 356708 673426 356720
rect 676030 356708 676036 356720
rect 673420 356680 676036 356708
rect 673420 356668 673426 356680
rect 676030 356668 676036 356680
rect 676088 356668 676094 356720
rect 672994 356192 673000 356244
rect 673052 356232 673058 356244
rect 676030 356232 676036 356244
rect 673052 356204 676036 356232
rect 673052 356192 673058 356204
rect 676030 356192 676036 356204
rect 676088 356192 676094 356244
rect 42150 355988 42156 356040
rect 42208 356028 42214 356040
rect 43162 356028 43168 356040
rect 42208 356000 43168 356028
rect 42208 355988 42214 356000
rect 43162 355988 43168 356000
rect 43220 355988 43226 356040
rect 674650 355036 674656 355088
rect 674708 355076 674714 355088
rect 676030 355076 676036 355088
rect 674708 355048 676036 355076
rect 674708 355036 674714 355048
rect 676030 355036 676036 355048
rect 676088 355036 676094 355088
rect 674650 354560 674656 354612
rect 674708 354600 674714 354612
rect 676030 354600 676036 354612
rect 674708 354572 676036 354600
rect 674708 354560 674714 354572
rect 676030 354560 676036 354572
rect 676088 354560 676094 354612
rect 27614 351160 27620 351212
rect 27672 351200 27678 351212
rect 46290 351200 46296 351212
rect 27672 351172 46296 351200
rect 27672 351160 27678 351172
rect 46290 351160 46296 351172
rect 46348 351160 46354 351212
rect 676214 351092 676220 351144
rect 676272 351132 676278 351144
rect 676858 351132 676864 351144
rect 676272 351104 676864 351132
rect 676272 351092 676278 351104
rect 676858 351092 676864 351104
rect 676916 351092 676922 351144
rect 674466 350888 674472 350940
rect 674524 350928 674530 350940
rect 676030 350928 676036 350940
rect 674524 350900 676036 350928
rect 674524 350888 674530 350900
rect 676030 350888 676036 350900
rect 676088 350888 676094 350940
rect 651558 350548 651564 350600
rect 651616 350588 651622 350600
rect 671522 350588 671528 350600
rect 651616 350560 671528 350588
rect 651616 350548 651622 350560
rect 671522 350548 671528 350560
rect 671580 350548 671586 350600
rect 673178 350548 673184 350600
rect 673236 350588 673242 350600
rect 676030 350588 676036 350600
rect 673236 350560 676036 350588
rect 673236 350548 673242 350560
rect 676030 350548 676036 350560
rect 676088 350548 676094 350600
rect 674558 349256 674564 349308
rect 674616 349296 674622 349308
rect 676030 349296 676036 349308
rect 674616 349268 676036 349296
rect 674616 349256 674622 349268
rect 676030 349256 676036 349268
rect 676088 349256 676094 349308
rect 673086 348848 673092 348900
rect 673144 348888 673150 348900
rect 676030 348888 676036 348900
rect 673144 348860 676036 348888
rect 673144 348848 673150 348860
rect 676030 348848 676036 348860
rect 676088 348848 676094 348900
rect 44910 347012 44916 347064
rect 44968 347052 44974 347064
rect 62114 347052 62120 347064
rect 44968 347024 62120 347052
rect 44968 347012 44974 347024
rect 62114 347012 62120 347024
rect 62172 347012 62178 347064
rect 671430 346400 671436 346452
rect 671488 346440 671494 346452
rect 676030 346440 676036 346452
rect 671488 346412 676036 346440
rect 671488 346400 671494 346412
rect 676030 346400 676036 346412
rect 676088 346400 676094 346452
rect 35710 344292 35716 344344
rect 35768 344332 35774 344344
rect 43714 344332 43720 344344
rect 35768 344304 43720 344332
rect 35768 344292 35774 344304
rect 43714 344292 43720 344304
rect 43772 344292 43778 344344
rect 35802 344156 35808 344208
rect 35860 344196 35866 344208
rect 55950 344196 55956 344208
rect 35860 344168 55956 344196
rect 35860 344156 35866 344168
rect 55950 344156 55956 344168
rect 56008 344156 56014 344208
rect 651650 338104 651656 338156
rect 651708 338144 651714 338156
rect 668762 338144 668768 338156
rect 651708 338116 668768 338144
rect 651708 338104 651714 338116
rect 668762 338104 668768 338116
rect 668820 338104 668826 338156
rect 46290 336744 46296 336796
rect 46348 336784 46354 336796
rect 62114 336784 62120 336796
rect 46348 336756 62120 336784
rect 46348 336744 46354 336756
rect 62114 336744 62120 336756
rect 62172 336744 62178 336796
rect 674466 336540 674472 336592
rect 674524 336580 674530 336592
rect 675478 336580 675484 336592
rect 674524 336552 675484 336580
rect 674524 336540 674530 336552
rect 675478 336540 675484 336552
rect 675536 336540 675542 336592
rect 674834 336268 674840 336320
rect 674892 336308 674898 336320
rect 675386 336308 675392 336320
rect 674892 336280 675392 336308
rect 674892 336268 674898 336280
rect 675386 336268 675392 336280
rect 675444 336268 675450 336320
rect 30374 333208 30380 333260
rect 30432 333248 30438 333260
rect 64138 333248 64144 333260
rect 30432 333220 64144 333248
rect 30432 333208 30438 333220
rect 64138 333208 64144 333220
rect 64196 333208 64202 333260
rect 674558 332596 674564 332648
rect 674616 332636 674622 332648
rect 675386 332636 675392 332648
rect 674616 332608 675392 332636
rect 674616 332596 674622 332608
rect 675386 332596 675392 332608
rect 675444 332596 675450 332648
rect 673086 331576 673092 331628
rect 673144 331616 673150 331628
rect 675386 331616 675392 331628
rect 673144 331588 675392 331616
rect 673144 331576 673150 331588
rect 675386 331576 675392 331588
rect 675444 331576 675450 331628
rect 674834 329468 674840 329520
rect 674892 329508 674898 329520
rect 675386 329508 675392 329520
rect 674892 329480 675392 329508
rect 674892 329468 674898 329480
rect 675386 329468 675392 329480
rect 675444 329468 675450 329520
rect 673178 328380 673184 328432
rect 673236 328420 673242 328432
rect 674834 328420 674840 328432
rect 673236 328392 674840 328420
rect 673236 328380 673242 328392
rect 674834 328380 674840 328392
rect 674892 328380 674898 328432
rect 675110 327632 675116 327684
rect 675168 327672 675174 327684
rect 675478 327672 675484 327684
rect 675168 327644 675484 327672
rect 675168 327632 675174 327644
rect 675478 327632 675484 327644
rect 675536 327632 675542 327684
rect 42058 326748 42064 326800
rect 42116 326788 42122 326800
rect 44174 326788 44180 326800
rect 42116 326760 44180 326788
rect 42116 326748 42122 326760
rect 44174 326748 44180 326760
rect 44232 326748 44238 326800
rect 675754 325796 675760 325848
rect 675812 325796 675818 325848
rect 675772 325644 675800 325796
rect 675754 325592 675760 325644
rect 675812 325592 675818 325644
rect 651558 324300 651564 324352
rect 651616 324340 651622 324352
rect 670234 324340 670240 324352
rect 651616 324312 670240 324340
rect 651616 324300 651622 324312
rect 670234 324300 670240 324312
rect 670292 324300 670298 324352
rect 42150 323280 42156 323332
rect 42208 323320 42214 323332
rect 42610 323320 42616 323332
rect 42208 323292 42616 323320
rect 42208 323280 42214 323292
rect 42610 323280 42616 323292
rect 42668 323280 42674 323332
rect 47670 322940 47676 322992
rect 47728 322980 47734 322992
rect 62114 322980 62120 322992
rect 47728 322952 62120 322980
rect 47728 322940 47734 322952
rect 62114 322940 62120 322952
rect 62172 322940 62178 322992
rect 42058 322872 42064 322924
rect 42116 322912 42122 322924
rect 44358 322912 44364 322924
rect 42116 322884 44364 322912
rect 42116 322872 42122 322884
rect 44358 322872 44364 322884
rect 44416 322872 44422 322924
rect 42610 321512 42616 321564
rect 42668 321552 42674 321564
rect 50430 321552 50436 321564
rect 42668 321524 50436 321552
rect 42668 321512 42674 321524
rect 50430 321512 50436 321524
rect 50488 321512 50494 321564
rect 42150 321444 42156 321496
rect 42208 321484 42214 321496
rect 44450 321484 44456 321496
rect 42208 321456 44456 321484
rect 42208 321444 42214 321456
rect 44450 321444 44456 321456
rect 44508 321444 44514 321496
rect 42150 319948 42156 320000
rect 42208 319988 42214 320000
rect 43070 319988 43076 320000
rect 42208 319960 43076 319988
rect 42208 319948 42214 319960
rect 43070 319948 43076 319960
rect 43128 319948 43134 320000
rect 42150 316684 42156 316736
rect 42208 316724 42214 316736
rect 42978 316724 42984 316736
rect 42208 316696 42984 316724
rect 42208 316684 42214 316696
rect 42978 316684 42984 316696
rect 43036 316684 43042 316736
rect 664530 313488 664536 313540
rect 664588 313528 664594 313540
rect 676214 313528 676220 313540
rect 664588 313500 676220 313528
rect 664588 313488 664594 313500
rect 676214 313488 676220 313500
rect 676272 313488 676278 313540
rect 663150 313352 663156 313404
rect 663208 313392 663214 313404
rect 676030 313392 676036 313404
rect 663208 313364 676036 313392
rect 663208 313352 663214 313364
rect 676030 313352 676036 313364
rect 676088 313352 676094 313404
rect 673270 312128 673276 312180
rect 673328 312168 673334 312180
rect 676214 312168 676220 312180
rect 673328 312140 676220 312168
rect 673328 312128 673334 312140
rect 676214 312128 676220 312140
rect 676272 312128 676278 312180
rect 659010 311992 659016 312044
rect 659068 312032 659074 312044
rect 676122 312032 676128 312044
rect 659068 312004 676128 312032
rect 659068 311992 659074 312004
rect 676122 311992 676128 312004
rect 676180 311992 676186 312044
rect 673362 311856 673368 311908
rect 673420 311896 673426 311908
rect 676214 311896 676220 311908
rect 673420 311868 676220 311896
rect 673420 311856 673426 311868
rect 676214 311856 676220 311868
rect 676272 311856 676278 311908
rect 672994 310632 673000 310684
rect 673052 310672 673058 310684
rect 676214 310672 676220 310684
rect 673052 310644 676220 310672
rect 673052 310632 673058 310644
rect 676214 310632 676220 310644
rect 676272 310632 676278 310684
rect 651558 310564 651564 310616
rect 651616 310604 651622 310616
rect 674098 310604 674104 310616
rect 651616 310576 674104 310604
rect 651616 310564 651622 310576
rect 674098 310564 674104 310576
rect 674156 310564 674162 310616
rect 46198 310496 46204 310548
rect 46256 310536 46262 310548
rect 62114 310536 62120 310548
rect 46256 310508 62120 310536
rect 46256 310496 46262 310508
rect 62114 310496 62120 310508
rect 62172 310496 62178 310548
rect 673270 310496 673276 310548
rect 673328 310536 673334 310548
rect 676122 310536 676128 310548
rect 673328 310508 676128 310536
rect 673328 310496 673334 310508
rect 676122 310496 676128 310508
rect 676180 310496 676186 310548
rect 674742 310224 674748 310276
rect 674800 310264 674806 310276
rect 676214 310264 676220 310276
rect 674800 310236 676220 310264
rect 674800 310224 674806 310236
rect 676214 310224 676220 310236
rect 676272 310224 676278 310276
rect 674650 310020 674656 310072
rect 674708 310060 674714 310072
rect 676030 310060 676036 310072
rect 674708 310032 676036 310060
rect 674708 310020 674714 310032
rect 676030 310020 676036 310032
rect 676088 310020 676094 310072
rect 674742 309408 674748 309460
rect 674800 309448 674806 309460
rect 676214 309448 676220 309460
rect 674800 309420 676220 309448
rect 674800 309408 674806 309420
rect 676214 309408 676220 309420
rect 676272 309408 676278 309460
rect 673178 303764 673184 303816
rect 673236 303804 673242 303816
rect 676214 303804 676220 303816
rect 673236 303776 676220 303804
rect 673236 303764 673242 303776
rect 676214 303764 676220 303776
rect 676272 303764 676278 303816
rect 673086 303696 673092 303748
rect 673144 303736 673150 303748
rect 676122 303736 676128 303748
rect 673144 303708 676128 303736
rect 673144 303696 673150 303708
rect 676122 303696 676128 303708
rect 676180 303696 676186 303748
rect 672994 303628 673000 303680
rect 673052 303668 673058 303680
rect 676306 303668 676312 303680
rect 673052 303640 676312 303668
rect 673052 303628 673058 303640
rect 676306 303628 676312 303640
rect 676364 303628 676370 303680
rect 674374 302200 674380 302252
rect 674432 302240 674438 302252
rect 683114 302240 683120 302252
rect 674432 302212 683120 302240
rect 674432 302200 674438 302212
rect 683114 302200 683120 302212
rect 683172 302200 683178 302252
rect 35802 301044 35808 301096
rect 35860 301084 35866 301096
rect 35860 301044 35894 301084
rect 35866 301016 35894 301044
rect 49050 301016 49056 301028
rect 35866 300988 49056 301016
rect 49050 300976 49056 300988
rect 49108 300976 49114 301028
rect 35802 300908 35808 300960
rect 35860 300948 35866 300960
rect 56042 300948 56048 300960
rect 35860 300920 56048 300948
rect 35860 300908 35866 300920
rect 56042 300908 56048 300920
rect 56100 300908 56106 300960
rect 43714 298120 43720 298172
rect 43772 298160 43778 298172
rect 62114 298160 62120 298172
rect 43772 298132 62120 298160
rect 43772 298120 43778 298132
rect 62114 298120 62120 298132
rect 62172 298120 62178 298172
rect 675202 298052 675208 298104
rect 675260 298092 675266 298104
rect 676858 298092 676864 298104
rect 675260 298064 676864 298092
rect 675260 298052 675266 298064
rect 676858 298052 676864 298064
rect 676916 298052 676922 298104
rect 675754 297984 675760 298036
rect 675812 298024 675818 298036
rect 678238 298024 678244 298036
rect 675812 297996 678244 298024
rect 675812 297984 675818 297996
rect 678238 297984 678244 297996
rect 678296 297984 678302 298036
rect 675110 297372 675116 297424
rect 675168 297412 675174 297424
rect 676490 297412 676496 297424
rect 675168 297384 676496 297412
rect 675168 297372 675174 297384
rect 676490 297372 676496 297384
rect 676548 297372 676554 297424
rect 675754 296148 675760 296200
rect 675812 296148 675818 296200
rect 675772 295996 675800 296148
rect 675754 295944 675760 295996
rect 675812 295944 675818 295996
rect 675202 295400 675208 295452
rect 675260 295440 675266 295452
rect 675386 295440 675392 295452
rect 675260 295412 675392 295440
rect 675260 295400 675266 295412
rect 675386 295400 675392 295412
rect 675444 295400 675450 295452
rect 675110 294080 675116 294092
rect 675036 294052 675116 294080
rect 675036 294024 675064 294052
rect 675110 294040 675116 294052
rect 675168 294040 675174 294092
rect 675018 293972 675024 294024
rect 675076 293972 675082 294024
rect 675018 291728 675024 291780
rect 675076 291768 675082 291780
rect 675386 291768 675392 291780
rect 675076 291740 675392 291768
rect 675076 291728 675082 291740
rect 675386 291728 675392 291740
rect 675444 291728 675450 291780
rect 672994 291048 673000 291100
rect 673052 291088 673058 291100
rect 675386 291088 675392 291100
rect 673052 291060 675392 291088
rect 673052 291048 673058 291060
rect 675386 291048 675392 291060
rect 675444 291048 675450 291100
rect 673086 287920 673092 287972
rect 673144 287960 673150 287972
rect 675386 287960 675392 287972
rect 673144 287932 675392 287960
rect 673144 287920 673150 287932
rect 675386 287920 675392 287932
rect 675444 287920 675450 287972
rect 673178 286560 673184 286612
rect 673236 286600 673242 286612
rect 675386 286600 675392 286612
rect 673236 286572 675392 286600
rect 673236 286560 673242 286572
rect 675386 286560 675392 286572
rect 675444 286560 675450 286612
rect 32398 284928 32404 284980
rect 32456 284968 32462 284980
rect 41874 284968 41880 284980
rect 32456 284940 41880 284968
rect 32456 284928 32462 284940
rect 41874 284928 41880 284940
rect 41932 284928 41938 284980
rect 43806 284316 43812 284368
rect 43864 284356 43870 284368
rect 62114 284356 62120 284368
rect 43864 284328 62120 284356
rect 43864 284316 43870 284328
rect 62114 284316 62120 284328
rect 62172 284316 62178 284368
rect 651558 284316 651564 284368
rect 651616 284356 651622 284368
rect 672810 284356 672816 284368
rect 651616 284328 672816 284356
rect 651616 284316 651622 284328
rect 672810 284316 672816 284328
rect 672868 284316 672874 284368
rect 41874 283772 41880 283824
rect 41932 283772 41938 283824
rect 41892 283620 41920 283772
rect 41874 283568 41880 283620
rect 41932 283568 41938 283620
rect 42150 280168 42156 280220
rect 42208 280208 42214 280220
rect 47578 280208 47584 280220
rect 42208 280180 47584 280208
rect 42208 280168 42214 280180
rect 47578 280168 47584 280180
rect 47636 280168 47642 280220
rect 42058 278604 42064 278656
rect 42116 278644 42122 278656
rect 44542 278644 44548 278656
rect 42116 278616 44548 278644
rect 42116 278604 42122 278616
rect 44542 278604 44548 278616
rect 44600 278604 44606 278656
rect 43438 278196 43444 278248
rect 43496 278236 43502 278248
rect 646038 278236 646044 278248
rect 43496 278208 646044 278236
rect 43496 278196 43502 278208
rect 646038 278196 646044 278208
rect 646096 278196 646102 278248
rect 53190 278128 53196 278180
rect 53248 278168 53254 278180
rect 656894 278168 656900 278180
rect 53248 278140 656900 278168
rect 53248 278128 53254 278140
rect 656894 278128 656900 278140
rect 656952 278128 656958 278180
rect 51810 278060 51816 278112
rect 51868 278100 51874 278112
rect 662414 278100 662420 278112
rect 51868 278072 662420 278100
rect 51868 278060 51874 278072
rect 662414 278060 662420 278072
rect 662472 278060 662478 278112
rect 43622 277992 43628 278044
rect 43680 278032 43686 278044
rect 658274 278032 658280 278044
rect 43680 278004 658280 278032
rect 43680 277992 43686 278004
rect 658274 277992 658280 278004
rect 658332 277992 658338 278044
rect 332502 277924 332508 277976
rect 332560 277964 332566 277976
rect 436646 277964 436652 277976
rect 332560 277936 436652 277964
rect 332560 277924 332566 277936
rect 436646 277924 436652 277936
rect 436704 277924 436710 277976
rect 333882 277856 333888 277908
rect 333940 277896 333946 277908
rect 440326 277896 440332 277908
rect 333940 277868 440332 277896
rect 333940 277856 333946 277868
rect 440326 277856 440332 277868
rect 440384 277856 440390 277908
rect 335078 277788 335084 277840
rect 335136 277828 335142 277840
rect 443822 277828 443828 277840
rect 335136 277800 443828 277828
rect 335136 277788 335142 277800
rect 443822 277788 443828 277800
rect 443880 277788 443886 277840
rect 336366 277720 336372 277772
rect 336424 277760 336430 277772
rect 447318 277760 447324 277772
rect 336424 277732 447324 277760
rect 336424 277720 336430 277732
rect 447318 277720 447324 277732
rect 447376 277720 447382 277772
rect 338022 277652 338028 277704
rect 338080 277692 338086 277704
rect 452470 277692 452476 277704
rect 338080 277664 452476 277692
rect 338080 277652 338086 277664
rect 452470 277652 452476 277664
rect 452528 277652 452534 277704
rect 339218 277584 339224 277636
rect 339276 277624 339282 277636
rect 454770 277624 454776 277636
rect 339276 277596 454776 277624
rect 339276 277584 339282 277596
rect 454770 277584 454776 277596
rect 454828 277584 454834 277636
rect 360102 277516 360108 277568
rect 360160 277556 360166 277568
rect 507946 277556 507952 277568
rect 360160 277528 507952 277556
rect 360160 277516 360166 277528
rect 507946 277516 507952 277528
rect 508004 277516 508010 277568
rect 391658 277448 391664 277500
rect 391716 277488 391722 277500
rect 594334 277488 594340 277500
rect 391716 277460 594340 277488
rect 391716 277448 391722 277460
rect 594334 277448 594340 277460
rect 594392 277448 594398 277500
rect 398742 277380 398748 277432
rect 398800 277420 398806 277432
rect 611998 277420 612004 277432
rect 398800 277392 612004 277420
rect 398800 277380 398806 277392
rect 611998 277380 612004 277392
rect 612056 277380 612062 277432
rect 353202 277312 353208 277364
rect 353260 277352 353266 277364
rect 492582 277352 492588 277364
rect 353260 277324 492588 277352
rect 353260 277312 353266 277324
rect 492582 277312 492588 277324
rect 492640 277312 492646 277364
rect 355962 277244 355968 277296
rect 356020 277284 356026 277296
rect 499758 277284 499764 277296
rect 356020 277256 499764 277284
rect 356020 277244 356026 277256
rect 499758 277244 499764 277256
rect 499816 277244 499822 277296
rect 358722 277176 358728 277228
rect 358780 277216 358786 277228
rect 506842 277216 506848 277228
rect 358780 277188 506848 277216
rect 358780 277176 358786 277188
rect 506842 277176 506848 277188
rect 506900 277176 506906 277228
rect 42150 277108 42156 277160
rect 42208 277148 42214 277160
rect 43162 277148 43168 277160
rect 42208 277120 43168 277148
rect 42208 277108 42214 277120
rect 43162 277108 43168 277120
rect 43220 277108 43226 277160
rect 380802 277108 380808 277160
rect 380860 277148 380866 277160
rect 563514 277148 563520 277160
rect 380860 277120 563520 277148
rect 380860 277108 380866 277120
rect 563514 277108 563520 277120
rect 563572 277108 563578 277160
rect 383470 277040 383476 277092
rect 383528 277080 383534 277092
rect 570690 277080 570696 277092
rect 383528 277052 570696 277080
rect 383528 277040 383534 277052
rect 570690 277040 570696 277052
rect 570748 277040 570754 277092
rect 383562 276972 383568 277024
rect 383620 277012 383626 277024
rect 571794 277012 571800 277024
rect 383620 276984 571800 277012
rect 383620 276972 383626 276984
rect 571794 276972 571800 276984
rect 571852 276972 571858 277024
rect 387242 276904 387248 276956
rect 387300 276944 387306 276956
rect 582466 276944 582472 276956
rect 387300 276916 582472 276944
rect 387300 276904 387306 276916
rect 582466 276904 582472 276916
rect 582524 276904 582530 276956
rect 389910 276836 389916 276888
rect 389968 276876 389974 276888
rect 589550 276876 589556 276888
rect 389968 276848 589556 276876
rect 389968 276836 389974 276848
rect 589550 276836 589556 276848
rect 589608 276836 589614 276888
rect 403894 276768 403900 276820
rect 403952 276808 403958 276820
rect 627362 276808 627368 276820
rect 403952 276780 627368 276808
rect 403952 276768 403958 276780
rect 627362 276768 627368 276780
rect 627420 276768 627426 276820
rect 42058 276700 42064 276752
rect 42116 276740 42122 276752
rect 42886 276740 42892 276752
rect 42116 276712 42892 276740
rect 42116 276700 42122 276712
rect 42886 276700 42892 276712
rect 42944 276700 42950 276752
rect 406654 276700 406660 276752
rect 406712 276740 406718 276752
rect 634446 276740 634452 276752
rect 406712 276712 634452 276740
rect 406712 276700 406718 276712
rect 634446 276700 634452 276712
rect 634504 276700 634510 276752
rect 409782 276632 409788 276684
rect 409840 276672 409846 276684
rect 641622 276672 641628 276684
rect 409840 276644 641628 276672
rect 409840 276632 409846 276644
rect 641622 276632 641628 276644
rect 641680 276632 641686 276684
rect 350442 276564 350448 276616
rect 350500 276604 350506 276616
rect 485498 276604 485504 276616
rect 350500 276576 485504 276604
rect 350500 276564 350506 276576
rect 485498 276564 485504 276576
rect 485556 276564 485562 276616
rect 349062 276496 349068 276548
rect 349120 276536 349126 276548
rect 478414 276536 478420 276548
rect 349120 276508 478420 276536
rect 349120 276496 349126 276508
rect 478414 276496 478420 276508
rect 478472 276496 478478 276548
rect 332410 276428 332416 276480
rect 332468 276468 332474 276480
rect 435910 276468 435916 276480
rect 332468 276440 435916 276468
rect 332468 276428 332474 276440
rect 435910 276428 435916 276440
rect 435968 276428 435974 276480
rect 329742 276360 329748 276412
rect 329800 276400 329806 276412
rect 428826 276400 428832 276412
rect 329800 276372 428832 276400
rect 329800 276360 329806 276372
rect 428826 276360 428832 276372
rect 428884 276360 428890 276412
rect 326706 276292 326712 276344
rect 326764 276332 326770 276344
rect 421650 276332 421656 276344
rect 326764 276304 421656 276332
rect 326764 276292 326770 276304
rect 421650 276292 421656 276304
rect 421708 276292 421714 276344
rect 324038 276224 324044 276276
rect 324096 276264 324102 276276
rect 414566 276264 414572 276276
rect 324096 276236 414572 276264
rect 324096 276224 324102 276236
rect 414566 276224 414572 276236
rect 414624 276224 414630 276276
rect 492646 276032 502334 276060
rect 146202 275952 146208 276004
rect 146260 275992 146266 276004
rect 195974 275992 195980 276004
rect 146260 275964 195980 275992
rect 146260 275952 146266 275964
rect 195974 275952 195980 275964
rect 196032 275952 196038 276004
rect 348970 275952 348976 276004
rect 349028 275992 349034 276004
rect 480806 275992 480812 276004
rect 349028 275964 480812 275992
rect 349028 275952 349034 275964
rect 480806 275952 480812 275964
rect 480864 275952 480870 276004
rect 487154 275952 487160 276004
rect 487212 275992 487218 276004
rect 487212 275964 489914 275992
rect 487212 275952 487218 275964
rect 163958 275884 163964 275936
rect 164016 275924 164022 275936
rect 216674 275924 216680 275936
rect 164016 275896 216680 275924
rect 164016 275884 164022 275896
rect 216674 275884 216680 275896
rect 216732 275884 216738 275936
rect 351822 275884 351828 275936
rect 351880 275924 351886 275936
rect 487890 275924 487896 275936
rect 351880 275896 487896 275924
rect 351880 275884 351886 275896
rect 487890 275884 487896 275896
rect 487948 275884 487954 275936
rect 489886 275924 489914 275964
rect 492646 275924 492674 276032
rect 489886 275896 492674 275924
rect 502306 275924 502334 276032
rect 583754 275952 583760 276004
rect 583812 275992 583818 276004
rect 600222 275992 600228 276004
rect 583812 275964 600228 275992
rect 583812 275952 583818 275964
rect 600222 275952 600228 275964
rect 600280 275952 600286 276004
rect 581270 275924 581276 275936
rect 502306 275896 581276 275924
rect 581270 275884 581276 275896
rect 581328 275884 581334 275936
rect 171042 275816 171048 275868
rect 171100 275856 171106 275868
rect 226978 275856 226984 275868
rect 171100 275828 226984 275856
rect 171100 275816 171106 275828
rect 226978 275816 226984 275828
rect 227036 275816 227042 275868
rect 354398 275816 354404 275868
rect 354456 275856 354462 275868
rect 494974 275856 494980 275868
rect 354456 275828 494980 275856
rect 354456 275816 354462 275828
rect 494974 275816 494980 275828
rect 495032 275816 495038 275868
rect 496722 275816 496728 275868
rect 496780 275856 496786 275868
rect 513926 275856 513932 275868
rect 496780 275828 513932 275856
rect 496780 275816 496786 275828
rect 513926 275816 513932 275828
rect 513984 275816 513990 275868
rect 581638 275816 581644 275868
rect 581696 275856 581702 275868
rect 599026 275856 599032 275868
rect 581696 275828 599032 275856
rect 581696 275816 581702 275828
rect 599026 275816 599032 275828
rect 599084 275816 599090 275868
rect 149790 275748 149796 275800
rect 149848 275788 149854 275800
rect 220630 275788 220636 275800
rect 149848 275760 220636 275788
rect 149848 275748 149854 275760
rect 220630 275748 220636 275760
rect 220688 275748 220694 275800
rect 258534 275748 258540 275800
rect 258592 275788 258598 275800
rect 264606 275788 264612 275800
rect 258592 275760 264612 275788
rect 258592 275748 258598 275760
rect 264606 275748 264612 275760
rect 264664 275748 264670 275800
rect 357342 275748 357348 275800
rect 357400 275788 357406 275800
rect 502058 275788 502064 275800
rect 357400 275760 502064 275788
rect 357400 275748 357406 275760
rect 502058 275748 502064 275760
rect 502116 275748 502122 275800
rect 502242 275748 502248 275800
rect 502300 275788 502306 275800
rect 584858 275788 584864 275800
rect 502300 275760 584864 275788
rect 502300 275748 502306 275760
rect 584858 275748 584864 275760
rect 584916 275748 584922 275800
rect 107194 275680 107200 275732
rect 107252 275720 107258 275732
rect 208302 275720 208308 275732
rect 107252 275692 208308 275720
rect 107252 275680 107258 275692
rect 208302 275680 208308 275692
rect 208360 275680 208366 275732
rect 214834 275680 214840 275732
rect 214892 275720 214898 275732
rect 227714 275720 227720 275732
rect 214892 275692 227720 275720
rect 214892 275680 214898 275692
rect 227714 275680 227720 275692
rect 227772 275680 227778 275732
rect 251450 275680 251456 275732
rect 251508 275720 251514 275732
rect 252370 275720 252376 275732
rect 251508 275692 252376 275720
rect 251508 275680 251514 275692
rect 252370 275680 252376 275692
rect 252428 275680 252434 275732
rect 362218 275680 362224 275732
rect 362276 275720 362282 275732
rect 509142 275720 509148 275732
rect 362276 275692 509148 275720
rect 362276 275680 362282 275692
rect 509142 275680 509148 275692
rect 509200 275680 509206 275732
rect 513466 275680 513472 275732
rect 513524 275720 513530 275732
rect 593138 275720 593144 275732
rect 513524 275692 593144 275720
rect 513524 275680 513530 275692
rect 593138 275680 593144 275692
rect 593196 275680 593202 275732
rect 100110 275612 100116 275664
rect 100168 275652 100174 275664
rect 205818 275652 205824 275664
rect 100168 275624 205824 275652
rect 100168 275612 100174 275624
rect 205818 275612 205824 275624
rect 205876 275612 205882 275664
rect 207750 275612 207756 275664
rect 207808 275652 207814 275664
rect 213454 275652 213460 275664
rect 207808 275624 213460 275652
rect 207808 275612 207814 275624
rect 213454 275612 213460 275624
rect 213512 275612 213518 275664
rect 223114 275612 223120 275664
rect 223172 275652 223178 275664
rect 241422 275652 241428 275664
rect 223172 275624 241428 275652
rect 223172 275612 223178 275624
rect 241422 275612 241428 275624
rect 241480 275612 241486 275664
rect 363506 275612 363512 275664
rect 363564 275652 363570 275664
rect 516226 275652 516232 275664
rect 363564 275624 516232 275652
rect 363564 275612 363570 275624
rect 516226 275612 516232 275624
rect 516284 275612 516290 275664
rect 521562 275612 521568 275664
rect 521620 275652 521626 275664
rect 596634 275652 596640 275664
rect 521620 275624 596640 275652
rect 521620 275612 521626 275624
rect 596634 275612 596640 275624
rect 596692 275612 596698 275664
rect 597830 275612 597836 275664
rect 597888 275652 597894 275664
rect 610802 275652 610808 275664
rect 597888 275624 610808 275652
rect 597888 275612 597894 275624
rect 610802 275612 610808 275624
rect 610860 275612 610866 275664
rect 90634 275544 90640 275596
rect 90692 275584 90698 275596
rect 201678 275584 201684 275596
rect 90692 275556 201684 275584
rect 90692 275544 90698 275556
rect 201678 275544 201684 275556
rect 201736 275544 201742 275596
rect 212442 275544 212448 275596
rect 212500 275584 212506 275596
rect 222470 275584 222476 275596
rect 212500 275556 222476 275584
rect 212500 275544 212506 275556
rect 222470 275544 222476 275556
rect 222528 275544 222534 275596
rect 224218 275544 224224 275596
rect 224276 275584 224282 275596
rect 243538 275584 243544 275596
rect 224276 275556 243544 275584
rect 224276 275544 224282 275556
rect 243538 275544 243544 275556
rect 243596 275544 243602 275596
rect 367002 275544 367008 275596
rect 367060 275584 367066 275596
rect 523402 275584 523408 275596
rect 367060 275556 523408 275584
rect 367060 275544 367066 275556
rect 523402 275544 523408 275556
rect 523460 275544 523466 275596
rect 523678 275544 523684 275596
rect 523736 275584 523742 275596
rect 591942 275584 591948 275596
rect 523736 275556 591948 275584
rect 523736 275544 523742 275556
rect 591942 275544 591948 275556
rect 592000 275544 592006 275596
rect 593414 275544 593420 275596
rect 593472 275584 593478 275596
rect 607306 275584 607312 275596
rect 593472 275556 607312 275584
rect 593472 275544 593478 275556
rect 607306 275544 607312 275556
rect 607364 275544 607370 275596
rect 83550 275476 83556 275528
rect 83608 275516 83614 275528
rect 199102 275516 199108 275528
rect 83608 275488 199108 275516
rect 83608 275476 83614 275488
rect 199102 275476 199108 275488
rect 199160 275476 199166 275528
rect 210050 275476 210056 275528
rect 210108 275516 210114 275528
rect 224954 275516 224960 275528
rect 210108 275488 224960 275516
rect 210108 275476 210114 275488
rect 224954 275476 224960 275488
rect 225012 275476 225018 275528
rect 227806 275476 227812 275528
rect 227864 275516 227870 275528
rect 249610 275516 249616 275528
rect 227864 275488 249616 275516
rect 227864 275476 227870 275488
rect 249610 275476 249616 275488
rect 249668 275476 249674 275528
rect 368382 275476 368388 275528
rect 368440 275516 368446 275528
rect 530486 275516 530492 275528
rect 368440 275488 530492 275516
rect 368440 275476 368446 275488
rect 530486 275476 530492 275488
rect 530544 275476 530550 275528
rect 543734 275476 543740 275528
rect 543792 275516 543798 275528
rect 595438 275516 595444 275528
rect 543792 275488 595444 275516
rect 543792 275476 543798 275488
rect 595438 275476 595444 275488
rect 595496 275476 595502 275528
rect 600038 275476 600044 275528
rect 600096 275516 600102 275528
rect 614390 275516 614396 275528
rect 600096 275488 614396 275516
rect 600096 275476 600102 275488
rect 614390 275476 614396 275488
rect 614448 275476 614454 275528
rect 81250 275408 81256 275460
rect 81308 275448 81314 275460
rect 197814 275448 197820 275460
rect 81308 275420 197820 275448
rect 81308 275408 81314 275420
rect 197814 275408 197820 275420
rect 197872 275408 197878 275460
rect 213638 275408 213644 275460
rect 213696 275448 213702 275460
rect 234614 275448 234620 275460
rect 213696 275420 234620 275448
rect 213696 275408 213702 275420
rect 234614 275408 234620 275420
rect 234672 275408 234678 275460
rect 239582 275408 239588 275460
rect 239640 275448 239646 275460
rect 249702 275448 249708 275460
rect 239640 275420 249708 275448
rect 239640 275408 239646 275420
rect 249702 275408 249708 275420
rect 249760 275408 249766 275460
rect 340598 275408 340604 275460
rect 340656 275448 340662 275460
rect 459554 275448 459560 275460
rect 340656 275420 459560 275448
rect 340656 275408 340662 275420
rect 459554 275408 459560 275420
rect 459612 275408 459618 275460
rect 459646 275408 459652 275460
rect 459704 275448 459710 275460
rect 626166 275448 626172 275460
rect 459704 275420 626172 275448
rect 459704 275408 459710 275420
rect 626166 275408 626172 275420
rect 626224 275408 626230 275460
rect 66990 275340 66996 275392
rect 67048 275380 67054 275392
rect 187694 275380 187700 275392
rect 67048 275352 187700 275380
rect 67048 275340 67054 275352
rect 187694 275340 187700 275352
rect 187752 275340 187758 275392
rect 208854 275340 208860 275392
rect 208912 275380 208918 275392
rect 233878 275380 233884 275392
rect 208912 275352 233884 275380
rect 208912 275340 208918 275352
rect 233878 275340 233884 275352
rect 233936 275340 233942 275392
rect 249058 275340 249064 275392
rect 249116 275380 249122 275392
rect 260742 275380 260748 275392
rect 249116 275352 260748 275380
rect 249116 275340 249122 275352
rect 260742 275340 260748 275352
rect 260800 275340 260806 275392
rect 336642 275340 336648 275392
rect 336700 275380 336706 275392
rect 448882 275380 448888 275392
rect 336700 275352 448888 275380
rect 336700 275340 336706 275352
rect 448882 275340 448888 275352
rect 448940 275340 448946 275392
rect 448974 275340 448980 275392
rect 449032 275380 449038 275392
rect 633342 275380 633348 275392
rect 449032 275352 633348 275380
rect 449032 275340 449038 275352
rect 633342 275340 633348 275352
rect 633400 275340 633406 275392
rect 71774 275272 71780 275324
rect 71832 275312 71838 275324
rect 194870 275312 194876 275324
rect 71832 275284 194876 275312
rect 71832 275272 71838 275284
rect 194870 275272 194876 275284
rect 194928 275272 194934 275324
rect 206554 275272 206560 275324
rect 206612 275312 206618 275324
rect 237374 275312 237380 275324
rect 206612 275284 237380 275312
rect 206612 275272 206618 275284
rect 237374 275272 237380 275284
rect 237432 275272 237438 275324
rect 240778 275272 240784 275324
rect 240836 275312 240842 275324
rect 258258 275312 258264 275324
rect 240836 275284 258264 275312
rect 240836 275272 240842 275284
rect 258258 275272 258264 275284
rect 258316 275272 258322 275324
rect 263226 275272 263232 275324
rect 263284 275312 263290 275324
rect 266538 275312 266544 275324
rect 263284 275284 266544 275312
rect 263284 275272 263290 275284
rect 266538 275272 266544 275284
rect 266596 275272 266602 275324
rect 388162 275272 388168 275324
rect 388220 275312 388226 275324
rect 402790 275312 402796 275324
rect 388220 275284 402796 275312
rect 388220 275272 388226 275284
rect 402790 275272 402796 275284
rect 402848 275272 402854 275324
rect 412542 275272 412548 275324
rect 412600 275312 412606 275324
rect 647510 275312 647516 275324
rect 412600 275284 647516 275312
rect 412600 275272 412606 275284
rect 647510 275272 647516 275284
rect 647568 275272 647574 275324
rect 128538 275204 128544 275256
rect 128596 275244 128602 275256
rect 131114 275244 131120 275256
rect 128596 275216 131120 275244
rect 128596 275204 128602 275216
rect 131114 275204 131120 275216
rect 131172 275204 131178 275256
rect 156874 275204 156880 275256
rect 156932 275244 156938 275256
rect 204898 275244 204904 275256
rect 156932 275216 204904 275244
rect 156932 275204 156938 275216
rect 204898 275204 204904 275216
rect 204956 275204 204962 275256
rect 234890 275204 234896 275256
rect 234948 275244 234954 275256
rect 235902 275244 235908 275256
rect 234948 275216 235908 275244
rect 234948 275204 234954 275216
rect 235902 275204 235908 275216
rect 235960 275204 235966 275256
rect 259730 275204 259736 275256
rect 259788 275244 259794 275256
rect 264974 275244 264980 275256
rect 259788 275216 264980 275244
rect 259788 275204 259794 275216
rect 264974 275204 264980 275216
rect 265032 275204 265038 275256
rect 346118 275204 346124 275256
rect 346176 275244 346182 275256
rect 473722 275244 473728 275256
rect 346176 275216 473728 275244
rect 346176 275204 346182 275216
rect 473722 275204 473728 275216
rect 473780 275204 473786 275256
rect 474182 275204 474188 275256
rect 474240 275244 474246 275256
rect 577774 275244 577780 275256
rect 474240 275216 577780 275244
rect 474240 275204 474246 275216
rect 577774 275204 577780 275216
rect 577832 275204 577838 275256
rect 139118 275136 139124 275188
rect 139176 275176 139182 275188
rect 185026 275176 185032 275188
rect 139176 275148 185032 275176
rect 139176 275136 139182 275148
rect 185026 275136 185032 275148
rect 185084 275136 185090 275188
rect 188798 275136 188804 275188
rect 188856 275176 188862 275188
rect 210418 275176 210424 275188
rect 188856 275148 210424 275176
rect 188856 275136 188862 275148
rect 210418 275136 210424 275148
rect 210476 275136 210482 275188
rect 343358 275136 343364 275188
rect 343416 275176 343422 275188
rect 466638 275176 466644 275188
rect 343416 275148 466644 275176
rect 343416 275136 343422 275148
rect 466638 275136 466644 275148
rect 466696 275136 466702 275188
rect 466730 275136 466736 275188
rect 466788 275176 466794 275188
rect 510338 275176 510344 275188
rect 466788 275148 510344 275176
rect 466788 275136 466794 275148
rect 510338 275136 510344 275148
rect 510396 275136 510402 275188
rect 178126 275068 178132 275120
rect 178184 275108 178190 275120
rect 221458 275108 221464 275120
rect 178184 275080 221464 275108
rect 178184 275068 178190 275080
rect 221458 275068 221464 275080
rect 221516 275068 221522 275120
rect 335170 275068 335176 275120
rect 335228 275108 335234 275120
rect 441798 275108 441804 275120
rect 335228 275080 441804 275108
rect 335228 275068 335234 275080
rect 441798 275068 441804 275080
rect 441856 275068 441862 275120
rect 185210 275000 185216 275052
rect 185268 275040 185274 275052
rect 214558 275040 214564 275052
rect 185268 275012 214564 275040
rect 185268 275000 185274 275012
rect 214558 275000 214564 275012
rect 214616 275000 214622 275052
rect 329650 275000 329656 275052
rect 329708 275040 329714 275052
rect 427630 275040 427636 275052
rect 329708 275012 427636 275040
rect 329708 275000 329714 275012
rect 427630 275000 427636 275012
rect 427688 275000 427694 275052
rect 427722 275000 427728 275052
rect 427780 275040 427786 275052
rect 458358 275040 458364 275052
rect 427780 275012 458364 275040
rect 427780 275000 427786 275012
rect 458358 275000 458364 275012
rect 458416 275000 458422 275052
rect 260926 274932 260932 274984
rect 260984 274972 260990 274984
rect 265066 274972 265072 274984
rect 260984 274944 265072 274972
rect 260984 274932 260990 274944
rect 265066 274932 265072 274944
rect 265124 274932 265130 274984
rect 375190 274932 375196 274984
rect 375248 274972 375254 274984
rect 434714 274972 434720 274984
rect 375248 274944 434720 274972
rect 375248 274932 375254 274944
rect 434714 274932 434720 274944
rect 434772 274932 434778 274984
rect 401778 274864 401784 274916
rect 401836 274904 401842 274916
rect 407482 274904 407488 274916
rect 401836 274876 407488 274904
rect 401836 274864 401842 274876
rect 407482 274864 407488 274876
rect 407540 274864 407546 274916
rect 409966 274864 409972 274916
rect 410024 274904 410030 274916
rect 419350 274904 419356 274916
rect 410024 274876 419356 274904
rect 410024 274864 410030 274876
rect 419350 274864 419356 274876
rect 419408 274864 419414 274916
rect 243170 274796 243176 274848
rect 243228 274836 243234 274848
rect 245838 274836 245844 274848
rect 243228 274808 245844 274836
rect 243228 274796 243234 274808
rect 245838 274796 245844 274808
rect 245896 274796 245902 274848
rect 250254 274796 250260 274848
rect 250312 274836 250318 274848
rect 254210 274836 254216 274848
rect 250312 274808 254216 274836
rect 250312 274796 250318 274808
rect 254210 274796 254216 274808
rect 254268 274796 254274 274848
rect 407022 274796 407028 274848
rect 407080 274836 407086 274848
rect 411070 274836 411076 274848
rect 407080 274808 411076 274836
rect 407080 274796 407086 274808
rect 411070 274796 411076 274808
rect 411128 274796 411134 274848
rect 458174 274796 458180 274848
rect 458232 274836 458238 274848
rect 461854 274836 461860 274848
rect 458232 274808 461860 274836
rect 458232 274796 458238 274808
rect 461854 274796 461860 274808
rect 461912 274796 461918 274848
rect 262122 274728 262128 274780
rect 262180 274768 262186 274780
rect 265894 274768 265900 274780
rect 262180 274740 265900 274768
rect 262180 274728 262186 274740
rect 265894 274728 265900 274740
rect 265952 274728 265958 274780
rect 401594 274728 401600 274780
rect 401652 274768 401658 274780
rect 406286 274768 406292 274780
rect 401652 274740 406292 274768
rect 401652 274728 401658 274740
rect 406286 274728 406292 274740
rect 406344 274728 406350 274780
rect 408586 274728 408592 274780
rect 408644 274768 408650 274780
rect 412266 274768 412272 274780
rect 408644 274740 412272 274768
rect 408644 274728 408650 274740
rect 412266 274728 412272 274740
rect 412324 274728 412330 274780
rect 516134 274728 516140 274780
rect 516192 274768 516198 274780
rect 516192 274740 518894 274768
rect 516192 274728 516198 274740
rect 74074 274660 74080 274712
rect 74132 274700 74138 274712
rect 76006 274700 76012 274712
rect 74132 274672 76012 274700
rect 74132 274660 74138 274672
rect 76006 274660 76012 274672
rect 76064 274660 76070 274712
rect 88334 274660 88340 274712
rect 88392 274700 88398 274712
rect 93118 274700 93124 274712
rect 88392 274672 93124 274700
rect 88392 274660 88398 274672
rect 93118 274660 93124 274672
rect 93176 274660 93182 274712
rect 160462 274660 160468 274712
rect 160520 274700 160526 274712
rect 161382 274700 161388 274712
rect 160520 274672 161388 274700
rect 160520 274660 160526 274672
rect 161382 274660 161388 274672
rect 161440 274660 161446 274712
rect 220722 274660 220728 274712
rect 220780 274700 220786 274712
rect 223574 274700 223580 274712
rect 220780 274672 223580 274700
rect 220780 274660 220786 274672
rect 223574 274660 223580 274672
rect 223632 274660 223638 274712
rect 225414 274660 225420 274712
rect 225472 274700 225478 274712
rect 229830 274700 229836 274712
rect 225472 274672 229836 274700
rect 225472 274660 225478 274672
rect 229830 274660 229836 274672
rect 229888 274660 229894 274712
rect 264422 274660 264428 274712
rect 264480 274700 264486 274712
rect 266722 274700 266728 274712
rect 264480 274672 266728 274700
rect 264480 274660 264486 274672
rect 266722 274660 266728 274672
rect 266780 274660 266786 274712
rect 266814 274660 266820 274712
rect 266872 274700 266878 274712
rect 267734 274700 267740 274712
rect 266872 274672 267740 274700
rect 266872 274660 266878 274672
rect 267734 274660 267740 274672
rect 267792 274660 267798 274712
rect 398834 274660 398840 274712
rect 398892 274700 398898 274712
rect 403986 274700 403992 274712
rect 398892 274672 403992 274700
rect 398892 274660 398898 274672
rect 403986 274660 403992 274672
rect 404044 274660 404050 274712
rect 404262 274660 404268 274712
rect 404320 274700 404326 274712
rect 409874 274700 409880 274712
rect 404320 274672 409880 274700
rect 404320 274660 404326 274672
rect 409874 274660 409880 274672
rect 409932 274660 409938 274712
rect 510522 274660 510528 274712
rect 510580 274700 510586 274712
rect 517422 274700 517428 274712
rect 510580 274672 517428 274700
rect 510580 274660 510586 274672
rect 517422 274660 517428 274672
rect 517480 274660 517486 274712
rect 518866 274700 518894 274740
rect 521010 274700 521016 274712
rect 518866 274672 521016 274700
rect 521010 274660 521016 274672
rect 521068 274660 521074 274712
rect 136818 274592 136824 274644
rect 136876 274632 136882 274644
rect 218238 274632 218244 274644
rect 136876 274604 218244 274632
rect 136876 274592 136882 274604
rect 218238 274592 218244 274604
rect 218296 274592 218302 274644
rect 297358 274592 297364 274644
rect 297416 274632 297422 274644
rect 319990 274632 319996 274644
rect 297416 274604 319996 274632
rect 297416 274592 297422 274604
rect 319990 274592 319996 274604
rect 320048 274592 320054 274644
rect 320082 274592 320088 274644
rect 320140 274632 320146 274644
rect 338942 274632 338948 274644
rect 320140 274604 338948 274632
rect 320140 274592 320146 274604
rect 338942 274592 338948 274604
rect 339000 274592 339006 274644
rect 348510 274592 348516 274644
rect 348568 274632 348574 274644
rect 479610 274632 479616 274644
rect 348568 274604 479616 274632
rect 348568 274592 348574 274604
rect 479610 274592 479616 274604
rect 479668 274592 479674 274644
rect 145006 274524 145012 274576
rect 145064 274564 145070 274576
rect 222194 274564 222200 274576
rect 145064 274536 222200 274564
rect 145064 274524 145070 274536
rect 222194 274524 222200 274536
rect 222252 274524 222258 274576
rect 309778 274524 309784 274576
rect 309836 274564 309842 274576
rect 333054 274564 333060 274576
rect 309836 274536 333060 274564
rect 309836 274524 309842 274536
rect 333054 274524 333060 274536
rect 333112 274524 333118 274576
rect 350350 274524 350356 274576
rect 350408 274564 350414 274576
rect 483198 274564 483204 274576
rect 350408 274536 483204 274564
rect 350408 274524 350414 274536
rect 483198 274524 483204 274536
rect 483256 274524 483262 274576
rect 137922 274456 137928 274508
rect 137980 274496 137986 274508
rect 219618 274496 219624 274508
rect 137980 274468 219624 274496
rect 137980 274456 137986 274468
rect 219618 274456 219624 274468
rect 219676 274456 219682 274508
rect 289630 274456 289636 274508
rect 289688 274496 289694 274508
rect 321186 274496 321192 274508
rect 289688 274468 321192 274496
rect 289688 274456 289694 274468
rect 321186 274456 321192 274468
rect 321244 274456 321250 274508
rect 351730 274456 351736 274508
rect 351788 274496 351794 274508
rect 486694 274496 486700 274508
rect 351788 274468 486700 274496
rect 351788 274456 351794 274468
rect 486694 274456 486700 274468
rect 486752 274456 486758 274508
rect 123754 274388 123760 274440
rect 123812 274428 123818 274440
rect 214098 274428 214104 274440
rect 123812 274400 214104 274428
rect 123812 274388 123818 274400
rect 214098 274388 214104 274400
rect 214156 274388 214162 274440
rect 291838 274388 291844 274440
rect 291896 274428 291902 274440
rect 311710 274428 311716 274440
rect 291896 274400 311716 274428
rect 291896 274388 291902 274400
rect 311710 274388 311716 274400
rect 311768 274388 311774 274440
rect 317782 274388 317788 274440
rect 317840 274428 317846 274440
rect 349614 274428 349620 274440
rect 317840 274400 349620 274428
rect 317840 274388 317846 274400
rect 349614 274388 349620 274400
rect 349672 274388 349678 274440
rect 353018 274388 353024 274440
rect 353076 274428 353082 274440
rect 490282 274428 490288 274440
rect 353076 274400 490288 274428
rect 353076 274388 353082 274400
rect 490282 274388 490288 274400
rect 490340 274388 490346 274440
rect 121362 274320 121368 274372
rect 121420 274360 121426 274372
rect 213086 274360 213092 274372
rect 121420 274332 213092 274360
rect 121420 274320 121426 274332
rect 213086 274320 213092 274332
rect 213144 274320 213150 274372
rect 295978 274320 295984 274372
rect 296036 274360 296042 274372
rect 329466 274360 329472 274372
rect 296036 274332 329472 274360
rect 296036 274320 296042 274332
rect 329466 274320 329472 274332
rect 329524 274320 329530 274372
rect 357250 274320 357256 274372
rect 357308 274360 357314 274372
rect 500862 274360 500868 274372
rect 357308 274332 500868 274360
rect 357308 274320 357314 274332
rect 500862 274320 500868 274332
rect 500920 274320 500926 274372
rect 42150 274252 42156 274304
rect 42208 274292 42214 274304
rect 42978 274292 42984 274304
rect 42208 274264 42984 274292
rect 42208 274252 42214 274264
rect 42978 274252 42984 274264
rect 43036 274252 43042 274304
rect 116670 274252 116676 274304
rect 116728 274292 116734 274304
rect 211338 274292 211344 274304
rect 116728 274264 211344 274292
rect 116728 274252 116734 274264
rect 211338 274252 211344 274264
rect 211396 274252 211402 274304
rect 237282 274252 237288 274304
rect 237340 274292 237346 274304
rect 256878 274292 256884 274304
rect 237340 274264 256884 274292
rect 237340 274252 237346 274264
rect 256878 274252 256884 274264
rect 256936 274252 256942 274304
rect 288342 274252 288348 274304
rect 288400 274292 288406 274304
rect 318794 274292 318800 274304
rect 288400 274264 318800 274292
rect 288400 274252 288406 274264
rect 318794 274252 318800 274264
rect 318852 274252 318858 274304
rect 319438 274252 319444 274304
rect 319496 274292 319502 274304
rect 353110 274292 353116 274304
rect 319496 274264 353116 274292
rect 319496 274252 319502 274264
rect 353110 274252 353116 274264
rect 353168 274252 353174 274304
rect 362586 274252 362592 274304
rect 362644 274292 362650 274304
rect 518618 274292 518624 274304
rect 362644 274264 518624 274292
rect 362644 274252 362650 274264
rect 518618 274252 518624 274264
rect 518676 274252 518682 274304
rect 111978 274184 111984 274236
rect 112036 274224 112042 274236
rect 208946 274224 208952 274236
rect 112036 274196 208952 274224
rect 112036 274184 112042 274196
rect 208946 274184 208952 274196
rect 209004 274184 209010 274236
rect 229002 274184 229008 274236
rect 229060 274224 229066 274236
rect 253474 274224 253480 274236
rect 229060 274196 253480 274224
rect 229060 274184 229066 274196
rect 253474 274184 253480 274196
rect 253532 274184 253538 274236
rect 293678 274184 293684 274236
rect 293736 274224 293742 274236
rect 335354 274224 335360 274236
rect 293736 274196 335360 274224
rect 293736 274184 293742 274196
rect 335354 274184 335360 274196
rect 335412 274184 335418 274236
rect 365622 274184 365628 274236
rect 365680 274224 365686 274236
rect 525702 274224 525708 274236
rect 365680 274196 525708 274224
rect 365680 274184 365686 274196
rect 525702 274184 525708 274196
rect 525760 274184 525766 274236
rect 97718 274116 97724 274168
rect 97776 274156 97782 274168
rect 203610 274156 203616 274168
rect 97776 274128 203616 274156
rect 97776 274116 97782 274128
rect 203610 274116 203616 274128
rect 203668 274116 203674 274168
rect 205358 274116 205364 274168
rect 205416 274156 205422 274168
rect 244550 274156 244556 274168
rect 205416 274128 244556 274156
rect 205416 274116 205422 274128
rect 244550 274116 244556 274128
rect 244608 274116 244614 274168
rect 298002 274116 298008 274168
rect 298060 274156 298066 274168
rect 346026 274156 346032 274168
rect 298060 274128 346032 274156
rect 298060 274116 298066 274128
rect 346026 274116 346032 274128
rect 346084 274116 346090 274168
rect 372522 274116 372528 274168
rect 372580 274156 372586 274168
rect 543458 274156 543464 274168
rect 372580 274128 543464 274156
rect 372580 274116 372586 274128
rect 543458 274116 543464 274128
rect 543516 274116 543522 274168
rect 94222 274048 94228 274100
rect 94280 274088 94286 274100
rect 201586 274088 201592 274100
rect 94280 274060 201592 274088
rect 94280 274048 94286 274060
rect 201586 274048 201592 274060
rect 201644 274048 201650 274100
rect 202966 274048 202972 274100
rect 203024 274088 203030 274100
rect 242894 274088 242900 274100
rect 203024 274060 242900 274088
rect 203024 274048 203030 274060
rect 242894 274048 242900 274060
rect 242952 274048 242958 274100
rect 279418 274048 279424 274100
rect 279476 274088 279482 274100
rect 288066 274088 288072 274100
rect 279476 274060 288072 274088
rect 279476 274048 279482 274060
rect 288066 274048 288072 274060
rect 288124 274048 288130 274100
rect 289722 274048 289728 274100
rect 289780 274088 289786 274100
rect 322382 274088 322388 274100
rect 289780 274060 322388 274088
rect 289780 274048 289786 274060
rect 322382 274048 322388 274060
rect 322440 274048 322446 274100
rect 323670 274048 323676 274100
rect 323728 274088 323734 274100
rect 374362 274088 374368 274100
rect 323728 274060 374368 274088
rect 323728 274048 323734 274060
rect 374362 274048 374368 274060
rect 374420 274048 374426 274100
rect 376662 274048 376668 274100
rect 376720 274088 376726 274100
rect 551738 274088 551744 274100
rect 376720 274060 551744 274088
rect 376720 274048 376726 274060
rect 551738 274048 551744 274060
rect 551796 274048 551802 274100
rect 84746 273980 84752 274032
rect 84804 274020 84810 274032
rect 198826 274020 198832 274032
rect 84804 273992 198832 274020
rect 84804 273980 84810 273992
rect 198826 273980 198832 273992
rect 198884 273980 198890 274032
rect 201770 273980 201776 274032
rect 201828 274020 201834 274032
rect 242986 274020 242992 274032
rect 201828 273992 242992 274020
rect 201828 273980 201834 273992
rect 242986 273980 242992 273992
rect 243044 273980 243050 274032
rect 243538 273980 243544 274032
rect 243596 274020 243602 274032
rect 251634 274020 251640 274032
rect 243596 273992 251640 274020
rect 243596 273980 243602 273992
rect 251634 273980 251640 273992
rect 251692 273980 251698 274032
rect 253842 273980 253848 274032
rect 253900 274020 253906 274032
rect 262766 274020 262772 274032
rect 253900 273992 262772 274020
rect 253900 273980 253906 273992
rect 262766 273980 262772 273992
rect 262824 273980 262830 274032
rect 275922 273980 275928 274032
rect 275980 274020 275986 274032
rect 285766 274020 285772 274032
rect 275980 273992 285772 274020
rect 275980 273980 275986 273992
rect 285766 273980 285772 273992
rect 285824 273980 285830 274032
rect 287698 273980 287704 274032
rect 287756 274020 287762 274032
rect 297542 274020 297548 274032
rect 287756 273992 297548 274020
rect 287756 273980 287762 273992
rect 297542 273980 297548 273992
rect 297600 273980 297606 274032
rect 303338 273980 303344 274032
rect 303396 274020 303402 274032
rect 360194 274020 360200 274032
rect 303396 273992 360200 274020
rect 303396 273980 303402 273992
rect 360194 273980 360200 273992
rect 360252 273980 360258 274032
rect 378042 273980 378048 274032
rect 378100 274020 378106 274032
rect 558822 274020 558828 274032
rect 378100 273992 558828 274020
rect 378100 273980 378106 273992
rect 558822 273980 558828 273992
rect 558880 273980 558886 274032
rect 72970 273912 72976 273964
rect 73028 273952 73034 273964
rect 194594 273952 194600 273964
rect 73028 273924 194600 273952
rect 73028 273912 73034 273924
rect 194594 273912 194600 273924
rect 194652 273912 194658 273964
rect 195882 273912 195888 273964
rect 195940 273952 195946 273964
rect 240226 273952 240232 273964
rect 195940 273924 240232 273952
rect 195940 273912 195946 273924
rect 240226 273912 240232 273924
rect 240284 273912 240290 273964
rect 277302 273912 277308 273964
rect 277360 273952 277366 273964
rect 289262 273952 289268 273964
rect 277360 273924 289268 273952
rect 277360 273912 277366 273924
rect 289262 273912 289268 273924
rect 289320 273912 289326 273964
rect 291102 273912 291108 273964
rect 291160 273952 291166 273964
rect 324774 273952 324780 273964
rect 291160 273924 324780 273952
rect 291160 273912 291166 273924
rect 324774 273912 324780 273924
rect 324832 273912 324838 273964
rect 326338 273912 326344 273964
rect 326396 273952 326402 273964
rect 385034 273952 385040 273964
rect 326396 273924 385040 273952
rect 326396 273912 326402 273924
rect 385034 273912 385040 273924
rect 385092 273912 385098 273964
rect 390370 273912 390376 273964
rect 390428 273952 390434 273964
rect 590746 273952 590752 273964
rect 390428 273924 590752 273952
rect 390428 273912 390434 273924
rect 590746 273912 590752 273924
rect 590804 273912 590810 273964
rect 155678 273844 155684 273896
rect 155736 273884 155742 273896
rect 225874 273884 225880 273896
rect 155736 273856 225880 273884
rect 155736 273844 155742 273856
rect 225874 273844 225880 273856
rect 225932 273844 225938 273896
rect 245562 273844 245568 273896
rect 245620 273884 245626 273896
rect 259638 273884 259644 273896
rect 245620 273856 259644 273884
rect 245620 273844 245626 273856
rect 259638 273844 259644 273856
rect 259696 273844 259702 273896
rect 307018 273844 307024 273896
rect 307076 273884 307082 273896
rect 325970 273884 325976 273896
rect 307076 273856 325976 273884
rect 307076 273844 307082 273856
rect 325970 273844 325976 273856
rect 326028 273844 326034 273896
rect 347682 273844 347688 273896
rect 347740 273884 347746 273896
rect 476114 273884 476120 273896
rect 347740 273856 476120 273884
rect 347740 273844 347746 273856
rect 476114 273844 476120 273856
rect 476172 273844 476178 273896
rect 132034 273776 132040 273828
rect 132092 273816 132098 273828
rect 196618 273816 196624 273828
rect 132092 273788 196624 273816
rect 132092 273776 132098 273788
rect 196618 273776 196624 273788
rect 196676 273776 196682 273828
rect 197078 273776 197084 273828
rect 197136 273816 197142 273828
rect 236638 273816 236644 273828
rect 197136 273788 236644 273816
rect 197136 273776 197142 273788
rect 236638 273776 236644 273788
rect 236696 273776 236702 273828
rect 305638 273776 305644 273828
rect 305696 273816 305702 273828
rect 315298 273816 315304 273828
rect 305696 273788 315304 273816
rect 305696 273776 305702 273788
rect 315298 273776 315304 273788
rect 315356 273776 315362 273828
rect 315390 273776 315396 273828
rect 315448 273816 315454 273828
rect 328270 273816 328276 273828
rect 315448 273788 328276 273816
rect 315448 273776 315454 273788
rect 328270 273776 328276 273788
rect 328328 273776 328334 273828
rect 346210 273776 346216 273828
rect 346268 273816 346274 273828
rect 472526 273816 472532 273828
rect 346268 273788 472532 273816
rect 346268 273776 346274 273788
rect 472526 273776 472532 273788
rect 472584 273776 472590 273828
rect 182910 273708 182916 273760
rect 182968 273748 182974 273760
rect 231118 273748 231124 273760
rect 182968 273720 231124 273748
rect 182968 273708 182974 273720
rect 231118 273708 231124 273720
rect 231176 273708 231182 273760
rect 311158 273708 311164 273760
rect 311216 273748 311222 273760
rect 323578 273748 323584 273760
rect 311216 273720 323584 273748
rect 311216 273708 311222 273720
rect 323578 273708 323584 273720
rect 323636 273708 323642 273760
rect 344554 273708 344560 273760
rect 344612 273748 344618 273760
rect 468938 273748 468944 273760
rect 344612 273720 468944 273748
rect 344612 273708 344618 273720
rect 468938 273708 468944 273720
rect 468996 273708 469002 273760
rect 194686 273640 194692 273692
rect 194744 273680 194750 273692
rect 240134 273680 240140 273692
rect 194744 273652 240140 273680
rect 194744 273640 194750 273652
rect 240134 273640 240140 273652
rect 240192 273640 240198 273692
rect 343450 273640 343456 273692
rect 343508 273680 343514 273692
rect 465442 273680 465448 273692
rect 343508 273652 465448 273680
rect 343508 273640 343514 273652
rect 465442 273640 465448 273652
rect 465500 273640 465506 273692
rect 204162 273572 204168 273624
rect 204220 273612 204226 273624
rect 239398 273612 239404 273624
rect 204220 273584 239404 273612
rect 204220 273572 204226 273584
rect 239398 273572 239404 273584
rect 239456 273572 239462 273624
rect 273162 273572 273168 273624
rect 273220 273612 273226 273624
rect 279786 273612 279792 273624
rect 273220 273584 279792 273612
rect 273220 273572 273226 273584
rect 279786 273572 279792 273584
rect 279844 273572 279850 273624
rect 341886 273572 341892 273624
rect 341944 273612 341950 273624
rect 458174 273612 458180 273624
rect 341944 273584 458180 273612
rect 341944 273572 341950 273584
rect 458174 273572 458180 273584
rect 458232 273572 458238 273624
rect 187694 273504 187700 273556
rect 187752 273544 187758 273556
rect 192386 273544 192392 273556
rect 187752 273516 192392 273544
rect 187752 273504 187758 273516
rect 192386 273504 192392 273516
rect 192444 273504 192450 273556
rect 327718 273504 327724 273556
rect 327776 273544 327782 273556
rect 416958 273544 416964 273556
rect 327776 273516 416964 273544
rect 327776 273504 327782 273516
rect 416958 273504 416964 273516
rect 417016 273504 417022 273556
rect 340690 273436 340696 273488
rect 340748 273476 340754 273488
rect 427722 273476 427728 273488
rect 340748 273448 427728 273476
rect 340748 273436 340754 273448
rect 427722 273436 427728 273448
rect 427780 273436 427786 273488
rect 322198 273368 322204 273420
rect 322256 273408 322262 273420
rect 367278 273408 367284 273420
rect 322256 273380 367284 273408
rect 322256 273368 322262 273380
rect 367278 273368 367284 273380
rect 367336 273368 367342 273420
rect 319530 273232 319536 273284
rect 319588 273272 319594 273284
rect 320082 273272 320088 273284
rect 319588 273244 320088 273272
rect 319588 273232 319594 273244
rect 320082 273232 320088 273244
rect 320140 273232 320146 273284
rect 148594 273164 148600 273216
rect 148652 273204 148658 273216
rect 222286 273204 222292 273216
rect 148652 273176 222292 273204
rect 148652 273164 148658 273176
rect 222286 273164 222292 273176
rect 222344 273164 222350 273216
rect 303522 273164 303528 273216
rect 303580 273204 303586 273216
rect 357894 273204 357900 273216
rect 303580 273176 357900 273204
rect 303580 273164 303586 273176
rect 357894 273164 357900 273176
rect 357952 273164 357958 273216
rect 368290 273164 368296 273216
rect 368348 273204 368354 273216
rect 532786 273204 532792 273216
rect 368348 273176 532792 273204
rect 368348 273164 368354 273176
rect 532786 273164 532792 273176
rect 532844 273164 532850 273216
rect 141510 273096 141516 273148
rect 141568 273136 141574 273148
rect 220814 273136 220820 273148
rect 141568 273108 220820 273136
rect 141568 273096 141574 273108
rect 220814 273096 220820 273108
rect 220872 273096 220878 273148
rect 306282 273096 306288 273148
rect 306340 273136 306346 273148
rect 364978 273136 364984 273148
rect 306340 273108 364984 273136
rect 306340 273096 306346 273108
rect 364978 273096 364984 273108
rect 365036 273096 365042 273148
rect 394418 273096 394424 273148
rect 394476 273136 394482 273148
rect 583754 273136 583760 273148
rect 394476 273108 583760 273136
rect 394476 273096 394482 273108
rect 583754 273096 583760 273108
rect 583812 273096 583818 273148
rect 42150 273028 42156 273080
rect 42208 273068 42214 273080
rect 44450 273068 44456 273080
rect 42208 273040 44456 273068
rect 42208 273028 42214 273040
rect 44450 273028 44456 273040
rect 44508 273028 44514 273080
rect 131114 273028 131120 273080
rect 131172 273068 131178 273080
rect 216030 273068 216036 273080
rect 131172 273040 216036 273068
rect 131172 273028 131178 273040
rect 216030 273028 216036 273040
rect 216088 273028 216094 273080
rect 313090 273028 313096 273080
rect 313148 273068 313154 273080
rect 383838 273068 383844 273080
rect 313148 273040 383844 273068
rect 313148 273028 313154 273040
rect 383838 273028 383844 273040
rect 383896 273028 383902 273080
rect 397270 273028 397276 273080
rect 397328 273068 397334 273080
rect 593414 273068 593420 273080
rect 397328 273040 593420 273068
rect 397328 273028 397334 273040
rect 593414 273028 593420 273040
rect 593472 273028 593478 273080
rect 127342 272960 127348 273012
rect 127400 273000 127406 273012
rect 215386 273000 215392 273012
rect 127400 272972 215392 273000
rect 127400 272960 127406 272972
rect 215386 272960 215392 272972
rect 215444 272960 215450 273012
rect 314470 272960 314476 273012
rect 314528 273000 314534 273012
rect 387426 273000 387432 273012
rect 314528 272972 387432 273000
rect 314528 272960 314534 272972
rect 387426 272960 387432 272972
rect 387484 272960 387490 273012
rect 398926 272960 398932 273012
rect 398984 273000 398990 273012
rect 600038 273000 600044 273012
rect 398984 272972 600044 273000
rect 398984 272960 398990 272972
rect 600038 272960 600044 272972
rect 600096 272960 600102 273012
rect 120258 272892 120264 272944
rect 120316 272932 120322 272944
rect 212626 272932 212632 272944
rect 120316 272904 212632 272932
rect 120316 272892 120322 272904
rect 212626 272892 212632 272904
rect 212684 272892 212690 272944
rect 315850 272892 315856 272944
rect 315908 272932 315914 272944
rect 390922 272932 390928 272944
rect 315908 272904 390928 272932
rect 315908 272892 315914 272904
rect 390922 272892 390928 272904
rect 390980 272892 390986 272944
rect 398650 272892 398656 272944
rect 398708 272932 398714 272944
rect 597830 272932 597836 272944
rect 398708 272904 597836 272932
rect 398708 272892 398714 272904
rect 597830 272892 597836 272904
rect 597888 272892 597894 272944
rect 113174 272824 113180 272876
rect 113232 272864 113238 272876
rect 209958 272864 209964 272876
rect 113232 272836 209964 272864
rect 113232 272824 113238 272836
rect 209958 272824 209964 272836
rect 210016 272824 210022 272876
rect 288434 272824 288440 272876
rect 288492 272864 288498 272876
rect 304626 272864 304632 272876
rect 288492 272836 304632 272864
rect 288492 272824 288498 272836
rect 304626 272824 304632 272836
rect 304684 272824 304690 272876
rect 317230 272824 317236 272876
rect 317288 272864 317294 272876
rect 394510 272864 394516 272876
rect 317288 272836 394516 272864
rect 317288 272824 317294 272836
rect 394510 272824 394516 272836
rect 394568 272824 394574 272876
rect 400306 272824 400312 272876
rect 400364 272864 400370 272876
rect 617978 272864 617984 272876
rect 400364 272836 617984 272864
rect 400364 272824 400370 272836
rect 617978 272824 617984 272836
rect 618036 272824 618042 272876
rect 108390 272756 108396 272808
rect 108448 272796 108454 272808
rect 207566 272796 207572 272808
rect 108448 272768 207572 272796
rect 108448 272756 108454 272768
rect 207566 272756 207572 272768
rect 207624 272756 207630 272808
rect 233694 272756 233700 272808
rect 233752 272796 233758 272808
rect 255498 272796 255504 272808
rect 233752 272768 255504 272796
rect 233752 272756 233758 272768
rect 255498 272756 255504 272768
rect 255556 272756 255562 272808
rect 282730 272756 282736 272808
rect 282788 272796 282794 272808
rect 305822 272796 305828 272808
rect 282788 272768 305828 272796
rect 282788 272756 282794 272768
rect 305822 272756 305828 272768
rect 305880 272756 305886 272808
rect 318610 272756 318616 272808
rect 318668 272796 318674 272808
rect 398006 272796 398012 272808
rect 318668 272768 398012 272796
rect 318668 272756 318674 272768
rect 398006 272756 398012 272768
rect 398064 272756 398070 272808
rect 401962 272756 401968 272808
rect 402020 272796 402026 272808
rect 621474 272796 621480 272808
rect 402020 272768 621480 272796
rect 402020 272756 402026 272768
rect 621474 272756 621480 272768
rect 621532 272756 621538 272808
rect 101306 272688 101312 272740
rect 101364 272728 101370 272740
rect 204806 272728 204812 272740
rect 101364 272700 204812 272728
rect 101364 272688 101370 272700
rect 204806 272688 204812 272700
rect 204864 272688 204870 272740
rect 222470 272688 222476 272740
rect 222528 272728 222534 272740
rect 247218 272728 247224 272740
rect 222528 272700 247224 272728
rect 222528 272688 222534 272700
rect 247218 272688 247224 272700
rect 247276 272688 247282 272740
rect 285582 272688 285588 272740
rect 285640 272728 285646 272740
rect 308214 272728 308220 272740
rect 285640 272700 308220 272728
rect 285640 272688 285646 272700
rect 308214 272688 308220 272700
rect 308272 272688 308278 272740
rect 321278 272688 321284 272740
rect 321336 272728 321342 272740
rect 401594 272728 401600 272740
rect 321336 272700 401600 272728
rect 321336 272688 321342 272700
rect 401594 272688 401600 272700
rect 401652 272688 401658 272740
rect 402974 272688 402980 272740
rect 403032 272728 403038 272740
rect 625062 272728 625068 272740
rect 403032 272700 625068 272728
rect 403032 272688 403038 272700
rect 625062 272688 625068 272700
rect 625120 272688 625126 272740
rect 89530 272620 89536 272672
rect 89588 272660 89594 272672
rect 200482 272660 200488 272672
rect 89588 272632 200488 272660
rect 89588 272620 89594 272632
rect 200482 272620 200488 272632
rect 200540 272620 200546 272672
rect 200574 272620 200580 272672
rect 200632 272660 200638 272672
rect 243078 272660 243084 272672
rect 200632 272632 243084 272660
rect 200632 272620 200638 272632
rect 243078 272620 243084 272632
rect 243136 272620 243142 272672
rect 285398 272620 285404 272672
rect 285456 272660 285462 272672
rect 312906 272660 312912 272672
rect 285456 272632 312912 272660
rect 285456 272620 285462 272632
rect 312906 272620 312912 272632
rect 312964 272620 312970 272672
rect 319898 272620 319904 272672
rect 319956 272660 319962 272672
rect 401686 272660 401692 272672
rect 319956 272632 401692 272660
rect 319956 272620 319962 272632
rect 401686 272620 401692 272632
rect 401744 272620 401750 272672
rect 405642 272620 405648 272672
rect 405700 272660 405706 272672
rect 632146 272660 632152 272672
rect 405700 272632 632152 272660
rect 405700 272620 405706 272632
rect 632146 272620 632152 272632
rect 632204 272620 632210 272672
rect 76006 272552 76012 272604
rect 76064 272592 76070 272604
rect 194778 272592 194784 272604
rect 76064 272564 194784 272592
rect 76064 272552 76070 272564
rect 194778 272552 194784 272564
rect 194836 272552 194842 272604
rect 198274 272552 198280 272604
rect 198332 272592 198338 272604
rect 241882 272592 241888 272604
rect 198332 272564 241888 272592
rect 198332 272552 198338 272564
rect 241882 272552 241888 272564
rect 241940 272552 241946 272604
rect 246758 272552 246764 272604
rect 246816 272592 246822 272604
rect 260098 272592 260104 272604
rect 246816 272564 260104 272592
rect 246816 272552 246822 272564
rect 260098 272552 260104 272564
rect 260156 272552 260162 272604
rect 285858 272552 285864 272604
rect 285916 272592 285922 272604
rect 314102 272592 314108 272604
rect 285916 272564 314108 272592
rect 285916 272552 285922 272564
rect 314102 272552 314108 272564
rect 314160 272552 314166 272604
rect 321370 272552 321376 272604
rect 321428 272592 321434 272604
rect 405182 272592 405188 272604
rect 321428 272564 405188 272592
rect 321428 272552 321434 272564
rect 405182 272552 405188 272564
rect 405240 272552 405246 272604
rect 408310 272552 408316 272604
rect 408368 272592 408374 272604
rect 639230 272592 639236 272604
rect 408368 272564 639236 272592
rect 408368 272552 408374 272564
rect 639230 272552 639236 272564
rect 639288 272552 639294 272604
rect 68186 272484 68192 272536
rect 68244 272524 68250 272536
rect 193214 272524 193220 272536
rect 68244 272496 193220 272524
rect 68244 272484 68250 272496
rect 193214 272484 193220 272496
rect 193272 272484 193278 272536
rect 193490 272484 193496 272536
rect 193548 272524 193554 272536
rect 240318 272524 240324 272536
rect 193548 272496 240324 272524
rect 193548 272484 193554 272496
rect 240318 272484 240324 272496
rect 240376 272484 240382 272536
rect 241974 272484 241980 272536
rect 242032 272524 242038 272536
rect 258350 272524 258356 272536
rect 242032 272496 258356 272524
rect 242032 272484 242038 272496
rect 258350 272484 258356 272496
rect 258408 272484 258414 272536
rect 274726 272484 274732 272536
rect 274784 272524 274790 272536
rect 284570 272524 284576 272536
rect 274784 272496 284576 272524
rect 274784 272484 274790 272496
rect 284570 272484 284576 272496
rect 284628 272484 284634 272536
rect 286778 272484 286784 272536
rect 286836 272524 286842 272536
rect 316494 272524 316500 272536
rect 286836 272496 316500 272524
rect 286836 272484 286842 272496
rect 316494 272484 316500 272496
rect 316552 272484 316558 272536
rect 321186 272484 321192 272536
rect 321244 272524 321250 272536
rect 408402 272524 408408 272536
rect 321244 272496 408408 272524
rect 321244 272484 321250 272496
rect 408402 272484 408408 272496
rect 408460 272484 408466 272536
rect 409598 272484 409604 272536
rect 409656 272524 409662 272536
rect 642726 272524 642732 272536
rect 409656 272496 642732 272524
rect 409656 272484 409662 272496
rect 642726 272484 642732 272496
rect 642784 272484 642790 272536
rect 159266 272416 159272 272468
rect 159324 272456 159330 272468
rect 226886 272456 226892 272468
rect 159324 272428 226892 272456
rect 159324 272416 159330 272428
rect 226886 272416 226892 272428
rect 226944 272416 226950 272468
rect 301498 272416 301504 272468
rect 301556 272456 301562 272468
rect 317690 272456 317696 272468
rect 301556 272428 317696 272456
rect 301556 272416 301562 272428
rect 317690 272416 317696 272428
rect 317748 272416 317754 272468
rect 358630 272416 358636 272468
rect 358688 272456 358694 272468
rect 504450 272456 504456 272468
rect 358688 272428 504456 272456
rect 358688 272416 358694 272428
rect 504450 272416 504456 272428
rect 504508 272416 504514 272468
rect 179322 272348 179328 272400
rect 179380 272388 179386 272400
rect 233786 272388 233792 272400
rect 179380 272360 233792 272388
rect 179380 272348 179386 272360
rect 233786 272348 233792 272360
rect 233844 272348 233850 272400
rect 363598 272348 363604 272400
rect 363656 272388 363662 272400
rect 392118 272388 392124 272400
rect 363656 272360 392124 272388
rect 363656 272348 363662 272360
rect 392118 272348 392124 272360
rect 392176 272348 392182 272400
rect 393130 272348 393136 272400
rect 393188 272388 393194 272400
rect 521562 272388 521568 272400
rect 393188 272360 521568 272388
rect 393188 272348 393194 272360
rect 521562 272348 521568 272360
rect 521620 272348 521626 272400
rect 191190 272280 191196 272332
rect 191248 272320 191254 272332
rect 239214 272320 239220 272332
rect 191248 272292 239220 272320
rect 191248 272280 191254 272292
rect 239214 272280 239220 272292
rect 239272 272280 239278 272332
rect 391750 272280 391756 272332
rect 391808 272320 391814 272332
rect 513466 272320 513472 272332
rect 391808 272292 513472 272320
rect 391808 272280 391814 272292
rect 513466 272280 513472 272292
rect 513524 272280 513530 272332
rect 153286 272212 153292 272264
rect 153344 272252 153350 272264
rect 192478 272252 192484 272264
rect 153344 272224 192484 272252
rect 153344 272212 153350 272224
rect 192478 272212 192484 272224
rect 192536 272212 192542 272264
rect 192570 272212 192576 272264
rect 192628 272252 192634 272264
rect 238846 272252 238852 272264
rect 192628 272224 238852 272252
rect 192628 272212 192634 272224
rect 238846 272212 238852 272224
rect 238904 272212 238910 272264
rect 322658 272212 322664 272264
rect 322716 272252 322722 272264
rect 408586 272252 408592 272264
rect 322716 272224 408592 272252
rect 322716 272212 322722 272224
rect 408586 272212 408592 272224
rect 408644 272212 408650 272264
rect 410426 272212 410432 272264
rect 410484 272252 410490 272264
rect 410484 272224 412634 272252
rect 410484 272212 410490 272224
rect 199470 272144 199476 272196
rect 199528 272184 199534 272196
rect 241606 272184 241612 272196
rect 199528 272156 241612 272184
rect 199528 272144 199534 272156
rect 241606 272144 241612 272156
rect 241664 272144 241670 272196
rect 325602 272144 325608 272196
rect 325660 272184 325666 272196
rect 409966 272184 409972 272196
rect 325660 272156 409972 272184
rect 325660 272144 325666 272156
rect 409966 272144 409972 272156
rect 410024 272144 410030 272196
rect 412606 272184 412634 272224
rect 422938 272212 422944 272264
rect 422996 272252 423002 272264
rect 431126 272252 431132 272264
rect 422996 272224 431132 272252
rect 422996 272212 423002 272224
rect 431126 272212 431132 272224
rect 431184 272212 431190 272264
rect 431218 272212 431224 272264
rect 431276 272252 431282 272264
rect 438210 272252 438216 272264
rect 431276 272224 438216 272252
rect 431276 272212 431282 272224
rect 438210 272212 438216 272224
rect 438268 272212 438274 272264
rect 424042 272184 424048 272196
rect 412606 272156 424048 272184
rect 424042 272144 424048 272156
rect 424100 272144 424106 272196
rect 322750 272076 322756 272128
rect 322808 272116 322814 272128
rect 404262 272116 404268 272128
rect 322808 272088 404268 272116
rect 322808 272076 322814 272088
rect 404262 272076 404268 272088
rect 404320 272076 404326 272128
rect 404354 272076 404360 272128
rect 404412 272116 404418 272128
rect 459646 272116 459652 272128
rect 404412 272088 459652 272116
rect 404412 272076 404418 272088
rect 459646 272076 459652 272088
rect 459704 272076 459710 272128
rect 349798 272008 349804 272060
rect 349856 272048 349862 272060
rect 422846 272048 422852 272060
rect 349856 272020 422852 272048
rect 349856 272008 349862 272020
rect 422846 272008 422852 272020
rect 422904 272008 422910 272060
rect 347038 271940 347044 271992
rect 347096 271980 347102 271992
rect 415762 271980 415768 271992
rect 347096 271952 415768 271980
rect 347096 271940 347102 271952
rect 415762 271940 415768 271952
rect 415820 271940 415826 271992
rect 273806 271872 273812 271924
rect 273864 271912 273870 271924
rect 282178 271912 282184 271924
rect 273864 271884 282184 271912
rect 273864 271872 273870 271884
rect 282178 271872 282184 271884
rect 282236 271872 282242 271924
rect 360838 271872 360844 271924
rect 360896 271912 360902 271924
rect 399202 271912 399208 271924
rect 360896 271884 399208 271912
rect 360896 271872 360902 271884
rect 399202 271872 399208 271884
rect 399260 271872 399266 271924
rect 403434 271872 403440 271924
rect 403492 271912 403498 271924
rect 404354 271912 404360 271924
rect 403492 271884 404360 271912
rect 403492 271872 403498 271884
rect 404354 271872 404360 271884
rect 404412 271872 404418 271924
rect 161566 271804 161572 271856
rect 161624 271844 161630 271856
rect 227806 271844 227812 271856
rect 161624 271816 227812 271844
rect 161624 271804 161630 271816
rect 227806 271804 227812 271816
rect 227864 271804 227870 271856
rect 295242 271804 295248 271856
rect 295300 271844 295306 271856
rect 336550 271844 336556 271856
rect 295300 271816 336556 271844
rect 295300 271804 295306 271816
rect 336550 271804 336556 271816
rect 336608 271804 336614 271856
rect 366910 271804 366916 271856
rect 366968 271844 366974 271856
rect 529290 271844 529296 271856
rect 366968 271816 529296 271844
rect 366968 271804 366974 271816
rect 529290 271804 529296 271816
rect 529348 271804 529354 271856
rect 142706 271736 142712 271788
rect 142764 271776 142770 271788
rect 162118 271776 162124 271788
rect 142764 271748 162124 271776
rect 142764 271736 142770 271748
rect 162118 271736 162124 271748
rect 162176 271736 162182 271788
rect 162762 271736 162768 271788
rect 162820 271776 162826 271788
rect 228266 271776 228272 271788
rect 162820 271748 228272 271776
rect 162820 271736 162826 271748
rect 228266 271736 228272 271748
rect 228324 271736 228330 271788
rect 296438 271736 296444 271788
rect 296496 271776 296502 271788
rect 340138 271776 340144 271788
rect 296496 271748 340144 271776
rect 296496 271736 296502 271748
rect 340138 271736 340144 271748
rect 340196 271736 340202 271788
rect 368106 271736 368112 271788
rect 368164 271776 368170 271788
rect 531590 271776 531596 271788
rect 368164 271748 531596 271776
rect 368164 271736 368170 271748
rect 531590 271736 531596 271748
rect 531648 271736 531654 271788
rect 93026 271668 93032 271720
rect 93084 271708 93090 271720
rect 153838 271708 153844 271720
rect 93084 271680 153844 271708
rect 93084 271668 93090 271680
rect 153838 271668 153844 271680
rect 153896 271668 153902 271720
rect 158070 271668 158076 271720
rect 158128 271708 158134 271720
rect 226426 271708 226432 271720
rect 158128 271680 226432 271708
rect 158128 271668 158134 271680
rect 226426 271668 226432 271680
rect 226484 271668 226490 271720
rect 300762 271668 300768 271720
rect 300820 271708 300826 271720
rect 350718 271708 350724 271720
rect 300820 271680 350724 271708
rect 300820 271668 300826 271680
rect 350718 271668 350724 271680
rect 350776 271668 350782 271720
rect 360010 271668 360016 271720
rect 360068 271708 360074 271720
rect 362218 271708 362224 271720
rect 360068 271680 362224 271708
rect 360068 271668 360074 271680
rect 362218 271668 362224 271680
rect 362276 271668 362282 271720
rect 369486 271668 369492 271720
rect 369544 271708 369550 271720
rect 535178 271708 535184 271720
rect 369544 271680 535184 271708
rect 369544 271668 369550 271680
rect 535178 271668 535184 271680
rect 535236 271668 535242 271720
rect 152182 271600 152188 271652
rect 152240 271640 152246 271652
rect 224494 271640 224500 271652
rect 152240 271612 224500 271640
rect 152240 271600 152246 271612
rect 224494 271600 224500 271612
rect 224552 271600 224558 271652
rect 303154 271600 303160 271652
rect 303212 271640 303218 271652
rect 358998 271640 359004 271652
rect 303212 271612 359004 271640
rect 303212 271600 303218 271612
rect 358998 271600 359004 271612
rect 359056 271600 359062 271652
rect 365530 271600 365536 271652
rect 365588 271640 365594 271652
rect 367002 271640 367008 271652
rect 365588 271612 367008 271640
rect 365588 271600 365594 271612
rect 367002 271600 367008 271612
rect 367060 271600 367066 271652
rect 370774 271600 370780 271652
rect 370832 271640 370838 271652
rect 538766 271640 538772 271652
rect 370832 271612 538772 271640
rect 370832 271600 370838 271612
rect 538766 271600 538772 271612
rect 538824 271600 538830 271652
rect 150986 271532 150992 271584
rect 151044 271572 151050 271584
rect 223666 271572 223672 271584
rect 151044 271544 223672 271572
rect 151044 271532 151050 271544
rect 223666 271532 223672 271544
rect 223724 271532 223730 271584
rect 241422 271532 241428 271584
rect 241480 271572 241486 271584
rect 251266 271572 251272 271584
rect 241480 271544 251272 271572
rect 241480 271532 241486 271544
rect 251266 271532 251272 271544
rect 251324 271532 251330 271584
rect 304442 271532 304448 271584
rect 304500 271572 304506 271584
rect 362310 271572 362316 271584
rect 304500 271544 362316 271572
rect 304500 271532 304506 271544
rect 362310 271532 362316 271544
rect 362368 271532 362374 271584
rect 362678 271532 362684 271584
rect 362736 271572 362742 271584
rect 363506 271572 363512 271584
rect 362736 271544 363512 271572
rect 362736 271532 362742 271544
rect 363506 271532 363512 271544
rect 363564 271532 363570 271584
rect 372154 271532 372160 271584
rect 372212 271572 372218 271584
rect 542262 271572 542268 271584
rect 372212 271544 542268 271572
rect 372212 271532 372218 271544
rect 542262 271532 542268 271544
rect 542320 271532 542326 271584
rect 78858 271464 78864 271516
rect 78916 271504 78922 271516
rect 152458 271504 152464 271516
rect 78916 271476 152464 271504
rect 78916 271464 78922 271476
rect 152458 271464 152464 271476
rect 152516 271464 152522 271516
rect 154482 271464 154488 271516
rect 154540 271504 154546 271516
rect 225046 271504 225052 271516
rect 154540 271476 225052 271504
rect 154540 271464 154546 271476
rect 225046 271464 225052 271476
rect 225104 271464 225110 271516
rect 233878 271464 233884 271516
rect 233936 271504 233942 271516
rect 246022 271504 246028 271516
rect 233936 271476 246028 271504
rect 233936 271464 233942 271476
rect 246022 271464 246028 271476
rect 246080 271464 246086 271516
rect 306190 271464 306196 271516
rect 306248 271504 306254 271516
rect 366082 271504 366088 271516
rect 306248 271476 366088 271504
rect 306248 271464 306254 271476
rect 366082 271464 366088 271476
rect 366140 271464 366146 271516
rect 373810 271464 373816 271516
rect 373868 271504 373874 271516
rect 547046 271504 547052 271516
rect 373868 271476 547052 271504
rect 373868 271464 373874 271476
rect 547046 271464 547052 271476
rect 547104 271464 547110 271516
rect 143902 271396 143908 271448
rect 143960 271436 143966 271448
rect 143960 271408 144316 271436
rect 143960 271396 143966 271408
rect 96614 271328 96620 271380
rect 96672 271368 96678 271380
rect 144178 271368 144184 271380
rect 96672 271340 144184 271368
rect 96672 271328 96678 271340
rect 144178 271328 144184 271340
rect 144236 271328 144242 271380
rect 144288 271368 144316 271408
rect 147398 271396 147404 271448
rect 147456 271436 147462 271448
rect 222470 271436 222476 271448
rect 147456 271408 222476 271436
rect 147456 271396 147462 271408
rect 222470 271396 222476 271408
rect 222528 271396 222534 271448
rect 224954 271396 224960 271448
rect 225012 271436 225018 271448
rect 245930 271436 245936 271448
rect 225012 271408 245936 271436
rect 225012 271396 225018 271408
rect 245930 271396 245936 271408
rect 245988 271396 245994 271448
rect 281534 271396 281540 271448
rect 281592 271436 281598 271448
rect 294046 271436 294052 271448
rect 281592 271408 294052 271436
rect 281592 271396 281598 271408
rect 294046 271396 294052 271408
rect 294104 271396 294110 271448
rect 307478 271396 307484 271448
rect 307536 271436 307542 271448
rect 369670 271436 369676 271448
rect 307536 271408 369676 271436
rect 307536 271396 307542 271408
rect 369670 271396 369676 271408
rect 369728 271396 369734 271448
rect 375282 271396 375288 271448
rect 375340 271436 375346 271448
rect 550542 271436 550548 271448
rect 375340 271408 550548 271436
rect 375340 271396 375346 271408
rect 550542 271396 550548 271408
rect 550600 271396 550606 271448
rect 220906 271368 220912 271380
rect 144288 271340 220912 271368
rect 220906 271328 220912 271340
rect 220964 271328 220970 271380
rect 231394 271328 231400 271380
rect 231452 271368 231458 271380
rect 254302 271368 254308 271380
rect 231452 271340 254308 271368
rect 231452 271328 231458 271340
rect 254302 271328 254308 271340
rect 254360 271328 254366 271380
rect 275646 271328 275652 271380
rect 275704 271368 275710 271380
rect 286502 271368 286508 271380
rect 275704 271340 286508 271368
rect 275704 271328 275710 271340
rect 286502 271328 286508 271340
rect 286560 271328 286566 271380
rect 296346 271368 296352 271380
rect 287532 271340 296352 271368
rect 124950 271260 124956 271312
rect 125008 271300 125014 271312
rect 214006 271300 214012 271312
rect 125008 271272 214012 271300
rect 125008 271260 125014 271272
rect 214006 271260 214012 271272
rect 214064 271260 214070 271312
rect 230198 271260 230204 271312
rect 230256 271300 230262 271312
rect 254026 271300 254032 271312
rect 230256 271272 254032 271300
rect 230256 271260 230262 271272
rect 254026 271260 254032 271272
rect 254084 271260 254090 271312
rect 254210 271260 254216 271312
rect 254268 271300 254274 271312
rect 261478 271300 261484 271312
rect 254268 271272 261484 271300
rect 254268 271260 254274 271272
rect 261478 271260 261484 271272
rect 261536 271260 261542 271312
rect 273346 271260 273352 271312
rect 273404 271300 273410 271312
rect 280982 271300 280988 271312
rect 273404 271272 280988 271300
rect 273404 271260 273410 271272
rect 280982 271260 280988 271272
rect 281040 271260 281046 271312
rect 114278 271192 114284 271244
rect 114336 271232 114342 271244
rect 209866 271232 209872 271244
rect 114336 271204 209872 271232
rect 114336 271192 114342 271204
rect 209866 271192 209872 271204
rect 209924 271192 209930 271244
rect 226610 271192 226616 271244
rect 226668 271232 226674 271244
rect 252646 271232 252652 271244
rect 226668 271204 252652 271232
rect 226668 271192 226674 271204
rect 252646 271192 252652 271204
rect 252704 271192 252710 271244
rect 256142 271192 256148 271244
rect 256200 271232 256206 271244
rect 263686 271232 263692 271244
rect 256200 271204 263692 271232
rect 256200 271192 256206 271204
rect 263686 271192 263692 271204
rect 263744 271192 263750 271244
rect 279142 271192 279148 271244
rect 279200 271232 279206 271244
rect 287532 271232 287560 271340
rect 296346 271328 296352 271340
rect 296404 271328 296410 271380
rect 307570 271328 307576 271380
rect 307628 271368 307634 271380
rect 370866 271368 370872 271380
rect 307628 271340 370872 271368
rect 307628 271328 307634 271340
rect 370866 271328 370872 271340
rect 370924 271328 370930 271380
rect 376570 271328 376576 271380
rect 376628 271368 376634 271380
rect 554130 271368 554136 271380
rect 376628 271340 554136 271368
rect 376628 271328 376634 271340
rect 554130 271328 554136 271340
rect 554188 271328 554194 271380
rect 287790 271260 287796 271312
rect 287848 271300 287854 271312
rect 303430 271300 303436 271312
rect 287848 271272 303436 271300
rect 287848 271260 287854 271272
rect 303430 271260 303436 271272
rect 303488 271260 303494 271312
rect 308950 271260 308956 271312
rect 309008 271300 309014 271312
rect 373258 271300 373264 271312
rect 309008 271272 373264 271300
rect 309008 271260 309014 271272
rect 373258 271260 373264 271272
rect 373316 271260 373322 271312
rect 377950 271260 377956 271312
rect 378008 271300 378014 271312
rect 557626 271300 557632 271312
rect 378008 271272 557632 271300
rect 378008 271260 378014 271272
rect 557626 271260 557632 271272
rect 557684 271260 557690 271312
rect 299934 271232 299940 271244
rect 279200 271204 287560 271232
rect 287624 271204 299940 271232
rect 279200 271192 279206 271204
rect 104894 271124 104900 271176
rect 104952 271164 104958 271176
rect 206278 271164 206284 271176
rect 104952 271136 206284 271164
rect 104952 271124 104958 271136
rect 206278 271124 206284 271136
rect 206336 271124 206342 271176
rect 223574 271124 223580 271176
rect 223632 271164 223638 271176
rect 250346 271164 250352 271176
rect 223632 271136 250352 271164
rect 223632 271124 223638 271136
rect 250346 271124 250352 271136
rect 250404 271124 250410 271176
rect 252922 271124 252928 271176
rect 252980 271164 252986 271176
rect 262306 271164 262312 271176
rect 252980 271136 262312 271164
rect 252980 271124 252986 271136
rect 262306 271124 262312 271136
rect 262364 271124 262370 271176
rect 280522 271124 280528 271176
rect 280580 271164 280586 271176
rect 287624 271164 287652 271204
rect 299934 271192 299940 271204
rect 299992 271192 299998 271244
rect 310330 271192 310336 271244
rect 310388 271232 310394 271244
rect 376754 271232 376760 271244
rect 310388 271204 376760 271232
rect 310388 271192 310394 271204
rect 376754 271192 376760 271204
rect 376812 271192 376818 271244
rect 379422 271192 379428 271244
rect 379480 271232 379486 271244
rect 561214 271232 561220 271244
rect 379480 271204 561220 271232
rect 379480 271192 379486 271204
rect 561214 271192 561220 271204
rect 561272 271192 561278 271244
rect 301130 271164 301136 271176
rect 280580 271136 287652 271164
rect 292546 271136 301136 271164
rect 280580 271124 280586 271136
rect 165154 271056 165160 271108
rect 165212 271096 165218 271108
rect 229278 271096 229284 271108
rect 165212 271068 229284 271096
rect 165212 271056 165218 271068
rect 229278 271056 229284 271068
rect 229336 271056 229342 271108
rect 168650 270988 168656 271040
rect 168708 271028 168714 271040
rect 230658 271028 230664 271040
rect 168708 271000 230664 271028
rect 168708 270988 168714 271000
rect 230658 270988 230664 271000
rect 230716 270988 230722 271040
rect 280982 270988 280988 271040
rect 281040 271028 281046 271040
rect 292546 271028 292574 271136
rect 301130 271124 301136 271136
rect 301188 271124 301194 271176
rect 311802 271124 311808 271176
rect 311860 271164 311866 271176
rect 380342 271164 380348 271176
rect 311860 271136 380348 271164
rect 311860 271124 311866 271136
rect 380342 271124 380348 271136
rect 380400 271124 380406 271176
rect 385954 271124 385960 271176
rect 386012 271164 386018 271176
rect 578878 271164 578884 271176
rect 386012 271136 578884 271164
rect 386012 271124 386018 271136
rect 578878 271124 578884 271136
rect 578936 271124 578942 271176
rect 312446 271056 312452 271108
rect 312504 271096 312510 271108
rect 343634 271096 343640 271108
rect 312504 271068 343640 271096
rect 312504 271056 312510 271068
rect 343634 271056 343640 271068
rect 343692 271056 343698 271108
rect 367002 271056 367008 271108
rect 367060 271096 367066 271108
rect 528094 271096 528100 271108
rect 367060 271068 528100 271096
rect 367060 271056 367066 271068
rect 528094 271056 528100 271068
rect 528152 271056 528158 271108
rect 281040 271000 292574 271028
rect 281040 270988 281046 271000
rect 333238 270988 333244 271040
rect 333296 271028 333302 271040
rect 354306 271028 354312 271040
rect 333296 271000 354312 271028
rect 333296 270988 333302 271000
rect 354306 270988 354312 271000
rect 354364 270988 354370 271040
rect 365438 270988 365444 271040
rect 365496 271028 365502 271040
rect 524506 271028 524512 271040
rect 365496 271000 524512 271028
rect 365496 270988 365502 271000
rect 524506 270988 524512 271000
rect 524564 270988 524570 271040
rect 172238 270920 172244 270972
rect 172296 270960 172302 270972
rect 232038 270960 232044 270972
rect 172296 270932 232044 270960
rect 172296 270920 172302 270932
rect 232038 270920 232044 270932
rect 232096 270920 232102 270972
rect 286962 270920 286968 270972
rect 287020 270960 287026 270972
rect 287790 270960 287796 270972
rect 287020 270932 287796 270960
rect 287020 270920 287026 270932
rect 287790 270920 287796 270932
rect 287848 270920 287854 270972
rect 327810 270920 327816 270972
rect 327868 270960 327874 270972
rect 347222 270960 347228 270972
rect 327868 270932 347228 270960
rect 327868 270920 327874 270932
rect 347222 270920 347228 270932
rect 347280 270920 347286 270972
rect 364150 270920 364156 270972
rect 364208 270960 364214 270972
rect 516134 270960 516140 270972
rect 364208 270932 516140 270960
rect 364208 270920 364214 270932
rect 516134 270920 516140 270932
rect 516192 270920 516198 270972
rect 175826 270852 175832 270904
rect 175884 270892 175890 270904
rect 233418 270892 233424 270904
rect 175884 270864 233424 270892
rect 175884 270852 175890 270864
rect 233418 270852 233424 270864
rect 233476 270852 233482 270904
rect 362770 270852 362776 270904
rect 362828 270892 362834 270904
rect 510522 270892 510528 270904
rect 362828 270864 510528 270892
rect 362828 270852 362834 270864
rect 510522 270852 510528 270864
rect 510580 270852 510586 270904
rect 189994 270784 190000 270836
rect 190052 270824 190058 270836
rect 235350 270824 235356 270836
rect 190052 270796 235356 270824
rect 190052 270784 190058 270796
rect 235350 270784 235356 270796
rect 235408 270784 235414 270836
rect 361482 270784 361488 270836
rect 361540 270824 361546 270836
rect 496722 270824 496728 270836
rect 361540 270796 496728 270824
rect 361540 270784 361546 270796
rect 496722 270784 496728 270796
rect 496780 270784 496786 270836
rect 221918 270716 221924 270768
rect 221976 270756 221982 270768
rect 238110 270756 238116 270768
rect 221976 270728 238116 270756
rect 221976 270716 221982 270728
rect 238110 270716 238116 270728
rect 238168 270716 238174 270768
rect 359918 270716 359924 270768
rect 359976 270756 359982 270768
rect 466730 270756 466736 270768
rect 359976 270728 466736 270756
rect 359976 270716 359982 270728
rect 466730 270716 466736 270728
rect 466788 270716 466794 270768
rect 329558 270648 329564 270700
rect 329616 270688 329622 270700
rect 429930 270688 429936 270700
rect 329616 270660 429936 270688
rect 329616 270648 329622 270660
rect 429930 270648 429936 270660
rect 429988 270648 429994 270700
rect 332318 270580 332324 270632
rect 332376 270620 332382 270632
rect 375190 270620 375196 270632
rect 332376 270592 375196 270620
rect 332376 270580 332382 270592
rect 375190 270580 375196 270592
rect 375248 270580 375254 270632
rect 70578 270444 70584 270496
rect 70636 270484 70642 270496
rect 71774 270484 71780 270496
rect 70636 270456 71780 270484
rect 70636 270444 70642 270456
rect 71774 270444 71780 270456
rect 71832 270444 71838 270496
rect 169846 270444 169852 270496
rect 169904 270484 169910 270496
rect 231486 270484 231492 270496
rect 169904 270456 231492 270484
rect 169904 270444 169910 270456
rect 231486 270444 231492 270456
rect 231544 270444 231550 270496
rect 296530 270444 296536 270496
rect 296588 270484 296594 270496
rect 342254 270484 342260 270496
rect 296588 270456 342260 270484
rect 296588 270444 296594 270456
rect 342254 270444 342260 270456
rect 342312 270444 342318 270496
rect 346394 270444 346400 270496
rect 346452 270484 346458 270496
rect 474734 270484 474740 270496
rect 346452 270456 474740 270484
rect 346452 270444 346458 270456
rect 474734 270444 474740 270456
rect 474792 270444 474798 270496
rect 166902 270376 166908 270428
rect 166960 270416 166966 270428
rect 230198 270416 230204 270428
rect 166960 270388 230204 270416
rect 166960 270376 166966 270388
rect 230198 270376 230204 270388
rect 230256 270376 230262 270428
rect 297450 270376 297456 270428
rect 297508 270416 297514 270428
rect 343818 270416 343824 270428
rect 297508 270388 343824 270416
rect 297508 270376 297514 270388
rect 343818 270376 343824 270388
rect 343876 270376 343882 270428
rect 354858 270376 354864 270428
rect 354916 270416 354922 270428
rect 496814 270416 496820 270428
rect 354916 270388 496820 270416
rect 354916 270376 354922 270388
rect 496814 270376 496820 270388
rect 496872 270376 496878 270428
rect 140682 270308 140688 270360
rect 140740 270348 140746 270360
rect 219986 270348 219992 270360
rect 140740 270320 219992 270348
rect 140740 270308 140746 270320
rect 219986 270308 219992 270320
rect 220044 270308 220050 270360
rect 220630 270308 220636 270360
rect 220688 270348 220694 270360
rect 224402 270348 224408 270360
rect 220688 270320 224408 270348
rect 220688 270308 220694 270320
rect 224402 270308 224408 270320
rect 224460 270308 224466 270360
rect 298738 270308 298744 270360
rect 298796 270348 298802 270360
rect 347774 270348 347780 270360
rect 298796 270320 347780 270348
rect 298796 270308 298802 270320
rect 347774 270308 347780 270320
rect 347832 270308 347838 270360
rect 360194 270308 360200 270360
rect 360252 270348 360258 270360
rect 510614 270348 510620 270360
rect 360252 270320 510620 270348
rect 360252 270308 360258 270320
rect 510614 270308 510620 270320
rect 510672 270308 510678 270360
rect 133782 270240 133788 270292
rect 133840 270280 133846 270292
rect 216950 270280 216956 270292
rect 133840 270252 216956 270280
rect 133840 270240 133846 270252
rect 216950 270240 216956 270252
rect 217008 270240 217014 270292
rect 300118 270240 300124 270292
rect 300176 270280 300182 270292
rect 351914 270280 351920 270292
rect 300176 270252 351920 270280
rect 300176 270240 300182 270252
rect 351914 270240 351920 270252
rect 351972 270240 351978 270292
rect 364242 270240 364248 270292
rect 364300 270280 364306 270292
rect 521654 270280 521660 270292
rect 364300 270252 521660 270280
rect 364300 270240 364306 270252
rect 521654 270240 521660 270252
rect 521712 270240 521718 270292
rect 129642 270172 129648 270224
rect 129700 270212 129706 270224
rect 215938 270212 215944 270224
rect 129700 270184 215944 270212
rect 129700 270172 129706 270184
rect 215938 270172 215944 270184
rect 215996 270172 216002 270224
rect 301406 270172 301412 270224
rect 301464 270212 301470 270224
rect 354674 270212 354680 270224
rect 301464 270184 354680 270212
rect 301464 270172 301470 270184
rect 354674 270172 354680 270184
rect 354732 270172 354738 270224
rect 369578 270172 369584 270224
rect 369636 270212 369642 270224
rect 535454 270212 535460 270224
rect 369636 270184 535460 270212
rect 369636 270172 369642 270184
rect 535454 270172 535460 270184
rect 535512 270172 535518 270224
rect 103698 270104 103704 270156
rect 103756 270144 103762 270156
rect 125962 270144 125968 270156
rect 103756 270116 125968 270144
rect 103756 270104 103762 270116
rect 125962 270104 125968 270116
rect 126020 270104 126026 270156
rect 126882 270104 126888 270156
rect 126940 270144 126946 270156
rect 214650 270144 214656 270156
rect 126940 270116 214656 270144
rect 126940 270104 126946 270116
rect 214650 270104 214656 270116
rect 214708 270104 214714 270156
rect 248046 270144 248052 270156
rect 238726 270116 248052 270144
rect 119062 270036 119068 270088
rect 119120 270076 119126 270088
rect 119120 270048 119752 270076
rect 119120 270036 119126 270048
rect 110782 269968 110788 270020
rect 110840 270008 110846 270020
rect 119614 270008 119620 270020
rect 110840 269980 119620 270008
rect 110840 269968 110846 269980
rect 119614 269968 119620 269980
rect 119672 269968 119678 270020
rect 119724 270008 119752 270048
rect 122742 270036 122748 270088
rect 122800 270076 122806 270088
rect 212902 270076 212908 270088
rect 122800 270048 212908 270076
rect 122800 270036 122806 270048
rect 212902 270036 212908 270048
rect 212960 270036 212966 270088
rect 234614 270036 234620 270088
rect 234672 270076 234678 270088
rect 238726 270076 238754 270116
rect 248046 270104 248052 270116
rect 248104 270104 248110 270156
rect 301866 270104 301872 270156
rect 301924 270144 301930 270156
rect 356054 270144 356060 270156
rect 301924 270116 356060 270144
rect 301924 270104 301930 270116
rect 356054 270104 356060 270116
rect 356112 270104 356118 270156
rect 373994 270104 374000 270156
rect 374052 270144 374058 270156
rect 547874 270144 547880 270156
rect 374052 270116 547880 270144
rect 374052 270104 374058 270116
rect 547874 270104 547880 270116
rect 547932 270104 547938 270156
rect 245286 270076 245292 270088
rect 234672 270048 238754 270076
rect 241992 270048 245292 270076
rect 234672 270036 234678 270048
rect 211890 270008 211896 270020
rect 119724 269980 211896 270008
rect 211890 269968 211896 269980
rect 211948 269968 211954 270020
rect 237374 269968 237380 270020
rect 237432 270008 237438 270020
rect 241992 270008 242020 270048
rect 245286 270036 245292 270048
rect 245344 270036 245350 270088
rect 248322 270036 248328 270088
rect 248380 270076 248386 270088
rect 260926 270076 260932 270088
rect 248380 270048 260932 270076
rect 248380 270036 248386 270048
rect 260926 270036 260932 270048
rect 260984 270036 260990 270088
rect 293402 270036 293408 270088
rect 293460 270076 293466 270088
rect 333974 270076 333980 270088
rect 293460 270048 333980 270076
rect 293460 270036 293466 270048
rect 333974 270036 333980 270048
rect 334032 270036 334038 270088
rect 339770 270036 339776 270088
rect 339828 270076 339834 270088
rect 456794 270076 456800 270088
rect 339828 270048 456800 270076
rect 339828 270036 339834 270048
rect 456794 270036 456800 270048
rect 456852 270036 456858 270088
rect 457990 270036 457996 270088
rect 458048 270076 458054 270088
rect 636194 270076 636200 270088
rect 458048 270048 636200 270076
rect 458048 270036 458054 270048
rect 636194 270036 636200 270048
rect 636252 270036 636258 270088
rect 237432 269980 242020 270008
rect 237432 269968 237438 269980
rect 244366 269968 244372 270020
rect 244424 270008 244430 270020
rect 259546 270008 259552 270020
rect 244424 269980 259552 270008
rect 244424 269968 244430 269980
rect 259546 269968 259552 269980
rect 259604 269968 259610 270020
rect 303338 269968 303344 270020
rect 303396 270008 303402 270020
rect 303522 270008 303528 270020
rect 303396 269980 303528 270008
rect 303396 269968 303402 269980
rect 303522 269968 303528 269980
rect 303580 269968 303586 270020
rect 304534 269968 304540 270020
rect 304592 270008 304598 270020
rect 362954 270008 362960 270020
rect 304592 269980 362960 270008
rect 304592 269968 304598 269980
rect 362954 269968 362960 269980
rect 363012 269968 363018 270020
rect 381630 269968 381636 270020
rect 381688 270008 381694 270020
rect 567194 270008 567200 270020
rect 381688 269980 567200 270008
rect 381688 269968 381694 269980
rect 567194 269968 567200 269980
rect 567252 269968 567258 270020
rect 85942 269900 85948 269952
rect 86000 269940 86006 269952
rect 110506 269940 110512 269952
rect 86000 269912 110512 269940
rect 86000 269900 86006 269912
rect 110506 269900 110512 269912
rect 110564 269900 110570 269952
rect 118602 269900 118608 269952
rect 118660 269940 118666 269952
rect 212350 269940 212356 269952
rect 118660 269912 212356 269940
rect 118660 269900 118666 269912
rect 212350 269900 212356 269912
rect 212408 269900 212414 269952
rect 236086 269900 236092 269952
rect 236144 269940 236150 269952
rect 256418 269940 256424 269952
rect 236144 269912 256424 269940
rect 236144 269900 236150 269912
rect 256418 269900 256424 269912
rect 256476 269900 256482 269952
rect 274266 269900 274272 269952
rect 274324 269940 274330 269952
rect 282914 269940 282920 269952
rect 274324 269912 282920 269940
rect 274324 269900 274330 269912
rect 282914 269900 282920 269912
rect 282972 269900 282978 269952
rect 283558 269900 283564 269952
rect 283616 269940 283622 269952
rect 292574 269940 292580 269952
rect 283616 269912 292580 269940
rect 283616 269900 283622 269912
rect 292574 269900 292580 269912
rect 292632 269900 292638 269952
rect 314286 269900 314292 269952
rect 314344 269940 314350 269952
rect 376938 269940 376944 269952
rect 314344 269912 376944 269940
rect 314344 269900 314350 269912
rect 376938 269900 376944 269912
rect 376996 269900 377002 269952
rect 380710 269900 380716 269952
rect 380768 269940 380774 269952
rect 565906 269940 565912 269952
rect 380768 269912 565912 269940
rect 380768 269900 380774 269912
rect 565906 269900 565912 269912
rect 565964 269900 565970 269952
rect 77202 269832 77208 269884
rect 77260 269872 77266 269884
rect 113174 269872 113180 269884
rect 77260 269844 113180 269872
rect 77260 269832 77266 269844
rect 113174 269832 113180 269844
rect 113232 269832 113238 269884
rect 115842 269832 115848 269884
rect 115900 269872 115906 269884
rect 210602 269872 210608 269884
rect 115900 269844 210608 269872
rect 115900 269832 115906 269844
rect 210602 269832 210608 269844
rect 210660 269832 210666 269884
rect 227714 269832 227720 269884
rect 227772 269872 227778 269884
rect 248414 269872 248420 269884
rect 227772 269844 248420 269872
rect 227772 269832 227778 269844
rect 248414 269832 248420 269844
rect 248472 269832 248478 269884
rect 276934 269832 276940 269884
rect 276992 269872 276998 269884
rect 289814 269872 289820 269884
rect 276992 269844 289820 269872
rect 276992 269832 276998 269844
rect 289814 269832 289820 269844
rect 289872 269832 289878 269884
rect 294782 269832 294788 269884
rect 294840 269872 294846 269884
rect 336734 269872 336740 269884
rect 294840 269844 336740 269872
rect 294840 269832 294846 269844
rect 336734 269832 336740 269844
rect 336792 269832 336798 269884
rect 337102 269832 337108 269884
rect 337160 269872 337166 269884
rect 449894 269872 449900 269884
rect 337160 269844 449900 269872
rect 337160 269832 337166 269844
rect 449894 269832 449900 269844
rect 449952 269832 449958 269884
rect 451366 269832 451372 269884
rect 451424 269872 451430 269884
rect 644474 269872 644480 269884
rect 451424 269844 644480 269872
rect 451424 269832 451430 269844
rect 644474 269832 644480 269844
rect 644532 269832 644538 269884
rect 110322 269764 110328 269816
rect 110380 269804 110386 269816
rect 208854 269804 208860 269816
rect 110380 269776 208860 269804
rect 110380 269764 110386 269776
rect 208854 269764 208860 269776
rect 208912 269764 208918 269816
rect 216674 269764 216680 269816
rect 216732 269804 216738 269816
rect 229462 269804 229468 269816
rect 216732 269776 229468 269804
rect 216732 269764 216738 269776
rect 229462 269764 229468 269776
rect 229520 269764 229526 269816
rect 229830 269764 229836 269816
rect 229888 269804 229894 269816
rect 252462 269804 252468 269816
rect 229888 269776 252468 269804
rect 229888 269764 229894 269776
rect 252462 269764 252468 269776
rect 252520 269764 252526 269816
rect 278682 269764 278688 269816
rect 278740 269804 278746 269816
rect 294138 269804 294144 269816
rect 278740 269776 294144 269804
rect 278740 269764 278746 269776
rect 294138 269764 294144 269776
rect 294196 269764 294202 269816
rect 319254 269764 319260 269816
rect 319312 269804 319318 269816
rect 388162 269804 388168 269816
rect 319312 269776 388168 269804
rect 319312 269764 319318 269776
rect 388162 269764 388168 269776
rect 388220 269764 388226 269816
rect 388714 269764 388720 269816
rect 388772 269804 388778 269816
rect 586514 269804 586520 269816
rect 388772 269776 586520 269804
rect 388772 269764 388778 269776
rect 586514 269764 586520 269776
rect 586572 269764 586578 269816
rect 173802 269696 173808 269748
rect 173860 269736 173866 269748
rect 232866 269736 232872 269748
rect 173860 269708 232872 269736
rect 173860 269696 173866 269708
rect 232866 269696 232872 269708
rect 232924 269696 232930 269748
rect 296070 269696 296076 269748
rect 296128 269736 296134 269748
rect 340874 269736 340880 269748
rect 296128 269708 340880 269736
rect 296128 269696 296134 269708
rect 340874 269696 340880 269708
rect 340932 269696 340938 269748
rect 345106 269696 345112 269748
rect 345164 269736 345170 269748
rect 470594 269736 470600 269748
rect 345164 269708 470600 269736
rect 345164 269696 345170 269708
rect 470594 269696 470600 269708
rect 470652 269696 470658 269748
rect 470686 269696 470692 269748
rect 470744 269736 470750 269748
rect 476298 269736 476304 269748
rect 470744 269708 476304 269736
rect 470744 269696 470750 269708
rect 476298 269696 476304 269708
rect 476356 269696 476362 269748
rect 176930 269628 176936 269680
rect 176988 269668 176994 269680
rect 234154 269668 234160 269680
rect 176988 269640 234160 269668
rect 176988 269628 176994 269640
rect 234154 269628 234160 269640
rect 234212 269628 234218 269680
rect 292574 269628 292580 269680
rect 292632 269668 292638 269680
rect 331214 269668 331220 269680
rect 292632 269640 331220 269668
rect 292632 269628 292638 269640
rect 331214 269628 331220 269640
rect 331272 269628 331278 269680
rect 343726 269628 343732 269680
rect 343784 269668 343790 269680
rect 467834 269668 467840 269680
rect 343784 269640 467840 269668
rect 343784 269628 343790 269640
rect 467834 269628 467840 269640
rect 467892 269628 467898 269680
rect 180702 269560 180708 269612
rect 180760 269600 180766 269612
rect 235534 269600 235540 269612
rect 180760 269572 235540 269600
rect 180760 269560 180766 269572
rect 235534 269560 235540 269572
rect 235592 269560 235598 269612
rect 292114 269560 292120 269612
rect 292172 269600 292178 269612
rect 329834 269600 329840 269612
rect 292172 269572 329840 269600
rect 292172 269560 292178 269572
rect 329834 269560 329840 269572
rect 329892 269560 329898 269612
rect 342438 269560 342444 269612
rect 342496 269600 342502 269612
rect 463694 269600 463700 269612
rect 342496 269572 463700 269600
rect 342496 269560 342502 269572
rect 463694 269560 463700 269572
rect 463752 269560 463758 269612
rect 135622 269492 135628 269544
rect 135680 269532 135686 269544
rect 184750 269532 184756 269544
rect 135680 269504 184756 269532
rect 135680 269492 135686 269504
rect 184750 269492 184756 269504
rect 184808 269492 184814 269544
rect 184842 269492 184848 269544
rect 184900 269532 184906 269544
rect 236914 269532 236920 269544
rect 184900 269504 236920 269532
rect 184900 269492 184906 269504
rect 236914 269492 236920 269504
rect 236972 269492 236978 269544
rect 290734 269492 290740 269544
rect 290792 269532 290798 269544
rect 327074 269532 327080 269544
rect 290792 269504 327080 269532
rect 290792 269492 290798 269504
rect 327074 269492 327080 269504
rect 327132 269492 327138 269544
rect 341058 269492 341064 269544
rect 341116 269532 341122 269544
rect 459738 269532 459744 269544
rect 341116 269504 459744 269532
rect 341116 269492 341122 269504
rect 459738 269492 459744 269504
rect 459796 269492 459802 269544
rect 187510 269424 187516 269476
rect 187568 269464 187574 269476
rect 238202 269464 238208 269476
rect 187568 269436 238208 269464
rect 187568 269424 187574 269436
rect 238202 269424 238208 269436
rect 238260 269424 238266 269476
rect 338390 269424 338396 269476
rect 338448 269464 338454 269476
rect 452654 269464 452660 269476
rect 338448 269436 452660 269464
rect 338448 269424 338454 269436
rect 452654 269424 452660 269436
rect 452712 269424 452718 269476
rect 335722 269356 335728 269408
rect 335780 269396 335786 269408
rect 445754 269396 445760 269408
rect 335780 269368 445760 269396
rect 335780 269356 335786 269368
rect 445754 269356 445760 269368
rect 445812 269356 445818 269408
rect 334342 269288 334348 269340
rect 334400 269328 334406 269340
rect 442994 269328 443000 269340
rect 334400 269300 443000 269328
rect 334400 269288 334406 269300
rect 442994 269288 443000 269300
rect 443052 269288 443058 269340
rect 353294 269220 353300 269272
rect 353352 269260 353358 269272
rect 380894 269260 380900 269272
rect 353352 269232 380900 269260
rect 353352 269220 353358 269232
rect 380894 269220 380900 269232
rect 380952 269220 380958 269272
rect 102502 269016 102508 269068
rect 102560 269056 102566 269068
rect 206186 269056 206192 269068
rect 102560 269028 206192 269056
rect 102560 269016 102566 269028
rect 206186 269016 206192 269028
rect 206244 269016 206250 269068
rect 249610 269016 249616 269068
rect 249668 269056 249674 269068
rect 253382 269056 253388 269068
rect 249668 269028 253388 269056
rect 249668 269016 249674 269028
rect 253382 269016 253388 269028
rect 253440 269016 253446 269068
rect 303706 269016 303712 269068
rect 303764 269056 303770 269068
rect 360378 269056 360384 269068
rect 303764 269028 360384 269056
rect 303764 269016 303770 269028
rect 360378 269016 360384 269028
rect 360436 269016 360442 269068
rect 361574 269016 361580 269068
rect 361632 269056 361638 269068
rect 514754 269056 514760 269068
rect 361632 269028 514760 269056
rect 361632 269016 361638 269028
rect 514754 269016 514760 269028
rect 514812 269016 514818 269068
rect 99282 268948 99288 269000
rect 99340 268988 99346 269000
rect 204438 268988 204444 269000
rect 99340 268960 204444 268988
rect 99340 268948 99346 268960
rect 204438 268948 204444 268960
rect 204496 268948 204502 269000
rect 249702 268948 249708 269000
rect 249760 268988 249766 269000
rect 257798 268988 257804 269000
rect 249760 268960 257804 268988
rect 249760 268948 249766 268960
rect 257798 268948 257804 268960
rect 257856 268948 257862 269000
rect 308858 268948 308864 269000
rect 308916 268988 308922 269000
rect 375374 268988 375380 269000
rect 308916 268960 375380 268988
rect 308916 268948 308922 268960
rect 375374 268948 375380 268960
rect 375432 268948 375438 269000
rect 391842 268948 391848 269000
rect 391900 268988 391906 269000
rect 543734 268988 543740 269000
rect 391900 268960 543740 268988
rect 391900 268948 391906 268960
rect 543734 268948 543740 268960
rect 543792 268948 543798 269000
rect 95418 268880 95424 268932
rect 95476 268920 95482 268932
rect 203518 268920 203524 268932
rect 95476 268892 203524 268920
rect 95476 268880 95482 268892
rect 203518 268880 203524 268892
rect 203576 268880 203582 268932
rect 306650 268880 306656 268932
rect 306708 268920 306714 268932
rect 368474 268920 368480 268932
rect 306708 268892 368480 268920
rect 306708 268880 306714 268892
rect 368474 268880 368480 268892
rect 368532 268880 368538 268932
rect 370866 268880 370872 268932
rect 370924 268920 370930 268932
rect 539594 268920 539600 268932
rect 370924 268892 539600 268920
rect 370924 268880 370930 268892
rect 539594 268880 539600 268892
rect 539652 268880 539658 268932
rect 92382 268812 92388 268864
rect 92440 268852 92446 268864
rect 202138 268852 202144 268864
rect 92440 268824 202144 268852
rect 92440 268812 92446 268824
rect 202138 268812 202144 268824
rect 202196 268812 202202 268864
rect 321002 268812 321008 268864
rect 321060 268852 321066 268864
rect 401778 268852 401784 268864
rect 321060 268824 401784 268852
rect 321060 268812 321066 268824
rect 401778 268812 401784 268824
rect 401836 268812 401842 268864
rect 404354 268812 404360 268864
rect 404412 268852 404418 268864
rect 587894 268852 587900 268864
rect 404412 268824 587900 268852
rect 404412 268812 404418 268824
rect 587894 268812 587900 268824
rect 587952 268812 587958 268864
rect 87138 268744 87144 268796
rect 87196 268784 87202 268796
rect 200390 268784 200396 268796
rect 87196 268756 200396 268784
rect 87196 268744 87202 268756
rect 200390 268744 200396 268756
rect 200448 268744 200454 268796
rect 204898 268744 204904 268796
rect 204956 268784 204962 268796
rect 226702 268784 226708 268796
rect 204956 268756 226708 268784
rect 204956 268744 204962 268756
rect 226702 268744 226708 268756
rect 226760 268744 226766 268796
rect 310422 268744 310428 268796
rect 310480 268784 310486 268796
rect 378134 268784 378140 268796
rect 310480 268756 378140 268784
rect 310480 268744 310486 268756
rect 378134 268744 378140 268756
rect 378192 268744 378198 268796
rect 393222 268744 393228 268796
rect 393280 268784 393286 268796
rect 581638 268784 581644 268796
rect 393280 268756 581644 268784
rect 393280 268744 393286 268756
rect 581638 268744 581644 268756
rect 581696 268744 581702 268796
rect 82722 268676 82728 268728
rect 82780 268716 82786 268728
rect 198550 268716 198556 268728
rect 82780 268688 198556 268716
rect 82780 268676 82786 268688
rect 198550 268676 198556 268688
rect 198608 268676 198614 268728
rect 218330 268676 218336 268728
rect 218388 268716 218394 268728
rect 242802 268716 242808 268728
rect 218388 268688 242808 268716
rect 218388 268676 218394 268688
rect 242802 268676 242808 268688
rect 242860 268676 242866 268728
rect 277394 268676 277400 268728
rect 277452 268716 277458 268728
rect 291194 268716 291200 268728
rect 277452 268688 291200 268716
rect 277452 268676 277458 268688
rect 291194 268676 291200 268688
rect 291252 268676 291258 268728
rect 312998 268676 313004 268728
rect 313056 268716 313062 268728
rect 385218 268716 385224 268728
rect 313056 268688 385224 268716
rect 313056 268676 313062 268688
rect 385218 268676 385224 268688
rect 385276 268676 385282 268728
rect 394050 268676 394056 268728
rect 394108 268716 394114 268728
rect 600314 268716 600320 268728
rect 394108 268688 600320 268716
rect 394108 268676 394114 268688
rect 600314 268676 600320 268688
rect 600372 268676 600378 268728
rect 80054 268608 80060 268660
rect 80112 268648 80118 268660
rect 197262 268648 197268 268660
rect 80112 268620 197268 268648
rect 80112 268608 80118 268620
rect 197262 268608 197268 268620
rect 197320 268608 197326 268660
rect 219526 268608 219532 268660
rect 219584 268648 219590 268660
rect 250254 268648 250260 268660
rect 219584 268620 250260 268648
rect 219584 268608 219590 268620
rect 250254 268608 250260 268620
rect 250312 268608 250318 268660
rect 280062 268608 280068 268660
rect 280120 268648 280126 268660
rect 298094 268648 298100 268660
rect 280120 268620 298100 268648
rect 280120 268608 280126 268620
rect 298094 268608 298100 268620
rect 298152 268608 298158 268660
rect 314378 268608 314384 268660
rect 314436 268648 314442 268660
rect 389174 268648 389180 268660
rect 314436 268620 389180 268648
rect 314436 268608 314442 268620
rect 389174 268608 389180 268620
rect 389232 268608 389238 268660
rect 394510 268608 394516 268660
rect 394568 268648 394574 268660
rect 601694 268648 601700 268660
rect 394568 268620 601700 268648
rect 394568 268608 394574 268620
rect 601694 268608 601700 268620
rect 601752 268608 601758 268660
rect 77662 268540 77668 268592
rect 77720 268580 77726 268592
rect 196802 268580 196808 268592
rect 77720 268552 196808 268580
rect 77720 268540 77726 268552
rect 196802 268540 196808 268552
rect 196860 268540 196866 268592
rect 217134 268540 217140 268592
rect 217192 268580 217198 268592
rect 249334 268580 249340 268592
rect 217192 268552 249340 268580
rect 217192 268540 217198 268552
rect 249334 268540 249340 268552
rect 249392 268540 249398 268592
rect 289906 268540 289912 268592
rect 289964 268580 289970 268592
rect 310514 268580 310520 268592
rect 289964 268552 310520 268580
rect 289964 268540 289970 268552
rect 310514 268540 310520 268552
rect 310572 268540 310578 268592
rect 315666 268540 315672 268592
rect 315724 268580 315730 268592
rect 393314 268580 393320 268592
rect 315724 268552 393320 268580
rect 315724 268540 315730 268552
rect 393314 268540 393320 268552
rect 393372 268540 393378 268592
rect 395798 268540 395804 268592
rect 395856 268580 395862 268592
rect 605834 268580 605840 268592
rect 395856 268552 605840 268580
rect 395856 268540 395862 268552
rect 605834 268540 605840 268552
rect 605892 268540 605898 268592
rect 75822 268472 75828 268524
rect 75880 268512 75886 268524
rect 195422 268512 195428 268524
rect 75880 268484 195428 268512
rect 75880 268472 75886 268484
rect 195422 268472 195428 268484
rect 195480 268472 195486 268524
rect 216582 268472 216588 268524
rect 216640 268512 216646 268524
rect 248874 268512 248880 268524
rect 216640 268484 248880 268512
rect 216640 268472 216646 268484
rect 248874 268472 248880 268484
rect 248932 268472 248938 268524
rect 283190 268472 283196 268524
rect 283248 268512 283254 268524
rect 306374 268512 306380 268524
rect 283248 268484 306380 268512
rect 283248 268472 283254 268484
rect 306374 268472 306380 268484
rect 306432 268472 306438 268524
rect 317046 268472 317052 268524
rect 317104 268512 317110 268524
rect 396074 268512 396080 268524
rect 317104 268484 396080 268512
rect 317104 268472 317110 268484
rect 396074 268472 396080 268484
rect 396132 268472 396138 268524
rect 397178 268472 397184 268524
rect 397236 268512 397242 268524
rect 608594 268512 608600 268524
rect 397236 268484 608600 268512
rect 397236 268472 397242 268484
rect 608594 268472 608600 268484
rect 608652 268472 608658 268524
rect 69382 268404 69388 268456
rect 69440 268444 69446 268456
rect 193674 268444 193680 268456
rect 69440 268416 193680 268444
rect 69440 268404 69446 268416
rect 193674 268404 193680 268416
rect 193732 268404 193738 268456
rect 213454 268404 213460 268456
rect 213512 268444 213518 268456
rect 245746 268444 245752 268456
rect 213512 268416 245752 268444
rect 213512 268404 213518 268416
rect 245746 268404 245752 268416
rect 245804 268404 245810 268456
rect 245838 268404 245844 268456
rect 245896 268444 245902 268456
rect 259178 268444 259184 268456
rect 245896 268416 259184 268444
rect 245896 268404 245902 268416
rect 259178 268404 259184 268416
rect 259236 268404 259242 268456
rect 281442 268404 281448 268456
rect 281500 268444 281506 268456
rect 302234 268444 302240 268456
rect 281500 268416 302240 268444
rect 281500 268404 281506 268416
rect 302234 268404 302240 268416
rect 302292 268404 302298 268456
rect 319714 268404 319720 268456
rect 319772 268444 319778 268456
rect 398834 268444 398840 268456
rect 319772 268416 398840 268444
rect 319772 268404 319778 268416
rect 398834 268404 398840 268416
rect 398892 268404 398898 268456
rect 399846 268404 399852 268456
rect 399904 268444 399910 268456
rect 615678 268444 615684 268456
rect 399904 268416 615684 268444
rect 399904 268404 399910 268416
rect 615678 268404 615684 268416
rect 615736 268404 615742 268456
rect 66162 268336 66168 268388
rect 66220 268376 66226 268388
rect 192110 268376 192116 268388
rect 66220 268348 192116 268376
rect 66220 268336 66226 268348
rect 192110 268336 192116 268348
rect 192168 268336 192174 268388
rect 211246 268336 211252 268388
rect 211304 268376 211310 268388
rect 247126 268376 247132 268388
rect 211304 268348 247132 268376
rect 211304 268336 211310 268348
rect 247126 268336 247132 268348
rect 247184 268336 247190 268388
rect 257982 268336 257988 268388
rect 258040 268376 258046 268388
rect 264514 268376 264520 268388
rect 258040 268348 264520 268376
rect 258040 268336 258046 268348
rect 264514 268336 264520 268348
rect 264572 268336 264578 268388
rect 284110 268336 284116 268388
rect 284168 268376 284174 268388
rect 309134 268376 309140 268388
rect 284168 268348 309140 268376
rect 284168 268336 284174 268348
rect 309134 268336 309140 268348
rect 309192 268336 309198 268388
rect 318334 268336 318340 268388
rect 318392 268376 318398 268388
rect 400214 268376 400220 268388
rect 318392 268348 400220 268376
rect 318392 268336 318398 268348
rect 400214 268336 400220 268348
rect 400272 268336 400278 268388
rect 401134 268336 401140 268388
rect 401192 268376 401198 268388
rect 619634 268376 619640 268388
rect 401192 268348 619640 268376
rect 401192 268336 401198 268348
rect 619634 268336 619640 268348
rect 619692 268336 619698 268388
rect 106182 268268 106188 268320
rect 106240 268308 106246 268320
rect 207474 268308 207480 268320
rect 106240 268280 207480 268308
rect 106240 268268 106246 268280
rect 207474 268268 207480 268280
rect 207532 268268 207538 268320
rect 307662 268268 307668 268320
rect 307720 268308 307726 268320
rect 371326 268308 371332 268320
rect 307720 268280 371332 268308
rect 307720 268268 307726 268280
rect 371326 268268 371332 268280
rect 371384 268268 371390 268320
rect 372706 268268 372712 268320
rect 372764 268308 372770 268320
rect 391934 268308 391940 268320
rect 372764 268280 391940 268308
rect 372764 268268 372770 268280
rect 391934 268268 391940 268280
rect 391992 268268 391998 268320
rect 131022 268200 131028 268252
rect 131080 268240 131086 268252
rect 216858 268240 216864 268252
rect 131080 268212 216864 268240
rect 131080 268200 131086 268212
rect 216858 268200 216864 268212
rect 216916 268200 216922 268252
rect 339402 268200 339408 268252
rect 339460 268240 339466 268252
rect 382274 268240 382280 268252
rect 339460 268212 382280 268240
rect 339460 268200 339466 268212
rect 382274 268200 382280 268212
rect 382332 268200 382338 268252
rect 388162 268200 388168 268252
rect 388220 268240 388226 268252
rect 502242 268240 502248 268252
rect 388220 268212 502248 268240
rect 388220 268200 388226 268212
rect 502242 268200 502248 268212
rect 502300 268200 502306 268252
rect 135162 268132 135168 268184
rect 135220 268172 135226 268184
rect 218146 268172 218152 268184
rect 135220 268144 218152 268172
rect 135220 268132 135226 268144
rect 218146 268132 218152 268144
rect 218204 268132 218210 268184
rect 386506 268132 386512 268184
rect 386564 268172 386570 268184
rect 487154 268172 487160 268184
rect 386564 268144 487160 268172
rect 386564 268132 386570 268144
rect 487154 268132 487160 268144
rect 487212 268132 487218 268184
rect 186406 268064 186412 268116
rect 186464 268104 186470 268116
rect 237282 268104 237288 268116
rect 186464 268076 237288 268104
rect 186464 268064 186470 268076
rect 237282 268064 237288 268076
rect 237340 268064 237346 268116
rect 331122 268064 331128 268116
rect 331180 268104 331186 268116
rect 419534 268104 419540 268116
rect 331180 268076 419540 268104
rect 331180 268064 331186 268076
rect 419534 268064 419540 268076
rect 419592 268064 419598 268116
rect 663058 268064 663064 268116
rect 663116 268104 663122 268116
rect 676214 268104 676220 268116
rect 663116 268076 676220 268104
rect 663116 268064 663122 268076
rect 676214 268064 676220 268076
rect 676272 268064 676278 268116
rect 185026 267996 185032 268048
rect 185084 268036 185090 268048
rect 220354 268036 220360 268048
rect 185084 268008 220360 268036
rect 185084 267996 185090 268008
rect 220354 267996 220360 268008
rect 220412 267996 220418 268048
rect 385126 267996 385132 268048
rect 385184 268036 385190 268048
rect 474182 268036 474188 268048
rect 385184 268008 474188 268036
rect 385184 267996 385190 268008
rect 474182 267996 474188 268008
rect 474240 267996 474246 268048
rect 195974 267928 195980 267980
rect 196032 267968 196038 267980
rect 223022 267968 223028 267980
rect 196032 267940 223028 267968
rect 196032 267928 196038 267940
rect 223022 267928 223028 267940
rect 223080 267928 223086 267980
rect 322382 267928 322388 267980
rect 322440 267968 322446 267980
rect 407022 267968 407028 267980
rect 322440 267940 407028 267968
rect 322440 267928 322446 267940
rect 407022 267928 407028 267940
rect 407080 267928 407086 267980
rect 661862 267928 661868 267980
rect 661920 267968 661926 267980
rect 676214 267968 676220 267980
rect 661920 267940 676220 267968
rect 661920 267928 661926 267940
rect 676214 267928 676220 267940
rect 676272 267928 676278 267980
rect 343634 267860 343640 267912
rect 343692 267900 343698 267912
rect 426434 267900 426440 267912
rect 343692 267872 426440 267900
rect 343692 267860 343698 267872
rect 426434 267860 426440 267872
rect 426492 267860 426498 267912
rect 371878 267792 371884 267844
rect 371936 267832 371942 267844
rect 394694 267832 394700 267844
rect 371936 267804 394700 267832
rect 371936 267792 371942 267804
rect 394694 267792 394700 267804
rect 394752 267792 394758 267844
rect 409874 267792 409880 267844
rect 409932 267832 409938 267844
rect 412634 267832 412640 267844
rect 409932 267804 412640 267832
rect 409932 267792 409938 267804
rect 412634 267792 412640 267804
rect 412692 267792 412698 267844
rect 365714 267724 365720 267776
rect 365772 267764 365778 267776
rect 387794 267764 387800 267776
rect 365772 267736 387800 267764
rect 365772 267724 365778 267736
rect 387794 267724 387800 267736
rect 387852 267724 387858 267776
rect 390462 267724 390468 267776
rect 390520 267764 390526 267776
rect 523678 267764 523684 267776
rect 390520 267736 523684 267764
rect 390520 267724 390526 267736
rect 523678 267724 523684 267736
rect 523736 267724 523742 267776
rect 660298 267724 660304 267776
rect 660356 267764 660362 267776
rect 676122 267764 676128 267776
rect 660356 267736 676128 267764
rect 660356 267724 660362 267736
rect 676122 267724 676128 267736
rect 676180 267724 676186 267776
rect 175182 267656 175188 267708
rect 175240 267696 175246 267708
rect 233786 267696 233792 267708
rect 175240 267668 233792 267696
rect 175240 267656 175246 267668
rect 233786 267656 233792 267668
rect 233844 267656 233850 267708
rect 276474 267656 276480 267708
rect 276532 267696 276538 267708
rect 277302 267696 277308 267708
rect 276532 267668 277308 267696
rect 276532 267656 276538 267668
rect 277302 267656 277308 267668
rect 277360 267656 277366 267708
rect 287606 267656 287612 267708
rect 287664 267696 287670 267708
rect 288342 267696 288348 267708
rect 287664 267668 288348 267696
rect 287664 267656 287670 267668
rect 288342 267656 288348 267668
rect 288400 267656 288406 267708
rect 289814 267656 289820 267708
rect 289872 267696 289878 267708
rect 291102 267696 291108 267708
rect 289872 267668 291108 267696
rect 289872 267656 289878 267668
rect 291102 267656 291108 267668
rect 291160 267656 291166 267708
rect 299198 267656 299204 267708
rect 299256 267696 299262 267708
rect 309318 267696 309324 267708
rect 299256 267668 309324 267696
rect 299256 267656 299262 267668
rect 309318 267656 309324 267668
rect 309376 267656 309382 267708
rect 311710 267656 311716 267708
rect 311768 267696 311774 267708
rect 311768 267668 319668 267696
rect 311768 267656 311774 267668
rect 162118 267588 162124 267640
rect 162176 267628 162182 267640
rect 221734 267628 221740 267640
rect 162176 267600 221740 267628
rect 162176 267588 162182 267600
rect 221734 267588 221740 267600
rect 221792 267588 221798 267640
rect 231118 267588 231124 267640
rect 231176 267628 231182 267640
rect 235994 267628 236000 267640
rect 231176 267600 236000 267628
rect 231176 267588 231182 267600
rect 235994 267588 236000 267600
rect 236052 267588 236058 267640
rect 300578 267588 300584 267640
rect 300636 267628 300642 267640
rect 319438 267628 319444 267640
rect 300636 267600 319444 267628
rect 300636 267588 300642 267600
rect 319438 267588 319444 267600
rect 319496 267588 319502 267640
rect 144178 267520 144184 267572
rect 144236 267560 144242 267572
rect 204346 267560 204352 267572
rect 144236 267532 204352 267560
rect 144236 267520 144242 267532
rect 204346 267520 204352 267532
rect 204404 267520 204410 267572
rect 284938 267520 284944 267572
rect 284996 267560 285002 267572
rect 291838 267560 291844 267572
rect 284996 267532 291844 267560
rect 284996 267520 285002 267532
rect 291838 267520 291844 267532
rect 291896 267520 291902 267572
rect 295150 267520 295156 267572
rect 295208 267560 295214 267572
rect 319530 267560 319536 267572
rect 295208 267532 319536 267560
rect 295208 267520 295214 267532
rect 319530 267520 319536 267532
rect 319588 267520 319594 267572
rect 168282 267452 168288 267504
rect 168340 267492 168346 267504
rect 231118 267492 231124 267504
rect 168340 267464 231124 267492
rect 168340 267452 168346 267464
rect 231118 267452 231124 267464
rect 231176 267452 231182 267504
rect 287146 267452 287152 267504
rect 287204 267492 287210 267504
rect 301498 267492 301504 267504
rect 287204 267464 301504 267492
rect 287204 267452 287210 267464
rect 301498 267452 301504 267464
rect 301556 267452 301562 267504
rect 306374 267452 306380 267504
rect 306432 267492 306438 267504
rect 311158 267492 311164 267504
rect 306432 267464 311164 267492
rect 306432 267452 306438 267464
rect 311158 267452 311164 267464
rect 311216 267452 311222 267504
rect 311250 267452 311256 267504
rect 311308 267492 311314 267504
rect 316034 267492 316040 267504
rect 311308 267464 316040 267492
rect 311308 267452 311314 267464
rect 316034 267452 316040 267464
rect 316092 267452 316098 267504
rect 319640 267492 319668 267668
rect 344646 267656 344652 267708
rect 344704 267696 344710 267708
rect 469214 267696 469220 267708
rect 344704 267668 469220 267696
rect 344704 267656 344710 267668
rect 469214 267656 469220 267668
rect 469272 267656 469278 267708
rect 324130 267588 324136 267640
rect 324188 267628 324194 267640
rect 347038 267628 347044 267640
rect 324188 267600 347044 267628
rect 324188 267588 324194 267600
rect 347038 267588 347044 267600
rect 347096 267588 347102 267640
rect 349982 267588 349988 267640
rect 350040 267628 350046 267640
rect 483382 267628 483388 267640
rect 350040 267600 483388 267628
rect 350040 267588 350046 267600
rect 483382 267588 483388 267600
rect 483440 267588 483446 267640
rect 326798 267520 326804 267572
rect 326856 267560 326862 267572
rect 349798 267560 349804 267572
rect 326856 267532 349804 267560
rect 326856 267520 326862 267532
rect 349798 267520 349804 267532
rect 349856 267520 349862 267572
rect 352650 267520 352656 267572
rect 352708 267560 352714 267572
rect 491386 267560 491392 267572
rect 352708 267532 491392 267560
rect 352708 267520 352714 267532
rect 491386 267520 491392 267532
rect 491444 267520 491450 267572
rect 339402 267492 339408 267504
rect 319640 267464 339408 267492
rect 339402 267452 339408 267464
rect 339460 267452 339466 267504
rect 355318 267452 355324 267504
rect 355376 267492 355382 267504
rect 498194 267492 498200 267504
rect 355376 267464 498200 267492
rect 355376 267452 355382 267464
rect 498194 267452 498200 267464
rect 498252 267452 498258 267504
rect 161382 267384 161388 267436
rect 161440 267424 161446 267436
rect 228450 267424 228456 267436
rect 161440 267396 228456 267424
rect 161440 267384 161446 267396
rect 228450 267384 228456 267396
rect 228508 267384 228514 267436
rect 236638 267384 236644 267436
rect 236696 267424 236702 267436
rect 241790 267424 241796 267436
rect 236696 267396 241796 267424
rect 236696 267384 236702 267396
rect 241790 267384 241796 267396
rect 241848 267384 241854 267436
rect 278314 267384 278320 267436
rect 278372 267424 278378 267436
rect 281534 267424 281540 267436
rect 278372 267396 281540 267424
rect 278372 267384 278378 267396
rect 281534 267384 281540 267396
rect 281592 267384 281598 267436
rect 283650 267384 283656 267436
rect 283708 267424 283714 267436
rect 285582 267424 285588 267436
rect 283708 267396 285588 267424
rect 283708 267384 283714 267396
rect 285582 267384 285588 267396
rect 285640 267384 285646 267436
rect 298278 267384 298284 267436
rect 298336 267424 298342 267436
rect 327810 267424 327816 267436
rect 298336 267396 327816 267424
rect 298336 267384 298342 267396
rect 327810 267384 327816 267396
rect 327868 267384 327874 267436
rect 357986 267384 357992 267436
rect 358044 267424 358050 267436
rect 505094 267424 505100 267436
rect 358044 267396 505100 267424
rect 358044 267384 358050 267396
rect 505094 267384 505100 267396
rect 505152 267384 505158 267436
rect 125962 267316 125968 267368
rect 126020 267356 126026 267368
rect 207014 267356 207020 267368
rect 126020 267328 207020 267356
rect 126020 267316 126026 267328
rect 207014 267316 207020 267328
rect 207072 267316 207078 267368
rect 276014 267316 276020 267368
rect 276072 267356 276078 267368
rect 279418 267356 279424 267368
rect 276072 267328 279424 267356
rect 276072 267316 276078 267328
rect 279418 267316 279424 267328
rect 279476 267316 279482 267368
rect 288066 267316 288072 267368
rect 288124 267356 288130 267368
rect 297358 267356 297364 267368
rect 288124 267328 297364 267356
rect 288124 267316 288130 267328
rect 297358 267316 297364 267328
rect 297416 267316 297422 267368
rect 300946 267316 300952 267368
rect 301004 267356 301010 267368
rect 333238 267356 333244 267368
rect 301004 267328 333244 267356
rect 301004 267316 301010 267328
rect 333238 267316 333244 267328
rect 333296 267316 333302 267368
rect 360654 267316 360660 267368
rect 360712 267356 360718 267368
rect 511994 267356 512000 267368
rect 360712 267328 512000 267356
rect 360712 267316 360718 267328
rect 511994 267316 512000 267328
rect 512052 267316 512058 267368
rect 113174 267248 113180 267300
rect 113232 267288 113238 267300
rect 196342 267288 196348 267300
rect 113232 267260 196348 267288
rect 113232 267248 113238 267260
rect 196342 267248 196348 267260
rect 196400 267248 196406 267300
rect 196618 267248 196624 267300
rect 196676 267288 196682 267300
rect 217686 267288 217692 267300
rect 196676 267260 217692 267288
rect 196676 267248 196682 267260
rect 217686 267248 217692 267260
rect 217744 267248 217750 267300
rect 238110 267248 238116 267300
rect 238168 267288 238174 267300
rect 251082 267288 251088 267300
rect 238168 267260 251088 267288
rect 238168 267248 238174 267260
rect 251082 267248 251088 267260
rect 251140 267248 251146 267300
rect 281810 267248 281816 267300
rect 281868 267288 281874 267300
rect 286962 267288 286968 267300
rect 281868 267260 286968 267288
rect 281868 267248 281874 267260
rect 286962 267248 286968 267260
rect 287020 267248 287026 267300
rect 288526 267248 288532 267300
rect 288584 267288 288590 267300
rect 289630 267288 289636 267300
rect 288584 267260 289636 267288
rect 288584 267248 288590 267260
rect 289630 267248 289636 267260
rect 289688 267248 289694 267300
rect 292942 267248 292948 267300
rect 293000 267288 293006 267300
rect 293000 267260 308076 267288
rect 293000 267248 293006 267260
rect 110506 267180 110512 267232
rect 110564 267220 110570 267232
rect 199930 267220 199936 267232
rect 110564 267192 199936 267220
rect 110564 267180 110570 267192
rect 199930 267180 199936 267192
rect 199988 267180 199994 267232
rect 221458 267180 221464 267232
rect 221516 267220 221522 267232
rect 235074 267220 235080 267232
rect 221516 267192 235080 267220
rect 221516 267180 221522 267192
rect 235074 267180 235080 267192
rect 235132 267180 235138 267232
rect 235902 267180 235908 267232
rect 235960 267220 235966 267232
rect 256050 267220 256056 267232
rect 235960 267192 256056 267220
rect 235960 267180 235966 267192
rect 256050 267180 256056 267192
rect 256108 267180 256114 267232
rect 272518 267180 272524 267232
rect 272576 267220 272582 267232
rect 277854 267220 277860 267232
rect 272576 267192 277860 267220
rect 272576 267180 272582 267192
rect 277854 267180 277860 267192
rect 277912 267180 277918 267232
rect 290274 267180 290280 267232
rect 290332 267220 290338 267232
rect 307018 267220 307024 267232
rect 290332 267192 307024 267220
rect 290332 267180 290338 267192
rect 307018 267180 307024 267192
rect 307076 267180 307082 267232
rect 308048 267220 308076 267260
rect 309318 267248 309324 267300
rect 309376 267288 309382 267300
rect 317782 267288 317788 267300
rect 309376 267260 317788 267288
rect 309376 267248 309382 267260
rect 317782 267248 317788 267260
rect 317840 267248 317846 267300
rect 317874 267248 317880 267300
rect 317932 267288 317938 267300
rect 360838 267288 360844 267300
rect 317932 267260 360844 267288
rect 317932 267248 317938 267260
rect 360838 267248 360844 267260
rect 360896 267248 360902 267300
rect 363322 267248 363328 267300
rect 363380 267288 363386 267300
rect 518894 267288 518900 267300
rect 363380 267260 518900 267288
rect 363380 267248 363386 267260
rect 518894 267248 518900 267260
rect 518952 267248 518958 267300
rect 309778 267220 309784 267232
rect 308048 267192 309784 267220
rect 309778 267180 309784 267192
rect 309836 267180 309842 267232
rect 313918 267180 313924 267232
rect 313976 267220 313982 267232
rect 316034 267220 316040 267232
rect 313976 267192 316040 267220
rect 313976 267180 313982 267192
rect 316034 267180 316040 267192
rect 316092 267180 316098 267232
rect 316126 267180 316132 267232
rect 316184 267220 316190 267232
rect 353294 267220 353300 267232
rect 316184 267192 353300 267220
rect 316184 267180 316190 267192
rect 353294 267180 353300 267192
rect 353352 267180 353358 267232
rect 363598 267220 363604 267232
rect 354646 267192 363604 267220
rect 119614 267112 119620 267164
rect 119672 267152 119678 267164
rect 209682 267152 209688 267164
rect 119672 267124 209688 267152
rect 119672 267112 119678 267124
rect 209682 267112 209688 267124
rect 209740 267112 209746 267164
rect 226978 267112 226984 267164
rect 227036 267152 227042 267164
rect 232406 267152 232412 267164
rect 227036 267124 232412 267152
rect 227036 267112 227042 267124
rect 232406 267112 232412 267124
rect 232464 267112 232470 267164
rect 233142 267112 233148 267164
rect 233200 267152 233206 267164
rect 255130 267152 255136 267164
rect 233200 267124 255136 267152
rect 233200 267112 233206 267124
rect 255130 267112 255136 267124
rect 255188 267112 255194 267164
rect 255222 267112 255228 267164
rect 255280 267152 255286 267164
rect 263594 267152 263600 267164
rect 255280 267124 263600 267152
rect 255280 267112 255286 267124
rect 263594 267112 263600 267124
rect 263652 267112 263658 267164
rect 286318 267112 286324 267164
rect 286376 267152 286382 267164
rect 305638 267152 305644 267164
rect 286376 267124 305644 267152
rect 286376 267112 286382 267124
rect 305638 267112 305644 267124
rect 305696 267112 305702 267164
rect 309244 267124 309456 267152
rect 93118 267044 93124 267096
rect 93176 267084 93182 267096
rect 201218 267084 201224 267096
rect 93176 267056 201224 267084
rect 93176 267044 93182 267056
rect 201218 267044 201224 267056
rect 201276 267044 201282 267096
rect 214558 267044 214564 267096
rect 214616 267084 214622 267096
rect 237742 267084 237748 267096
rect 214616 267056 237748 267084
rect 214616 267044 214622 267056
rect 237742 267044 237748 267056
rect 237800 267044 237806 267096
rect 238662 267044 238668 267096
rect 238720 267084 238726 267096
rect 257338 267084 257344 267096
rect 238720 267056 257344 267084
rect 238720 267044 238726 267056
rect 257338 267044 257344 267056
rect 257396 267044 257402 267096
rect 289446 267044 289452 267096
rect 289504 267084 289510 267096
rect 306374 267084 306380 267096
rect 289504 267056 306380 267084
rect 289504 267044 289510 267056
rect 306374 267044 306380 267056
rect 306432 267044 306438 267096
rect 71774 266976 71780 267028
rect 71832 267016 71838 267028
rect 194134 267016 194140 267028
rect 71832 266988 194140 267016
rect 71832 266976 71838 266988
rect 194134 266976 194140 266988
rect 194192 266976 194198 267028
rect 210418 266976 210424 267028
rect 210476 267016 210482 267028
rect 239122 267016 239128 267028
rect 210476 266988 239128 267016
rect 210476 266976 210482 266988
rect 239122 266976 239128 266988
rect 239180 266976 239186 267028
rect 252370 266976 252376 267028
rect 252428 267016 252434 267028
rect 262214 267016 262220 267028
rect 252428 266988 262220 267016
rect 252428 266976 252434 266988
rect 262214 266976 262220 266988
rect 262272 266976 262278 267028
rect 272426 266976 272432 267028
rect 272484 267016 272490 267028
rect 277762 267016 277768 267028
rect 272484 266988 277768 267016
rect 272484 266976 272490 266988
rect 277762 266976 277768 266988
rect 277820 266976 277826 267028
rect 279602 266976 279608 267028
rect 279660 267016 279666 267028
rect 287698 267016 287704 267028
rect 279660 266988 287704 267016
rect 279660 266976 279666 266988
rect 287698 266976 287704 266988
rect 287756 266976 287762 267028
rect 291194 266976 291200 267028
rect 291252 267016 291258 267028
rect 309244 267016 309272 267124
rect 309428 267084 309456 267124
rect 315206 267112 315212 267164
rect 315264 267152 315270 267164
rect 354646 267152 354674 267192
rect 363598 267180 363604 267192
rect 363656 267180 363662 267232
rect 365714 267220 365720 267232
rect 364306 267192 365720 267220
rect 315264 267124 354674 267152
rect 315264 267112 315270 267124
rect 356238 267112 356244 267164
rect 356296 267152 356302 267164
rect 357250 267152 357256 267164
rect 356296 267124 357256 267152
rect 356296 267112 356302 267124
rect 357250 267112 357256 267124
rect 357308 267112 357314 267164
rect 358906 267112 358912 267164
rect 358964 267152 358970 267164
rect 360102 267152 360108 267164
rect 358964 267124 360108 267152
rect 358964 267112 358970 267124
rect 360102 267112 360108 267124
rect 360160 267112 360166 267164
rect 362034 267112 362040 267164
rect 362092 267152 362098 267164
rect 362678 267152 362684 267164
rect 362092 267124 362684 267152
rect 362092 267112 362098 267124
rect 362678 267112 362684 267124
rect 362736 267112 362742 267164
rect 315390 267084 315396 267096
rect 309428 267056 315396 267084
rect 315390 267044 315396 267056
rect 315448 267044 315454 267096
rect 316034 267044 316040 267096
rect 316092 267084 316098 267096
rect 364306 267084 364334 267192
rect 365714 267180 365720 267192
rect 365772 267180 365778 267232
rect 365990 267180 365996 267232
rect 366048 267220 366054 267232
rect 525794 267220 525800 267232
rect 366048 267192 525800 267220
rect 366048 267180 366054 267192
rect 525794 267180 525800 267192
rect 525852 267180 525858 267232
rect 368658 267112 368664 267164
rect 368716 267152 368722 267164
rect 532878 267152 532884 267164
rect 368716 267124 532884 267152
rect 368716 267112 368722 267124
rect 532878 267112 532884 267124
rect 532936 267112 532942 267164
rect 316092 267056 364334 267084
rect 316092 267044 316098 267056
rect 371326 267044 371332 267096
rect 371384 267084 371390 267096
rect 540974 267084 540980 267096
rect 371384 267056 540980 267084
rect 371384 267044 371390 267056
rect 540974 267044 540980 267056
rect 541032 267044 541038 267096
rect 312446 267016 312452 267028
rect 291252 266988 309272 267016
rect 309428 266988 312452 267016
rect 291252 266976 291258 266988
rect 182082 266908 182088 266960
rect 182140 266948 182146 266960
rect 236454 266948 236460 266960
rect 182140 266920 236460 266948
rect 182140 266908 182146 266920
rect 236454 266908 236460 266920
rect 236512 266908 236518 266960
rect 153838 266840 153844 266892
rect 153896 266880 153902 266892
rect 203058 266880 203064 266892
rect 153896 266852 203064 266880
rect 153896 266840 153902 266852
rect 203058 266840 203064 266852
rect 203116 266840 203122 266892
rect 152458 266772 152464 266824
rect 152516 266812 152522 266824
rect 197722 266812 197728 266824
rect 152516 266784 197728 266812
rect 152516 266772 152522 266784
rect 197722 266772 197728 266784
rect 197780 266772 197786 266824
rect 296990 266772 296996 266824
rect 297048 266812 297054 266824
rect 309428 266812 309456 266988
rect 312446 266976 312452 266988
rect 312504 266976 312510 267028
rect 316586 266976 316592 267028
rect 316644 267016 316650 267028
rect 371878 267016 371884 267028
rect 316644 266988 371884 267016
rect 316644 266976 316650 266988
rect 371878 266976 371884 266988
rect 371936 266976 371942 267028
rect 375374 266976 375380 267028
rect 375432 267016 375438 267028
rect 376662 267016 376668 267028
rect 375432 266988 376668 267016
rect 375432 266976 375438 266988
rect 376662 266976 376668 266988
rect 376720 266976 376726 267028
rect 382458 266976 382464 267028
rect 382516 267016 382522 267028
rect 383470 267016 383476 267028
rect 382516 266988 383476 267016
rect 382516 266976 382522 266988
rect 383470 266976 383476 266988
rect 383528 266976 383534 267028
rect 397638 266976 397644 267028
rect 397696 267016 397702 267028
rect 398650 267016 398656 267028
rect 397696 266988 398656 267016
rect 397696 266976 397702 266988
rect 398650 266976 398656 266988
rect 398708 266976 398714 267028
rect 399018 266976 399024 267028
rect 399076 267016 399082 267028
rect 409874 267016 409880 267028
rect 399076 266988 409880 267016
rect 399076 266976 399082 266988
rect 409874 266976 409880 266988
rect 409932 266976 409938 267028
rect 417418 266976 417424 267028
rect 417476 267016 417482 267028
rect 643094 267016 643100 267028
rect 417476 266988 643100 267016
rect 417476 266976 417482 266988
rect 643094 266976 643100 266988
rect 643152 266976 643158 267028
rect 673914 266976 673920 267028
rect 673972 267016 673978 267028
rect 676030 267016 676036 267028
rect 673972 266988 676036 267016
rect 673972 266976 673978 266988
rect 676030 266976 676036 266988
rect 676088 266976 676094 267028
rect 322198 266948 322204 266960
rect 297048 266784 309456 266812
rect 311176 266920 322204 266948
rect 297048 266772 297054 266784
rect 184750 266704 184756 266756
rect 184808 266744 184814 266756
rect 219066 266744 219072 266756
rect 184808 266716 219072 266744
rect 184808 266704 184814 266716
rect 219066 266704 219072 266716
rect 219124 266704 219130 266756
rect 282270 266704 282276 266756
rect 282328 266744 282334 266756
rect 288434 266744 288440 266756
rect 282328 266716 288440 266744
rect 282328 266704 282334 266716
rect 288434 266704 288440 266716
rect 288492 266704 288498 266756
rect 192478 266636 192484 266688
rect 192536 266676 192542 266688
rect 225782 266676 225788 266688
rect 192536 266648 225788 266676
rect 192536 266636 192542 266648
rect 225782 266636 225788 266648
rect 225840 266636 225846 266688
rect 305914 266636 305920 266688
rect 305972 266676 305978 266688
rect 311176 266676 311204 266920
rect 322198 266908 322204 266920
rect 322256 266908 322262 266960
rect 324590 266908 324596 266960
rect 324648 266948 324654 266960
rect 327718 266948 327724 266960
rect 324648 266920 327724 266948
rect 324648 266908 324654 266920
rect 327718 266908 327724 266920
rect 327776 266908 327782 266960
rect 328178 266908 328184 266960
rect 328236 266948 328242 266960
rect 343634 266948 343640 266960
rect 328236 266920 343640 266948
rect 328236 266908 328242 266920
rect 343634 266908 343640 266920
rect 343692 266908 343698 266960
rect 347314 266908 347320 266960
rect 347372 266948 347378 266960
rect 470686 266948 470692 266960
rect 347372 266920 470692 266948
rect 347372 266908 347378 266920
rect 470686 266908 470692 266920
rect 470744 266908 470750 266960
rect 323670 266880 323676 266892
rect 305972 266648 311204 266676
rect 311268 266852 323676 266880
rect 305972 266636 305978 266648
rect 271598 266568 271604 266620
rect 271656 266608 271662 266620
rect 276290 266608 276296 266620
rect 271656 266580 276296 266608
rect 271656 266568 271662 266580
rect 276290 266568 276296 266580
rect 276348 266568 276354 266620
rect 277854 266568 277860 266620
rect 277912 266608 277918 266620
rect 283558 266608 283564 266620
rect 277912 266580 283564 266608
rect 277912 266568 277918 266580
rect 283558 266568 283564 266580
rect 283616 266568 283622 266620
rect 308582 266568 308588 266620
rect 308640 266608 308646 266620
rect 311268 266608 311296 266852
rect 323670 266840 323676 266852
rect 323728 266840 323734 266892
rect 341978 266840 341984 266892
rect 342036 266880 342042 266892
rect 462314 266880 462320 266892
rect 342036 266852 462320 266880
rect 342036 266840 342042 266852
rect 462314 266840 462320 266852
rect 462372 266840 462378 266892
rect 339310 266772 339316 266824
rect 339368 266812 339374 266824
rect 455414 266812 455420 266824
rect 339368 266784 455420 266812
rect 339368 266772 339374 266784
rect 455414 266772 455420 266784
rect 455472 266772 455478 266824
rect 312538 266704 312544 266756
rect 312596 266744 312602 266756
rect 312596 266716 316034 266744
rect 312596 266704 312602 266716
rect 316006 266676 316034 266716
rect 335262 266704 335268 266756
rect 335320 266744 335326 266756
rect 444374 266744 444380 266756
rect 335320 266716 444380 266744
rect 335320 266704 335326 266716
rect 444374 266704 444380 266716
rect 444432 266704 444438 266756
rect 326338 266676 326344 266688
rect 316006 266648 326344 266676
rect 326338 266636 326344 266648
rect 326396 266636 326402 266688
rect 329926 266636 329932 266688
rect 329984 266676 329990 266688
rect 329984 266648 331260 266676
rect 329984 266636 329990 266648
rect 308640 266580 311296 266608
rect 308640 266568 308646 266580
rect 325970 266568 325976 266620
rect 326028 266608 326034 266620
rect 331122 266608 331128 266620
rect 326028 266580 331128 266608
rect 326028 266568 326034 266580
rect 331122 266568 331128 266580
rect 331180 266568 331186 266620
rect 331232 266608 331260 266648
rect 332594 266636 332600 266688
rect 332652 266676 332658 266688
rect 431218 266676 431224 266688
rect 332652 266648 431224 266676
rect 332652 266636 332658 266648
rect 431218 266636 431224 266648
rect 431276 266636 431282 266688
rect 422938 266608 422944 266620
rect 331232 266580 422944 266608
rect 422938 266568 422944 266580
rect 422996 266568 423002 266620
rect 673362 266568 673368 266620
rect 673420 266608 673426 266620
rect 676214 266608 676220 266620
rect 673420 266580 676220 266608
rect 673420 266568 673426 266580
rect 676214 266568 676220 266580
rect 676272 266568 676278 266620
rect 271138 266500 271144 266552
rect 271196 266540 271202 266552
rect 274634 266540 274640 266552
rect 271196 266512 274640 266540
rect 271196 266500 271202 266512
rect 274634 266500 274640 266512
rect 274692 266500 274698 266552
rect 323210 266500 323216 266552
rect 323268 266540 323274 266552
rect 399018 266540 399024 266552
rect 323268 266512 399024 266540
rect 323268 266500 323274 266512
rect 399018 266500 399024 266512
rect 399076 266500 399082 266552
rect 408466 266512 409828 266540
rect 239398 266432 239404 266484
rect 239456 266472 239462 266484
rect 244458 266472 244464 266484
rect 239456 266444 244464 266472
rect 239456 266432 239462 266444
rect 244458 266432 244464 266444
rect 244516 266432 244522 266484
rect 270678 266432 270684 266484
rect 270736 266472 270742 266484
rect 273254 266472 273260 266484
rect 270736 266444 273260 266472
rect 270736 266432 270742 266444
rect 273254 266432 273260 266444
rect 273312 266432 273318 266484
rect 291654 266432 291660 266484
rect 291712 266472 291718 266484
rect 295978 266472 295984 266484
rect 291712 266444 295984 266472
rect 291712 266432 291718 266444
rect 295978 266432 295984 266444
rect 296036 266432 296042 266484
rect 304994 266432 305000 266484
rect 305052 266472 305058 266484
rect 306282 266472 306288 266484
rect 305052 266444 306288 266472
rect 305052 266432 305058 266444
rect 306282 266432 306288 266444
rect 306340 266432 306346 266484
rect 309870 266432 309876 266484
rect 309928 266472 309934 266484
rect 314286 266472 314292 266484
rect 309928 266444 314292 266472
rect 309928 266432 309934 266444
rect 314286 266432 314292 266444
rect 314344 266432 314350 266484
rect 320174 266432 320180 266484
rect 320232 266472 320238 266484
rect 321370 266472 321376 266484
rect 320232 266444 321376 266472
rect 320232 266432 320238 266444
rect 321370 266432 321376 266444
rect 321428 266432 321434 266484
rect 328638 266432 328644 266484
rect 328696 266472 328702 266484
rect 329650 266472 329656 266484
rect 328696 266444 329656 266472
rect 328696 266432 328702 266444
rect 329650 266432 329656 266444
rect 329708 266432 329714 266484
rect 408466 266472 408494 266512
rect 329852 266444 408494 266472
rect 233878 266364 233884 266416
rect 233936 266404 233942 266416
rect 234614 266404 234620 266416
rect 233936 266376 234620 266404
rect 233936 266364 233942 266376
rect 234614 266364 234620 266376
rect 234672 266364 234678 266416
rect 235350 266364 235356 266416
rect 235408 266404 235414 266416
rect 238662 266404 238668 266416
rect 235408 266376 238668 266404
rect 235408 266364 235414 266376
rect 238662 266364 238668 266376
rect 238720 266364 238726 266416
rect 242802 266364 242808 266416
rect 242860 266404 242866 266416
rect 249794 266404 249800 266416
rect 242860 266376 249800 266404
rect 242860 266364 242866 266376
rect 249794 266364 249800 266376
rect 249852 266364 249858 266416
rect 270310 266364 270316 266416
rect 270368 266404 270374 266416
rect 272058 266404 272064 266416
rect 270368 266376 272064 266404
rect 270368 266364 270374 266376
rect 272058 266364 272064 266376
rect 272116 266364 272122 266416
rect 284478 266364 284484 266416
rect 284536 266404 284542 266416
rect 289906 266404 289912 266416
rect 284536 266376 289912 266404
rect 284536 266364 284542 266376
rect 289906 266364 289912 266376
rect 289964 266364 289970 266416
rect 294322 266364 294328 266416
rect 294380 266404 294386 266416
rect 295242 266404 295248 266416
rect 294380 266376 295248 266404
rect 294380 266364 294386 266376
rect 295242 266364 295248 266376
rect 295300 266364 295306 266416
rect 295610 266364 295616 266416
rect 295668 266404 295674 266416
rect 296438 266404 296444 266416
rect 295668 266376 296444 266404
rect 295668 266364 295674 266376
rect 296438 266364 296444 266376
rect 296496 266364 296502 266416
rect 299658 266364 299664 266416
rect 299716 266404 299722 266416
rect 300762 266404 300768 266416
rect 299716 266376 300768 266404
rect 299716 266364 299722 266376
rect 300762 266364 300768 266376
rect 300820 266364 300826 266416
rect 302326 266364 302332 266416
rect 302384 266404 302390 266416
rect 303430 266404 303436 266416
rect 302384 266376 303436 266404
rect 302384 266364 302390 266376
rect 303430 266364 303436 266376
rect 303488 266364 303494 266416
rect 305454 266364 305460 266416
rect 305512 266404 305518 266416
rect 306190 266404 306196 266416
rect 305512 266376 306196 266404
rect 305512 266364 305518 266376
rect 306190 266364 306196 266376
rect 306248 266364 306254 266416
rect 306742 266364 306748 266416
rect 306800 266404 306806 266416
rect 307478 266404 307484 266416
rect 306800 266376 307484 266404
rect 306800 266364 306806 266376
rect 307478 266364 307484 266376
rect 307536 266364 307542 266416
rect 308122 266364 308128 266416
rect 308180 266404 308186 266416
rect 308950 266404 308956 266416
rect 308180 266376 308956 266404
rect 308180 266364 308186 266376
rect 308950 266364 308956 266376
rect 309008 266364 309014 266416
rect 309410 266364 309416 266416
rect 309468 266404 309474 266416
rect 310330 266404 310336 266416
rect 309468 266376 310336 266404
rect 309468 266364 309474 266376
rect 310330 266364 310336 266376
rect 310388 266364 310394 266416
rect 310790 266364 310796 266416
rect 310848 266404 310854 266416
rect 311802 266404 311808 266416
rect 310848 266376 311808 266404
rect 310848 266364 310854 266376
rect 311802 266364 311808 266376
rect 311860 266364 311866 266416
rect 312078 266364 312084 266416
rect 312136 266404 312142 266416
rect 313090 266404 313096 266416
rect 312136 266376 313096 266404
rect 312136 266364 312142 266376
rect 313090 266364 313096 266376
rect 313148 266364 313154 266416
rect 313458 266364 313464 266416
rect 313516 266404 313522 266416
rect 314470 266404 314476 266416
rect 313516 266376 314476 266404
rect 313516 266364 313522 266376
rect 314470 266364 314476 266376
rect 314528 266364 314534 266416
rect 314838 266364 314844 266416
rect 314896 266404 314902 266416
rect 315850 266404 315856 266416
rect 314896 266376 315856 266404
rect 314896 266364 314902 266376
rect 315850 266364 315856 266376
rect 315908 266364 315914 266416
rect 316126 266364 316132 266416
rect 316184 266404 316190 266416
rect 317230 266404 317236 266416
rect 316184 266376 317236 266404
rect 316184 266364 316190 266376
rect 317230 266364 317236 266376
rect 317288 266364 317294 266416
rect 317506 266364 317512 266416
rect 317564 266404 317570 266416
rect 318610 266404 318616 266416
rect 317564 266376 318616 266404
rect 317564 266364 317570 266376
rect 318610 266364 318616 266376
rect 318668 266364 318674 266416
rect 318794 266364 318800 266416
rect 318852 266404 318858 266416
rect 319898 266404 319904 266416
rect 318852 266376 319904 266404
rect 318852 266364 318858 266376
rect 319898 266364 319904 266376
rect 319956 266364 319962 266416
rect 320542 266364 320548 266416
rect 320600 266404 320606 266416
rect 321278 266404 321284 266416
rect 320600 266376 321284 266404
rect 320600 266364 320606 266376
rect 321278 266364 321284 266376
rect 321336 266364 321342 266416
rect 321922 266364 321928 266416
rect 321980 266404 321986 266416
rect 322750 266404 322756 266416
rect 321980 266376 322756 266404
rect 321980 266364 321986 266376
rect 322750 266364 322756 266376
rect 322808 266364 322814 266416
rect 327258 266364 327264 266416
rect 327316 266404 327322 266416
rect 327316 266376 328960 266404
rect 327316 266364 327322 266376
rect 328932 266336 328960 266376
rect 329006 266364 329012 266416
rect 329064 266404 329070 266416
rect 329742 266404 329748 266416
rect 329064 266376 329748 266404
rect 329064 266364 329070 266376
rect 329742 266364 329748 266376
rect 329800 266364 329806 266416
rect 329852 266336 329880 266444
rect 408770 266432 408776 266484
rect 408828 266472 408834 266484
rect 409690 266472 409696 266484
rect 408828 266444 409696 266472
rect 408828 266432 408834 266444
rect 409690 266432 409696 266444
rect 409748 266432 409754 266484
rect 409800 266472 409828 266512
rect 410058 266500 410064 266552
rect 410116 266540 410122 266552
rect 417418 266540 417424 266552
rect 410116 266512 417424 266540
rect 410116 266500 410122 266512
rect 417418 266500 417424 266512
rect 417476 266500 417482 266552
rect 410426 266472 410432 266484
rect 409800 266444 410432 266472
rect 410426 266432 410432 266444
rect 410484 266432 410490 266484
rect 411438 266432 411444 266484
rect 411496 266472 411502 266484
rect 412542 266472 412548 266484
rect 411496 266444 412548 266472
rect 411496 266432 411502 266444
rect 412542 266432 412548 266444
rect 412600 266432 412606 266484
rect 673270 266432 673276 266484
rect 673328 266472 673334 266484
rect 676214 266472 676220 266484
rect 673328 266444 676220 266472
rect 673328 266432 673334 266444
rect 676214 266432 676220 266444
rect 676272 266432 676278 266484
rect 331306 266364 331312 266416
rect 331364 266404 331370 266416
rect 332318 266404 332324 266416
rect 331364 266376 332324 266404
rect 331364 266364 331370 266376
rect 332318 266364 332324 266376
rect 332376 266364 332382 266416
rect 333974 266364 333980 266416
rect 334032 266404 334038 266416
rect 335170 266404 335176 266416
rect 334032 266376 335176 266404
rect 334032 266364 334038 266376
rect 335170 266364 335176 266376
rect 335228 266364 335234 266416
rect 340138 266364 340144 266416
rect 340196 266404 340202 266416
rect 340690 266404 340696 266416
rect 340196 266376 340696 266404
rect 340196 266364 340202 266376
rect 340690 266364 340696 266376
rect 340748 266364 340754 266416
rect 342806 266364 342812 266416
rect 342864 266404 342870 266416
rect 343450 266404 343456 266416
rect 342864 266376 343456 266404
rect 342864 266364 342870 266376
rect 343450 266364 343456 266376
rect 343508 266364 343514 266416
rect 345474 266364 345480 266416
rect 345532 266404 345538 266416
rect 346210 266404 346216 266416
rect 345532 266376 346216 266404
rect 345532 266364 345538 266376
rect 346210 266364 346216 266376
rect 346268 266364 346274 266416
rect 346854 266364 346860 266416
rect 346912 266404 346918 266416
rect 347682 266404 347688 266416
rect 346912 266376 347688 266404
rect 346912 266364 346918 266376
rect 347682 266364 347688 266376
rect 347740 266364 347746 266416
rect 347774 266364 347780 266416
rect 347832 266404 347838 266416
rect 349062 266404 349068 266416
rect 347832 266376 349068 266404
rect 347832 266364 347838 266376
rect 349062 266364 349068 266376
rect 349120 266364 349126 266416
rect 349522 266364 349528 266416
rect 349580 266404 349586 266416
rect 350350 266404 350356 266416
rect 349580 266376 350356 266404
rect 349580 266364 349586 266376
rect 350350 266364 350356 266376
rect 350408 266364 350414 266416
rect 350902 266364 350908 266416
rect 350960 266404 350966 266416
rect 351730 266404 351736 266416
rect 350960 266376 351736 266404
rect 350960 266364 350966 266376
rect 351730 266364 351736 266376
rect 351788 266364 351794 266416
rect 352190 266364 352196 266416
rect 352248 266404 352254 266416
rect 353018 266404 353024 266416
rect 352248 266376 353024 266404
rect 352248 266364 352254 266376
rect 353018 266364 353024 266376
rect 353076 266364 353082 266416
rect 356606 266364 356612 266416
rect 356664 266404 356670 266416
rect 357342 266404 357348 266416
rect 356664 266376 357348 266404
rect 356664 266364 356670 266376
rect 357342 266364 357348 266376
rect 357400 266364 357406 266416
rect 357526 266364 357532 266416
rect 357584 266404 357590 266416
rect 358630 266404 358636 266416
rect 357584 266376 358636 266404
rect 357584 266364 357590 266376
rect 358630 266364 358636 266376
rect 358688 266364 358694 266416
rect 359366 266364 359372 266416
rect 359424 266404 359430 266416
rect 360010 266404 360016 266416
rect 359424 266376 360016 266404
rect 359424 266364 359430 266376
rect 360010 266364 360016 266376
rect 360068 266364 360074 266416
rect 362402 266364 362408 266416
rect 362460 266404 362466 266416
rect 362770 266404 362776 266416
rect 362460 266376 362776 266404
rect 362460 266364 362466 266376
rect 362770 266364 362776 266376
rect 362828 266364 362834 266416
rect 364702 266364 364708 266416
rect 364760 266404 364766 266416
rect 365530 266404 365536 266416
rect 364760 266376 365536 266404
rect 364760 266364 364766 266376
rect 365530 266364 365536 266376
rect 365588 266364 365594 266416
rect 366450 266364 366456 266416
rect 366508 266404 366514 266416
rect 367002 266404 367008 266416
rect 366508 266376 367008 266404
rect 366508 266364 366514 266376
rect 367002 266364 367008 266376
rect 367060 266364 367066 266416
rect 367370 266364 367376 266416
rect 367428 266404 367434 266416
rect 368382 266404 368388 266416
rect 367428 266376 368388 266404
rect 367428 266364 367434 266376
rect 368382 266364 368388 266376
rect 368440 266364 368446 266416
rect 370038 266364 370044 266416
rect 370096 266404 370102 266416
rect 371050 266404 371056 266416
rect 370096 266376 371056 266404
rect 370096 266364 370102 266376
rect 371050 266364 371056 266376
rect 371108 266364 371114 266416
rect 376478 266364 376484 266416
rect 376536 266404 376542 266416
rect 376662 266404 376668 266416
rect 376536 266376 376668 266404
rect 376536 266364 376542 266376
rect 376662 266364 376668 266376
rect 376720 266364 376726 266416
rect 378870 266364 378876 266416
rect 378928 266404 378934 266416
rect 379422 266404 379428 266416
rect 378928 266376 379428 266404
rect 378928 266364 378934 266376
rect 379422 266364 379428 266376
rect 379480 266364 379486 266416
rect 379790 266364 379796 266416
rect 379848 266404 379854 266416
rect 380802 266404 380808 266416
rect 379848 266376 380808 266404
rect 379848 266364 379854 266376
rect 380802 266364 380808 266376
rect 380860 266364 380866 266416
rect 382918 266364 382924 266416
rect 382976 266404 382982 266416
rect 383562 266404 383568 266416
rect 382976 266376 383568 266404
rect 382976 266364 382982 266376
rect 383562 266364 383568 266376
rect 383620 266364 383626 266416
rect 390922 266364 390928 266416
rect 390980 266404 390986 266416
rect 391750 266404 391756 266416
rect 390980 266376 391756 266404
rect 390980 266364 390986 266376
rect 391750 266364 391756 266376
rect 391808 266364 391814 266416
rect 392302 266364 392308 266416
rect 392360 266404 392366 266416
rect 393130 266404 393136 266416
rect 392360 266376 393136 266404
rect 392360 266364 392366 266376
rect 393130 266364 393136 266376
rect 393188 266364 393194 266416
rect 393590 266364 393596 266416
rect 393648 266404 393654 266416
rect 394418 266404 394424 266416
rect 393648 266376 394424 266404
rect 393648 266364 393654 266376
rect 394418 266364 394424 266376
rect 394476 266364 394482 266416
rect 396258 266364 396264 266416
rect 396316 266404 396322 266416
rect 397270 266404 397276 266416
rect 396316 266376 397276 266404
rect 396316 266364 396322 266376
rect 397270 266364 397276 266376
rect 397328 266364 397334 266416
rect 398098 266364 398104 266416
rect 398156 266404 398162 266416
rect 398742 266404 398748 266416
rect 398156 266376 398748 266404
rect 398156 266364 398162 266376
rect 398742 266364 398748 266376
rect 398800 266364 398806 266416
rect 409230 266364 409236 266416
rect 409288 266404 409294 266416
rect 409782 266404 409788 266416
rect 409288 266376 409788 266404
rect 409288 266364 409294 266376
rect 409782 266364 409788 266376
rect 409840 266364 409846 266416
rect 410518 266364 410524 266416
rect 410576 266404 410582 266416
rect 451366 266404 451372 266416
rect 410576 266376 451372 266404
rect 410576 266364 410582 266376
rect 451366 266364 451372 266376
rect 451424 266364 451430 266416
rect 328932 266308 329880 266336
rect 354398 266296 354404 266348
rect 354456 266336 354462 266348
rect 495434 266336 495440 266348
rect 354456 266308 495440 266336
rect 354456 266296 354462 266308
rect 495434 266296 495440 266308
rect 495492 266296 495498 266348
rect 357066 266228 357072 266280
rect 357124 266268 357130 266280
rect 502334 266268 502340 266280
rect 357124 266240 502340 266268
rect 357124 266228 357130 266240
rect 502334 266228 502340 266240
rect 502392 266228 502398 266280
rect 373166 266160 373172 266212
rect 373224 266200 373230 266212
rect 545114 266200 545120 266212
rect 373224 266172 545120 266200
rect 373224 266160 373230 266172
rect 545114 266160 545120 266172
rect 545172 266160 545178 266212
rect 374454 266092 374460 266144
rect 374512 266132 374518 266144
rect 549254 266132 549260 266144
rect 374512 266104 549260 266132
rect 374512 266092 374518 266104
rect 549254 266092 549260 266104
rect 549312 266092 549318 266144
rect 375834 266024 375840 266076
rect 375892 266064 375898 266076
rect 552014 266064 552020 266076
rect 375892 266036 552020 266064
rect 375892 266024 375898 266036
rect 552014 266024 552020 266036
rect 552072 266024 552078 266076
rect 674006 266024 674012 266076
rect 674064 266064 674070 266076
rect 676214 266064 676220 266076
rect 674064 266036 676220 266064
rect 674064 266024 674070 266036
rect 676214 266024 676220 266036
rect 676272 266024 676278 266076
rect 377122 265956 377128 266008
rect 377180 265996 377186 266008
rect 556154 265996 556160 266008
rect 377180 265968 556160 265996
rect 377180 265956 377186 265968
rect 556154 265956 556160 265968
rect 556212 265956 556218 266008
rect 378502 265888 378508 265940
rect 378560 265928 378566 265940
rect 558914 265928 558920 265940
rect 378560 265900 558920 265928
rect 378560 265888 378566 265900
rect 558914 265888 558920 265900
rect 558972 265888 558978 265940
rect 380250 265820 380256 265872
rect 380308 265860 380314 265872
rect 564434 265860 564440 265872
rect 380308 265832 564440 265860
rect 380308 265820 380314 265832
rect 564434 265820 564440 265832
rect 564492 265820 564498 265872
rect 674650 265820 674656 265872
rect 674708 265860 674714 265872
rect 676030 265860 676036 265872
rect 674708 265832 676036 265860
rect 674708 265820 674714 265832
rect 676030 265820 676036 265832
rect 676088 265820 676094 265872
rect 381170 265752 381176 265804
rect 381228 265792 381234 265804
rect 565998 265792 566004 265804
rect 381228 265764 566004 265792
rect 381228 265752 381234 265764
rect 565998 265752 566004 265764
rect 566056 265752 566062 265804
rect 384298 265684 384304 265736
rect 384356 265724 384362 265736
rect 574278 265724 574284 265736
rect 384356 265696 574284 265724
rect 384356 265684 384362 265696
rect 574278 265684 574284 265696
rect 574336 265684 574342 265736
rect 28350 265616 28356 265668
rect 28408 265656 28414 265668
rect 46290 265656 46296 265668
rect 28408 265628 46296 265656
rect 28408 265616 28414 265628
rect 46290 265616 46296 265628
rect 46348 265616 46354 265668
rect 383838 265616 383844 265668
rect 383896 265656 383902 265668
rect 574094 265656 574100 265668
rect 383896 265628 574100 265656
rect 383896 265616 383902 265628
rect 574094 265616 574100 265628
rect 574152 265616 574158 265668
rect 194778 265548 194784 265600
rect 194836 265588 194842 265600
rect 195606 265588 195612 265600
rect 194836 265560 195612 265588
rect 194836 265548 194842 265560
rect 195606 265548 195612 265560
rect 195664 265548 195670 265600
rect 201586 265548 201592 265600
rect 201644 265588 201650 265600
rect 202230 265588 202236 265600
rect 201644 265560 202236 265588
rect 201644 265548 201650 265560
rect 202230 265548 202236 265560
rect 202288 265548 202294 265600
rect 209866 265548 209872 265600
rect 209924 265588 209930 265600
rect 210694 265588 210700 265600
rect 209924 265560 210700 265588
rect 209924 265548 209930 265560
rect 210694 265548 210700 265560
rect 210752 265548 210758 265600
rect 214006 265548 214012 265600
rect 214064 265588 214070 265600
rect 214742 265588 214748 265600
rect 214064 265560 214748 265588
rect 214064 265548 214070 265560
rect 214742 265548 214748 265560
rect 214800 265548 214806 265600
rect 222286 265548 222292 265600
rect 222344 265588 222350 265600
rect 223206 265588 223212 265600
rect 222344 265560 223212 265588
rect 222344 265548 222350 265560
rect 223206 265548 223212 265560
rect 223264 265548 223270 265600
rect 238846 265548 238852 265600
rect 238904 265588 238910 265600
rect 239674 265588 239680 265600
rect 238904 265560 239680 265588
rect 238904 265548 238910 265560
rect 239674 265548 239680 265560
rect 239732 265548 239738 265600
rect 240134 265548 240140 265600
rect 240192 265588 240198 265600
rect 240502 265588 240508 265600
rect 240192 265560 240508 265588
rect 240192 265548 240198 265560
rect 240502 265548 240508 265560
rect 240560 265548 240566 265600
rect 241606 265548 241612 265600
rect 241664 265588 241670 265600
rect 242342 265588 242348 265600
rect 241664 265560 242348 265588
rect 241664 265548 241670 265560
rect 242342 265548 242348 265560
rect 242400 265548 242406 265600
rect 242986 265548 242992 265600
rect 243044 265588 243050 265600
rect 243262 265588 243268 265600
rect 243044 265560 243268 265588
rect 243044 265548 243050 265560
rect 243262 265548 243268 265560
rect 243320 265548 243326 265600
rect 266354 265548 266360 265600
rect 266412 265588 266418 265600
rect 267274 265588 267280 265600
rect 266412 265560 267280 265588
rect 266412 265548 266418 265560
rect 267274 265548 267280 265560
rect 267332 265548 267338 265600
rect 351730 265548 351736 265600
rect 351788 265588 351794 265600
rect 488534 265588 488540 265600
rect 351788 265560 488540 265588
rect 351788 265548 351794 265560
rect 488534 265548 488540 265560
rect 488592 265548 488598 265600
rect 194594 265480 194600 265532
rect 194652 265520 194658 265532
rect 194962 265520 194968 265532
rect 194652 265492 194968 265520
rect 194652 265480 194658 265492
rect 194962 265480 194968 265492
rect 195020 265480 195026 265532
rect 240226 265480 240232 265532
rect 240284 265520 240290 265532
rect 241054 265520 241060 265532
rect 240284 265492 241060 265520
rect 240284 265480 240290 265492
rect 241054 265480 241060 265492
rect 241112 265480 241118 265532
rect 242894 265480 242900 265532
rect 242952 265520 242958 265532
rect 243630 265520 243636 265532
rect 242952 265492 243636 265520
rect 242952 265480 242958 265492
rect 243630 265480 243636 265492
rect 243688 265480 243694 265532
rect 349062 265480 349068 265532
rect 349120 265520 349126 265532
rect 481634 265520 481640 265532
rect 349120 265492 481640 265520
rect 349120 265480 349126 265492
rect 481634 265480 481640 265492
rect 481692 265480 481698 265532
rect 333054 265412 333060 265464
rect 333112 265452 333118 265464
rect 438854 265452 438860 265464
rect 333112 265424 438860 265452
rect 333112 265412 333118 265424
rect 438854 265412 438860 265424
rect 438912 265412 438918 265464
rect 330846 265344 330852 265396
rect 330904 265384 330910 265396
rect 433334 265384 433340 265396
rect 330904 265356 433340 265384
rect 330904 265344 330910 265356
rect 433334 265344 433340 265356
rect 433392 265344 433398 265396
rect 330386 265276 330392 265328
rect 330444 265316 330450 265328
rect 431954 265316 431960 265328
rect 330444 265288 431960 265316
rect 330444 265276 330450 265288
rect 431954 265276 431960 265288
rect 432012 265276 432018 265328
rect 327718 265208 327724 265260
rect 327776 265248 327782 265260
rect 425054 265248 425060 265260
rect 327776 265220 425060 265248
rect 327776 265208 327782 265220
rect 425054 265208 425060 265220
rect 425112 265208 425118 265260
rect 325050 265140 325056 265192
rect 325108 265180 325114 265192
rect 418154 265180 418160 265192
rect 325108 265152 418160 265180
rect 325108 265140 325114 265152
rect 418154 265140 418160 265152
rect 418212 265140 418218 265192
rect 245838 264936 245844 264988
rect 245896 264976 245902 264988
rect 246390 264976 246396 264988
rect 245896 264948 246396 264976
rect 245896 264936 245902 264948
rect 246390 264936 246396 264948
rect 246448 264936 246454 264988
rect 673362 264936 673368 264988
rect 673420 264976 673426 264988
rect 676214 264976 676220 264988
rect 673420 264948 676220 264976
rect 673420 264936 673426 264948
rect 676214 264936 676220 264948
rect 676272 264936 676278 264988
rect 337470 264528 337476 264580
rect 337528 264568 337534 264580
rect 451274 264568 451280 264580
rect 337528 264540 451280 264568
rect 337528 264528 337534 264540
rect 451274 264528 451280 264540
rect 451332 264528 451338 264580
rect 353846 264460 353852 264512
rect 353904 264500 353910 264512
rect 492674 264500 492680 264512
rect 353904 264472 492680 264500
rect 353904 264460 353910 264472
rect 492674 264460 492680 264472
rect 492732 264460 492738 264512
rect 384942 264392 384948 264444
rect 385000 264432 385006 264444
rect 575474 264432 575480 264444
rect 385000 264404 575480 264432
rect 385000 264392 385006 264404
rect 575474 264392 575480 264404
rect 575532 264392 575538 264444
rect 387610 264324 387616 264376
rect 387668 264364 387674 264376
rect 582558 264364 582564 264376
rect 387668 264336 582564 264364
rect 387668 264324 387674 264336
rect 582558 264324 582564 264336
rect 582616 264324 582622 264376
rect 393038 264256 393044 264308
rect 393096 264296 393102 264308
rect 597554 264296 597560 264308
rect 393096 264268 597560 264296
rect 393096 264256 393102 264268
rect 597554 264256 597560 264268
rect 597612 264256 597618 264308
rect 45002 264188 45008 264240
rect 45060 264228 45066 264240
rect 662506 264228 662512 264240
rect 45060 264200 662512 264228
rect 45060 264188 45066 264200
rect 662506 264188 662512 264200
rect 662564 264188 662570 264240
rect 399754 264120 399760 264172
rect 399812 264120 399818 264172
rect 401226 264120 401232 264172
rect 401284 264160 401290 264172
rect 607398 264160 607404 264172
rect 401284 264132 607404 264160
rect 401284 264120 401290 264132
rect 607398 264120 607404 264132
rect 607456 264120 607462 264172
rect 399772 264092 399800 264120
rect 615494 264092 615500 264104
rect 399772 264064 615500 264092
rect 615494 264052 615500 264064
rect 615552 264052 615558 264104
rect 673270 263576 673276 263628
rect 673328 263616 673334 263628
rect 676214 263616 676220 263628
rect 673328 263588 676220 263616
rect 673328 263576 673334 263588
rect 676214 263576 676220 263588
rect 676272 263576 676278 263628
rect 675018 262624 675024 262676
rect 675076 262664 675082 262676
rect 676030 262664 676036 262676
rect 675076 262636 676036 262664
rect 675076 262624 675082 262636
rect 676030 262624 676036 262636
rect 676088 262624 676094 262676
rect 415302 262216 415308 262268
rect 415360 262256 415366 262268
rect 572714 262256 572720 262268
rect 415360 262228 572720 262256
rect 415360 262216 415366 262228
rect 572714 262216 572720 262228
rect 572772 262216 572778 262268
rect 675202 262216 675208 262268
rect 675260 262256 675266 262268
rect 676030 262256 676036 262268
rect 675260 262228 676036 262256
rect 675260 262216 675266 262228
rect 676030 262216 676036 262228
rect 676088 262216 676094 262268
rect 674466 261944 674472 261996
rect 674524 261984 674530 261996
rect 676214 261984 676220 261996
rect 674524 261956 676220 261984
rect 674524 261944 674530 261956
rect 676214 261944 676220 261956
rect 676272 261944 676278 261996
rect 674742 261536 674748 261588
rect 674800 261576 674806 261588
rect 676214 261576 676220 261588
rect 674800 261548 676220 261576
rect 674800 261536 674806 261548
rect 676214 261536 676220 261548
rect 676272 261536 676278 261588
rect 672994 260856 673000 260908
rect 673052 260896 673058 260908
rect 676214 260896 676220 260908
rect 673052 260868 676220 260896
rect 673052 260856 673058 260868
rect 676214 260856 676220 260868
rect 676272 260856 676278 260908
rect 674558 259904 674564 259956
rect 674616 259944 674622 259956
rect 676214 259944 676220 259956
rect 674616 259916 676220 259944
rect 674616 259904 674622 259916
rect 676214 259904 676220 259916
rect 676272 259904 676278 259956
rect 675478 259360 675484 259412
rect 675536 259400 675542 259412
rect 676306 259400 676312 259412
rect 675536 259372 676312 259400
rect 675536 259360 675542 259372
rect 676306 259360 676312 259372
rect 676364 259360 676370 259412
rect 185210 258340 185216 258392
rect 185268 258380 185274 258392
rect 189074 258380 189080 258392
rect 185268 258352 189080 258380
rect 185268 258340 185274 258352
rect 189074 258340 189080 258352
rect 189132 258340 189138 258392
rect 673178 258136 673184 258188
rect 673236 258176 673242 258188
rect 676214 258176 676220 258188
rect 673236 258148 676220 258176
rect 673236 258136 673242 258148
rect 676214 258136 676220 258148
rect 676272 258136 676278 258188
rect 414198 258068 414204 258120
rect 414256 258108 414262 258120
rect 571518 258108 571524 258120
rect 414256 258080 571524 258108
rect 414256 258068 414262 258080
rect 571518 258068 571524 258080
rect 571576 258068 571582 258120
rect 673086 258068 673092 258120
rect 673144 258108 673150 258120
rect 676122 258108 676128 258120
rect 673144 258080 676128 258108
rect 673144 258068 673150 258080
rect 676122 258068 676128 258080
rect 676180 258068 676186 258120
rect 31570 258000 31576 258052
rect 31628 258040 31634 258052
rect 44358 258040 44364 258052
rect 31628 258012 44364 258040
rect 31628 258000 31634 258012
rect 44358 258000 44364 258012
rect 44416 258000 44422 258052
rect 31478 257864 31484 257916
rect 31536 257904 31542 257916
rect 44910 257904 44916 257916
rect 31536 257876 44916 257904
rect 31536 257864 31542 257876
rect 44910 257864 44916 257876
rect 44968 257864 44974 257916
rect 31662 257728 31668 257780
rect 31720 257768 31726 257780
rect 47670 257768 47676 257780
rect 31720 257740 47676 257768
rect 31720 257728 31726 257740
rect 47670 257728 47676 257740
rect 47728 257728 47734 257780
rect 671614 256708 671620 256760
rect 671672 256748 671678 256760
rect 683114 256748 683120 256760
rect 671672 256720 683120 256748
rect 671672 256708 671678 256720
rect 683114 256708 683120 256720
rect 683172 256708 683178 256760
rect 415302 255280 415308 255332
rect 415360 255320 415366 255332
rect 571426 255320 571432 255332
rect 415360 255292 571432 255320
rect 415360 255280 415366 255292
rect 571426 255280 571432 255292
rect 571484 255280 571490 255332
rect 414382 252560 414388 252612
rect 414440 252600 414446 252612
rect 574738 252600 574744 252612
rect 414440 252572 574744 252600
rect 414440 252560 414446 252572
rect 574738 252560 574744 252572
rect 574796 252560 574802 252612
rect 674650 251676 674656 251728
rect 674708 251716 674714 251728
rect 675018 251716 675024 251728
rect 674708 251688 675024 251716
rect 674708 251676 674714 251688
rect 675018 251676 675024 251688
rect 675076 251676 675082 251728
rect 675018 251540 675024 251592
rect 675076 251580 675082 251592
rect 675478 251580 675484 251592
rect 675076 251552 675484 251580
rect 675076 251540 675082 251552
rect 675478 251540 675484 251552
rect 675536 251540 675542 251592
rect 675386 251200 675392 251252
rect 675444 251200 675450 251252
rect 675404 250980 675432 251200
rect 675386 250928 675392 250980
rect 675444 250928 675450 250980
rect 674742 250180 674748 250232
rect 674800 250220 674806 250232
rect 675478 250220 675484 250232
rect 674800 250192 675484 250220
rect 674800 250180 674806 250192
rect 675478 250180 675484 250192
rect 675536 250180 675542 250232
rect 675018 249704 675024 249756
rect 675076 249744 675082 249756
rect 675386 249744 675392 249756
rect 675076 249716 675392 249744
rect 675076 249704 675082 249716
rect 675386 249704 675392 249716
rect 675444 249704 675450 249756
rect 674650 249568 674656 249620
rect 674708 249608 674714 249620
rect 675018 249608 675024 249620
rect 674708 249580 675024 249608
rect 674708 249568 674714 249580
rect 675018 249568 675024 249580
rect 675076 249568 675082 249620
rect 675202 248480 675208 248532
rect 675260 248480 675266 248532
rect 414198 248412 414204 248464
rect 414256 248452 414262 248464
rect 438210 248452 438216 248464
rect 414256 248424 438216 248452
rect 414256 248412 414262 248424
rect 438210 248412 438216 248424
rect 438268 248412 438274 248464
rect 675220 248328 675248 248480
rect 675202 248276 675208 248328
rect 675260 248276 675266 248328
rect 675018 247868 675024 247920
rect 675076 247908 675082 247920
rect 675478 247908 675484 247920
rect 675076 247880 675484 247908
rect 675076 247868 675082 247880
rect 675478 247868 675484 247880
rect 675536 247868 675542 247920
rect 672994 246984 673000 247036
rect 673052 247024 673058 247036
rect 675386 247024 675392 247036
rect 673052 246996 675392 247024
rect 673052 246984 673058 246996
rect 675386 246984 675392 246996
rect 675444 246984 675450 247036
rect 35802 245624 35808 245676
rect 35860 245664 35866 245676
rect 117958 245664 117964 245676
rect 35860 245636 117964 245664
rect 35860 245624 35866 245636
rect 117958 245624 117964 245636
rect 118016 245624 118022 245676
rect 415302 245624 415308 245676
rect 415360 245664 415366 245676
rect 438118 245664 438124 245676
rect 415360 245636 438124 245664
rect 415360 245624 415366 245636
rect 438118 245624 438124 245636
rect 438176 245624 438182 245676
rect 674742 243856 674748 243908
rect 674800 243896 674806 243908
rect 675110 243896 675116 243908
rect 674800 243868 675116 243896
rect 674800 243856 674806 243868
rect 675110 243856 675116 243868
rect 675168 243856 675174 243908
rect 675202 243856 675208 243908
rect 675260 243896 675266 243908
rect 675260 243868 675340 243896
rect 675260 243856 675266 243868
rect 675312 243636 675340 243868
rect 675294 243584 675300 243636
rect 675352 243584 675358 243636
rect 414382 242904 414388 242956
rect 414440 242944 414446 242956
rect 621658 242944 621664 242956
rect 414440 242916 621664 242944
rect 414440 242904 414446 242916
rect 621658 242904 621664 242916
rect 621716 242904 621722 242956
rect 32398 242292 32404 242344
rect 32456 242332 32462 242344
rect 41966 242332 41972 242344
rect 32456 242304 41972 242332
rect 32456 242292 32462 242304
rect 41966 242292 41972 242304
rect 42024 242292 42030 242344
rect 31110 242224 31116 242276
rect 31168 242264 31174 242276
rect 42426 242264 42432 242276
rect 31168 242236 42432 242264
rect 31168 242224 31174 242236
rect 42426 242224 42432 242236
rect 42484 242224 42490 242276
rect 31018 242156 31024 242208
rect 31076 242196 31082 242208
rect 42702 242196 42708 242208
rect 31076 242168 42708 242196
rect 31076 242156 31082 242168
rect 42702 242156 42708 242168
rect 42760 242156 42766 242208
rect 674558 242156 674564 242208
rect 674616 242196 674622 242208
rect 675386 242196 675392 242208
rect 674616 242168 675392 242196
rect 674616 242156 674622 242168
rect 675386 242156 675392 242168
rect 675444 242156 675450 242208
rect 673086 241612 673092 241664
rect 673144 241652 673150 241664
rect 675294 241652 675300 241664
rect 673144 241624 675300 241652
rect 673144 241612 673150 241624
rect 675294 241612 675300 241624
rect 675352 241612 675358 241664
rect 174998 241544 175004 241596
rect 175056 241544 175062 241596
rect 155862 240796 155868 240848
rect 155920 240836 155926 240848
rect 175016 240836 175044 241544
rect 673178 241068 673184 241120
rect 673236 241108 673242 241120
rect 675294 241108 675300 241120
rect 673236 241080 675300 241108
rect 673236 241068 673242 241080
rect 675294 241068 675300 241080
rect 675352 241068 675358 241120
rect 155920 240808 175044 240836
rect 155920 240796 155926 240808
rect 42426 240048 42432 240100
rect 42484 240088 42490 240100
rect 42794 240088 42800 240100
rect 42484 240060 42800 240088
rect 42484 240048 42490 240060
rect 42794 240048 42800 240060
rect 42852 240048 42858 240100
rect 42150 239980 42156 240032
rect 42208 240020 42214 240032
rect 44174 240020 44180 240032
rect 42208 239992 44180 240020
rect 42208 239980 42214 239992
rect 44174 239980 44180 239992
rect 44232 239980 44238 240032
rect 414934 238756 414940 238808
rect 414992 238796 414998 238808
rect 428458 238796 428464 238808
rect 414992 238768 428464 238796
rect 414992 238756 414998 238768
rect 428458 238756 428464 238768
rect 428516 238756 428522 238808
rect 674742 238756 674748 238808
rect 674800 238796 674806 238808
rect 674800 238768 675340 238796
rect 674800 238756 674806 238768
rect 675312 238728 675340 238768
rect 675386 238728 675392 238740
rect 675312 238700 675392 238728
rect 675386 238688 675392 238700
rect 675444 238688 675450 238740
rect 438210 238008 438216 238060
rect 438268 238048 438274 238060
rect 574094 238048 574100 238060
rect 438268 238020 574100 238048
rect 438268 238008 438274 238020
rect 574094 238008 574100 238020
rect 574152 238008 574158 238060
rect 184934 237396 184940 237448
rect 184992 237436 184998 237448
rect 189074 237436 189080 237448
rect 184992 237408 189080 237436
rect 184992 237396 184998 237408
rect 189074 237396 189080 237408
rect 189132 237396 189138 237448
rect 153102 235968 153108 236020
rect 153160 236008 153166 236020
rect 155862 236008 155868 236020
rect 153160 235980 155868 236008
rect 153160 235968 153166 235980
rect 155862 235968 155868 235980
rect 155920 235968 155926 236020
rect 42150 235356 42156 235408
rect 42208 235396 42214 235408
rect 44634 235396 44640 235408
rect 42208 235368 44640 235396
rect 42208 235356 42214 235368
rect 44634 235356 44640 235368
rect 44692 235356 44698 235408
rect 42150 234540 42156 234592
rect 42208 234580 42214 234592
rect 44542 234580 44548 234592
rect 42208 234552 44548 234580
rect 42208 234540 42214 234552
rect 44542 234540 44548 234552
rect 44600 234540 44606 234592
rect 42150 233996 42156 234048
rect 42208 234036 42214 234048
rect 44910 234036 44916 234048
rect 42208 234008 44916 234036
rect 42208 233996 42214 234008
rect 44910 233996 44916 234008
rect 44968 233996 44974 234048
rect 130378 233860 130384 233912
rect 130436 233900 130442 233912
rect 153102 233900 153108 233912
rect 130436 233872 153108 233900
rect 130436 233860 130442 233872
rect 153102 233860 153108 233872
rect 153160 233860 153166 233912
rect 438118 233860 438124 233912
rect 438176 233900 438182 233912
rect 572806 233900 572812 233912
rect 438176 233872 572812 233900
rect 438176 233860 438182 233872
rect 572806 233860 572812 233872
rect 572864 233860 572870 233912
rect 42150 233248 42156 233300
rect 42208 233288 42214 233300
rect 43162 233288 43168 233300
rect 42208 233260 43168 233288
rect 42208 233248 42214 233260
rect 43162 233248 43168 233260
rect 43220 233248 43226 233300
rect 415302 233248 415308 233300
rect 415360 233288 415366 233300
rect 427078 233288 427084 233300
rect 415360 233260 427084 233288
rect 415360 233248 415366 233260
rect 427078 233248 427084 233260
rect 427136 233248 427142 233300
rect 177114 232500 177120 232552
rect 177172 232540 177178 232552
rect 184842 232540 184848 232552
rect 177172 232512 184848 232540
rect 177172 232500 177178 232512
rect 184842 232500 184848 232512
rect 184900 232500 184906 232552
rect 414198 232500 414204 232552
rect 414256 232540 414262 232552
rect 639598 232540 639604 232552
rect 414256 232512 639604 232540
rect 414256 232500 414262 232512
rect 639598 232500 639604 232512
rect 639656 232500 639662 232552
rect 427078 232432 427084 232484
rect 427136 232472 427142 232484
rect 639138 232472 639144 232484
rect 427136 232444 639144 232472
rect 427136 232432 427142 232444
rect 639138 232432 639144 232444
rect 639196 232432 639202 232484
rect 428458 231752 428464 231804
rect 428516 231792 428522 231804
rect 639046 231792 639052 231804
rect 428516 231764 639052 231792
rect 428516 231752 428522 231764
rect 639046 231752 639052 231764
rect 639104 231752 639110 231804
rect 190362 231684 190368 231736
rect 190420 231724 190426 231736
rect 604454 231724 604460 231736
rect 190420 231696 604460 231724
rect 190420 231684 190426 231696
rect 604454 231684 604460 231696
rect 604512 231684 604518 231736
rect 191098 231616 191104 231668
rect 191156 231656 191162 231668
rect 663794 231656 663800 231668
rect 191156 231628 663800 231656
rect 191156 231616 191162 231628
rect 663794 231616 663800 231628
rect 663852 231616 663858 231668
rect 65150 231548 65156 231600
rect 65208 231588 65214 231600
rect 177114 231588 177120 231600
rect 65208 231560 177120 231588
rect 65208 231548 65214 231560
rect 177114 231548 177120 231560
rect 177172 231548 177178 231600
rect 189718 231548 189724 231600
rect 189776 231588 189782 231600
rect 663886 231588 663892 231600
rect 189776 231560 663892 231588
rect 189776 231548 189782 231560
rect 663886 231548 663892 231560
rect 663944 231548 663950 231600
rect 55858 231480 55864 231532
rect 55916 231520 55922 231532
rect 649350 231520 649356 231532
rect 55916 231492 649356 231520
rect 55916 231480 55922 231492
rect 649350 231480 649356 231492
rect 649408 231480 649414 231532
rect 64138 231412 64144 231464
rect 64196 231452 64202 231464
rect 661034 231452 661040 231464
rect 64196 231424 661040 231452
rect 64196 231412 64202 231424
rect 661034 231412 661040 231424
rect 661092 231412 661098 231464
rect 54478 231344 54484 231396
rect 54536 231384 54542 231396
rect 654134 231384 654140 231396
rect 54536 231356 654140 231384
rect 54536 231344 54542 231356
rect 654134 231344 654140 231356
rect 654192 231344 654198 231396
rect 50338 231276 50344 231328
rect 50396 231316 50402 231328
rect 650638 231316 650644 231328
rect 50396 231288 650644 231316
rect 50396 231276 50402 231288
rect 650638 231276 650644 231288
rect 650696 231276 650702 231328
rect 51718 231208 51724 231260
rect 51776 231248 51782 231260
rect 652754 231248 652760 231260
rect 51776 231220 652760 231248
rect 51776 231208 51782 231220
rect 652754 231208 652760 231220
rect 652812 231208 652818 231260
rect 53098 231140 53104 231192
rect 53156 231180 53162 231192
rect 655514 231180 655520 231192
rect 53156 231152 655520 231180
rect 53156 231140 53162 231152
rect 655514 231140 655520 231152
rect 655572 231140 655578 231192
rect 42150 231072 42156 231124
rect 42208 231112 42214 231124
rect 43254 231112 43260 231124
rect 42208 231084 43260 231112
rect 42208 231072 42214 231084
rect 43254 231072 43260 231084
rect 43312 231072 43318 231124
rect 43898 231072 43904 231124
rect 43956 231112 43962 231124
rect 662598 231112 662604 231124
rect 43956 231084 662604 231112
rect 43956 231072 43962 231084
rect 662598 231072 662604 231084
rect 662656 231072 662662 231124
rect 42150 230528 42156 230580
rect 42208 230568 42214 230580
rect 42426 230568 42432 230580
rect 42208 230540 42432 230568
rect 42208 230528 42214 230540
rect 42426 230528 42432 230540
rect 42484 230528 42490 230580
rect 271248 230472 271552 230500
rect 179322 230392 179328 230444
rect 179380 230432 179386 230444
rect 246114 230432 246120 230444
rect 179380 230404 246120 230432
rect 179380 230392 179386 230404
rect 246114 230392 246120 230404
rect 246172 230392 246178 230444
rect 262214 230392 262220 230444
rect 262272 230432 262278 230444
rect 263226 230432 263232 230444
rect 262272 230404 263232 230432
rect 262272 230392 262278 230404
rect 263226 230392 263232 230404
rect 263284 230392 263290 230444
rect 263594 230392 263600 230444
rect 263652 230432 263658 230444
rect 263778 230432 263784 230444
rect 263652 230404 263784 230432
rect 263652 230392 263658 230404
rect 263778 230392 263784 230404
rect 263836 230392 263842 230444
rect 175182 230324 175188 230376
rect 175240 230364 175246 230376
rect 244642 230364 244648 230376
rect 175240 230336 244648 230364
rect 175240 230324 175246 230336
rect 244642 230324 244648 230336
rect 244700 230324 244706 230376
rect 246942 230324 246948 230376
rect 247000 230364 247006 230376
rect 271248 230364 271276 230472
rect 271524 230432 271552 230472
rect 333606 230460 333612 230512
rect 333664 230500 333670 230512
rect 333664 230472 334020 230500
rect 333664 230460 333670 230472
rect 274634 230432 274640 230444
rect 271524 230404 274640 230432
rect 274634 230392 274640 230404
rect 274692 230392 274698 230444
rect 276750 230392 276756 230444
rect 276808 230432 276814 230444
rect 277762 230432 277768 230444
rect 276808 230404 277768 230432
rect 276808 230392 276814 230404
rect 277762 230392 277768 230404
rect 277820 230392 277826 230444
rect 285306 230432 285312 230444
rect 277964 230404 285312 230432
rect 247000 230336 271276 230364
rect 247000 230324 247006 230336
rect 271322 230324 271328 230376
rect 271380 230364 271386 230376
rect 272794 230364 272800 230376
rect 271380 230336 272800 230364
rect 271380 230324 271386 230336
rect 272794 230324 272800 230336
rect 272852 230324 272858 230376
rect 169662 230256 169668 230308
rect 169720 230296 169726 230308
rect 241790 230296 241796 230308
rect 169720 230268 241796 230296
rect 169720 230256 169726 230268
rect 241790 230256 241796 230268
rect 241848 230256 241854 230308
rect 244182 230256 244188 230308
rect 244240 230296 244246 230308
rect 274266 230296 274272 230308
rect 244240 230268 274272 230296
rect 244240 230256 244246 230268
rect 274266 230256 274272 230268
rect 274324 230256 274330 230308
rect 274542 230256 274548 230308
rect 274600 230296 274606 230308
rect 277964 230296 277992 230404
rect 285306 230392 285312 230404
rect 285364 230392 285370 230444
rect 288342 230392 288348 230444
rect 288400 230432 288406 230444
rect 292758 230432 292764 230444
rect 288400 230404 292764 230432
rect 288400 230392 288406 230404
rect 292758 230392 292764 230404
rect 292816 230392 292822 230444
rect 299934 230392 299940 230444
rect 299992 230432 299998 230444
rect 303982 230432 303988 230444
rect 299992 230404 303988 230432
rect 299992 230392 299998 230404
rect 303982 230392 303988 230404
rect 304040 230392 304046 230444
rect 314930 230392 314936 230444
rect 314988 230432 314994 230444
rect 315942 230432 315948 230444
rect 314988 230404 315948 230432
rect 314988 230392 314994 230404
rect 315942 230392 315948 230404
rect 316000 230392 316006 230444
rect 318794 230392 318800 230444
rect 318852 230432 318858 230444
rect 326338 230432 326344 230444
rect 318852 230404 326344 230432
rect 318852 230392 318858 230404
rect 326338 230392 326344 230404
rect 326396 230392 326402 230444
rect 331306 230392 331312 230444
rect 331364 230432 331370 230444
rect 332226 230432 332232 230444
rect 331364 230404 332232 230432
rect 331364 230392 331370 230404
rect 332226 230392 332232 230404
rect 332284 230392 332290 230444
rect 333054 230392 333060 230444
rect 333112 230432 333118 230444
rect 333882 230432 333888 230444
rect 333112 230404 333888 230432
rect 333112 230392 333118 230404
rect 333882 230392 333888 230404
rect 333940 230392 333946 230444
rect 333992 230432 334020 230472
rect 385126 230460 385132 230512
rect 385184 230500 385190 230512
rect 507946 230500 507952 230512
rect 385184 230472 507952 230500
rect 385184 230460 385190 230472
rect 507946 230460 507952 230472
rect 508004 230460 508010 230512
rect 604454 230460 604460 230512
rect 604512 230500 604518 230512
rect 605742 230500 605748 230512
rect 604512 230472 605748 230500
rect 604512 230460 604518 230472
rect 605742 230460 605748 230472
rect 605800 230500 605806 230512
rect 636838 230500 636844 230512
rect 605800 230472 636844 230500
rect 605800 230460 605806 230472
rect 636838 230460 636844 230472
rect 636896 230460 636902 230512
rect 371878 230432 371884 230444
rect 333992 230404 371884 230432
rect 371878 230392 371884 230404
rect 371936 230392 371942 230444
rect 380710 230432 380716 230444
rect 373966 230404 380716 230432
rect 279418 230324 279424 230376
rect 279476 230364 279482 230376
rect 283190 230364 283196 230376
rect 279476 230336 283196 230364
rect 279476 230324 279482 230336
rect 283190 230324 283196 230336
rect 283248 230324 283254 230376
rect 287422 230364 287428 230376
rect 283300 230336 287428 230364
rect 274600 230268 277992 230296
rect 274600 230256 274606 230268
rect 278038 230256 278044 230308
rect 278096 230296 278102 230308
rect 283300 230296 283328 230336
rect 287422 230324 287428 230336
rect 287480 230324 287486 230376
rect 305638 230324 305644 230376
rect 305696 230364 305702 230376
rect 306190 230364 306196 230376
rect 305696 230336 306196 230364
rect 305696 230324 305702 230336
rect 306190 230324 306196 230336
rect 306248 230324 306254 230376
rect 307018 230324 307024 230376
rect 307076 230364 307082 230376
rect 307570 230364 307576 230376
rect 307076 230336 307576 230364
rect 307076 230324 307082 230336
rect 307570 230324 307576 230336
rect 307628 230324 307634 230376
rect 312078 230324 312084 230376
rect 312136 230364 312142 230376
rect 313182 230364 313188 230376
rect 312136 230336 313188 230364
rect 312136 230324 312142 230336
rect 313182 230324 313188 230336
rect 313240 230324 313246 230376
rect 314562 230324 314568 230376
rect 314620 230364 314626 230376
rect 314620 230336 316034 230364
rect 314620 230324 314626 230336
rect 278096 230268 283328 230296
rect 278096 230256 278102 230268
rect 286962 230256 286968 230308
rect 287020 230296 287026 230308
rect 291746 230296 291752 230308
rect 287020 230268 291752 230296
rect 287020 230256 287026 230268
rect 291746 230256 291752 230268
rect 291804 230256 291810 230308
rect 316006 230296 316034 230336
rect 316310 230324 316316 230376
rect 316368 230364 316374 230376
rect 317322 230364 317328 230376
rect 316368 230336 317328 230364
rect 316368 230324 316374 230336
rect 317322 230324 317328 230336
rect 317380 230324 317386 230376
rect 317782 230324 317788 230376
rect 317840 230364 317846 230376
rect 318702 230364 318708 230376
rect 317840 230336 318708 230364
rect 317840 230324 317846 230336
rect 318702 230324 318708 230336
rect 318760 230324 318766 230376
rect 319254 230324 319260 230376
rect 319312 230364 319318 230376
rect 319898 230364 319904 230376
rect 319312 230336 319904 230364
rect 319312 230324 319318 230336
rect 319898 230324 319904 230336
rect 319956 230324 319962 230376
rect 320634 230324 320640 230376
rect 320692 230364 320698 230376
rect 321370 230364 321376 230376
rect 320692 230336 321376 230364
rect 320692 230324 320698 230336
rect 321370 230324 321376 230336
rect 321428 230324 321434 230376
rect 321646 230324 321652 230376
rect 321704 230364 321710 230376
rect 338758 230364 338764 230376
rect 321704 230336 338764 230364
rect 321704 230324 321710 230336
rect 338758 230324 338764 230336
rect 338816 230324 338822 230376
rect 341978 230324 341984 230376
rect 342036 230364 342042 230376
rect 373966 230364 373994 230404
rect 380710 230392 380716 230404
rect 380768 230392 380774 230444
rect 393682 230392 393688 230444
rect 393740 230432 393746 230444
rect 400674 230432 400680 230444
rect 393740 230404 400680 230432
rect 393740 230392 393746 230404
rect 400674 230392 400680 230404
rect 400732 230392 400738 230444
rect 401870 230392 401876 230444
rect 401928 230432 401934 230444
rect 456150 230432 456156 230444
rect 401928 230404 456156 230432
rect 401928 230392 401934 230404
rect 456150 230392 456156 230404
rect 456208 230392 456214 230444
rect 342036 230336 373994 230364
rect 342036 230324 342042 230336
rect 374086 230324 374092 230376
rect 374144 230364 374150 230376
rect 377398 230364 377404 230376
rect 374144 230336 377404 230364
rect 374144 230324 374150 230336
rect 377398 230324 377404 230336
rect 377456 230324 377462 230376
rect 390830 230324 390836 230376
rect 390888 230364 390894 230376
rect 391842 230364 391848 230376
rect 390888 230336 391848 230364
rect 390888 230324 390894 230336
rect 391842 230324 391848 230336
rect 391900 230324 391906 230376
rect 393314 230324 393320 230376
rect 393372 230364 393378 230376
rect 394602 230364 394608 230376
rect 393372 230336 394608 230364
rect 393372 230324 393378 230336
rect 394602 230324 394608 230336
rect 394660 230324 394666 230376
rect 397638 230324 397644 230376
rect 397696 230364 397702 230376
rect 398558 230364 398564 230376
rect 397696 230336 398564 230364
rect 397696 230324 397702 230336
rect 398558 230324 398564 230336
rect 398616 230324 398622 230376
rect 399018 230324 399024 230376
rect 399076 230364 399082 230376
rect 400122 230364 400128 230376
rect 399076 230336 400128 230364
rect 399076 230324 399082 230336
rect 400122 230324 400128 230336
rect 400180 230324 400186 230376
rect 403342 230324 403348 230376
rect 403400 230364 403406 230376
rect 404170 230364 404176 230376
rect 403400 230336 404176 230364
rect 403400 230324 403406 230336
rect 404170 230324 404176 230336
rect 404228 230324 404234 230376
rect 404354 230324 404360 230376
rect 404412 230364 404418 230376
rect 406654 230364 406660 230376
rect 404412 230336 406660 230364
rect 404412 230324 404418 230336
rect 406654 230324 406660 230336
rect 406712 230324 406718 230376
rect 406838 230324 406844 230376
rect 406896 230364 406902 230376
rect 410978 230364 410984 230376
rect 406896 230336 410984 230364
rect 406896 230324 406902 230336
rect 410978 230324 410984 230336
rect 411036 230324 411042 230376
rect 411162 230324 411168 230376
rect 411220 230364 411226 230376
rect 461578 230364 461584 230376
rect 411220 230336 461584 230364
rect 411220 230324 411226 230336
rect 461578 230324 461584 230336
rect 461636 230324 461642 230376
rect 319346 230296 319352 230308
rect 316006 230268 319352 230296
rect 319346 230256 319352 230268
rect 319404 230256 319410 230308
rect 339126 230256 339132 230308
rect 339184 230296 339190 230308
rect 378226 230296 378232 230308
rect 339184 230268 378232 230296
rect 339184 230256 339190 230268
rect 378226 230256 378232 230268
rect 378284 230256 378290 230308
rect 395430 230256 395436 230308
rect 395488 230296 395494 230308
rect 396718 230296 396724 230308
rect 395488 230268 396724 230296
rect 395488 230256 395494 230268
rect 396718 230256 396724 230268
rect 396776 230256 396782 230308
rect 398650 230256 398656 230308
rect 398708 230296 398714 230308
rect 400858 230296 400864 230308
rect 398708 230268 400864 230296
rect 398708 230256 398714 230268
rect 400858 230256 400864 230268
rect 400916 230256 400922 230308
rect 402974 230256 402980 230308
rect 403032 230296 403038 230308
rect 404262 230296 404268 230308
rect 403032 230268 404268 230296
rect 403032 230256 403038 230268
rect 404262 230256 404268 230268
rect 404320 230256 404326 230308
rect 404722 230256 404728 230308
rect 404780 230296 404786 230308
rect 409782 230296 409788 230308
rect 404780 230268 409788 230296
rect 404780 230256 404786 230268
rect 409782 230256 409788 230268
rect 409840 230256 409846 230308
rect 467098 230296 467104 230308
rect 409892 230268 467104 230296
rect 136358 230188 136364 230240
rect 136416 230228 136422 230240
rect 213270 230228 213276 230240
rect 136416 230200 213276 230228
rect 136416 230188 136422 230200
rect 213270 230188 213276 230200
rect 213328 230188 213334 230240
rect 219250 230188 219256 230240
rect 219308 230228 219314 230240
rect 262214 230228 262220 230240
rect 219308 230200 262220 230228
rect 219308 230188 219314 230200
rect 262214 230188 262220 230200
rect 262272 230188 262278 230240
rect 262766 230188 262772 230240
rect 262824 230228 262830 230240
rect 269942 230228 269948 230240
rect 262824 230200 269948 230228
rect 262824 230188 262830 230200
rect 269942 230188 269948 230200
rect 270000 230188 270006 230240
rect 276658 230188 276664 230240
rect 276716 230228 276722 230240
rect 287054 230228 287060 230240
rect 276716 230200 287060 230228
rect 276716 230188 276722 230200
rect 287054 230188 287060 230200
rect 287112 230188 287118 230240
rect 311710 230188 311716 230240
rect 311768 230228 311774 230240
rect 315298 230228 315304 230240
rect 311768 230200 315304 230228
rect 311768 230188 311774 230200
rect 315298 230188 315304 230200
rect 315356 230188 315362 230240
rect 320266 230188 320272 230240
rect 320324 230228 320330 230240
rect 337378 230228 337384 230240
rect 320324 230200 337384 230228
rect 320324 230188 320330 230200
rect 337378 230188 337384 230200
rect 337436 230188 337442 230240
rect 347682 230188 347688 230240
rect 347740 230228 347746 230240
rect 386414 230228 386420 230240
rect 347740 230200 386420 230228
rect 347740 230188 347746 230200
rect 386414 230188 386420 230200
rect 386472 230188 386478 230240
rect 398098 230188 398104 230240
rect 398156 230228 398162 230240
rect 403066 230228 403072 230240
rect 398156 230200 403072 230228
rect 398156 230188 398162 230200
rect 403066 230188 403072 230200
rect 403124 230188 403130 230240
rect 406194 230188 406200 230240
rect 406252 230228 406258 230240
rect 409892 230228 409920 230268
rect 467098 230256 467104 230268
rect 467156 230256 467162 230308
rect 406252 230200 409920 230228
rect 406252 230188 406258 230200
rect 409966 230188 409972 230240
rect 410024 230228 410030 230240
rect 469214 230228 469220 230240
rect 410024 230200 469220 230228
rect 410024 230188 410030 230200
rect 469214 230188 469220 230200
rect 469272 230188 469278 230240
rect 155862 230120 155868 230172
rect 155920 230160 155926 230172
rect 236086 230160 236092 230172
rect 155920 230132 236092 230160
rect 155920 230120 155926 230132
rect 236086 230120 236092 230132
rect 236144 230120 236150 230172
rect 240042 230120 240048 230172
rect 240100 230160 240106 230172
rect 271782 230160 271788 230172
rect 240100 230132 271788 230160
rect 240100 230120 240106 230132
rect 271782 230120 271788 230132
rect 271840 230120 271846 230172
rect 275278 230120 275284 230172
rect 275336 230160 275342 230172
rect 277670 230160 277676 230172
rect 275336 230132 277676 230160
rect 275336 230120 275342 230132
rect 277670 230120 277676 230132
rect 277728 230120 277734 230172
rect 277762 230120 277768 230172
rect 277820 230160 277826 230172
rect 286042 230160 286048 230172
rect 277820 230132 286048 230160
rect 277820 230120 277826 230132
rect 286042 230120 286048 230132
rect 286100 230120 286106 230172
rect 317414 230120 317420 230172
rect 317472 230160 317478 230172
rect 334618 230160 334624 230172
rect 317472 230132 334624 230160
rect 317472 230120 317478 230132
rect 334618 230120 334624 230132
rect 334676 230120 334682 230172
rect 336642 230120 336648 230172
rect 336700 230160 336706 230172
rect 376018 230160 376024 230172
rect 336700 230132 376024 230160
rect 336700 230120 336706 230132
rect 376018 230120 376024 230132
rect 376076 230120 376082 230172
rect 378318 230120 378324 230172
rect 378376 230160 378382 230172
rect 443638 230160 443644 230172
rect 378376 230132 443644 230160
rect 378376 230120 378382 230132
rect 443638 230120 443644 230132
rect 443696 230120 443702 230172
rect 146202 230052 146208 230104
rect 146260 230092 146266 230104
rect 231854 230092 231860 230104
rect 146260 230064 231860 230092
rect 146260 230052 146266 230064
rect 231854 230052 231860 230064
rect 231912 230052 231918 230104
rect 233142 230052 233148 230104
rect 233200 230092 233206 230104
rect 233200 230064 267734 230092
rect 233200 230052 233206 230064
rect 139302 229984 139308 230036
rect 139360 230024 139366 230036
rect 229002 230024 229008 230036
rect 139360 229996 229008 230024
rect 139360 229984 139366 229996
rect 229002 229984 229008 229996
rect 229060 229984 229066 230036
rect 234522 229984 234528 230036
rect 234580 230024 234586 230036
rect 262766 230024 262772 230036
rect 234580 229996 262772 230024
rect 234580 229984 234586 229996
rect 262766 229984 262772 229996
rect 262824 229984 262830 230036
rect 267706 230024 267734 230064
rect 271138 230052 271144 230104
rect 271196 230092 271202 230104
rect 277118 230092 277124 230104
rect 271196 230064 277124 230092
rect 271196 230052 271202 230064
rect 277118 230052 277124 230064
rect 277176 230052 277182 230104
rect 277210 230052 277216 230104
rect 277268 230092 277274 230104
rect 282454 230092 282460 230104
rect 277268 230064 282460 230092
rect 277268 230052 277274 230064
rect 282454 230052 282460 230064
rect 282512 230052 282518 230104
rect 315850 230052 315856 230104
rect 315908 230092 315914 230104
rect 322198 230092 322204 230104
rect 315908 230064 322204 230092
rect 315908 230052 315914 230064
rect 322198 230052 322204 230064
rect 322256 230052 322262 230104
rect 323762 230052 323768 230104
rect 323820 230092 323826 230104
rect 364518 230092 364524 230104
rect 323820 230064 364524 230092
rect 323820 230052 323826 230064
rect 364518 230052 364524 230064
rect 364576 230052 364582 230104
rect 387978 230052 387984 230104
rect 388036 230092 388042 230104
rect 515398 230092 515404 230104
rect 388036 230064 515404 230092
rect 388036 230052 388042 230064
rect 515398 230052 515404 230064
rect 515456 230052 515462 230104
rect 268930 230024 268936 230036
rect 267706 229996 268936 230024
rect 268930 229984 268936 229996
rect 268988 229984 268994 230036
rect 270402 229984 270408 230036
rect 270460 230024 270466 230036
rect 283834 230024 283840 230036
rect 270460 229996 283840 230024
rect 270460 229984 270466 229996
rect 283834 229984 283840 229996
rect 283892 229984 283898 230036
rect 285490 229984 285496 230036
rect 285548 230024 285554 230036
rect 290642 230024 290648 230036
rect 285548 229996 290648 230024
rect 285548 229984 285554 229996
rect 290642 229984 290648 229996
rect 290700 229984 290706 230036
rect 312354 229984 312360 230036
rect 312412 230024 312418 230036
rect 337010 230024 337016 230036
rect 312412 229996 337016 230024
rect 312412 229984 312418 229996
rect 337010 229984 337016 229996
rect 337068 229984 337074 230036
rect 343726 229984 343732 230036
rect 343784 230024 343790 230036
rect 385678 230024 385684 230036
rect 343784 229996 385684 230024
rect 343784 229984 343790 229996
rect 385678 229984 385684 229996
rect 385736 229984 385742 230036
rect 387610 229984 387616 230036
rect 387668 230024 387674 230036
rect 399478 230024 399484 230036
rect 387668 229996 399484 230024
rect 387668 229984 387674 229996
rect 399478 229984 399484 229996
rect 399536 229984 399542 230036
rect 400858 229984 400864 230036
rect 400916 230024 400922 230036
rect 407758 230024 407764 230036
rect 400916 229996 407764 230024
rect 400916 229984 400922 229996
rect 407758 229984 407764 229996
rect 407816 229984 407822 230036
rect 408310 229984 408316 230036
rect 408368 230024 408374 230036
rect 408368 229996 411944 230024
rect 408368 229984 408374 229996
rect 132402 229916 132408 229968
rect 132460 229956 132466 229968
rect 226150 229956 226156 229968
rect 132460 229928 226156 229956
rect 132460 229916 132466 229928
rect 226150 229916 226156 229928
rect 226208 229916 226214 229968
rect 226242 229916 226248 229968
rect 226300 229956 226306 229968
rect 259914 229956 259920 229968
rect 226300 229928 259920 229956
rect 226300 229916 226306 229928
rect 259914 229916 259920 229928
rect 259972 229916 259978 229968
rect 260098 229916 260104 229968
rect 260156 229956 260162 229968
rect 262858 229956 262864 229968
rect 260156 229928 262864 229956
rect 260156 229916 260162 229928
rect 262858 229916 262864 229928
rect 262916 229916 262922 229968
rect 270310 229916 270316 229968
rect 270368 229956 270374 229968
rect 284570 229956 284576 229968
rect 270368 229928 284576 229956
rect 270368 229916 270374 229928
rect 284570 229916 284576 229928
rect 284628 229916 284634 229968
rect 285582 229916 285588 229968
rect 285640 229956 285646 229968
rect 291378 229956 291384 229968
rect 285640 229928 291384 229956
rect 285640 229916 285646 229928
rect 291378 229916 291384 229928
rect 291436 229916 291442 229968
rect 313826 229916 313832 229968
rect 313884 229956 313890 229968
rect 341242 229956 341248 229968
rect 313884 229928 341248 229956
rect 313884 229916 313890 229928
rect 341242 229916 341248 229928
rect 341300 229916 341306 229968
rect 345566 229916 345572 229968
rect 345624 229956 345630 229968
rect 354766 229956 354772 229968
rect 345624 229928 354772 229956
rect 345624 229916 345630 229928
rect 354766 229916 354772 229928
rect 354824 229916 354830 229968
rect 356238 229916 356244 229968
rect 356296 229956 356302 229968
rect 357066 229956 357072 229968
rect 356296 229928 357072 229956
rect 356296 229916 356302 229928
rect 357066 229916 357072 229928
rect 357124 229916 357130 229968
rect 359090 229916 359096 229968
rect 359148 229956 359154 229968
rect 360102 229956 360108 229968
rect 359148 229928 360108 229956
rect 359148 229916 359154 229928
rect 360102 229916 360108 229928
rect 360160 229916 360166 229968
rect 360562 229916 360568 229968
rect 360620 229956 360626 229968
rect 361298 229956 361304 229968
rect 360620 229928 361304 229956
rect 360620 229916 360626 229928
rect 361298 229916 361304 229928
rect 361356 229916 361362 229968
rect 361942 229916 361948 229968
rect 362000 229956 362006 229968
rect 362678 229956 362684 229968
rect 362000 229928 362684 229956
rect 362000 229916 362006 229928
rect 362678 229916 362684 229928
rect 362736 229916 362742 229968
rect 364242 229916 364248 229968
rect 364300 229956 364306 229968
rect 407022 229956 407028 229968
rect 364300 229928 407028 229956
rect 364300 229916 364306 229928
rect 407022 229916 407028 229928
rect 407080 229916 407086 229968
rect 409322 229916 409328 229968
rect 409380 229956 409386 229968
rect 411916 229956 411944 229996
rect 411990 229984 411996 230036
rect 412048 230024 412054 230036
rect 539594 230024 539600 230036
rect 412048 229996 539600 230024
rect 412048 229984 412054 229996
rect 539594 229984 539600 229996
rect 539652 229984 539658 230036
rect 547138 229956 547144 229968
rect 409380 229928 411668 229956
rect 411916 229928 547144 229956
rect 409380 229916 409386 229928
rect 42150 229848 42156 229900
rect 42208 229888 42214 229900
rect 43070 229888 43076 229900
rect 42208 229860 43076 229888
rect 42208 229848 42214 229860
rect 43070 229848 43076 229860
rect 43128 229848 43134 229900
rect 91738 229848 91744 229900
rect 91796 229888 91802 229900
rect 206186 229888 206192 229900
rect 91796 229860 206192 229888
rect 91796 229848 91802 229860
rect 206186 229848 206192 229860
rect 206244 229848 206250 229900
rect 212442 229848 212448 229900
rect 212500 229888 212506 229900
rect 260374 229888 260380 229900
rect 212500 229860 260380 229888
rect 212500 229848 212506 229860
rect 260374 229848 260380 229860
rect 260432 229848 260438 229900
rect 263502 229848 263508 229900
rect 263560 229888 263566 229900
rect 281718 229888 281724 229900
rect 263560 229860 281724 229888
rect 263560 229848 263566 229860
rect 281718 229848 281724 229860
rect 281776 229848 281782 229900
rect 284110 229848 284116 229900
rect 284168 229888 284174 229900
rect 290274 229888 290280 229900
rect 284168 229860 290280 229888
rect 284168 229848 284174 229860
rect 290274 229848 290280 229860
rect 290332 229848 290338 229900
rect 304902 229848 304908 229900
rect 304960 229888 304966 229900
rect 311618 229888 311624 229900
rect 304960 229860 311624 229888
rect 304960 229848 304966 229860
rect 311618 229848 311624 229860
rect 311676 229848 311682 229900
rect 316678 229848 316684 229900
rect 316736 229888 316742 229900
rect 346486 229888 346492 229900
rect 316736 229860 346492 229888
rect 316736 229848 316742 229860
rect 346486 229848 346492 229860
rect 346544 229848 346550 229900
rect 352006 229848 352012 229900
rect 352064 229888 352070 229900
rect 398098 229888 398104 229900
rect 352064 229860 398104 229888
rect 352064 229848 352070 229860
rect 398098 229848 398104 229860
rect 398156 229848 398162 229900
rect 399754 229848 399760 229900
rect 399812 229888 399818 229900
rect 407850 229888 407856 229900
rect 399812 229860 407856 229888
rect 399812 229848 399818 229860
rect 407850 229848 407856 229860
rect 407908 229848 407914 229900
rect 410426 229848 410432 229900
rect 410484 229888 410490 229900
rect 411640 229888 411668 229928
rect 547138 229916 547144 229928
rect 547196 229916 547202 229968
rect 551278 229888 551284 229900
rect 410484 229860 411576 229888
rect 411640 229860 551284 229888
rect 410484 229848 410490 229860
rect 82814 229780 82820 229832
rect 82872 229820 82878 229832
rect 203334 229820 203340 229832
rect 82872 229792 203340 229820
rect 82872 229780 82878 229792
rect 203334 229780 203340 229792
rect 203392 229780 203398 229832
rect 203518 229780 203524 229832
rect 203576 229820 203582 229832
rect 204714 229820 204720 229832
rect 203576 229792 204720 229820
rect 203576 229780 203582 229792
rect 204714 229780 204720 229792
rect 204772 229780 204778 229832
rect 206738 229780 206744 229832
rect 206796 229820 206802 229832
rect 257522 229820 257528 229832
rect 206796 229792 257528 229820
rect 206796 229780 206802 229792
rect 257522 229780 257528 229792
rect 257580 229780 257586 229832
rect 259362 229780 259368 229832
rect 259420 229820 259426 229832
rect 280338 229820 280344 229832
rect 259420 229792 280344 229820
rect 259420 229780 259426 229792
rect 280338 229780 280344 229792
rect 280396 229780 280402 229832
rect 281350 229780 281356 229832
rect 281408 229820 281414 229832
rect 289906 229820 289912 229832
rect 281408 229792 289912 229820
rect 281408 229780 281414 229792
rect 289906 229780 289912 229792
rect 289964 229780 289970 229832
rect 298830 229780 298836 229832
rect 298888 229820 298894 229832
rect 302510 229820 302516 229832
rect 298888 229792 302516 229820
rect 298888 229780 298894 229792
rect 302510 229780 302516 229792
rect 302568 229780 302574 229832
rect 303522 229780 303528 229832
rect 303580 229820 303586 229832
rect 312538 229820 312544 229832
rect 303580 229792 312544 229820
rect 303580 229780 303586 229792
rect 312538 229780 312544 229792
rect 312596 229780 312602 229832
rect 318058 229780 318064 229832
rect 318116 229820 318122 229832
rect 350902 229820 350908 229832
rect 318116 229792 350908 229820
rect 318116 229780 318122 229792
rect 350902 229780 350908 229792
rect 350960 229780 350966 229832
rect 362310 229780 362316 229832
rect 362368 229820 362374 229832
rect 364150 229820 364156 229832
rect 362368 229792 364156 229820
rect 362368 229780 362374 229792
rect 364150 229780 364156 229792
rect 364208 229780 364214 229832
rect 364242 229780 364248 229832
rect 364300 229820 364306 229832
rect 407390 229820 407396 229832
rect 364300 229792 407396 229820
rect 364300 229780 364306 229792
rect 407390 229780 407396 229792
rect 407448 229780 407454 229832
rect 407684 229792 409000 229820
rect 73798 229712 73804 229764
rect 73856 229752 73862 229764
rect 200482 229752 200488 229764
rect 73856 229724 200488 229752
rect 73856 229712 73862 229724
rect 200482 229712 200488 229724
rect 200540 229712 200546 229764
rect 200666 229712 200672 229764
rect 200724 229752 200730 229764
rect 254670 229752 254676 229764
rect 200724 229724 254676 229752
rect 200724 229712 200730 229724
rect 254670 229712 254676 229724
rect 254728 229712 254734 229764
rect 255222 229712 255228 229764
rect 255280 229752 255286 229764
rect 278498 229752 278504 229764
rect 255280 229724 278504 229752
rect 255280 229712 255286 229724
rect 278498 229712 278504 229724
rect 278556 229712 278562 229764
rect 278682 229712 278688 229764
rect 278740 229752 278746 229764
rect 288526 229752 288532 229764
rect 278740 229724 288532 229752
rect 278740 229712 278746 229724
rect 288526 229712 288532 229724
rect 288584 229712 288590 229764
rect 302050 229712 302056 229764
rect 302108 229752 302114 229764
rect 311158 229752 311164 229764
rect 302108 229724 311164 229752
rect 302108 229712 302114 229724
rect 311158 229712 311164 229724
rect 311216 229712 311222 229764
rect 326338 229712 326344 229764
rect 326396 229752 326402 229764
rect 334710 229752 334716 229764
rect 326396 229724 334716 229752
rect 326396 229712 326402 229724
rect 334710 229712 334716 229724
rect 334768 229712 334774 229764
rect 344830 229712 344836 229764
rect 344888 229752 344894 229764
rect 406378 229752 406384 229764
rect 344888 229724 406384 229752
rect 344888 229712 344894 229724
rect 406378 229712 406384 229724
rect 406436 229712 406442 229764
rect 406654 229712 406660 229764
rect 406712 229752 406718 229764
rect 407684 229752 407712 229792
rect 406712 229724 407712 229752
rect 408972 229752 409000 229792
rect 409046 229780 409052 229832
rect 409104 229820 409110 229832
rect 411070 229820 411076 229832
rect 409104 229792 411076 229820
rect 409104 229780 409110 229792
rect 411070 229780 411076 229792
rect 411128 229780 411134 229832
rect 411548 229820 411576 229860
rect 551278 229848 551284 229860
rect 551336 229848 551342 229900
rect 563698 229820 563704 229832
rect 411548 229792 563704 229820
rect 563698 229780 563704 229792
rect 563756 229780 563762 229832
rect 411162 229752 411168 229764
rect 408972 229724 411168 229752
rect 406712 229712 406718 229724
rect 411162 229712 411168 229724
rect 411220 229712 411226 229764
rect 411530 229712 411536 229764
rect 411588 229752 411594 229764
rect 570598 229752 570604 229764
rect 411588 229724 570604 229752
rect 411588 229712 411594 229724
rect 570598 229712 570604 229724
rect 570656 229712 570662 229764
rect 140038 229644 140044 229696
rect 140096 229684 140102 229696
rect 205818 229684 205824 229696
rect 140096 229656 205824 229684
rect 140096 229644 140102 229656
rect 205818 229644 205824 229656
rect 205876 229644 205882 229696
rect 227530 229644 227536 229696
rect 227588 229684 227594 229696
rect 227588 229656 259776 229684
rect 227588 229644 227594 229656
rect 151814 229576 151820 229628
rect 151872 229616 151878 229628
rect 218974 229616 218980 229628
rect 151872 229588 218980 229616
rect 151872 229576 151878 229588
rect 218974 229576 218980 229588
rect 219032 229576 219038 229628
rect 248322 229576 248328 229628
rect 248380 229616 248386 229628
rect 248380 229588 258074 229616
rect 248380 229576 248386 229588
rect 149698 229508 149704 229560
rect 149756 229548 149762 229560
rect 216122 229548 216128 229560
rect 149756 229520 216128 229548
rect 149756 229508 149762 229520
rect 216122 229508 216128 229520
rect 216180 229508 216186 229560
rect 244918 229508 244924 229560
rect 244976 229548 244982 229560
rect 254302 229548 254308 229560
rect 244976 229520 254308 229548
rect 244976 229508 244982 229520
rect 254302 229508 254308 229520
rect 254360 229508 254366 229560
rect 146386 229440 146392 229492
rect 146444 229480 146450 229492
rect 209038 229480 209044 229492
rect 146444 229452 209044 229480
rect 146444 229440 146450 229452
rect 209038 229440 209044 229452
rect 209096 229440 209102 229492
rect 258046 229480 258074 229588
rect 259748 229548 259776 229656
rect 259914 229644 259920 229696
rect 259972 229684 259978 229696
rect 266078 229684 266084 229696
rect 259972 229656 266084 229684
rect 259972 229644 259978 229656
rect 266078 229644 266084 229656
rect 266136 229644 266142 229696
rect 268378 229644 268384 229696
rect 268436 229684 268442 229696
rect 277210 229684 277216 229696
rect 268436 229656 277216 229684
rect 268436 229644 268442 229656
rect 277210 229644 277216 229656
rect 277268 229644 277274 229696
rect 280062 229644 280068 229696
rect 280120 229684 280126 229696
rect 288894 229684 288900 229696
rect 280120 229656 288900 229684
rect 280120 229644 280126 229656
rect 288894 229644 288900 229656
rect 288952 229644 288958 229696
rect 323118 229644 323124 229696
rect 323176 229684 323182 229696
rect 340138 229684 340144 229696
rect 323176 229656 340144 229684
rect 323176 229644 323182 229656
rect 340138 229644 340144 229656
rect 340196 229644 340202 229696
rect 340874 229644 340880 229696
rect 340932 229684 340938 229696
rect 380250 229684 380256 229696
rect 340932 229656 380256 229684
rect 340932 229644 340938 229656
rect 380250 229644 380256 229656
rect 380308 229644 380314 229696
rect 400766 229644 400772 229696
rect 400824 229684 400830 229696
rect 453298 229684 453304 229696
rect 400824 229656 453304 229684
rect 400824 229644 400830 229656
rect 453298 229644 453304 229656
rect 453356 229644 453362 229696
rect 275646 229616 275652 229628
rect 267706 229588 275652 229616
rect 267090 229548 267096 229560
rect 259748 229520 267096 229548
rect 267090 229508 267096 229520
rect 267148 229508 267154 229560
rect 267706 229480 267734 229588
rect 275646 229576 275652 229588
rect 275704 229576 275710 229628
rect 277302 229576 277308 229628
rect 277360 229616 277366 229628
rect 277486 229616 277492 229628
rect 277360 229588 277492 229616
rect 277360 229576 277366 229588
rect 277486 229576 277492 229588
rect 277544 229576 277550 229628
rect 277670 229576 277676 229628
rect 277728 229616 277734 229628
rect 285674 229616 285680 229628
rect 277728 229588 285680 229616
rect 277728 229576 277734 229588
rect 285674 229576 285680 229588
rect 285732 229576 285738 229628
rect 313458 229576 313464 229628
rect 313516 229616 313522 229628
rect 314562 229616 314568 229628
rect 313516 229588 314568 229616
rect 313516 229576 313522 229588
rect 314562 229576 314568 229588
rect 314620 229576 314626 229628
rect 331674 229576 331680 229628
rect 331732 229616 331738 229628
rect 332410 229616 332416 229628
rect 331732 229588 332416 229616
rect 331732 229576 331738 229588
rect 332410 229576 332416 229588
rect 332468 229576 332474 229628
rect 341518 229616 341524 229628
rect 332520 229588 341524 229616
rect 270126 229508 270132 229560
rect 270184 229548 270190 229560
rect 271414 229548 271420 229560
rect 270184 229520 271420 229548
rect 270184 229508 270190 229520
rect 271414 229508 271420 229520
rect 271472 229508 271478 229560
rect 272978 229508 272984 229560
rect 273036 229548 273042 229560
rect 281074 229548 281080 229560
rect 273036 229520 281080 229548
rect 273036 229508 273042 229520
rect 281074 229508 281080 229520
rect 281132 229508 281138 229560
rect 300670 229508 300676 229560
rect 300728 229548 300734 229560
rect 305546 229548 305552 229560
rect 300728 229520 305552 229548
rect 300728 229508 300734 229520
rect 305546 229508 305552 229520
rect 305604 229508 305610 229560
rect 327350 229508 327356 229560
rect 327408 229548 327414 229560
rect 332520 229548 332548 229588
rect 341518 229576 341524 229588
rect 341576 229576 341582 229628
rect 350534 229576 350540 229628
rect 350592 229616 350598 229628
rect 387794 229616 387800 229628
rect 350592 229588 387800 229616
rect 350592 229576 350598 229588
rect 387794 229576 387800 229588
rect 387852 229576 387858 229628
rect 398098 229576 398104 229628
rect 398156 229616 398162 229628
rect 404354 229616 404360 229628
rect 398156 229588 404360 229616
rect 398156 229576 398162 229588
rect 404354 229576 404360 229588
rect 404412 229576 404418 229628
rect 407850 229576 407856 229628
rect 407908 229616 407914 229628
rect 449158 229616 449164 229628
rect 407908 229588 449164 229616
rect 407908 229576 407914 229588
rect 449158 229576 449164 229588
rect 449216 229576 449222 229628
rect 327408 229520 332548 229548
rect 327408 229508 327414 229520
rect 332686 229508 332692 229560
rect 332744 229548 332750 229560
rect 333790 229548 333796 229560
rect 332744 229520 333796 229548
rect 332744 229508 332750 229520
rect 333790 229508 333796 229520
rect 333848 229508 333854 229560
rect 338022 229508 338028 229560
rect 338080 229548 338086 229560
rect 352558 229548 352564 229560
rect 338080 229520 352564 229548
rect 338080 229508 338086 229520
rect 352558 229508 352564 229520
rect 352616 229508 352622 229560
rect 354858 229508 354864 229560
rect 354916 229548 354922 229560
rect 364242 229548 364248 229560
rect 354916 229520 364248 229548
rect 354916 229508 354922 229520
rect 364242 229508 364248 229520
rect 364300 229508 364306 229560
rect 366542 229508 366548 229560
rect 366600 229548 366606 229560
rect 409874 229548 409880 229560
rect 366600 229520 409880 229548
rect 366600 229508 366606 229520
rect 409874 229508 409880 229520
rect 409932 229508 409938 229560
rect 411898 229508 411904 229560
rect 411956 229548 411962 229560
rect 422294 229548 422300 229560
rect 411956 229520 422300 229548
rect 411956 229508 411962 229520
rect 422294 229508 422300 229520
rect 422352 229508 422358 229560
rect 258046 229452 267734 229480
rect 273898 229440 273904 229492
rect 273956 229480 273962 229492
rect 282822 229480 282828 229492
rect 273956 229452 282828 229480
rect 273956 229440 273962 229452
rect 282822 229440 282828 229452
rect 282880 229440 282886 229492
rect 339494 229440 339500 229492
rect 339552 229480 339558 229492
rect 353938 229480 353944 229492
rect 339552 229452 353944 229480
rect 339552 229440 339558 229452
rect 353938 229440 353944 229452
rect 353996 229440 354002 229492
rect 355502 229440 355508 229492
rect 355560 229480 355566 229492
rect 379514 229480 379520 229492
rect 355560 229452 379520 229480
rect 355560 229440 355566 229452
rect 379514 229440 379520 229452
rect 379572 229440 379578 229492
rect 382090 229440 382096 229492
rect 382148 229480 382154 229492
rect 393406 229480 393412 229492
rect 382148 229452 393412 229480
rect 382148 229440 382154 229452
rect 393406 229440 393412 229452
rect 393464 229440 393470 229492
rect 401502 229440 401508 229492
rect 401560 229480 401566 229492
rect 404998 229480 405004 229492
rect 401560 229452 405004 229480
rect 401560 229440 401566 229452
rect 404998 229440 405004 229452
rect 405056 229440 405062 229492
rect 407758 229440 407764 229492
rect 407816 229480 407822 229492
rect 438946 229480 438952 229492
rect 407816 229452 438952 229480
rect 407816 229440 407822 229452
rect 438946 229440 438952 229452
rect 439004 229440 439010 229492
rect 186958 229372 186964 229424
rect 187016 229412 187022 229424
rect 248966 229412 248972 229424
rect 187016 229384 248972 229412
rect 187016 229372 187022 229384
rect 248966 229372 248972 229384
rect 249024 229372 249030 229424
rect 275370 229372 275376 229424
rect 275428 229412 275434 229424
rect 284202 229412 284208 229424
rect 275428 229384 284208 229412
rect 275428 229372 275434 229384
rect 284202 229372 284208 229384
rect 284260 229372 284266 229424
rect 298462 229372 298468 229424
rect 298520 229412 298526 229424
rect 301130 229412 301136 229424
rect 298520 229384 301136 229412
rect 298520 229372 298526 229384
rect 301130 229372 301136 229384
rect 301188 229372 301194 229424
rect 310606 229372 310612 229424
rect 310664 229412 310670 229424
rect 314470 229412 314476 229424
rect 310664 229384 314476 229412
rect 310664 229372 310670 229384
rect 314470 229372 314476 229384
rect 314528 229372 314534 229424
rect 334526 229372 334532 229424
rect 334584 229412 334590 229424
rect 342898 229412 342904 229424
rect 334584 229384 342904 229412
rect 334584 229372 334590 229384
rect 342898 229372 342904 229384
rect 342956 229372 342962 229424
rect 361206 229372 361212 229424
rect 361264 229412 361270 229424
rect 382458 229412 382464 229424
rect 361264 229384 382464 229412
rect 361264 229372 361270 229384
rect 382458 229372 382464 229384
rect 382516 229372 382522 229424
rect 392210 229372 392216 229424
rect 392268 229412 392274 229424
rect 431954 229412 431960 229424
rect 392268 229384 431960 229412
rect 392268 229372 392274 229384
rect 431954 229372 431960 229384
rect 432012 229372 432018 229424
rect 162854 229304 162860 229356
rect 162912 229344 162918 229356
rect 223298 229344 223304 229356
rect 162912 229316 223304 229344
rect 162912 229304 162918 229316
rect 223298 229304 223304 229316
rect 223356 229304 223362 229356
rect 277486 229304 277492 229356
rect 277544 229344 277550 229356
rect 286686 229344 286692 229356
rect 277544 229316 286692 229344
rect 277544 229304 277550 229316
rect 286686 229304 286692 229316
rect 286744 229304 286750 229356
rect 296714 229304 296720 229356
rect 296772 229344 296778 229356
rect 300118 229344 300124 229356
rect 296772 229316 300124 229344
rect 296772 229304 296778 229316
rect 300118 229304 300124 229316
rect 300176 229304 300182 229356
rect 315206 229304 315212 229356
rect 315264 229344 315270 229356
rect 315264 229316 335354 229344
rect 315264 229304 315270 229316
rect 180794 229236 180800 229288
rect 180852 229276 180858 229288
rect 238938 229276 238944 229288
rect 180852 229248 238944 229276
rect 180852 229236 180858 229248
rect 238938 229236 238944 229248
rect 238996 229236 239002 229288
rect 271230 229236 271236 229288
rect 271288 229276 271294 229288
rect 279970 229276 279976 229288
rect 271288 229248 279976 229276
rect 271288 229236 271294 229248
rect 279970 229236 279976 229248
rect 280028 229236 280034 229288
rect 281442 229236 281448 229288
rect 281500 229276 281506 229288
rect 288158 229276 288164 229288
rect 281500 229248 288164 229276
rect 281500 229236 281506 229248
rect 288158 229236 288164 229248
rect 288216 229236 288222 229288
rect 296346 229236 296352 229288
rect 296404 229276 296410 229288
rect 298462 229276 298468 229288
rect 296404 229248 298468 229276
rect 296404 229236 296410 229248
rect 298462 229236 298468 229248
rect 298520 229236 298526 229288
rect 313090 229236 313096 229288
rect 313148 229276 313154 229288
rect 318058 229276 318064 229288
rect 313148 229248 318064 229276
rect 313148 229236 313154 229248
rect 318058 229236 318064 229248
rect 318116 229236 318122 229288
rect 335326 229276 335354 229316
rect 342346 229304 342352 229356
rect 342404 229344 342410 229356
rect 343266 229344 343272 229356
rect 342404 229316 343272 229344
rect 342404 229304 342410 229316
rect 343266 229304 343272 229316
rect 343324 229304 343330 229356
rect 363414 229304 363420 229356
rect 363472 229344 363478 229356
rect 364150 229344 364156 229356
rect 363472 229316 364156 229344
rect 363472 229304 363478 229316
rect 364150 229304 364156 229316
rect 364208 229304 364214 229356
rect 371970 229304 371976 229356
rect 372028 229344 372034 229356
rect 398098 229344 398104 229356
rect 372028 229316 398104 229344
rect 372028 229304 372034 229316
rect 398098 229304 398104 229316
rect 398156 229304 398162 229356
rect 407206 229304 407212 229356
rect 407264 229344 407270 229356
rect 411990 229344 411996 229356
rect 407264 229316 411996 229344
rect 407264 229304 407270 229316
rect 411990 229304 411996 229316
rect 412048 229304 412054 229356
rect 343818 229276 343824 229288
rect 335326 229248 343824 229276
rect 343818 229236 343824 229248
rect 343876 229236 343882 229288
rect 357710 229236 357716 229288
rect 357768 229276 357774 229288
rect 376110 229276 376116 229288
rect 357768 229248 376116 229276
rect 357768 229236 357774 229248
rect 376110 229236 376116 229248
rect 376168 229236 376174 229288
rect 379698 229236 379704 229288
rect 379756 229276 379762 229288
rect 379756 229248 383608 229276
rect 379756 229236 379762 229248
rect 255958 229168 255964 229220
rect 256016 229208 256022 229220
rect 260006 229208 260012 229220
rect 256016 229180 260012 229208
rect 256016 229168 256022 229180
rect 260006 229168 260012 229180
rect 260064 229168 260070 229220
rect 282822 229168 282828 229220
rect 282880 229208 282886 229220
rect 289262 229208 289268 229220
rect 282880 229180 289268 229208
rect 282880 229168 282886 229180
rect 289262 229168 289268 229180
rect 289320 229168 289326 229220
rect 295242 229168 295248 229220
rect 295300 229208 295306 229220
rect 296898 229208 296904 229220
rect 295300 229180 296904 229208
rect 295300 229168 295306 229180
rect 296898 229168 296904 229180
rect 296956 229168 296962 229220
rect 297450 229168 297456 229220
rect 297508 229208 297514 229220
rect 299474 229208 299480 229220
rect 297508 229180 299480 229208
rect 297508 229168 297514 229180
rect 299474 229168 299480 229180
rect 299532 229168 299538 229220
rect 324866 229168 324872 229220
rect 324924 229208 324930 229220
rect 325510 229208 325516 229220
rect 324924 229180 325516 229208
rect 324924 229168 324930 229180
rect 325510 229168 325516 229180
rect 325568 229168 325574 229220
rect 328454 229168 328460 229220
rect 328512 229208 328518 229220
rect 329558 229208 329564 229220
rect 328512 229180 329564 229208
rect 328512 229168 328518 229180
rect 329558 229168 329564 229180
rect 329616 229168 329622 229220
rect 369394 229168 369400 229220
rect 369452 229208 369458 229220
rect 382090 229208 382096 229220
rect 369452 229180 382096 229208
rect 369452 229168 369458 229180
rect 382090 229168 382096 229180
rect 382148 229168 382154 229220
rect 382274 229168 382280 229220
rect 382332 229208 382338 229220
rect 383470 229208 383476 229220
rect 382332 229180 383476 229208
rect 382332 229168 382338 229180
rect 383470 229168 383476 229180
rect 383528 229168 383534 229220
rect 383580 229208 383608 229248
rect 384390 229236 384396 229288
rect 384448 229276 384454 229288
rect 411254 229276 411260 229288
rect 384448 229248 411260 229276
rect 384448 229236 384454 229248
rect 411254 229236 411260 229248
rect 411312 229236 411318 229288
rect 386598 229208 386604 229220
rect 383580 229180 386604 229208
rect 386598 229168 386604 229180
rect 386656 229168 386662 229220
rect 386874 229168 386880 229220
rect 386932 229208 386938 229220
rect 388438 229208 388444 229220
rect 386932 229180 388444 229208
rect 386932 229168 386938 229180
rect 388438 229168 388444 229180
rect 388496 229168 388502 229220
rect 390094 229168 390100 229220
rect 390152 229208 390158 229220
rect 395338 229208 395344 229220
rect 390152 229180 395344 229208
rect 390152 229168 390158 229180
rect 395338 229168 395344 229180
rect 395396 229168 395402 229220
rect 395430 229168 395436 229220
rect 395488 229208 395494 229220
rect 407298 229208 407304 229220
rect 395488 229180 407304 229208
rect 395488 229168 395494 229180
rect 407298 229168 407304 229180
rect 407356 229168 407362 229220
rect 407390 229168 407396 229220
rect 407448 229208 407454 229220
rect 407758 229208 407764 229220
rect 407448 229180 407764 229208
rect 407448 229168 407454 229180
rect 407758 229168 407764 229180
rect 407816 229168 407822 229220
rect 410058 229168 410064 229220
rect 410116 229208 410122 229220
rect 416222 229208 416228 229220
rect 410116 229180 416228 229208
rect 410116 229168 410122 229180
rect 416222 229168 416228 229180
rect 416280 229168 416286 229220
rect 62114 229100 62120 229152
rect 62172 229140 62178 229152
rect 65150 229140 65156 229152
rect 62172 229112 65156 229140
rect 62172 229100 62178 229112
rect 65150 229100 65156 229112
rect 65208 229100 65214 229152
rect 257338 229100 257344 229152
rect 257396 229140 257402 229152
rect 258902 229140 258908 229152
rect 257396 229112 258908 229140
rect 257396 229100 257402 229112
rect 258902 229100 258908 229112
rect 258960 229100 258966 229152
rect 284202 229100 284208 229152
rect 284260 229140 284266 229152
rect 289538 229140 289544 229152
rect 284260 229112 289544 229140
rect 284260 229100 284266 229112
rect 289538 229100 289544 229112
rect 289596 229100 289602 229152
rect 292574 229100 292580 229152
rect 292632 229140 292638 229152
rect 293862 229140 293868 229152
rect 292632 229112 293868 229140
rect 292632 229100 292638 229112
rect 293862 229100 293868 229112
rect 293920 229100 293926 229152
rect 298094 229100 298100 229152
rect 298152 229140 298158 229152
rect 299382 229140 299388 229152
rect 298152 229112 299388 229140
rect 298152 229100 298158 229112
rect 299382 229100 299388 229112
rect 299440 229100 299446 229152
rect 299566 229100 299572 229152
rect 299624 229140 299630 229152
rect 300486 229140 300492 229152
rect 299624 229112 300492 229140
rect 299624 229100 299630 229112
rect 300486 229100 300492 229112
rect 300544 229100 300550 229152
rect 323486 229100 323492 229152
rect 323544 229140 323550 229152
rect 324222 229140 324228 229152
rect 323544 229112 324228 229140
rect 323544 229100 323550 229112
rect 324222 229100 324228 229112
rect 324280 229100 324286 229152
rect 324498 229100 324504 229152
rect 324556 229140 324562 229152
rect 325326 229140 325332 229152
rect 324556 229112 325332 229140
rect 324556 229100 324562 229112
rect 325326 229100 325332 229112
rect 325384 229100 325390 229152
rect 328822 229100 328828 229152
rect 328880 229140 328886 229152
rect 329650 229140 329656 229152
rect 328880 229112 329656 229140
rect 328880 229100 328886 229112
rect 329650 229100 329656 229112
rect 329708 229100 329714 229152
rect 329834 229100 329840 229152
rect 329892 229140 329898 229152
rect 331030 229140 331036 229152
rect 329892 229112 331036 229140
rect 329892 229100 329898 229112
rect 331030 229100 331036 229112
rect 331088 229100 331094 229152
rect 381170 229100 381176 229152
rect 381228 229140 381234 229152
rect 382182 229140 382188 229152
rect 381228 229112 382188 229140
rect 381228 229100 381234 229112
rect 382182 229100 382188 229112
rect 382240 229100 382246 229152
rect 382642 229100 382648 229152
rect 382700 229140 382706 229152
rect 383378 229140 383384 229152
rect 382700 229112 383384 229140
rect 382700 229100 382706 229112
rect 383378 229100 383384 229112
rect 383436 229100 383442 229152
rect 383654 229100 383660 229152
rect 383712 229140 383718 229152
rect 384942 229140 384948 229152
rect 383712 229112 384948 229140
rect 383712 229100 383718 229112
rect 384942 229100 384948 229112
rect 385000 229100 385006 229152
rect 385494 229100 385500 229152
rect 385552 229140 385558 229152
rect 386322 229140 386328 229152
rect 385552 229112 386328 229140
rect 385552 229100 385558 229112
rect 386322 229100 386328 229112
rect 386380 229100 386386 229152
rect 386506 229100 386512 229152
rect 386564 229140 386570 229152
rect 387702 229140 387708 229152
rect 386564 229112 387708 229140
rect 386564 229100 386570 229112
rect 387702 229100 387708 229112
rect 387760 229100 387766 229152
rect 405090 229100 405096 229152
rect 405148 229140 405154 229152
rect 409966 229140 409972 229152
rect 405148 229112 409972 229140
rect 405148 229100 405154 229112
rect 409966 229100 409972 229112
rect 410024 229100 410030 229152
rect 410886 229100 410892 229152
rect 410944 229140 410950 229152
rect 421006 229140 421012 229152
rect 410944 229112 421012 229140
rect 410944 229100 410950 229112
rect 421006 229100 421012 229112
rect 421064 229100 421070 229152
rect 120810 229032 120816 229084
rect 120868 229072 120874 229084
rect 220814 229072 220820 229084
rect 120868 229044 220820 229072
rect 120868 229032 120874 229044
rect 220814 229032 220820 229044
rect 220872 229032 220878 229084
rect 365162 229032 365168 229084
rect 365220 229072 365226 229084
rect 460934 229072 460940 229084
rect 365220 229044 460940 229072
rect 365220 229032 365226 229044
rect 460934 229032 460940 229044
rect 460992 229032 460998 229084
rect 117222 228964 117228 229016
rect 117280 229004 117286 229016
rect 219342 229004 219348 229016
rect 117280 228976 219348 229004
rect 117280 228964 117286 228976
rect 219342 228964 219348 228976
rect 219400 228964 219406 229016
rect 332042 228964 332048 229016
rect 332100 229004 332106 229016
rect 370222 229004 370228 229016
rect 332100 228976 370228 229004
rect 332100 228964 332106 228976
rect 370222 228964 370228 228976
rect 370280 228964 370286 229016
rect 373350 228964 373356 229016
rect 373408 229004 373414 229016
rect 480254 229004 480260 229016
rect 373408 228976 480260 229004
rect 373408 228964 373414 228976
rect 480254 228964 480260 228976
rect 480312 228964 480318 229016
rect 114186 228896 114192 228948
rect 114244 228936 114250 228948
rect 217962 228936 217968 228948
rect 114244 228908 217968 228936
rect 114244 228896 114250 228908
rect 217962 228896 217968 228908
rect 218020 228896 218026 228948
rect 224034 228896 224040 228948
rect 224092 228936 224098 228948
rect 234706 228936 234712 228948
rect 224092 228908 234712 228936
rect 224092 228896 224098 228908
rect 234706 228896 234712 228908
rect 234764 228896 234770 228948
rect 329190 228896 329196 228948
rect 329248 228936 329254 228948
rect 371326 228936 371332 228948
rect 329248 228908 371332 228936
rect 329248 228896 329254 228908
rect 371326 228896 371332 228908
rect 371384 228896 371390 228948
rect 375098 228896 375104 228948
rect 375156 228936 375162 228948
rect 483474 228936 483480 228948
rect 375156 228908 483480 228936
rect 375156 228896 375162 228908
rect 483474 228896 483480 228908
rect 483532 228896 483538 228948
rect 110690 228828 110696 228880
rect 110748 228868 110754 228880
rect 216490 228868 216496 228880
rect 110748 228840 216496 228868
rect 110748 228828 110754 228840
rect 216490 228828 216496 228840
rect 216548 228828 216554 228880
rect 227714 228828 227720 228880
rect 227772 228868 227778 228880
rect 240410 228868 240416 228880
rect 227772 228840 240416 228868
rect 227772 228828 227778 228840
rect 240410 228828 240416 228840
rect 240468 228828 240474 228880
rect 327718 228828 327724 228880
rect 327776 228868 327782 228880
rect 372706 228868 372712 228880
rect 327776 228840 372712 228868
rect 327776 228828 327782 228840
rect 372706 228828 372712 228840
rect 372764 228828 372770 228880
rect 376570 228828 376576 228880
rect 376628 228868 376634 228880
rect 487706 228868 487712 228880
rect 376628 228840 487712 228868
rect 376628 228828 376634 228840
rect 487706 228828 487712 228840
rect 487764 228828 487770 228880
rect 107470 228760 107476 228812
rect 107528 228800 107534 228812
rect 215110 228800 215116 228812
rect 107528 228772 215116 228800
rect 107528 228760 107534 228772
rect 215110 228760 215116 228772
rect 215168 228760 215174 228812
rect 216674 228760 216680 228812
rect 216732 228800 216738 228812
rect 224678 228800 224684 228812
rect 216732 228772 224684 228800
rect 216732 228760 216738 228772
rect 224678 228760 224684 228772
rect 224736 228760 224742 228812
rect 230290 228760 230296 228812
rect 230348 228800 230354 228812
rect 230348 228772 230612 228800
rect 230348 228760 230354 228772
rect 103974 228692 103980 228744
rect 104032 228732 104038 228744
rect 213638 228732 213644 228744
rect 104032 228704 213644 228732
rect 104032 228692 104038 228704
rect 213638 228692 213644 228704
rect 213696 228692 213702 228744
rect 222102 228692 222108 228744
rect 222160 228732 222166 228744
rect 230382 228732 230388 228744
rect 222160 228704 230388 228732
rect 222160 228692 222166 228704
rect 230382 228692 230388 228704
rect 230440 228692 230446 228744
rect 230584 228732 230612 228772
rect 233510 228760 233516 228812
rect 233568 228800 233574 228812
rect 268194 228800 268200 228812
rect 233568 228772 268200 228800
rect 233568 228760 233574 228772
rect 268194 228760 268200 228772
rect 268252 228760 268258 228812
rect 330570 228760 330576 228812
rect 330628 228800 330634 228812
rect 375282 228800 375288 228812
rect 330628 228772 375288 228800
rect 330628 228760 330634 228772
rect 375282 228760 375288 228772
rect 375340 228760 375346 228812
rect 377950 228760 377956 228812
rect 378008 228800 378014 228812
rect 491294 228800 491300 228812
rect 378008 228772 491300 228800
rect 378008 228760 378014 228772
rect 491294 228760 491300 228772
rect 491352 228760 491358 228812
rect 266722 228732 266728 228744
rect 230584 228704 266728 228732
rect 266722 228692 266728 228704
rect 266780 228692 266786 228744
rect 328086 228692 328092 228744
rect 328144 228732 328150 228744
rect 374086 228732 374092 228744
rect 328144 228704 374092 228732
rect 328144 228692 328150 228704
rect 374086 228692 374092 228704
rect 374144 228692 374150 228744
rect 391934 228692 391940 228744
rect 391992 228732 391998 228744
rect 523034 228732 523040 228744
rect 391992 228704 523040 228732
rect 391992 228692 391998 228704
rect 523034 228692 523040 228704
rect 523092 228692 523098 228744
rect 100662 228624 100668 228676
rect 100720 228664 100726 228676
rect 212258 228664 212264 228676
rect 100720 228636 212264 228664
rect 100720 228624 100726 228636
rect 212258 228624 212264 228636
rect 212316 228624 212322 228676
rect 215110 228624 215116 228676
rect 215168 228664 215174 228676
rect 260742 228664 260748 228676
rect 215168 228636 260748 228664
rect 215168 228624 215174 228636
rect 260742 228624 260748 228636
rect 260800 228624 260806 228676
rect 334894 228624 334900 228676
rect 334952 228664 334958 228676
rect 389266 228664 389272 228676
rect 334952 228636 389272 228664
rect 334952 228624 334958 228636
rect 389266 228624 389272 228636
rect 389324 228624 389330 228676
rect 392946 228624 392952 228676
rect 393004 228664 393010 228676
rect 526346 228664 526352 228676
rect 393004 228636 526352 228664
rect 393004 228624 393010 228636
rect 526346 228624 526352 228636
rect 526404 228624 526410 228676
rect 97258 228556 97264 228608
rect 97316 228596 97322 228608
rect 210786 228596 210792 228608
rect 97316 228568 210792 228596
rect 97316 228556 97322 228568
rect 210786 228556 210792 228568
rect 210844 228556 210850 228608
rect 213822 228556 213828 228608
rect 213880 228596 213886 228608
rect 258534 228596 258540 228608
rect 213880 228568 258540 228596
rect 213880 228556 213886 228568
rect 258534 228556 258540 228568
rect 258592 228556 258598 228608
rect 336274 228556 336280 228608
rect 336332 228596 336338 228608
rect 392578 228596 392584 228608
rect 336332 228568 392584 228596
rect 336332 228556 336338 228568
rect 392578 228556 392584 228568
rect 392636 228556 392642 228608
rect 397270 228556 397276 228608
rect 397328 228596 397334 228608
rect 536834 228596 536840 228608
rect 397328 228568 536840 228596
rect 397328 228556 397334 228568
rect 536834 228556 536840 228568
rect 536892 228556 536898 228608
rect 93762 228488 93768 228540
rect 93820 228528 93826 228540
rect 209406 228528 209412 228540
rect 93820 228500 209412 228528
rect 93820 228488 93826 228500
rect 209406 228488 209412 228500
rect 209464 228488 209470 228540
rect 209866 228488 209872 228540
rect 209924 228528 209930 228540
rect 257154 228528 257160 228540
rect 209924 228500 257160 228528
rect 209924 228488 209930 228500
rect 257154 228488 257160 228500
rect 257212 228488 257218 228540
rect 306650 228488 306656 228540
rect 306708 228528 306714 228540
rect 323670 228528 323676 228540
rect 306708 228500 323676 228528
rect 306708 228488 306714 228500
rect 323670 228488 323676 228500
rect 323728 228488 323734 228540
rect 337746 228488 337752 228540
rect 337804 228528 337810 228540
rect 396166 228528 396172 228540
rect 337804 228500 396172 228528
rect 337804 228488 337810 228500
rect 396166 228488 396172 228500
rect 396224 228488 396230 228540
rect 398282 228488 398288 228540
rect 398340 228528 398346 228540
rect 538214 228528 538220 228540
rect 398340 228500 538220 228528
rect 398340 228488 398346 228500
rect 538214 228488 538220 228500
rect 538272 228488 538278 228540
rect 56318 228420 56324 228472
rect 56376 228460 56382 228472
rect 193306 228460 193312 228472
rect 56376 228432 193312 228460
rect 56376 228420 56382 228432
rect 193306 228420 193312 228432
rect 193364 228420 193370 228472
rect 194962 228420 194968 228472
rect 195020 228460 195026 228472
rect 252186 228460 252192 228472
rect 195020 228432 252192 228460
rect 195020 228420 195026 228432
rect 252186 228420 252192 228432
rect 252244 228420 252250 228472
rect 276382 228460 276388 228472
rect 258046 228432 276388 228460
rect 53650 228352 53656 228404
rect 53708 228392 53714 228404
rect 192294 228392 192300 228404
rect 53708 228364 192300 228392
rect 53708 228352 53714 228364
rect 192294 228352 192300 228364
rect 192352 228352 192358 228404
rect 194134 228352 194140 228404
rect 194192 228392 194198 228404
rect 252830 228392 252836 228404
rect 194192 228364 252836 228392
rect 194192 228352 194198 228364
rect 252830 228352 252836 228364
rect 252888 228352 252894 228404
rect 127526 228284 127532 228336
rect 127584 228324 127590 228336
rect 223666 228324 223672 228336
rect 127584 228296 223672 228324
rect 127584 228284 127590 228296
rect 223666 228284 223672 228296
rect 223724 228284 223730 228336
rect 252002 228284 252008 228336
rect 252060 228324 252066 228336
rect 258046 228324 258074 228432
rect 276382 228420 276388 228432
rect 276440 228420 276446 228472
rect 309870 228420 309876 228472
rect 309928 228460 309934 228472
rect 327810 228460 327816 228472
rect 309928 228432 327816 228460
rect 309928 228420 309934 228432
rect 327810 228420 327816 228432
rect 327868 228420 327874 228472
rect 345198 228420 345204 228472
rect 345256 228460 345262 228472
rect 408494 228460 408500 228472
rect 345256 228432 408500 228460
rect 345256 228420 345262 228432
rect 408494 228420 408500 228432
rect 408552 228420 408558 228472
rect 409782 228420 409788 228472
rect 409840 228460 409846 228472
rect 553394 228460 553400 228472
rect 409840 228432 553400 228460
rect 409840 228420 409846 228432
rect 553394 228420 553400 228432
rect 553452 228420 553458 228472
rect 260558 228352 260564 228404
rect 260616 228392 260622 228404
rect 279602 228392 279608 228404
rect 260616 228364 279608 228392
rect 260616 228352 260622 228364
rect 279602 228352 279608 228364
rect 279660 228352 279666 228404
rect 294230 228392 294236 228404
rect 294064 228364 294236 228392
rect 252060 228296 258074 228324
rect 252060 228284 252066 228296
rect 131022 228216 131028 228268
rect 131080 228256 131086 228268
rect 225046 228256 225052 228268
rect 131080 228228 225052 228256
rect 131080 228216 131086 228228
rect 225046 228216 225052 228228
rect 225104 228216 225110 228268
rect 294064 228200 294092 228364
rect 294230 228352 294236 228364
rect 294288 228352 294294 228404
rect 308122 228352 308128 228404
rect 308180 228392 308186 228404
rect 327074 228392 327080 228404
rect 308180 228364 327080 228392
rect 308180 228352 308186 228364
rect 327074 228352 327080 228364
rect 327132 228352 327138 228404
rect 346302 228352 346308 228404
rect 346360 228392 346366 228404
rect 409966 228392 409972 228404
rect 346360 228364 409972 228392
rect 346360 228352 346366 228364
rect 409966 228352 409972 228364
rect 410024 228352 410030 228404
rect 410794 228352 410800 228404
rect 410852 228392 410858 228404
rect 568574 228392 568580 228404
rect 410852 228364 568580 228392
rect 410852 228352 410858 228364
rect 568574 228352 568580 228364
rect 568632 228352 568638 228404
rect 353386 228284 353392 228336
rect 353444 228324 353450 228336
rect 433334 228324 433340 228336
rect 353444 228296 433340 228324
rect 353444 228284 353450 228296
rect 433334 228284 433340 228296
rect 433392 228284 433398 228336
rect 349154 228216 349160 228268
rect 349212 228256 349218 228268
rect 422202 228256 422208 228268
rect 349212 228228 422208 228256
rect 349212 228216 349218 228228
rect 422202 228216 422208 228228
rect 422260 228216 422266 228268
rect 422294 228216 422300 228268
rect 422352 228256 422358 228268
rect 485130 228256 485136 228268
rect 422352 228228 485136 228256
rect 422352 228216 422358 228228
rect 485130 228216 485136 228228
rect 485188 228216 485194 228268
rect 137738 228148 137744 228200
rect 137796 228188 137802 228200
rect 227898 228188 227904 228200
rect 137796 228160 227904 228188
rect 137796 228148 137802 228160
rect 227898 228148 227904 228160
rect 227956 228148 227962 228200
rect 294046 228148 294052 228200
rect 294104 228148 294110 228200
rect 340598 228148 340604 228200
rect 340656 228188 340662 228200
rect 402974 228188 402980 228200
rect 340656 228160 402980 228188
rect 340656 228148 340662 228160
rect 402974 228148 402980 228160
rect 403032 228148 403038 228200
rect 404354 228148 404360 228200
rect 404412 228188 404418 228200
rect 476114 228188 476120 228200
rect 404412 228160 476120 228188
rect 404412 228148 404418 228160
rect 476114 228148 476120 228160
rect 476172 228148 476178 228200
rect 144362 228080 144368 228132
rect 144420 228120 144426 228132
rect 230750 228120 230756 228132
rect 144420 228092 230756 228120
rect 144420 228080 144426 228092
rect 230750 228080 230756 228092
rect 230808 228080 230814 228132
rect 334158 228080 334164 228132
rect 334216 228120 334222 228132
rect 378502 228120 378508 228132
rect 334216 228092 378508 228120
rect 334216 228080 334222 228092
rect 378502 228080 378508 228092
rect 378560 228080 378566 228132
rect 380710 228080 380716 228132
rect 380768 228120 380774 228132
rect 406010 228120 406016 228132
rect 380768 228092 406016 228120
rect 380768 228080 380774 228092
rect 406010 228080 406016 228092
rect 406068 228080 406074 228132
rect 407022 228080 407028 228132
rect 407080 228120 407086 228132
rect 454034 228120 454040 228132
rect 407080 228092 454040 228120
rect 407080 228080 407086 228092
rect 454034 228080 454040 228092
rect 454092 228080 454098 228132
rect 154482 228012 154488 228064
rect 154540 228052 154546 228064
rect 235074 228052 235080 228064
rect 154540 228024 235080 228052
rect 154540 228012 154546 228024
rect 235074 228012 235080 228024
rect 235132 228012 235138 228064
rect 343450 228012 343456 228064
rect 343508 228052 343514 228064
rect 387150 228052 387156 228064
rect 343508 228024 387156 228052
rect 343508 228012 343514 228024
rect 387150 228012 387156 228024
rect 387208 228012 387214 228064
rect 387794 228012 387800 228064
rect 387852 228052 387858 228064
rect 426434 228052 426440 228064
rect 387852 228024 426440 228052
rect 387852 228012 387858 228024
rect 426434 228012 426440 228024
rect 426492 228012 426498 228064
rect 161290 227944 161296 227996
rect 161348 227984 161354 227996
rect 237926 227984 237932 227996
rect 161348 227956 237932 227984
rect 161348 227944 161354 227956
rect 237926 227944 237932 227956
rect 237984 227944 237990 227996
rect 386414 227944 386420 227996
rect 386472 227984 386478 227996
rect 419534 227984 419540 227996
rect 386472 227956 419540 227984
rect 386472 227944 386478 227956
rect 419534 227944 419540 227956
rect 419592 227944 419598 227996
rect 171042 227876 171048 227928
rect 171100 227916 171106 227928
rect 242158 227916 242164 227928
rect 171100 227888 242164 227916
rect 171100 227876 171106 227888
rect 242158 227876 242164 227888
rect 242216 227876 242222 227928
rect 378226 227876 378232 227928
rect 378284 227916 378290 227928
rect 399386 227916 399392 227928
rect 378284 227888 399392 227916
rect 378284 227876 378290 227888
rect 399386 227876 399392 227888
rect 399444 227876 399450 227928
rect 403066 227876 403072 227928
rect 403124 227916 403130 227928
rect 429654 227916 429660 227928
rect 403124 227888 429660 227916
rect 403124 227876 403130 227888
rect 429654 227876 429660 227888
rect 429712 227876 429718 227928
rect 375466 227808 375472 227860
rect 375524 227848 375530 227860
rect 380986 227848 380992 227860
rect 375524 227820 380992 227848
rect 375524 227808 375530 227820
rect 380986 227808 380992 227820
rect 381044 227808 381050 227860
rect 77938 227740 77944 227792
rect 77996 227780 78002 227792
rect 82814 227780 82820 227792
rect 77996 227752 82820 227780
rect 77996 227740 78002 227752
rect 82814 227740 82820 227752
rect 82872 227740 82878 227792
rect 84654 227740 84660 227792
rect 84712 227780 84718 227792
rect 91738 227780 91744 227792
rect 84712 227752 91744 227780
rect 84712 227740 84718 227752
rect 91738 227740 91744 227752
rect 91796 227740 91802 227792
rect 377306 227740 377312 227792
rect 377364 227780 377370 227792
rect 380342 227780 380348 227792
rect 377364 227752 380348 227780
rect 377364 227740 377370 227752
rect 380342 227740 380348 227752
rect 380400 227740 380406 227792
rect 160370 227672 160376 227724
rect 160428 227712 160434 227724
rect 238570 227712 238576 227724
rect 160428 227684 238576 227712
rect 160428 227672 160434 227684
rect 238570 227672 238576 227684
rect 238628 227672 238634 227724
rect 364426 227672 364432 227724
rect 364484 227712 364490 227724
rect 457346 227712 457352 227724
rect 364484 227684 457352 227712
rect 364484 227672 364490 227684
rect 457346 227672 457352 227684
rect 457404 227672 457410 227724
rect 157058 227604 157064 227656
rect 157116 227644 157122 227656
rect 237190 227644 237196 227656
rect 157116 227616 237196 227644
rect 157116 227604 157122 227616
rect 237190 227604 237196 227616
rect 237248 227604 237254 227656
rect 358722 227604 358728 227656
rect 358780 227644 358786 227656
rect 444374 227644 444380 227656
rect 358780 227616 444380 227644
rect 358780 227604 358786 227616
rect 444374 227604 444380 227616
rect 444432 227604 444438 227656
rect 449158 227604 449164 227656
rect 449216 227644 449222 227656
rect 542998 227644 543004 227656
rect 449216 227616 543004 227644
rect 449216 227604 449222 227616
rect 542998 227604 543004 227616
rect 543056 227604 543062 227656
rect 153654 227536 153660 227588
rect 153712 227576 153718 227588
rect 235718 227576 235724 227588
rect 153712 227548 235724 227576
rect 153712 227536 153718 227548
rect 235718 227536 235724 227548
rect 235776 227536 235782 227588
rect 365898 227536 365904 227588
rect 365956 227576 365962 227588
rect 461210 227576 461216 227588
rect 365956 227548 461216 227576
rect 365956 227536 365962 227548
rect 461210 227536 461216 227548
rect 461268 227536 461274 227588
rect 461578 227536 461584 227588
rect 461636 227576 461642 227588
rect 552658 227576 552664 227588
rect 461636 227548 552664 227576
rect 461636 227536 461642 227548
rect 552658 227536 552664 227548
rect 552716 227536 552722 227588
rect 108206 227468 108212 227520
rect 108264 227508 108270 227520
rect 149698 227508 149704 227520
rect 108264 227480 149704 227508
rect 108264 227468 108270 227480
rect 149698 227468 149704 227480
rect 149756 227468 149762 227520
rect 150342 227468 150348 227520
rect 150400 227508 150406 227520
rect 234338 227508 234344 227520
rect 150400 227480 234344 227508
rect 150400 227468 150406 227480
rect 234338 227468 234344 227480
rect 234396 227468 234402 227520
rect 367278 227468 367284 227520
rect 367336 227508 367342 227520
rect 464154 227508 464160 227520
rect 367336 227480 464160 227508
rect 367336 227468 367342 227480
rect 464154 227468 464160 227480
rect 464212 227468 464218 227520
rect 147582 227400 147588 227452
rect 147640 227440 147646 227452
rect 232222 227440 232228 227452
rect 147640 227412 232228 227440
rect 147640 227400 147646 227412
rect 232222 227400 232228 227412
rect 232280 227400 232286 227452
rect 309502 227400 309508 227452
rect 309560 227440 309566 227452
rect 330386 227440 330392 227452
rect 309560 227412 330392 227440
rect 309560 227400 309566 227412
rect 330386 227400 330392 227412
rect 330444 227400 330450 227452
rect 368750 227400 368756 227452
rect 368808 227440 368814 227452
rect 467834 227440 467840 227452
rect 368808 227412 467840 227440
rect 368808 227400 368814 227412
rect 467834 227400 467840 227412
rect 467892 227400 467898 227452
rect 469214 227400 469220 227452
rect 469272 227440 469278 227452
rect 555418 227440 555424 227452
rect 469272 227412 555424 227440
rect 469272 227400 469278 227412
rect 555418 227400 555424 227412
rect 555476 227400 555482 227452
rect 91370 227332 91376 227384
rect 91428 227372 91434 227384
rect 146386 227372 146392 227384
rect 91428 227344 146392 227372
rect 91428 227332 91434 227344
rect 146386 227332 146392 227344
rect 146444 227332 146450 227384
rect 146938 227332 146944 227384
rect 146996 227372 147002 227384
rect 232866 227372 232872 227384
rect 146996 227344 232872 227372
rect 146996 227332 147002 227344
rect 232866 227332 232872 227344
rect 232924 227332 232930 227384
rect 315574 227332 315580 227384
rect 315632 227372 315638 227384
rect 341334 227372 341340 227384
rect 315632 227344 341340 227372
rect 315632 227332 315638 227344
rect 341334 227332 341340 227344
rect 341392 227332 341398 227384
rect 370130 227332 370136 227384
rect 370188 227372 370194 227384
rect 470870 227372 470876 227384
rect 370188 227344 470876 227372
rect 370188 227332 370194 227344
rect 470870 227332 470876 227344
rect 470928 227332 470934 227384
rect 143442 227264 143448 227316
rect 143500 227304 143506 227316
rect 231486 227304 231492 227316
rect 143500 227276 231492 227304
rect 143500 227264 143506 227276
rect 231486 227264 231492 227276
rect 231544 227264 231550 227316
rect 312722 227264 312728 227316
rect 312780 227304 312786 227316
rect 333974 227304 333980 227316
rect 312780 227276 333980 227304
rect 312780 227264 312786 227276
rect 333974 227264 333980 227276
rect 334032 227264 334038 227316
rect 335170 227264 335176 227316
rect 335228 227304 335234 227316
rect 363138 227304 363144 227316
rect 335228 227276 363144 227304
rect 335228 227264 335234 227276
rect 363138 227264 363144 227276
rect 363196 227264 363202 227316
rect 371602 227264 371608 227316
rect 371660 227304 371666 227316
rect 474182 227304 474188 227316
rect 371660 227276 474188 227304
rect 371660 227264 371666 227276
rect 474182 227264 474188 227276
rect 474240 227264 474246 227316
rect 141050 227196 141056 227248
rect 141108 227236 141114 227248
rect 229370 227236 229376 227248
rect 141108 227208 229376 227236
rect 141108 227196 141114 227208
rect 229370 227196 229376 227208
rect 229428 227196 229434 227248
rect 232774 227196 232780 227248
rect 232832 227236 232838 227248
rect 247494 227236 247500 227248
rect 232832 227208 247500 227236
rect 232832 227196 232838 227208
rect 247494 227196 247500 227208
rect 247552 227196 247558 227248
rect 318426 227196 318432 227248
rect 318484 227236 318490 227248
rect 348050 227236 348056 227248
rect 318484 227208 348056 227236
rect 318484 227196 318490 227208
rect 348050 227196 348056 227208
rect 348108 227196 348114 227248
rect 372982 227196 372988 227248
rect 373040 227236 373046 227248
rect 477586 227236 477592 227248
rect 373040 227208 477592 227236
rect 373040 227196 373046 227208
rect 477586 227196 477592 227208
rect 477644 227196 477650 227248
rect 478138 227196 478144 227248
rect 478196 227236 478202 227248
rect 500218 227236 500224 227248
rect 478196 227208 500224 227236
rect 478196 227196 478202 227208
rect 500218 227196 500224 227208
rect 500276 227196 500282 227248
rect 82722 227128 82728 227180
rect 82780 227168 82786 227180
rect 140038 227168 140044 227180
rect 82780 227140 140044 227168
rect 82780 227128 82786 227140
rect 140038 227128 140044 227140
rect 140096 227128 140102 227180
rect 140130 227128 140136 227180
rect 140188 227168 140194 227180
rect 230014 227168 230020 227180
rect 140188 227140 230020 227168
rect 140188 227128 140194 227140
rect 230014 227128 230020 227140
rect 230072 227128 230078 227180
rect 237374 227128 237380 227180
rect 237432 227168 237438 227180
rect 256050 227168 256056 227180
rect 237432 227140 256056 227168
rect 237432 227128 237438 227140
rect 256050 227128 256056 227140
rect 256108 227128 256114 227180
rect 258810 227128 258816 227180
rect 258868 227168 258874 227180
rect 279234 227168 279240 227180
rect 258868 227140 279240 227168
rect 258868 227128 258874 227140
rect 279234 227128 279240 227140
rect 279292 227128 279298 227180
rect 321278 227128 321284 227180
rect 321336 227168 321342 227180
rect 354766 227168 354772 227180
rect 321336 227140 354772 227168
rect 321336 227128 321342 227140
rect 354766 227128 354772 227140
rect 354824 227128 354830 227180
rect 374454 227128 374460 227180
rect 374512 227168 374518 227180
rect 480898 227168 480904 227180
rect 374512 227140 480904 227168
rect 374512 227128 374518 227140
rect 480898 227128 480904 227140
rect 480956 227128 480962 227180
rect 134242 227060 134248 227112
rect 134300 227100 134306 227112
rect 226518 227100 226524 227112
rect 134300 227072 226524 227100
rect 134300 227060 134306 227072
rect 226518 227060 226524 227072
rect 226576 227060 226582 227112
rect 234706 227060 234712 227112
rect 234764 227100 234770 227112
rect 253198 227100 253204 227112
rect 234764 227072 253204 227100
rect 234764 227060 234770 227072
rect 253198 227060 253204 227072
rect 253256 227060 253262 227112
rect 255130 227060 255136 227112
rect 255188 227100 255194 227112
rect 277854 227100 277860 227112
rect 255188 227072 277860 227100
rect 255188 227060 255194 227072
rect 277854 227060 277860 227072
rect 277912 227060 277918 227112
rect 329466 227060 329472 227112
rect 329524 227100 329530 227112
rect 365254 227100 365260 227112
rect 329524 227072 365260 227100
rect 329524 227060 329530 227072
rect 365254 227060 365260 227072
rect 365312 227060 365318 227112
rect 374822 227060 374828 227112
rect 374880 227100 374886 227112
rect 483106 227100 483112 227112
rect 374880 227072 483112 227100
rect 374880 227060 374886 227072
rect 483106 227060 483112 227072
rect 483164 227060 483170 227112
rect 124122 226992 124128 227044
rect 124180 227032 124186 227044
rect 222194 227032 222200 227044
rect 124180 227004 222200 227032
rect 124180 226992 124186 227004
rect 222194 226992 222200 227004
rect 222252 226992 222258 227044
rect 237006 226992 237012 227044
rect 237064 227032 237070 227044
rect 269574 227032 269580 227044
rect 237064 227004 269580 227032
rect 237064 226992 237070 227004
rect 269574 226992 269580 227004
rect 269632 226992 269638 227044
rect 305270 226992 305276 227044
rect 305328 227032 305334 227044
rect 320266 227032 320272 227044
rect 305328 227004 320272 227032
rect 305328 226992 305334 227004
rect 320266 226992 320272 227004
rect 320324 226992 320330 227044
rect 325602 226992 325608 227044
rect 325660 227032 325666 227044
rect 360286 227032 360292 227044
rect 325660 227004 360292 227032
rect 325660 226992 325666 227004
rect 360286 226992 360292 227004
rect 360344 226992 360350 227044
rect 409690 226992 409696 227044
rect 409748 227032 409754 227044
rect 565906 227032 565912 227044
rect 409748 227004 565912 227032
rect 409748 226992 409754 227004
rect 565906 226992 565912 227004
rect 565964 226992 565970 227044
rect 125042 226924 125048 226976
rect 125100 226964 125106 226976
rect 162854 226964 162860 226976
rect 125100 226936 162860 226964
rect 125100 226924 125106 226936
rect 162854 226924 162860 226936
rect 162912 226924 162918 226976
rect 163682 226924 163688 226976
rect 163740 226964 163746 226976
rect 239766 226964 239772 226976
rect 163740 226936 239772 226964
rect 163740 226924 163746 226936
rect 239766 226924 239772 226936
rect 239824 226924 239830 226976
rect 293954 226924 293960 226976
rect 294012 226964 294018 226976
rect 294598 226964 294604 226976
rect 294012 226936 294604 226964
rect 294012 226924 294018 226936
rect 294598 226924 294604 226936
rect 294656 226924 294662 226976
rect 363046 226924 363052 226976
rect 363104 226964 363110 226976
rect 454126 226964 454132 226976
rect 363104 226936 454132 226964
rect 363104 226924 363110 226936
rect 454126 226924 454132 226936
rect 454184 226924 454190 226976
rect 166902 226856 166908 226908
rect 166960 226896 166966 226908
rect 241422 226896 241428 226908
rect 166960 226868 241428 226896
rect 166960 226856 166966 226868
rect 241422 226856 241428 226868
rect 241480 226856 241486 226908
rect 361574 226856 361580 226908
rect 361632 226896 361638 226908
rect 450630 226896 450636 226908
rect 361632 226868 450636 226896
rect 361632 226856 361638 226868
rect 450630 226856 450636 226868
rect 450688 226856 450694 226908
rect 164602 226788 164608 226840
rect 164660 226828 164666 226840
rect 239306 226828 239312 226840
rect 164660 226800 239312 226828
rect 164660 226788 164666 226800
rect 239306 226788 239312 226800
rect 239364 226788 239370 226840
rect 360194 226788 360200 226840
rect 360252 226828 360258 226840
rect 447318 226828 447324 226840
rect 360252 226800 447324 226828
rect 360252 226788 360258 226800
rect 447318 226788 447324 226800
rect 447376 226788 447382 226840
rect 173802 226720 173808 226772
rect 173860 226760 173866 226772
rect 244274 226760 244280 226772
rect 173860 226732 244280 226760
rect 173860 226720 173866 226732
rect 244274 226720 244280 226732
rect 244332 226720 244338 226772
rect 357342 226720 357348 226772
rect 357400 226760 357406 226772
rect 440602 226760 440608 226772
rect 357400 226732 440608 226760
rect 357400 226720 357406 226732
rect 440602 226720 440608 226732
rect 440660 226720 440666 226772
rect 42150 226652 42156 226704
rect 42208 226692 42214 226704
rect 44358 226692 44364 226704
rect 42208 226664 44364 226692
rect 42208 226652 42214 226664
rect 44358 226652 44364 226664
rect 44416 226652 44422 226704
rect 174630 226652 174636 226704
rect 174688 226692 174694 226704
rect 243630 226692 243636 226704
rect 174688 226664 243636 226692
rect 174688 226652 174694 226664
rect 243630 226652 243636 226664
rect 243688 226652 243694 226704
rect 355870 226652 355876 226704
rect 355928 226692 355934 226704
rect 437474 226692 437480 226704
rect 355928 226664 437480 226692
rect 355928 226652 355934 226664
rect 437474 226652 437480 226664
rect 437532 226652 437538 226704
rect 177206 226584 177212 226636
rect 177264 226624 177270 226636
rect 245746 226624 245752 226636
rect 177264 226596 245752 226624
rect 177264 226584 177270 226596
rect 245746 226584 245752 226596
rect 245804 226584 245810 226636
rect 354490 226584 354496 226636
rect 354548 226624 354554 226636
rect 433794 226624 433800 226636
rect 354548 226596 433800 226624
rect 354548 226584 354554 226596
rect 433794 226584 433800 226596
rect 433852 226584 433858 226636
rect 190270 226516 190276 226568
rect 190328 226556 190334 226568
rect 251450 226556 251456 226568
rect 190328 226528 251456 226556
rect 190328 226516 190334 226528
rect 251450 226516 251456 226528
rect 251508 226516 251514 226568
rect 351638 226516 351644 226568
rect 351696 226556 351702 226568
rect 427078 226556 427084 226568
rect 351696 226528 427084 226556
rect 351696 226516 351702 226528
rect 427078 226516 427084 226528
rect 427136 226516 427142 226568
rect 124858 226312 124864 226364
rect 124916 226352 124922 226364
rect 130378 226352 130384 226364
rect 124916 226324 130384 226352
rect 124916 226312 124922 226324
rect 130378 226312 130384 226324
rect 130436 226312 130442 226364
rect 116578 226244 116584 226296
rect 116636 226284 116642 226296
rect 220078 226284 220084 226296
rect 116636 226256 220084 226284
rect 116636 226244 116642 226256
rect 220078 226244 220084 226256
rect 220136 226244 220142 226296
rect 364058 226244 364064 226296
rect 364116 226284 364122 226296
rect 455690 226284 455696 226296
rect 364116 226256 455696 226284
rect 364116 226244 364122 226256
rect 455690 226244 455696 226256
rect 455748 226244 455754 226296
rect 456150 226244 456156 226296
rect 456208 226284 456214 226296
rect 548150 226284 548156 226296
rect 456208 226256 548156 226284
rect 456208 226244 456214 226256
rect 548150 226244 548156 226256
rect 548208 226244 548214 226296
rect 42150 226176 42156 226228
rect 42208 226216 42214 226228
rect 42978 226216 42984 226228
rect 42208 226188 42984 226216
rect 42208 226176 42214 226188
rect 42978 226176 42984 226188
rect 43036 226176 43042 226228
rect 112990 226176 112996 226228
rect 113048 226216 113054 226228
rect 218606 226216 218612 226228
rect 113048 226188 218612 226216
rect 113048 226176 113054 226188
rect 218606 226176 218612 226188
rect 218664 226176 218670 226228
rect 223114 226176 223120 226228
rect 223172 226216 223178 226228
rect 233234 226216 233240 226228
rect 223172 226188 233240 226216
rect 223172 226176 223178 226188
rect 233234 226176 233240 226188
rect 233292 226176 233298 226228
rect 365530 226176 365536 226228
rect 365588 226216 365594 226228
rect 459554 226216 459560 226228
rect 365588 226188 459560 226216
rect 365588 226176 365594 226188
rect 459554 226176 459560 226188
rect 459612 226176 459618 226228
rect 109862 226108 109868 226160
rect 109920 226148 109926 226160
rect 217226 226148 217232 226160
rect 109920 226120 217232 226148
rect 109920 226108 109926 226120
rect 217226 226108 217232 226120
rect 217284 226108 217290 226160
rect 218054 226108 218060 226160
rect 218112 226148 218118 226160
rect 227254 226148 227260 226160
rect 218112 226120 227260 226148
rect 218112 226108 218118 226120
rect 227254 226108 227260 226120
rect 227312 226108 227318 226160
rect 227346 226108 227352 226160
rect 227404 226148 227410 226160
rect 237558 226148 237564 226160
rect 227404 226120 237564 226148
rect 227404 226108 227410 226120
rect 237558 226108 237564 226120
rect 237616 226108 237622 226160
rect 366910 226108 366916 226160
rect 366968 226148 366974 226160
rect 462406 226148 462412 226160
rect 366968 226120 462412 226148
rect 366968 226108 366974 226120
rect 462406 226108 462412 226120
rect 462464 226108 462470 226160
rect 106550 226040 106556 226092
rect 106608 226080 106614 226092
rect 215754 226080 215760 226092
rect 106608 226052 215760 226080
rect 106608 226040 106614 226052
rect 215754 226040 215760 226052
rect 215812 226040 215818 226092
rect 224954 226040 224960 226092
rect 225012 226080 225018 226092
rect 251818 226080 251824 226092
rect 225012 226052 251824 226080
rect 225012 226040 225018 226052
rect 251818 226040 251824 226052
rect 251876 226040 251882 226092
rect 253842 226040 253848 226092
rect 253900 226080 253906 226092
rect 276474 226080 276480 226092
rect 253900 226052 276480 226080
rect 253900 226040 253906 226052
rect 276474 226040 276480 226052
rect 276532 226040 276538 226092
rect 335906 226040 335912 226092
rect 335964 226080 335970 226092
rect 367646 226080 367652 226092
rect 335964 226052 367652 226080
rect 335964 226040 335970 226052
rect 367646 226040 367652 226052
rect 367704 226040 367710 226092
rect 368382 226040 368388 226092
rect 368440 226080 368446 226092
rect 465074 226080 465080 226092
rect 368440 226052 465080 226080
rect 368440 226040 368446 226052
rect 465074 226040 465080 226052
rect 465132 226040 465138 226092
rect 103238 225972 103244 226024
rect 103296 226012 103302 226024
rect 214374 226012 214380 226024
rect 103296 225984 214380 226012
rect 103296 225972 103302 225984
rect 214374 225972 214380 225984
rect 214432 225972 214438 226024
rect 220630 225972 220636 226024
rect 220688 226012 220694 226024
rect 264238 226012 264244 226024
rect 220688 225984 264244 226012
rect 220688 225972 220694 225984
rect 264238 225972 264244 225984
rect 264296 225972 264302 226024
rect 322750 225972 322756 226024
rect 322808 226012 322814 226024
rect 358170 226012 358176 226024
rect 322808 225984 358176 226012
rect 322808 225972 322814 225984
rect 358170 225972 358176 225984
rect 358228 225972 358234 226024
rect 369762 225972 369768 226024
rect 369820 226012 369826 226024
rect 469214 226012 469220 226024
rect 369820 225984 469220 226012
rect 369820 225972 369826 225984
rect 469214 225972 469220 225984
rect 469272 225972 469278 226024
rect 99834 225904 99840 225956
rect 99892 225944 99898 225956
rect 212902 225944 212908 225956
rect 99892 225916 212908 225944
rect 99892 225904 99898 225916
rect 212902 225904 212908 225916
rect 212960 225904 212966 225956
rect 215294 225904 215300 225956
rect 215352 225944 215358 225956
rect 261386 225944 261392 225956
rect 215352 225916 261392 225944
rect 215352 225904 215358 225916
rect 261386 225904 261392 225916
rect 261444 225904 261450 225956
rect 326982 225904 326988 225956
rect 327040 225944 327046 225956
rect 362954 225944 362960 225956
rect 327040 225916 362960 225944
rect 327040 225904 327046 225916
rect 362954 225904 362960 225916
rect 363012 225904 363018 225956
rect 371234 225904 371240 225956
rect 371292 225944 371298 225956
rect 471974 225944 471980 225956
rect 371292 225916 471980 225944
rect 371292 225904 371298 225916
rect 471974 225904 471980 225916
rect 472032 225904 472038 225956
rect 96522 225836 96528 225888
rect 96580 225876 96586 225888
rect 211522 225876 211528 225888
rect 96580 225848 211528 225876
rect 96580 225836 96586 225848
rect 211522 225836 211528 225848
rect 211580 225836 211586 225888
rect 211706 225836 211712 225888
rect 211764 225876 211770 225888
rect 258994 225876 259000 225888
rect 211764 225848 259000 225876
rect 211764 225836 211770 225848
rect 258994 225836 259000 225848
rect 259052 225836 259058 225888
rect 356974 225836 356980 225888
rect 357032 225876 357038 225888
rect 438854 225876 438860 225888
rect 357032 225848 438860 225876
rect 357032 225836 357038 225848
rect 438854 225836 438860 225848
rect 438912 225836 438918 225888
rect 438946 225836 438952 225888
rect 439004 225876 439010 225888
rect 540422 225876 540428 225888
rect 439004 225848 540428 225876
rect 439004 225836 439010 225848
rect 540422 225836 540428 225848
rect 540480 225836 540486 225888
rect 86310 225768 86316 225820
rect 86368 225808 86374 225820
rect 207198 225808 207204 225820
rect 86368 225780 207204 225808
rect 86368 225768 86374 225780
rect 207198 225768 207204 225780
rect 207256 225768 207262 225820
rect 208302 225768 208308 225820
rect 208360 225808 208366 225820
rect 257890 225808 257896 225820
rect 208360 225780 257896 225808
rect 208360 225768 208366 225780
rect 257890 225768 257896 225780
rect 257948 225768 257954 225820
rect 324130 225768 324136 225820
rect 324188 225808 324194 225820
rect 361574 225808 361580 225820
rect 324188 225780 361580 225808
rect 324188 225768 324194 225780
rect 361574 225768 361580 225780
rect 361632 225768 361638 225820
rect 372614 225768 372620 225820
rect 372672 225808 372678 225820
rect 476206 225808 476212 225820
rect 372672 225780 476212 225808
rect 372672 225768 372678 225780
rect 476206 225768 476212 225780
rect 476264 225768 476270 225820
rect 76282 225700 76288 225752
rect 76340 225740 76346 225752
rect 202966 225740 202972 225752
rect 76340 225712 202972 225740
rect 76340 225700 76346 225712
rect 202966 225700 202972 225712
rect 203024 225700 203030 225752
rect 206830 225700 206836 225752
rect 206888 225740 206894 225752
rect 256786 225740 256792 225752
rect 206888 225712 256792 225740
rect 206888 225700 206894 225712
rect 256786 225700 256792 225712
rect 256844 225700 256850 225752
rect 303798 225700 303804 225752
rect 303856 225740 303862 225752
rect 317414 225740 317420 225752
rect 303856 225712 317420 225740
rect 303856 225700 303862 225712
rect 317414 225700 317420 225712
rect 317472 225700 317478 225752
rect 343082 225700 343088 225752
rect 343140 225740 343146 225752
rect 407114 225740 407120 225752
rect 343140 225712 407120 225740
rect 343140 225700 343146 225712
rect 407114 225700 407120 225712
rect 407172 225700 407178 225752
rect 407298 225700 407304 225752
rect 407356 225740 407362 225752
rect 531406 225740 531412 225752
rect 407356 225712 531412 225740
rect 407356 225700 407362 225712
rect 531406 225700 531412 225712
rect 531464 225700 531470 225752
rect 539594 225700 539600 225752
rect 539652 225740 539658 225752
rect 560846 225740 560852 225752
rect 539652 225712 560852 225740
rect 539652 225700 539658 225712
rect 560846 225700 560852 225712
rect 560904 225700 560910 225752
rect 56042 225632 56048 225684
rect 56100 225672 56106 225684
rect 194410 225672 194416 225684
rect 56100 225644 194416 225672
rect 56100 225632 56106 225644
rect 194410 225632 194416 225644
rect 194468 225632 194474 225684
rect 199010 225632 199016 225684
rect 199068 225672 199074 225684
rect 200666 225672 200672 225684
rect 199068 225644 200672 225672
rect 199068 225632 199074 225644
rect 200666 225632 200672 225644
rect 200724 225632 200730 225684
rect 203242 225632 203248 225684
rect 203300 225672 203306 225684
rect 255314 225672 255320 225684
rect 203300 225644 255320 225672
rect 203300 225632 203306 225644
rect 255314 225632 255320 225644
rect 255372 225632 255378 225684
rect 263410 225632 263416 225684
rect 263468 225672 263474 225684
rect 280982 225672 280988 225684
rect 263468 225644 280988 225672
rect 263468 225632 263474 225644
rect 280982 225632 280988 225644
rect 281040 225632 281046 225684
rect 302418 225632 302424 225684
rect 302476 225672 302482 225684
rect 313550 225672 313556 225684
rect 302476 225644 313556 225672
rect 302476 225632 302482 225644
rect 313550 225632 313556 225644
rect 313608 225632 313614 225684
rect 314470 225632 314476 225684
rect 314528 225672 314534 225684
rect 331214 225672 331220 225684
rect 314528 225644 331220 225672
rect 314528 225632 314534 225644
rect 331214 225632 331220 225644
rect 331272 225632 331278 225684
rect 341610 225632 341616 225684
rect 341668 225672 341674 225684
rect 403526 225672 403532 225684
rect 341668 225644 403532 225672
rect 341668 225632 341674 225644
rect 403526 225632 403532 225644
rect 403584 225632 403590 225684
rect 403618 225632 403624 225684
rect 403676 225672 403682 225684
rect 552014 225672 552020 225684
rect 403676 225644 552020 225672
rect 403676 225632 403682 225644
rect 552014 225632 552020 225644
rect 552072 225632 552078 225684
rect 52730 225564 52736 225616
rect 52788 225604 52794 225616
rect 192662 225604 192668 225616
rect 52788 225576 192668 225604
rect 52788 225564 52794 225576
rect 192662 225564 192668 225576
rect 192720 225564 192726 225616
rect 201402 225564 201408 225616
rect 201460 225604 201466 225616
rect 255038 225604 255044 225616
rect 201460 225576 255044 225604
rect 201460 225564 201466 225576
rect 255038 225564 255044 225576
rect 255096 225564 255102 225616
rect 257062 225564 257068 225616
rect 257120 225604 257126 225616
rect 278130 225604 278136 225616
rect 257120 225576 278136 225604
rect 257120 225564 257126 225576
rect 278130 225564 278136 225576
rect 278188 225564 278194 225616
rect 310974 225564 310980 225616
rect 311032 225604 311038 225616
rect 334066 225604 334072 225616
rect 311032 225576 334072 225604
rect 311032 225564 311038 225576
rect 334066 225564 334072 225576
rect 334124 225564 334130 225616
rect 344462 225564 344468 225616
rect 344520 225604 344526 225616
rect 410242 225604 410248 225616
rect 344520 225576 410248 225604
rect 344520 225564 344526 225576
rect 410242 225564 410248 225576
rect 410300 225564 410306 225616
rect 410978 225564 410984 225616
rect 411036 225604 411042 225616
rect 559190 225604 559196 225616
rect 411036 225576 559196 225604
rect 411036 225564 411042 225576
rect 559190 225564 559196 225576
rect 559248 225564 559254 225616
rect 119890 225496 119896 225548
rect 119948 225536 119954 225548
rect 221182 225536 221188 225548
rect 119948 225508 221188 225536
rect 119948 225496 119954 225508
rect 221182 225496 221188 225508
rect 221240 225496 221246 225548
rect 362862 225496 362868 225548
rect 362920 225536 362926 225548
rect 452654 225536 452660 225548
rect 362920 225508 452660 225536
rect 362920 225496 362926 225508
rect 452654 225496 452660 225508
rect 452712 225496 452718 225548
rect 123386 225428 123392 225480
rect 123444 225468 123450 225480
rect 222930 225468 222936 225480
rect 123444 225440 222936 225468
rect 123444 225428 123450 225440
rect 222930 225428 222936 225440
rect 222988 225428 222994 225480
rect 359826 225428 359832 225480
rect 359884 225468 359890 225480
rect 445754 225468 445760 225480
rect 359884 225440 445760 225468
rect 359884 225428 359890 225440
rect 445754 225428 445760 225440
rect 445812 225428 445818 225480
rect 126790 225360 126796 225412
rect 126848 225400 126854 225412
rect 224310 225400 224316 225412
rect 126848 225372 224316 225400
rect 126848 225360 126854 225372
rect 224310 225360 224316 225372
rect 224368 225360 224374 225412
rect 358354 225360 358360 225412
rect 358412 225400 358418 225412
rect 441614 225400 441620 225412
rect 358412 225372 441620 225400
rect 358412 225360 358418 225372
rect 441614 225360 441620 225372
rect 441672 225360 441678 225412
rect 130102 225292 130108 225344
rect 130160 225332 130166 225344
rect 225782 225332 225788 225344
rect 130160 225304 225788 225332
rect 130160 225292 130166 225304
rect 225782 225292 225788 225304
rect 225840 225292 225846 225344
rect 348786 225292 348792 225344
rect 348844 225332 348850 225344
rect 420362 225332 420368 225344
rect 348844 225304 420368 225332
rect 348844 225292 348850 225304
rect 420362 225292 420368 225304
rect 420420 225292 420426 225344
rect 133506 225224 133512 225276
rect 133564 225264 133570 225276
rect 227162 225264 227168 225276
rect 133564 225236 227168 225264
rect 133564 225224 133570 225236
rect 227162 225224 227168 225236
rect 227220 225224 227226 225276
rect 345934 225224 345940 225276
rect 345992 225264 345998 225276
rect 414014 225264 414020 225276
rect 345992 225236 414020 225264
rect 345992 225224 345998 225236
rect 414014 225224 414020 225236
rect 414072 225224 414078 225276
rect 170490 225156 170496 225208
rect 170548 225196 170554 225208
rect 242894 225196 242900 225208
rect 170548 225168 242900 225196
rect 170548 225156 170554 225168
rect 242894 225156 242900 225168
rect 242952 225156 242958 225208
rect 339034 225156 339040 225208
rect 339092 225196 339098 225208
rect 382274 225196 382280 225208
rect 339092 225168 382280 225196
rect 339092 225156 339098 225168
rect 382274 225156 382280 225168
rect 382332 225156 382338 225208
rect 382458 225156 382464 225208
rect 382516 225196 382522 225208
rect 448974 225196 448980 225208
rect 382516 225168 448980 225196
rect 382516 225156 382522 225168
rect 448974 225156 448980 225168
rect 449032 225156 449038 225208
rect 180610 225088 180616 225140
rect 180668 225128 180674 225140
rect 247126 225128 247132 225140
rect 180668 225100 247132 225128
rect 180668 225088 180674 225100
rect 247126 225088 247132 225100
rect 247184 225088 247190 225140
rect 340230 225088 340236 225140
rect 340288 225128 340294 225140
rect 385494 225128 385500 225140
rect 340288 225100 385500 225128
rect 340288 225088 340294 225100
rect 385494 225088 385500 225100
rect 385552 225088 385558 225140
rect 386598 225088 386604 225140
rect 386656 225128 386662 225140
rect 434714 225128 434720 225140
rect 386656 225100 434720 225128
rect 386656 225088 386662 225100
rect 434714 225088 434720 225100
rect 434772 225088 434778 225140
rect 192846 224952 192852 225004
rect 192904 224992 192910 225004
rect 197630 224992 197636 225004
rect 192904 224964 197636 224992
rect 192904 224952 192910 224964
rect 197630 224952 197636 224964
rect 197688 224952 197694 225004
rect 162762 224884 162768 224936
rect 162820 224924 162826 224936
rect 238202 224924 238208 224936
rect 162820 224896 238208 224924
rect 162820 224884 162826 224896
rect 238202 224884 238208 224896
rect 238260 224884 238266 224936
rect 368014 224884 368020 224936
rect 368072 224924 368078 224936
rect 468294 224924 468300 224936
rect 368072 224896 468300 224924
rect 368072 224884 368078 224896
rect 468294 224884 468300 224896
rect 468352 224884 468358 224936
rect 159542 224816 159548 224868
rect 159600 224856 159606 224868
rect 236822 224856 236828 224868
rect 159600 224828 236828 224856
rect 159600 224816 159606 224828
rect 236822 224816 236828 224828
rect 236880 224816 236886 224868
rect 377398 224816 377404 224868
rect 377456 224856 377462 224868
rect 479242 224856 479248 224868
rect 377456 224828 479248 224856
rect 377456 224816 377462 224828
rect 479242 224816 479248 224828
rect 479300 224816 479306 224868
rect 155770 224748 155776 224800
rect 155828 224788 155834 224800
rect 235350 224788 235356 224800
rect 155828 224760 235356 224788
rect 155828 224748 155834 224760
rect 235350 224748 235356 224760
rect 235408 224748 235414 224800
rect 370866 224748 370872 224800
rect 370924 224788 370930 224800
rect 475010 224788 475016 224800
rect 370924 224760 475016 224788
rect 370924 224748 370930 224760
rect 475010 224748 475016 224760
rect 475068 224748 475074 224800
rect 114922 224680 114928 224732
rect 114980 224720 114986 224732
rect 151814 224720 151820 224732
rect 114980 224692 151820 224720
rect 114980 224680 114986 224692
rect 151814 224680 151820 224692
rect 151872 224680 151878 224732
rect 152918 224680 152924 224732
rect 152976 224720 152982 224732
rect 233970 224720 233976 224732
rect 152976 224692 233976 224720
rect 152976 224680 152982 224692
rect 233970 224680 233976 224692
rect 234028 224680 234034 224732
rect 372246 224680 372252 224732
rect 372304 224720 372310 224732
rect 478966 224720 478972 224732
rect 372304 224692 478972 224720
rect 372304 224680 372310 224692
rect 478966 224680 478972 224692
rect 479024 224680 479030 224732
rect 149422 224612 149428 224664
rect 149480 224652 149486 224664
rect 232314 224652 232320 224664
rect 149480 224624 232320 224652
rect 149480 224612 149486 224624
rect 232314 224612 232320 224624
rect 232372 224612 232378 224664
rect 373718 224612 373724 224664
rect 373776 224652 373782 224664
rect 481818 224652 481824 224664
rect 373776 224624 481824 224652
rect 373776 224612 373782 224624
rect 481818 224612 481824 224624
rect 481876 224612 481882 224664
rect 146110 224544 146116 224596
rect 146168 224584 146174 224596
rect 231118 224584 231124 224596
rect 146168 224556 231124 224584
rect 146168 224544 146174 224556
rect 231118 224544 231124 224556
rect 231176 224544 231182 224596
rect 335538 224544 335544 224596
rect 335596 224584 335602 224596
rect 377306 224584 377312 224596
rect 335596 224556 377312 224584
rect 335596 224544 335602 224556
rect 377306 224544 377312 224556
rect 377364 224544 377370 224596
rect 388714 224544 388720 224596
rect 388772 224584 388778 224596
rect 516226 224584 516232 224596
rect 388772 224556 516232 224584
rect 388772 224544 388778 224556
rect 516226 224544 516232 224556
rect 516284 224544 516290 224596
rect 142706 224476 142712 224528
rect 142764 224516 142770 224528
rect 229646 224516 229652 224528
rect 142764 224488 229652 224516
rect 142764 224476 142770 224488
rect 229646 224476 229652 224488
rect 229704 224476 229710 224528
rect 332318 224476 332324 224528
rect 332376 224516 332382 224528
rect 372614 224516 372620 224528
rect 332376 224488 372620 224516
rect 332376 224476 332382 224488
rect 372614 224476 372620 224488
rect 372672 224476 372678 224528
rect 389726 224476 389732 224528
rect 389784 224516 389790 224528
rect 518894 224516 518900 224528
rect 389784 224488 518900 224516
rect 389784 224476 389790 224488
rect 518894 224476 518900 224488
rect 518952 224476 518958 224528
rect 139210 224408 139216 224460
rect 139268 224448 139274 224460
rect 228266 224448 228272 224460
rect 139268 224420 228272 224448
rect 139268 224408 139274 224420
rect 228266 224408 228272 224420
rect 228324 224408 228330 224460
rect 234614 224408 234620 224460
rect 234672 224448 234678 224460
rect 250346 224448 250352 224460
rect 234672 224420 250352 224448
rect 234672 224408 234678 224420
rect 250346 224408 250352 224420
rect 250404 224408 250410 224460
rect 268930 224408 268936 224460
rect 268988 224448 268994 224460
rect 283558 224448 283564 224460
rect 268988 224420 283564 224448
rect 268988 224408 268994 224420
rect 283558 224408 283564 224420
rect 283616 224408 283622 224460
rect 333698 224408 333704 224460
rect 333756 224448 333762 224460
rect 378042 224448 378048 224460
rect 333756 224420 378048 224448
rect 333756 224408 333762 224420
rect 378042 224408 378048 224420
rect 378100 224408 378106 224460
rect 400030 224408 400036 224460
rect 400088 224448 400094 224460
rect 543182 224448 543188 224460
rect 400088 224420 543188 224448
rect 400088 224408 400094 224420
rect 543182 224408 543188 224420
rect 543240 224408 543246 224460
rect 135990 224340 135996 224392
rect 136048 224380 136054 224392
rect 226794 224380 226800 224392
rect 136048 224352 226800 224380
rect 136048 224340 136054 224352
rect 226794 224340 226800 224352
rect 226852 224340 226858 224392
rect 246850 224340 246856 224392
rect 246908 224380 246914 224392
rect 273622 224380 273628 224392
rect 246908 224352 273628 224380
rect 246908 224340 246914 224352
rect 273622 224340 273628 224352
rect 273680 224340 273686 224392
rect 307754 224340 307760 224392
rect 307812 224380 307818 224392
rect 325694 224380 325700 224392
rect 307812 224352 325700 224380
rect 307812 224340 307818 224352
rect 325694 224340 325700 224352
rect 325752 224340 325758 224392
rect 339862 224340 339868 224392
rect 339920 224380 339926 224392
rect 386414 224380 386420 224392
rect 339920 224352 386420 224380
rect 339920 224340 339926 224352
rect 386414 224340 386420 224352
rect 386472 224340 386478 224392
rect 402238 224340 402244 224392
rect 402296 224380 402302 224392
rect 548518 224380 548524 224392
rect 402296 224352 548524 224380
rect 402296 224340 402302 224352
rect 548518 224340 548524 224352
rect 548576 224340 548582 224392
rect 101490 224272 101496 224324
rect 101548 224312 101554 224324
rect 136358 224312 136364 224324
rect 101548 224284 136364 224312
rect 101548 224272 101554 224284
rect 136358 224272 136364 224284
rect 136416 224272 136422 224324
rect 136542 224272 136548 224324
rect 136600 224312 136606 224324
rect 228634 224312 228640 224324
rect 136600 224284 228640 224312
rect 136600 224272 136606 224284
rect 228634 224272 228640 224284
rect 228692 224272 228698 224324
rect 232406 224272 232412 224324
rect 232464 224312 232470 224324
rect 243262 224312 243268 224324
rect 232464 224284 243268 224312
rect 232464 224272 232470 224284
rect 243262 224272 243268 224284
rect 243320 224272 243326 224324
rect 243630 224272 243636 224324
rect 243688 224312 243694 224324
rect 272242 224312 272248 224324
rect 243688 224284 272248 224312
rect 243688 224272 243694 224284
rect 272242 224272 272248 224284
rect 272300 224272 272306 224324
rect 309226 224272 309232 224324
rect 309284 224312 309290 224324
rect 328730 224312 328736 224324
rect 309284 224284 328736 224312
rect 309284 224272 309290 224284
rect 328730 224272 328736 224284
rect 328788 224272 328794 224324
rect 341426 224272 341432 224324
rect 341484 224312 341490 224324
rect 401870 224312 401876 224324
rect 341484 224284 401876 224312
rect 341484 224272 341490 224284
rect 401870 224272 401876 224284
rect 401928 224272 401934 224324
rect 405458 224272 405464 224324
rect 405516 224312 405522 224324
rect 556154 224312 556160 224324
rect 405516 224284 556160 224312
rect 405516 224272 405522 224284
rect 556154 224272 556160 224284
rect 556212 224272 556218 224324
rect 88150 224204 88156 224256
rect 88208 224244 88214 224256
rect 207566 224244 207572 224256
rect 88208 224216 207572 224244
rect 88208 224204 88214 224216
rect 207566 224204 207572 224216
rect 207624 224204 207630 224256
rect 239950 224204 239956 224256
rect 240008 224244 240014 224256
rect 271046 224244 271052 224256
rect 240008 224216 271052 224244
rect 240008 224204 240014 224216
rect 271046 224204 271052 224216
rect 271104 224204 271110 224256
rect 292574 224204 292580 224256
rect 292632 224244 292638 224256
rect 293494 224244 293500 224256
rect 292632 224216 293500 224244
rect 292632 224204 292638 224216
rect 293494 224204 293500 224216
rect 293552 224204 293558 224256
rect 311342 224204 311348 224256
rect 311400 224244 311406 224256
rect 331306 224244 331312 224256
rect 311400 224216 331312 224244
rect 311400 224204 311406 224216
rect 331306 224204 331312 224216
rect 331364 224204 331370 224256
rect 344094 224204 344100 224256
rect 344152 224244 344158 224256
rect 408586 224244 408592 224256
rect 344152 224216 408592 224244
rect 344152 224204 344158 224216
rect 408586 224204 408592 224216
rect 408644 224204 408650 224256
rect 408678 224204 408684 224256
rect 408736 224244 408742 224256
rect 563606 224244 563612 224256
rect 408736 224216 563612 224244
rect 408736 224204 408742 224216
rect 563606 224204 563612 224216
rect 563664 224204 563670 224256
rect 166258 224136 166264 224188
rect 166316 224176 166322 224188
rect 239674 224176 239680 224188
rect 166316 224148 239680 224176
rect 166316 224136 166322 224148
rect 239674 224136 239680 224148
rect 239732 224136 239738 224188
rect 342714 224136 342720 224188
rect 342772 224176 342778 224188
rect 405826 224176 405832 224188
rect 342772 224148 405832 224176
rect 342772 224136 342778 224148
rect 405826 224136 405832 224148
rect 405884 224136 405890 224188
rect 411254 224136 411260 224188
rect 411312 224176 411318 224188
rect 506474 224176 506480 224188
rect 411312 224148 506480 224176
rect 411312 224136 411318 224148
rect 506474 224136 506480 224148
rect 506532 224136 506538 224188
rect 169570 224068 169576 224120
rect 169628 224108 169634 224120
rect 241054 224108 241060 224120
rect 169628 224080 241060 224108
rect 169628 224068 169634 224080
rect 241054 224068 241060 224080
rect 241112 224068 241118 224120
rect 338390 224068 338396 224120
rect 338448 224108 338454 224120
rect 380710 224108 380716 224120
rect 338448 224080 380716 224108
rect 338448 224068 338454 224080
rect 380710 224068 380716 224080
rect 380768 224068 380774 224120
rect 393406 224068 393412 224120
rect 393464 224108 393470 224120
rect 472066 224108 472072 224120
rect 393464 224080 472072 224108
rect 393464 224068 393470 224080
rect 472066 224068 472072 224080
rect 472124 224068 472130 224120
rect 172974 224000 172980 224052
rect 173032 224040 173038 224052
rect 242526 224040 242532 224052
rect 173032 224012 242532 224040
rect 173032 224000 173038 224012
rect 242526 224000 242532 224012
rect 242584 224000 242590 224052
rect 349798 224000 349804 224052
rect 349856 224040 349862 224052
rect 422386 224040 422392 224052
rect 349856 224012 422392 224040
rect 349856 224000 349862 224012
rect 422386 224000 422392 224012
rect 422444 224000 422450 224052
rect 176470 223932 176476 223984
rect 176528 223972 176534 223984
rect 243906 223972 243912 223984
rect 176528 223944 243912 223972
rect 176528 223932 176534 223944
rect 243906 223932 243912 223944
rect 243964 223932 243970 223984
rect 347314 223932 347320 223984
rect 347372 223972 347378 223984
rect 417050 223972 417056 223984
rect 347372 223944 417056 223972
rect 347372 223932 347378 223944
rect 417050 223932 417056 223944
rect 417108 223932 417114 223984
rect 179690 223864 179696 223916
rect 179748 223904 179754 223916
rect 245378 223904 245384 223916
rect 179748 223876 245384 223904
rect 179748 223864 179754 223876
rect 245378 223864 245384 223876
rect 245436 223864 245442 223916
rect 348418 223864 348424 223916
rect 348476 223904 348482 223916
rect 418706 223904 418712 223916
rect 348476 223876 418712 223904
rect 348476 223864 348482 223876
rect 418706 223864 418712 223876
rect 418764 223864 418770 223916
rect 183186 223796 183192 223848
rect 183244 223836 183250 223848
rect 246758 223836 246764 223848
rect 183244 223808 246764 223836
rect 183244 223796 183250 223808
rect 246758 223796 246764 223808
rect 246816 223796 246822 223848
rect 346946 223796 346952 223848
rect 347004 223836 347010 223848
rect 415486 223836 415492 223848
rect 347004 223808 415492 223836
rect 347004 223796 347010 223808
rect 415486 223796 415492 223808
rect 415544 223796 415550 223848
rect 186222 223728 186228 223780
rect 186280 223768 186286 223780
rect 248230 223768 248236 223780
rect 186280 223740 248236 223768
rect 186280 223728 186286 223740
rect 248230 223728 248236 223740
rect 248288 223728 248294 223780
rect 354858 223728 354864 223780
rect 354916 223768 354922 223780
rect 411990 223768 411996 223780
rect 354916 223740 411996 223768
rect 354916 223728 354922 223740
rect 411990 223728 411996 223740
rect 412048 223728 412054 223780
rect 337286 223660 337292 223712
rect 337344 223700 337350 223712
rect 378778 223700 378784 223712
rect 337344 223672 378784 223700
rect 337344 223660 337350 223672
rect 378778 223660 378784 223672
rect 378836 223660 378842 223712
rect 409874 223660 409880 223712
rect 409932 223700 409938 223712
rect 465166 223700 465172 223712
rect 409932 223672 465172 223700
rect 409932 223660 409938 223672
rect 465166 223660 465172 223672
rect 465224 223660 465230 223712
rect 62022 223632 62028 223644
rect 59372 223604 62028 223632
rect 56594 223524 56600 223576
rect 56652 223564 56658 223576
rect 59372 223564 59400 223604
rect 62022 223592 62028 223604
rect 62080 223592 62086 223644
rect 56652 223536 59400 223564
rect 56652 223524 56658 223536
rect 125870 223524 125876 223576
rect 125928 223564 125934 223576
rect 222562 223564 222568 223576
rect 125928 223536 222568 223564
rect 125928 223524 125934 223536
rect 222562 223524 222568 223536
rect 222620 223524 222626 223576
rect 359458 223524 359464 223576
rect 359516 223564 359522 223576
rect 448606 223564 448612 223576
rect 359516 223536 448612 223564
rect 359516 223524 359522 223536
rect 448606 223524 448612 223536
rect 448664 223524 448670 223576
rect 115750 223456 115756 223508
rect 115808 223496 115814 223508
rect 115808 223468 210556 223496
rect 115808 223456 115814 223468
rect 108850 223388 108856 223440
rect 108908 223428 108914 223440
rect 108908 223400 210464 223428
rect 108908 223388 108914 223400
rect 105722 223320 105728 223372
rect 105780 223360 105786 223372
rect 209590 223360 209596 223372
rect 105780 223332 209596 223360
rect 105780 223320 105786 223332
rect 209590 223320 209596 223332
rect 209648 223320 209654 223372
rect 209700 223332 210004 223360
rect 101950 223252 101956 223304
rect 102008 223292 102014 223304
rect 209700 223292 209728 223332
rect 102008 223264 209728 223292
rect 102008 223252 102014 223264
rect 95602 223184 95608 223236
rect 95660 223224 95666 223236
rect 209682 223224 209688 223236
rect 95660 223196 209688 223224
rect 95660 223184 95666 223196
rect 209682 223184 209688 223196
rect 209740 223184 209746 223236
rect 209976 223224 210004 223332
rect 210436 223292 210464 223400
rect 210528 223360 210556 223468
rect 213914 223456 213920 223508
rect 213972 223496 213978 223508
rect 221826 223496 221832 223508
rect 213972 223468 221832 223496
rect 213972 223456 213978 223468
rect 221826 223456 221832 223468
rect 221884 223456 221890 223508
rect 361114 223456 361120 223508
rect 361172 223496 361178 223508
rect 451458 223496 451464 223508
rect 361172 223468 451464 223496
rect 361172 223456 361178 223468
rect 451458 223456 451464 223468
rect 451516 223456 451522 223508
rect 352282 223388 352288 223440
rect 352340 223428 352346 223440
rect 431310 223428 431316 223440
rect 352340 223400 431316 223428
rect 352340 223388 352346 223400
rect 431310 223388 431316 223400
rect 431368 223388 431374 223440
rect 431954 223388 431960 223440
rect 432012 223428 432018 223440
rect 525058 223428 525064 223440
rect 432012 223400 525064 223428
rect 432012 223388 432018 223400
rect 525058 223388 525064 223400
rect 525116 223388 525122 223440
rect 218238 223360 218244 223372
rect 210528 223332 218244 223360
rect 218238 223320 218244 223332
rect 218296 223320 218302 223372
rect 389082 223320 389088 223372
rect 389140 223360 389146 223372
rect 395706 223360 395712 223372
rect 389140 223332 395712 223360
rect 389140 223320 389146 223332
rect 395706 223320 395712 223332
rect 395764 223320 395770 223372
rect 523126 223360 523132 223372
rect 395908 223332 523132 223360
rect 215386 223292 215392 223304
rect 210436 223264 215392 223292
rect 215386 223252 215392 223264
rect 215444 223252 215450 223304
rect 212534 223224 212540 223236
rect 209976 223196 212540 223224
rect 212534 223184 212540 223196
rect 212592 223184 212598 223236
rect 319254 223184 319260 223236
rect 319312 223224 319318 223236
rect 350626 223224 350632 223236
rect 319312 223196 350632 223224
rect 319312 223184 319318 223196
rect 350626 223184 350632 223196
rect 350684 223184 350690 223236
rect 391566 223184 391572 223236
rect 391624 223224 391630 223236
rect 391624 223196 393314 223224
rect 391624 223184 391630 223196
rect 82170 223116 82176 223168
rect 82228 223156 82234 223168
rect 203978 223156 203984 223168
rect 82228 223128 203984 223156
rect 82228 223116 82234 223128
rect 203978 223116 203984 223128
rect 204036 223116 204042 223168
rect 209590 223116 209596 223168
rect 209648 223156 209654 223168
rect 214006 223156 214012 223168
rect 209648 223128 214012 223156
rect 209648 223116 209654 223128
rect 214006 223116 214012 223128
rect 214064 223116 214070 223168
rect 250346 223116 250352 223168
rect 250404 223156 250410 223168
rect 275094 223156 275100 223168
rect 250404 223128 275100 223156
rect 250404 223116 250410 223128
rect 275094 223116 275100 223128
rect 275152 223116 275158 223168
rect 311618 223116 311624 223168
rect 311676 223156 311682 223168
rect 318886 223156 318892 223168
rect 311676 223128 318892 223156
rect 311676 223116 311682 223128
rect 318886 223116 318892 223128
rect 318944 223116 318950 223168
rect 330938 223116 330944 223168
rect 330996 223156 331002 223168
rect 367002 223156 367008 223168
rect 330996 223128 367008 223156
rect 330996 223116 331002 223128
rect 367002 223116 367008 223128
rect 367060 223116 367066 223168
rect 385862 223116 385868 223168
rect 385920 223156 385926 223168
rect 387794 223156 387800 223168
rect 385920 223128 387800 223156
rect 385920 223116 385926 223128
rect 387794 223116 387800 223128
rect 387852 223116 387858 223168
rect 393286 223156 393314 223196
rect 395908 223156 395936 223332
rect 523126 223320 523132 223332
rect 523184 223320 523190 223372
rect 398282 223252 398288 223304
rect 398340 223292 398346 223304
rect 530578 223292 530584 223304
rect 398340 223264 530584 223292
rect 398340 223252 398346 223264
rect 530578 223252 530584 223264
rect 530636 223252 530642 223304
rect 395982 223184 395988 223236
rect 396040 223224 396046 223236
rect 533062 223224 533068 223236
rect 396040 223196 533068 223224
rect 396040 223184 396046 223196
rect 533062 223184 533068 223196
rect 533120 223184 533126 223236
rect 393286 223128 395936 223156
rect 397914 223116 397920 223168
rect 397972 223156 397978 223168
rect 538306 223156 538312 223168
rect 397972 223128 538312 223156
rect 397972 223116 397978 223128
rect 538306 223116 538312 223128
rect 538364 223116 538370 223168
rect 75362 223048 75368 223100
rect 75420 223088 75426 223100
rect 201126 223088 201132 223100
rect 75420 223060 201132 223088
rect 75420 223048 75426 223060
rect 201126 223048 201132 223060
rect 201184 223048 201190 223100
rect 204898 223048 204904 223100
rect 204956 223088 204962 223100
rect 256418 223088 256424 223100
rect 204956 223060 256424 223088
rect 204956 223048 204962 223060
rect 256418 223048 256424 223060
rect 256476 223048 256482 223100
rect 314194 223048 314200 223100
rect 314252 223088 314258 223100
rect 338114 223088 338120 223100
rect 314252 223060 338120 223088
rect 314252 223048 314258 223060
rect 338114 223048 338120 223060
rect 338172 223048 338178 223100
rect 348142 223048 348148 223100
rect 348200 223088 348206 223100
rect 421190 223088 421196 223100
rect 348200 223060 421196 223088
rect 348200 223048 348206 223060
rect 421190 223048 421196 223060
rect 421248 223048 421254 223100
rect 421282 223048 421288 223100
rect 421340 223088 421346 223100
rect 569310 223088 569316 223100
rect 421340 223060 569316 223088
rect 421340 223048 421346 223060
rect 569310 223048 569316 223060
rect 569368 223048 569374 223100
rect 69014 222980 69020 223032
rect 69072 223020 69078 223032
rect 69072 222992 194180 223020
rect 69072 222980 69078 222992
rect 68738 222912 68744 222964
rect 68796 222952 68802 222964
rect 193950 222952 193956 222964
rect 68796 222924 193956 222952
rect 68796 222912 68802 222924
rect 193950 222912 193956 222924
rect 194008 222912 194014 222964
rect 194152 222952 194180 222992
rect 198182 222980 198188 223032
rect 198240 223020 198246 223032
rect 253566 223020 253572 223032
rect 198240 222992 253572 223020
rect 198240 222980 198246 222992
rect 253566 222980 253572 222992
rect 253624 222980 253630 223032
rect 306374 222980 306380 223032
rect 306432 223020 306438 223032
rect 321922 223020 321928 223032
rect 306432 222992 321928 223020
rect 306432 222980 306438 222992
rect 321922 222980 321928 222992
rect 321980 222980 321986 223032
rect 326614 222980 326620 223032
rect 326672 223020 326678 223032
rect 371234 223020 371240 223032
rect 326672 222992 371240 223020
rect 326672 222980 326678 222992
rect 371234 222980 371240 222992
rect 371292 222980 371298 223032
rect 379790 222980 379796 223032
rect 379848 223020 379854 223032
rect 389174 223020 389180 223032
rect 379848 222992 389180 223020
rect 379848 222980 379854 222992
rect 389174 222980 389180 222992
rect 389232 222980 389238 223032
rect 394786 222980 394792 223032
rect 394844 223020 394850 223032
rect 398282 223020 398288 223032
rect 394844 222992 398288 223020
rect 394844 222980 394850 222992
rect 398282 222980 398288 222992
rect 398340 222980 398346 223032
rect 404630 222980 404636 223032
rect 404688 223020 404694 223032
rect 553670 223020 553676 223032
rect 404688 222992 553676 223020
rect 404688 222980 404694 222992
rect 553670 222980 553676 222992
rect 553728 222980 553734 223032
rect 198366 222952 198372 222964
rect 194152 222924 198372 222952
rect 198366 222912 198372 222924
rect 198424 222912 198430 222964
rect 199930 222912 199936 222964
rect 199988 222952 199994 222964
rect 253934 222952 253940 222964
rect 199988 222924 253940 222952
rect 199988 222912 199994 222924
rect 253934 222912 253940 222924
rect 253992 222912 253998 222964
rect 265526 222912 265532 222964
rect 265584 222952 265590 222964
rect 282086 222952 282092 222964
rect 265584 222924 282092 222952
rect 265584 222912 265590 222924
rect 282086 222912 282092 222924
rect 282144 222912 282150 222964
rect 317046 222912 317052 222964
rect 317104 222952 317110 222964
rect 345014 222952 345020 222964
rect 317104 222924 345020 222952
rect 317104 222912 317110 222924
rect 345014 222912 345020 222924
rect 345072 222912 345078 222964
rect 346670 222912 346676 222964
rect 346728 222952 346734 222964
rect 415302 222952 415308 222964
rect 346728 222924 415308 222952
rect 346728 222912 346734 222924
rect 415302 222912 415308 222924
rect 415360 222912 415366 222964
rect 416222 222912 416228 222964
rect 416280 222952 416286 222964
rect 567194 222952 567200 222964
rect 416280 222924 567200 222952
rect 416280 222912 416286 222924
rect 567194 222912 567200 222924
rect 567252 222912 567258 222964
rect 65334 222844 65340 222896
rect 65392 222884 65398 222896
rect 196894 222884 196900 222896
rect 65392 222856 196900 222884
rect 65392 222844 65398 222856
rect 196894 222844 196900 222856
rect 196952 222844 196958 222896
rect 200758 222844 200764 222896
rect 200816 222884 200822 222896
rect 255682 222884 255688 222896
rect 200816 222856 255688 222884
rect 200816 222844 200822 222856
rect 255682 222844 255688 222856
rect 255740 222844 255746 222896
rect 262122 222844 262128 222896
rect 262180 222884 262186 222896
rect 280706 222884 280712 222896
rect 262180 222856 280712 222884
rect 262180 222844 262186 222856
rect 280706 222844 280712 222856
rect 280764 222844 280770 222896
rect 308490 222844 308496 222896
rect 308548 222884 308554 222896
rect 324498 222884 324504 222896
rect 308548 222856 324504 222884
rect 308548 222844 308554 222856
rect 324498 222844 324504 222856
rect 324556 222844 324562 222896
rect 337654 222844 337660 222896
rect 337712 222884 337718 222896
rect 390646 222884 390652 222896
rect 337712 222856 390652 222884
rect 337712 222844 337718 222856
rect 390646 222844 390652 222856
rect 390704 222844 390710 222896
rect 407574 222844 407580 222896
rect 407632 222884 407638 222896
rect 560938 222884 560944 222896
rect 407632 222856 560944 222884
rect 407632 222844 407638 222856
rect 560938 222844 560944 222856
rect 560996 222844 561002 222896
rect 132310 222776 132316 222828
rect 132368 222816 132374 222828
rect 225414 222816 225420 222828
rect 132368 222788 225420 222816
rect 132368 222776 132374 222788
rect 225414 222776 225420 222788
rect 225472 222776 225478 222828
rect 357986 222776 357992 222828
rect 358044 222816 358050 222828
rect 444742 222816 444748 222828
rect 358044 222788 444748 222816
rect 358044 222776 358050 222788
rect 444742 222776 444748 222788
rect 444800 222776 444806 222828
rect 177850 222708 177856 222760
rect 177908 222748 177914 222760
rect 245010 222748 245016 222760
rect 177908 222720 245016 222748
rect 177908 222708 177914 222720
rect 245010 222708 245016 222720
rect 245068 222708 245074 222760
rect 356606 222708 356612 222760
rect 356664 222748 356670 222760
rect 441706 222748 441712 222760
rect 356664 222720 441712 222748
rect 356664 222708 356670 222720
rect 441706 222708 441712 222720
rect 441764 222708 441770 222760
rect 162026 222640 162032 222692
rect 162084 222680 162090 222692
rect 180794 222680 180800 222692
rect 162084 222652 180800 222680
rect 162084 222640 162090 222652
rect 180794 222640 180800 222652
rect 180852 222640 180858 222692
rect 181346 222640 181352 222692
rect 181404 222680 181410 222692
rect 246482 222680 246488 222692
rect 181404 222652 246488 222680
rect 181404 222640 181410 222652
rect 246482 222640 246488 222652
rect 246540 222640 246546 222692
rect 355134 222640 355140 222692
rect 355192 222680 355198 222692
rect 438026 222680 438032 222692
rect 355192 222652 438032 222680
rect 355192 222640 355198 222652
rect 438026 222640 438032 222652
rect 438084 222640 438090 222692
rect 187326 222572 187332 222624
rect 187384 222612 187390 222624
rect 249978 222612 249984 222624
rect 187384 222584 249984 222612
rect 187384 222572 187390 222584
rect 249978 222572 249984 222584
rect 250036 222572 250042 222624
rect 353754 222572 353760 222624
rect 353812 222612 353818 222624
rect 434806 222612 434812 222624
rect 353812 222584 434812 222612
rect 353812 222572 353818 222584
rect 434806 222572 434812 222584
rect 434864 222572 434870 222624
rect 184750 222504 184756 222556
rect 184808 222544 184814 222556
rect 247862 222544 247868 222556
rect 184808 222516 247868 222544
rect 184808 222504 184814 222516
rect 247862 222504 247868 222516
rect 247920 222504 247926 222556
rect 352650 222504 352656 222556
rect 352708 222544 352714 222556
rect 429286 222544 429292 222556
rect 352708 222516 429292 222544
rect 352708 222504 352714 222516
rect 429286 222504 429292 222516
rect 429344 222504 429350 222556
rect 665818 222504 665824 222556
rect 665876 222544 665882 222556
rect 675938 222544 675944 222556
rect 665876 222516 675944 222544
rect 665876 222504 665882 222516
rect 675938 222504 675944 222516
rect 675996 222504 676002 222556
rect 188154 222436 188160 222488
rect 188212 222476 188218 222488
rect 249334 222476 249340 222488
rect 188212 222448 249340 222476
rect 188212 222436 188218 222448
rect 249334 222436 249340 222448
rect 249392 222436 249398 222488
rect 351178 222436 351184 222488
rect 351236 222476 351242 222488
rect 427906 222476 427912 222488
rect 351236 222448 427912 222476
rect 351236 222436 351242 222448
rect 427906 222436 427912 222448
rect 427964 222436 427970 222488
rect 428642 222436 428648 222488
rect 428700 222476 428706 222488
rect 488534 222476 488540 222488
rect 428700 222448 488540 222476
rect 428700 222436 428706 222448
rect 488534 222436 488540 222448
rect 488592 222436 488598 222488
rect 191558 222368 191564 222420
rect 191616 222408 191622 222420
rect 250714 222408 250720 222420
rect 191616 222380 250720 222408
rect 191616 222368 191622 222380
rect 250714 222368 250720 222380
rect 250772 222368 250778 222420
rect 349430 222368 349436 222420
rect 349488 222408 349494 222420
rect 425054 222408 425060 222420
rect 349488 222380 425060 222408
rect 349488 222368 349494 222380
rect 425054 222368 425060 222380
rect 425112 222368 425118 222420
rect 664438 222368 664444 222420
rect 664496 222408 664502 222420
rect 676030 222408 676036 222420
rect 664496 222380 676036 222408
rect 664496 222368 664502 222380
rect 676030 222368 676036 222380
rect 676088 222368 676094 222420
rect 196526 222300 196532 222352
rect 196584 222340 196590 222352
rect 252278 222340 252284 222352
rect 196584 222312 252284 222340
rect 196584 222300 196590 222312
rect 252278 222300 252284 222312
rect 252336 222300 252342 222352
rect 193950 222232 193956 222284
rect 194008 222272 194014 222284
rect 198274 222272 198280 222284
rect 194008 222244 198280 222272
rect 194008 222232 194014 222244
rect 198274 222232 198280 222244
rect 198332 222232 198338 222284
rect 673914 222232 673920 222284
rect 673972 222272 673978 222284
rect 676030 222272 676036 222284
rect 673972 222244 676036 222272
rect 673972 222232 673978 222244
rect 676030 222232 676036 222244
rect 676088 222232 676094 222284
rect 660390 222164 660396 222216
rect 660448 222204 660454 222216
rect 675846 222204 675852 222216
rect 660448 222176 675852 222204
rect 660448 222164 660454 222176
rect 675846 222164 675852 222176
rect 675904 222164 675910 222216
rect 122466 222096 122472 222148
rect 122524 222136 122530 222148
rect 220998 222136 221004 222148
rect 122524 222108 221004 222136
rect 122524 222096 122530 222108
rect 220998 222096 221004 222108
rect 221056 222096 221062 222148
rect 228450 222096 228456 222148
rect 228508 222136 228514 222148
rect 266446 222136 266452 222148
rect 228508 222108 266452 222136
rect 228508 222096 228514 222108
rect 266446 222096 266452 222108
rect 266504 222096 266510 222148
rect 311158 222096 311164 222148
rect 311216 222136 311222 222148
rect 311986 222136 311992 222148
rect 311216 222108 311992 222136
rect 311216 222096 311222 222108
rect 311986 222096 311992 222108
rect 312044 222096 312050 222148
rect 312538 222096 312544 222148
rect 312596 222136 312602 222148
rect 315298 222136 315304 222148
rect 312596 222108 315304 222136
rect 312596 222096 312602 222108
rect 315298 222096 315304 222108
rect 315356 222096 315362 222148
rect 318702 222096 318708 222148
rect 318760 222136 318766 222148
rect 349154 222136 349160 222148
rect 318760 222108 349160 222136
rect 318760 222096 318766 222108
rect 349154 222096 349160 222108
rect 349212 222096 349218 222148
rect 362678 222096 362684 222148
rect 362736 222136 362742 222148
rect 453206 222136 453212 222148
rect 362736 222108 453212 222136
rect 362736 222096 362742 222108
rect 453206 222096 453212 222108
rect 453264 222096 453270 222148
rect 453298 222096 453304 222148
rect 453356 222136 453362 222148
rect 545206 222136 545212 222148
rect 453356 222108 545212 222136
rect 453356 222096 453362 222108
rect 545206 222096 545212 222108
rect 545264 222096 545270 222148
rect 574738 222096 574744 222148
rect 574796 222136 574802 222148
rect 575474 222136 575480 222148
rect 574796 222108 575480 222136
rect 574796 222096 574802 222108
rect 575474 222096 575480 222108
rect 575532 222096 575538 222148
rect 119154 222028 119160 222080
rect 119212 222068 119218 222080
rect 219618 222068 219624 222080
rect 119212 222040 219624 222068
rect 119212 222028 119218 222040
rect 219618 222028 219624 222040
rect 219676 222028 219682 222080
rect 226794 222028 226800 222080
rect 226852 222068 226858 222080
rect 265250 222068 265256 222080
rect 226852 222040 265256 222068
rect 226852 222028 226858 222040
rect 265250 222028 265256 222040
rect 265308 222028 265314 222080
rect 321370 222028 321376 222080
rect 321428 222068 321434 222080
rect 356054 222068 356060 222080
rect 321428 222040 356060 222068
rect 321428 222028 321434 222040
rect 356054 222028 356060 222040
rect 356112 222028 356118 222080
rect 364150 222028 364156 222080
rect 364208 222068 364214 222080
rect 456794 222068 456800 222080
rect 364208 222040 456800 222068
rect 364208 222028 364214 222040
rect 456794 222028 456800 222040
rect 456852 222028 456858 222080
rect 100754 221960 100760 222012
rect 100812 222000 100818 222012
rect 204346 222000 204352 222012
rect 100812 221972 204352 222000
rect 100812 221960 100818 221972
rect 204346 221960 204352 221972
rect 204404 221960 204410 222012
rect 223482 221960 223488 222012
rect 223540 222000 223546 222012
rect 263686 222000 263692 222012
rect 223540 221972 263692 222000
rect 223540 221960 223546 221972
rect 263686 221960 263692 221972
rect 263744 221960 263750 222012
rect 321186 221960 321192 222012
rect 321244 222000 321250 222012
rect 357526 222000 357532 222012
rect 321244 221972 357532 222000
rect 321244 221960 321250 221972
rect 357526 221960 357532 221972
rect 357584 221960 357590 222012
rect 363966 221960 363972 222012
rect 364024 222000 364030 222012
rect 458358 222000 458364 222012
rect 364024 221972 458364 222000
rect 364024 221960 364030 221972
rect 458358 221960 458364 221972
rect 458416 221960 458422 222012
rect 112438 221892 112444 221944
rect 112496 221932 112502 221944
rect 216858 221932 216864 221944
rect 112496 221904 216864 221932
rect 112496 221892 112502 221904
rect 216858 221892 216864 221904
rect 216916 221892 216922 221944
rect 224862 221892 224868 221944
rect 224920 221932 224926 221944
rect 265158 221932 265164 221944
rect 224920 221904 265164 221932
rect 224920 221892 224926 221904
rect 265158 221892 265164 221904
rect 265216 221892 265222 221944
rect 322290 221892 322296 221944
rect 322348 221932 322354 221944
rect 359090 221932 359096 221944
rect 322348 221904 359096 221932
rect 322348 221892 322354 221904
rect 359090 221892 359096 221904
rect 359148 221892 359154 221944
rect 365070 221892 365076 221944
rect 365128 221932 365134 221944
rect 460014 221932 460020 221944
rect 365128 221904 460020 221932
rect 365128 221892 365134 221904
rect 460014 221892 460020 221904
rect 460072 221892 460078 221944
rect 88886 221824 88892 221876
rect 88944 221864 88950 221876
rect 88944 221836 205312 221864
rect 88944 221824 88950 221836
rect 85482 221756 85488 221808
rect 85540 221796 85546 221808
rect 205174 221796 205180 221808
rect 85540 221768 205180 221796
rect 85540 221756 85546 221768
rect 205174 221756 205180 221768
rect 205232 221756 205238 221808
rect 83826 221688 83832 221740
rect 83884 221728 83890 221740
rect 204806 221728 204812 221740
rect 83884 221700 204812 221728
rect 83884 221688 83890 221700
rect 204806 221688 204812 221700
rect 204864 221688 204870 221740
rect 205284 221728 205312 221836
rect 205542 221824 205548 221876
rect 205600 221864 205606 221876
rect 206738 221864 206744 221876
rect 205600 221836 206744 221864
rect 205600 221824 205606 221836
rect 206738 221824 206744 221836
rect 206796 221824 206802 221876
rect 220078 221824 220084 221876
rect 220136 221864 220142 221876
rect 262306 221864 262312 221876
rect 220136 221836 262312 221864
rect 220136 221824 220142 221836
rect 262306 221824 262312 221836
rect 262364 221824 262370 221876
rect 322658 221824 322664 221876
rect 322716 221864 322722 221876
rect 360746 221864 360752 221876
rect 322716 221836 360752 221864
rect 322716 221824 322722 221836
rect 360746 221824 360752 221836
rect 360804 221824 360810 221876
rect 366450 221824 366456 221876
rect 366508 221864 366514 221876
rect 463694 221864 463700 221876
rect 366508 221836 463700 221864
rect 366508 221824 366514 221836
rect 463694 221824 463700 221836
rect 463752 221824 463758 221876
rect 674650 221824 674656 221876
rect 674708 221864 674714 221876
rect 676030 221864 676036 221876
rect 674708 221836 676036 221864
rect 674708 221824 674714 221836
rect 676030 221824 676036 221836
rect 676088 221824 676094 221876
rect 206922 221756 206928 221808
rect 206980 221796 206986 221808
rect 217318 221796 217324 221808
rect 206980 221768 217324 221796
rect 206980 221756 206986 221768
rect 217318 221756 217324 221768
rect 217376 221756 217382 221808
rect 218422 221756 218428 221808
rect 218480 221796 218486 221808
rect 261846 221796 261852 221808
rect 218480 221768 261852 221796
rect 218480 221756 218486 221768
rect 261846 221756 261852 221768
rect 261904 221756 261910 221808
rect 324222 221756 324228 221808
rect 324280 221796 324286 221808
rect 362402 221796 362408 221808
rect 324280 221768 362408 221796
rect 324280 221756 324286 221768
rect 362402 221756 362408 221768
rect 362460 221756 362466 221808
rect 367922 221756 367928 221808
rect 367980 221796 367986 221808
rect 466730 221796 466736 221808
rect 367980 221768 466736 221796
rect 367980 221756 367986 221768
rect 466730 221756 466736 221768
rect 466788 221756 466794 221808
rect 467098 221756 467104 221808
rect 467156 221796 467162 221808
rect 557810 221796 557816 221808
rect 467156 221768 557816 221796
rect 467156 221756 467162 221768
rect 557810 221756 557816 221768
rect 557868 221756 557874 221808
rect 206646 221728 206652 221740
rect 205284 221700 206652 221728
rect 206646 221688 206652 221700
rect 206704 221688 206710 221740
rect 208210 221688 208216 221740
rect 208268 221728 208274 221740
rect 220170 221728 220176 221740
rect 208268 221700 220176 221728
rect 208268 221688 208274 221700
rect 220170 221688 220176 221700
rect 220228 221688 220234 221740
rect 221734 221688 221740 221740
rect 221792 221728 221798 221740
rect 263778 221728 263784 221740
rect 221792 221700 263784 221728
rect 221792 221688 221798 221700
rect 263778 221688 263784 221700
rect 263836 221688 263842 221740
rect 325510 221688 325516 221740
rect 325568 221728 325574 221740
rect 365806 221728 365812 221740
rect 325568 221700 365812 221728
rect 325568 221688 325574 221700
rect 365806 221688 365812 221700
rect 365864 221688 365870 221740
rect 369302 221688 369308 221740
rect 369360 221728 369366 221740
rect 470134 221728 470140 221740
rect 369360 221700 470140 221728
rect 369360 221688 369366 221700
rect 470134 221688 470140 221700
rect 470192 221688 470198 221740
rect 80422 221620 80428 221672
rect 80480 221660 80486 221672
rect 203426 221660 203432 221672
rect 80480 221632 203432 221660
rect 80480 221620 80486 221632
rect 203426 221620 203432 221632
rect 203484 221620 203490 221672
rect 204162 221620 204168 221672
rect 204220 221660 204226 221672
rect 214466 221660 214472 221672
rect 204220 221632 214472 221660
rect 204220 221620 204226 221632
rect 214466 221620 214472 221632
rect 214524 221620 214530 221672
rect 216582 221620 216588 221672
rect 216640 221660 216646 221672
rect 261018 221660 261024 221672
rect 216640 221632 261024 221660
rect 216640 221620 216646 221632
rect 261018 221620 261024 221632
rect 261076 221620 261082 221672
rect 326522 221620 326528 221672
rect 326580 221660 326586 221672
rect 369118 221660 369124 221672
rect 326580 221632 369124 221660
rect 326580 221620 326586 221632
rect 369118 221620 369124 221632
rect 369176 221620 369182 221672
rect 370774 221620 370780 221672
rect 370832 221660 370838 221672
rect 473538 221660 473544 221672
rect 370832 221632 473544 221660
rect 370832 221620 370838 221632
rect 473538 221620 473544 221632
rect 473596 221620 473602 221672
rect 77018 221552 77024 221604
rect 77076 221592 77082 221604
rect 201954 221592 201960 221604
rect 77076 221564 201960 221592
rect 77076 221552 77082 221564
rect 201954 221552 201960 221564
rect 202012 221552 202018 221604
rect 202414 221552 202420 221604
rect 202472 221592 202478 221604
rect 210142 221592 210148 221604
rect 202472 221564 210148 221592
rect 202472 221552 202478 221564
rect 210142 221552 210148 221564
rect 210200 221552 210206 221604
rect 213362 221552 213368 221604
rect 213420 221592 213426 221604
rect 259638 221592 259644 221604
rect 213420 221564 259644 221592
rect 213420 221552 213426 221564
rect 259638 221552 259644 221564
rect 259696 221552 259702 221604
rect 325418 221552 325424 221604
rect 325476 221592 325482 221604
rect 367462 221592 367468 221604
rect 325476 221564 367468 221592
rect 325476 221552 325482 221564
rect 367462 221552 367468 221564
rect 367520 221552 367526 221604
rect 400122 221552 400128 221604
rect 400180 221592 400186 221604
rect 541066 221592 541072 221604
rect 400180 221564 541072 221592
rect 400180 221552 400186 221564
rect 541066 221552 541072 221564
rect 541124 221552 541130 221604
rect 547138 221552 547144 221604
rect 547196 221592 547202 221604
rect 561766 221592 561772 221604
rect 547196 221564 561772 221592
rect 547196 221552 547202 221564
rect 561766 221552 561772 221564
rect 561824 221552 561830 221604
rect 63402 221484 63408 221536
rect 63460 221524 63466 221536
rect 196250 221524 196256 221536
rect 63460 221496 196256 221524
rect 63460 221484 63466 221496
rect 196250 221484 196256 221496
rect 196308 221484 196314 221536
rect 197262 221484 197268 221536
rect 197320 221524 197326 221536
rect 244918 221524 244924 221536
rect 197320 221496 244924 221524
rect 197320 221484 197326 221496
rect 244918 221484 244924 221496
rect 244976 221484 244982 221536
rect 245286 221484 245292 221536
rect 245344 221524 245350 221536
rect 273438 221524 273444 221536
rect 245344 221496 273444 221524
rect 245344 221484 245350 221496
rect 273438 221484 273444 221496
rect 273496 221484 273502 221536
rect 275554 221484 275560 221536
rect 275612 221524 275618 221536
rect 286134 221524 286140 221536
rect 275612 221496 286140 221524
rect 275612 221484 275618 221496
rect 286134 221484 286140 221496
rect 286192 221484 286198 221536
rect 319438 221484 319444 221536
rect 319496 221524 319502 221536
rect 352374 221524 352380 221536
rect 319496 221496 352380 221524
rect 319496 221484 319502 221496
rect 352374 221484 352380 221496
rect 352432 221484 352438 221536
rect 352558 221484 352564 221536
rect 352616 221524 352622 221536
rect 397730 221524 397736 221536
rect 352616 221496 397736 221524
rect 352616 221484 352622 221496
rect 397730 221484 397736 221496
rect 397788 221484 397794 221536
rect 404170 221484 404176 221536
rect 404228 221524 404234 221536
rect 550818 221524 550824 221536
rect 404228 221496 550824 221524
rect 404228 221484 404234 221496
rect 550818 221484 550824 221496
rect 550876 221484 550882 221536
rect 551278 221484 551284 221536
rect 551336 221524 551342 221536
rect 565446 221524 565452 221536
rect 551336 221496 565452 221524
rect 551336 221484 551342 221496
rect 565446 221484 565452 221496
rect 565504 221484 565510 221536
rect 674006 221484 674012 221536
rect 674064 221524 674070 221536
rect 676030 221524 676036 221536
rect 674064 221496 676036 221524
rect 674064 221484 674070 221496
rect 676030 221484 676036 221496
rect 676088 221484 676094 221536
rect 28718 221416 28724 221468
rect 28776 221456 28782 221468
rect 43714 221456 43720 221468
rect 28776 221428 43720 221456
rect 28776 221416 28782 221428
rect 43714 221416 43720 221428
rect 43772 221416 43778 221468
rect 60274 221416 60280 221468
rect 60332 221456 60338 221468
rect 194870 221456 194876 221468
rect 60332 221428 194876 221456
rect 60332 221416 60338 221428
rect 194870 221416 194876 221428
rect 194928 221416 194934 221468
rect 209682 221416 209688 221468
rect 209740 221456 209746 221468
rect 258258 221456 258264 221468
rect 209740 221428 258264 221456
rect 209740 221416 209746 221428
rect 258258 221416 258264 221428
rect 258316 221416 258322 221468
rect 272242 221416 272248 221468
rect 272300 221456 272306 221468
rect 284662 221456 284668 221468
rect 272300 221428 284668 221456
rect 272300 221416 272306 221428
rect 284662 221416 284668 221428
rect 284720 221416 284726 221468
rect 301222 221416 301228 221468
rect 301280 221456 301286 221468
rect 310514 221456 310520 221468
rect 301280 221428 310520 221456
rect 301280 221416 301286 221428
rect 310514 221416 310520 221428
rect 310572 221416 310578 221468
rect 319806 221416 319812 221468
rect 319864 221456 319870 221468
rect 354030 221456 354036 221468
rect 319864 221428 354036 221456
rect 319864 221416 319870 221428
rect 354030 221416 354036 221428
rect 354088 221416 354094 221468
rect 401134 221456 401140 221468
rect 354646 221428 401140 221456
rect 129274 221348 129280 221400
rect 129332 221388 129338 221400
rect 223758 221388 223764 221400
rect 129332 221360 223764 221388
rect 129332 221348 129338 221360
rect 223758 221348 223764 221360
rect 223816 221348 223822 221400
rect 231670 221348 231676 221400
rect 231728 221388 231734 221400
rect 267826 221388 267832 221400
rect 231728 221360 267832 221388
rect 231728 221348 231734 221360
rect 267826 221348 267832 221360
rect 267884 221348 267890 221400
rect 317322 221348 317328 221400
rect 317380 221388 317386 221400
rect 345566 221388 345572 221400
rect 317380 221360 345572 221388
rect 317380 221348 317386 221360
rect 345566 221348 345572 221360
rect 345624 221348 345630 221400
rect 151078 221280 151084 221332
rect 151136 221320 151142 221332
rect 233418 221320 233424 221332
rect 151136 221292 233424 221320
rect 151136 221280 151142 221292
rect 233418 221280 233424 221292
rect 233476 221280 233482 221332
rect 235258 221280 235264 221332
rect 235316 221320 235322 221332
rect 269206 221320 269212 221332
rect 235316 221292 269212 221320
rect 235316 221280 235322 221292
rect 269206 221280 269212 221292
rect 269264 221280 269270 221332
rect 315942 221280 315948 221332
rect 316000 221320 316006 221332
rect 342254 221320 342260 221332
rect 316000 221292 342260 221320
rect 316000 221280 316006 221292
rect 342254 221280 342260 221292
rect 342312 221280 342318 221332
rect 353938 221280 353944 221332
rect 353996 221320 354002 221332
rect 354646 221320 354674 221428
rect 401134 221416 401140 221428
rect 401192 221416 401198 221468
rect 406746 221416 406752 221468
rect 406804 221456 406810 221468
rect 558454 221456 558460 221468
rect 406804 221428 558460 221456
rect 406804 221416 406810 221428
rect 558454 221416 558460 221428
rect 558512 221416 558518 221468
rect 361298 221348 361304 221400
rect 361356 221388 361362 221400
rect 449894 221388 449900 221400
rect 361356 221360 449900 221388
rect 361356 221348 361362 221360
rect 449894 221348 449900 221360
rect 449952 221348 449958 221400
rect 353996 221292 354674 221320
rect 353996 221280 354002 221292
rect 360102 221280 360108 221332
rect 360160 221320 360166 221332
rect 446582 221320 446588 221332
rect 360160 221292 446588 221320
rect 360160 221280 360166 221292
rect 446582 221280 446588 221292
rect 446640 221280 446646 221332
rect 157794 221212 157800 221264
rect 157852 221252 157858 221264
rect 236178 221252 236184 221264
rect 157852 221224 236184 221252
rect 157852 221212 157858 221224
rect 236178 221212 236184 221224
rect 236236 221212 236242 221264
rect 238570 221212 238576 221264
rect 238628 221252 238634 221264
rect 270678 221252 270684 221264
rect 238628 221224 270684 221252
rect 238628 221212 238634 221224
rect 270678 221212 270684 221224
rect 270736 221212 270742 221264
rect 314562 221212 314568 221264
rect 314620 221252 314626 221264
rect 338850 221252 338856 221264
rect 314620 221224 338856 221252
rect 314620 221212 314626 221224
rect 338850 221212 338856 221224
rect 338908 221212 338914 221264
rect 357066 221212 357072 221264
rect 357124 221252 357130 221264
rect 439774 221252 439780 221264
rect 357124 221224 439780 221252
rect 357124 221212 357130 221224
rect 439774 221212 439780 221224
rect 439832 221212 439838 221264
rect 443638 221212 443644 221264
rect 443696 221252 443702 221264
rect 491938 221252 491944 221264
rect 443696 221224 491944 221252
rect 443696 221212 443702 221224
rect 491938 221212 491944 221224
rect 491996 221212 492002 221264
rect 167914 221144 167920 221196
rect 167972 221184 167978 221196
rect 240502 221184 240508 221196
rect 167972 221156 240508 221184
rect 167972 221144 167978 221156
rect 240502 221144 240508 221156
rect 240560 221144 240566 221196
rect 241974 221144 241980 221196
rect 242032 221184 242038 221196
rect 271966 221184 271972 221196
rect 242032 221156 271972 221184
rect 242032 221144 242038 221156
rect 271966 221144 271972 221156
rect 272024 221144 272030 221196
rect 313182 221144 313188 221196
rect 313240 221184 313246 221196
rect 335538 221184 335544 221196
rect 313240 221156 335544 221184
rect 313240 221144 313246 221156
rect 335538 221144 335544 221156
rect 335596 221144 335602 221196
rect 351546 221144 351552 221196
rect 351604 221184 351610 221196
rect 425514 221184 425520 221196
rect 351604 221156 425520 221184
rect 351604 221144 351610 221156
rect 425514 221144 425520 221156
rect 425572 221144 425578 221196
rect 183922 221076 183928 221128
rect 183980 221116 183986 221128
rect 248598 221116 248604 221128
rect 183980 221088 248604 221116
rect 183980 221076 183986 221088
rect 248598 221076 248604 221088
rect 248656 221076 248662 221128
rect 248690 221076 248696 221128
rect 248748 221116 248754 221128
rect 274818 221116 274824 221128
rect 248748 221088 274824 221116
rect 248748 221076 248754 221088
rect 274818 221076 274824 221088
rect 274876 221076 274882 221128
rect 376110 221076 376116 221128
rect 376168 221116 376174 221128
rect 443178 221116 443184 221128
rect 376168 221088 443184 221116
rect 376168 221076 376174 221088
rect 443178 221076 443184 221088
rect 443236 221076 443242 221128
rect 189810 221008 189816 221060
rect 189868 221048 189874 221060
rect 249426 221048 249432 221060
rect 189868 221020 249432 221048
rect 189868 221008 189874 221020
rect 249426 221008 249432 221020
rect 249484 221008 249490 221060
rect 343266 221008 343272 221060
rect 343324 221048 343330 221060
rect 407850 221048 407856 221060
rect 343324 221020 407856 221048
rect 343324 221008 343330 221020
rect 407850 221008 407856 221020
rect 407908 221008 407914 221060
rect 407942 221008 407948 221060
rect 408000 221048 408006 221060
rect 436462 221048 436468 221060
rect 408000 221020 436468 221048
rect 408000 221008 408006 221020
rect 436462 221008 436468 221020
rect 436520 221008 436526 221060
rect 192938 220940 192944 220992
rect 192996 220980 193002 220992
rect 250806 220980 250812 220992
rect 192996 220952 250812 220980
rect 192996 220940 193002 220952
rect 250806 220940 250812 220952
rect 250864 220940 250870 220992
rect 385678 220940 385684 220992
rect 385736 220980 385742 220992
rect 411254 220980 411260 220992
rect 385736 220952 411260 220980
rect 385736 220940 385742 220952
rect 411254 220940 411260 220952
rect 411312 220940 411318 220992
rect 195146 220872 195152 220924
rect 195204 220912 195210 220924
rect 211614 220912 211620 220924
rect 195204 220884 211620 220912
rect 195204 220872 195210 220884
rect 211614 220872 211620 220884
rect 211672 220872 211678 220924
rect 380250 220872 380256 220924
rect 380308 220912 380314 220924
rect 404446 220912 404452 220924
rect 380308 220884 404452 220912
rect 380308 220872 380314 220884
rect 404446 220872 404452 220884
rect 404504 220872 404510 220924
rect 269592 220816 270448 220844
rect 61102 220736 61108 220788
rect 61160 220776 61166 220788
rect 64138 220776 64144 220788
rect 61160 220748 64144 220776
rect 61160 220736 61166 220748
rect 64138 220736 64144 220748
rect 64196 220736 64202 220788
rect 71222 220736 71228 220788
rect 71280 220776 71286 220788
rect 73798 220776 73804 220788
rect 71280 220748 73804 220776
rect 71280 220736 71286 220748
rect 73798 220736 73804 220748
rect 73856 220736 73862 220788
rect 131758 220736 131764 220788
rect 131816 220776 131822 220788
rect 132402 220776 132408 220788
rect 131816 220748 132408 220776
rect 131816 220736 131822 220748
rect 132402 220736 132408 220748
rect 132460 220736 132466 220788
rect 138474 220736 138480 220788
rect 138532 220776 138538 220788
rect 139302 220776 139308 220788
rect 138532 220748 139308 220776
rect 138532 220736 138538 220748
rect 139302 220736 139308 220748
rect 139360 220736 139366 220788
rect 141878 220736 141884 220788
rect 141936 220776 141942 220788
rect 222102 220776 222108 220788
rect 141936 220748 222108 220776
rect 141936 220736 141942 220748
rect 222102 220736 222108 220748
rect 222160 220736 222166 220788
rect 232682 220736 232688 220788
rect 232740 220776 232746 220788
rect 233142 220776 233148 220788
rect 232740 220748 233148 220776
rect 232740 220736 232746 220748
rect 233142 220736 233148 220748
rect 233200 220736 233206 220788
rect 239398 220736 239404 220788
rect 239456 220776 239462 220788
rect 240042 220776 240048 220788
rect 239456 220748 240048 220776
rect 239456 220736 239462 220748
rect 240042 220736 240048 220748
rect 240100 220736 240106 220788
rect 241146 220736 241152 220788
rect 241204 220776 241210 220788
rect 269592 220776 269620 220816
rect 241204 220748 269620 220776
rect 241204 220736 241210 220748
rect 269666 220736 269672 220788
rect 269724 220776 269730 220788
rect 270310 220776 270316 220788
rect 269724 220748 270316 220776
rect 269724 220736 269730 220748
rect 270310 220736 270316 220748
rect 270368 220736 270374 220788
rect 270420 220776 270448 220816
rect 305546 220804 305552 220856
rect 305604 220844 305610 220856
rect 308582 220844 308588 220856
rect 305604 220816 308588 220844
rect 305604 220804 305610 220816
rect 308582 220804 308588 220816
rect 308640 220804 308646 220856
rect 563698 220804 563704 220856
rect 563756 220844 563762 220856
rect 567930 220844 567936 220856
rect 563756 220816 567936 220844
rect 563756 220804 563762 220816
rect 567930 220804 567936 220816
rect 567988 220804 567994 220856
rect 271322 220776 271328 220788
rect 270420 220748 271328 220776
rect 271322 220736 271328 220748
rect 271380 220736 271386 220788
rect 273898 220736 273904 220788
rect 273956 220776 273962 220788
rect 274542 220776 274548 220788
rect 273956 220748 274548 220776
rect 273956 220736 273962 220748
rect 274542 220736 274548 220748
rect 274600 220736 274606 220788
rect 278130 220736 278136 220788
rect 278188 220776 278194 220788
rect 278682 220776 278688 220788
rect 278188 220748 278688 220776
rect 278188 220736 278194 220748
rect 278682 220736 278688 220748
rect 278740 220736 278746 220788
rect 282362 220736 282368 220788
rect 282420 220776 282426 220788
rect 282822 220776 282828 220788
rect 282420 220748 282828 220776
rect 282420 220736 282426 220748
rect 282822 220736 282828 220748
rect 282880 220736 282886 220788
rect 283190 220736 283196 220788
rect 283248 220776 283254 220788
rect 284110 220776 284116 220788
rect 283248 220748 284116 220776
rect 283248 220736 283254 220748
rect 284110 220736 284116 220748
rect 284168 220736 284174 220788
rect 286502 220736 286508 220788
rect 286560 220776 286566 220788
rect 286962 220776 286968 220788
rect 286560 220748 286968 220776
rect 286560 220736 286566 220748
rect 286962 220736 286968 220748
rect 287020 220736 287026 220788
rect 287330 220736 287336 220788
rect 287388 220776 287394 220788
rect 290642 220776 290648 220788
rect 287388 220748 290648 220776
rect 287388 220736 287394 220748
rect 290642 220736 290648 220748
rect 290700 220736 290706 220788
rect 290734 220736 290740 220788
rect 290792 220776 290798 220788
rect 292206 220776 292212 220788
rect 290792 220748 292212 220776
rect 290792 220736 290798 220748
rect 292206 220736 292212 220748
rect 292264 220736 292270 220788
rect 292482 220736 292488 220788
rect 292540 220776 292546 220788
rect 293218 220776 293224 220788
rect 292540 220748 293224 220776
rect 292540 220736 292546 220748
rect 293218 220736 293224 220748
rect 293276 220736 293282 220788
rect 294966 220736 294972 220788
rect 295024 220776 295030 220788
rect 295518 220776 295524 220788
rect 295024 220748 295524 220776
rect 295024 220736 295030 220748
rect 295518 220736 295524 220748
rect 295576 220736 295582 220788
rect 298002 220736 298008 220788
rect 298060 220776 298066 220788
rect 302234 220776 302240 220788
rect 298060 220748 302240 220776
rect 298060 220736 298066 220748
rect 302234 220736 302240 220748
rect 302292 220736 302298 220788
rect 325326 220736 325332 220788
rect 325384 220776 325390 220788
rect 363230 220776 363236 220788
rect 325384 220748 363236 220776
rect 325384 220736 325390 220748
rect 363230 220736 363236 220748
rect 363288 220736 363294 220788
rect 367002 220736 367008 220788
rect 367060 220776 367066 220788
rect 380894 220776 380900 220788
rect 367060 220748 380900 220776
rect 367060 220736 367066 220748
rect 380894 220736 380900 220748
rect 380952 220736 380958 220788
rect 387794 220736 387800 220788
rect 387852 220776 387858 220788
rect 509878 220776 509884 220788
rect 387852 220748 509884 220776
rect 387852 220736 387858 220748
rect 509878 220736 509884 220748
rect 509936 220736 509942 220788
rect 576394 220776 576400 220788
rect 518866 220748 576400 220776
rect 134978 220668 134984 220720
rect 135036 220708 135042 220720
rect 135036 220680 210464 220708
rect 135036 220668 135042 220680
rect 128170 220600 128176 220652
rect 128228 220640 128234 220652
rect 210436 220640 210464 220680
rect 214190 220668 214196 220720
rect 214248 220708 214254 220720
rect 215294 220708 215300 220720
rect 214248 220680 215300 220708
rect 214248 220668 214254 220680
rect 215294 220668 215300 220680
rect 215352 220668 215358 220720
rect 237742 220668 237748 220720
rect 237800 220708 237806 220720
rect 270126 220708 270132 220720
rect 237800 220680 270132 220708
rect 237800 220668 237806 220680
rect 270126 220668 270132 220680
rect 270184 220668 270190 220720
rect 274450 220668 274456 220720
rect 274508 220708 274514 220720
rect 276658 220708 276664 220720
rect 274508 220680 276664 220708
rect 274508 220668 274514 220680
rect 276658 220668 276664 220680
rect 276716 220668 276722 220720
rect 289078 220668 289084 220720
rect 289136 220708 289142 220720
rect 291838 220708 291844 220720
rect 289136 220680 291844 220708
rect 289136 220668 289142 220680
rect 291838 220668 291844 220680
rect 291896 220668 291902 220720
rect 303062 220668 303068 220720
rect 303120 220708 303126 220720
rect 311158 220708 311164 220720
rect 303120 220680 311164 220708
rect 303120 220668 303126 220680
rect 311158 220668 311164 220680
rect 311216 220668 311222 220720
rect 326246 220668 326252 220720
rect 326304 220708 326310 220720
rect 366634 220708 366640 220720
rect 326304 220680 366640 220708
rect 326304 220668 326310 220680
rect 366634 220668 366640 220680
rect 366692 220668 366698 220720
rect 367646 220668 367652 220720
rect 367704 220708 367710 220720
rect 390554 220708 390560 220720
rect 367704 220680 390560 220708
rect 367704 220668 367710 220680
rect 390554 220668 390560 220680
rect 390612 220668 390618 220720
rect 395706 220668 395712 220720
rect 395764 220708 395770 220720
rect 517514 220708 517520 220720
rect 395764 220680 517520 220708
rect 395764 220668 395770 220680
rect 517514 220668 517520 220680
rect 517572 220708 517578 220720
rect 518866 220708 518894 220748
rect 576394 220736 576400 220748
rect 576452 220736 576458 220788
rect 517572 220680 518894 220708
rect 517572 220668 517578 220680
rect 522574 220668 522580 220720
rect 522632 220708 522638 220720
rect 577314 220708 577320 220720
rect 522632 220680 577320 220708
rect 522632 220668 522638 220680
rect 577314 220668 577320 220680
rect 577372 220668 577378 220720
rect 673362 220668 673368 220720
rect 673420 220708 673426 220720
rect 676030 220708 676036 220720
rect 673420 220680 676036 220708
rect 673420 220668 673426 220680
rect 676030 220668 676036 220680
rect 676088 220668 676094 220720
rect 218054 220640 218060 220652
rect 128228 220612 206416 220640
rect 210436 220612 218060 220640
rect 128228 220600 128234 220612
rect 118326 220532 118332 220584
rect 118384 220572 118390 220584
rect 206388 220572 206416 220612
rect 218054 220600 218060 220612
rect 218112 220600 218118 220652
rect 235902 220600 235908 220652
rect 235960 220640 235966 220652
rect 270034 220640 270040 220652
rect 235960 220612 270040 220640
rect 235960 220600 235966 220612
rect 270034 220600 270040 220612
rect 270092 220600 270098 220652
rect 273070 220600 273076 220652
rect 273128 220640 273134 220652
rect 276750 220640 276756 220652
rect 273128 220612 276756 220640
rect 273128 220600 273134 220612
rect 276750 220600 276756 220612
rect 276808 220600 276814 220652
rect 291470 220600 291476 220652
rect 291528 220640 291534 220652
rect 294046 220640 294052 220652
rect 291528 220612 294052 220640
rect 291528 220600 291534 220612
rect 294046 220600 294052 220612
rect 294104 220600 294110 220652
rect 303430 220600 303436 220652
rect 303488 220640 303494 220652
rect 312814 220640 312820 220652
rect 303488 220612 312820 220640
rect 303488 220600 303494 220612
rect 312814 220600 312820 220612
rect 312872 220600 312878 220652
rect 329558 220600 329564 220652
rect 329616 220640 329622 220652
rect 371694 220640 371700 220652
rect 329616 220612 371700 220640
rect 329616 220600 329622 220612
rect 371694 220600 371700 220612
rect 371752 220600 371758 220652
rect 371878 220600 371884 220652
rect 371936 220640 371942 220652
rect 385954 220640 385960 220652
rect 371936 220612 385960 220640
rect 371936 220600 371942 220612
rect 385954 220600 385960 220612
rect 386012 220600 386018 220652
rect 388438 220600 388444 220652
rect 388496 220640 388502 220652
rect 512822 220640 512828 220652
rect 388496 220612 512828 220640
rect 388496 220600 388502 220612
rect 512822 220600 512828 220612
rect 512880 220600 512886 220652
rect 545758 220600 545764 220652
rect 545816 220640 545822 220652
rect 576486 220640 576492 220652
rect 545816 220612 576492 220640
rect 545816 220600 545822 220612
rect 576486 220600 576492 220612
rect 576544 220600 576550 220652
rect 216674 220572 216680 220584
rect 118384 220544 206324 220572
rect 206388 220544 216680 220572
rect 118384 220532 118390 220544
rect 121270 220464 121276 220516
rect 121328 220504 121334 220516
rect 206186 220504 206192 220516
rect 121328 220476 206192 220504
rect 121328 220464 121334 220476
rect 206186 220464 206192 220476
rect 206244 220464 206250 220516
rect 206296 220504 206324 220544
rect 216674 220532 216680 220544
rect 216732 220532 216738 220584
rect 229370 220532 229376 220584
rect 229428 220572 229434 220584
rect 262582 220572 262588 220584
rect 229428 220544 262588 220572
rect 229428 220532 229434 220544
rect 262582 220532 262588 220544
rect 262640 220532 262646 220584
rect 262950 220532 262956 220584
rect 263008 220572 263014 220584
rect 263502 220572 263508 220584
rect 263008 220544 263508 220572
rect 263008 220532 263014 220544
rect 263502 220532 263508 220544
rect 263560 220532 263566 220584
rect 299382 220532 299388 220584
rect 299440 220572 299446 220584
rect 303614 220572 303620 220584
rect 299440 220544 303620 220572
rect 299440 220532 299446 220544
rect 303614 220532 303620 220544
rect 303672 220532 303678 220584
rect 304810 220532 304816 220584
rect 304868 220572 304874 220584
rect 316126 220572 316132 220584
rect 304868 220544 316132 220572
rect 304868 220532 304874 220544
rect 316126 220532 316132 220544
rect 316184 220532 316190 220584
rect 329650 220532 329656 220584
rect 329708 220572 329714 220584
rect 373350 220572 373356 220584
rect 329708 220544 373356 220572
rect 329708 220532 329714 220544
rect 373350 220532 373356 220544
rect 373408 220532 373414 220584
rect 394694 220572 394700 220584
rect 389146 220544 394700 220572
rect 208210 220504 208216 220516
rect 206296 220476 208216 220504
rect 208210 220464 208216 220476
rect 208268 220464 208274 220516
rect 224954 220504 224960 220516
rect 219406 220476 224960 220504
rect 111610 220396 111616 220448
rect 111668 220436 111674 220448
rect 206922 220436 206928 220448
rect 111668 220408 206928 220436
rect 111668 220396 111674 220408
rect 206922 220396 206928 220408
rect 206980 220396 206986 220448
rect 145190 220328 145196 220380
rect 145248 220368 145254 220380
rect 146202 220368 146208 220380
rect 145248 220340 146208 220368
rect 145248 220328 145254 220340
rect 146202 220328 146208 220340
rect 146260 220328 146266 220380
rect 155310 220328 155316 220380
rect 155368 220368 155374 220380
rect 155862 220368 155868 220380
rect 155368 220340 155868 220368
rect 155368 220328 155374 220340
rect 155862 220328 155868 220340
rect 155920 220328 155926 220380
rect 168742 220328 168748 220380
rect 168800 220368 168806 220380
rect 169662 220368 169668 220380
rect 168800 220340 169668 220368
rect 168800 220328 168806 220340
rect 169662 220328 169668 220340
rect 169720 220328 169726 220380
rect 178862 220328 178868 220380
rect 178920 220368 178926 220380
rect 179322 220368 179328 220380
rect 178920 220340 179328 220368
rect 178920 220328 178926 220340
rect 179322 220328 179328 220340
rect 179380 220328 179386 220380
rect 192294 220328 192300 220380
rect 192352 220368 192358 220380
rect 219406 220368 219434 220476
rect 224954 220464 224960 220476
rect 225012 220464 225018 220516
rect 231026 220464 231032 220516
rect 231084 220504 231090 220516
rect 268286 220504 268292 220516
rect 231084 220476 268292 220504
rect 231084 220464 231090 220476
rect 268286 220464 268292 220476
rect 268344 220464 268350 220516
rect 299290 220464 299296 220516
rect 299348 220504 299354 220516
rect 305270 220504 305276 220516
rect 299348 220476 305276 220504
rect 299348 220464 299354 220476
rect 305270 220464 305276 220476
rect 305328 220464 305334 220516
rect 306190 220464 306196 220516
rect 306248 220504 306254 220516
rect 317874 220504 317880 220516
rect 306248 220476 317880 220504
rect 306248 220464 306254 220476
rect 317874 220464 317880 220476
rect 317932 220464 317938 220516
rect 319346 220464 319352 220516
rect 319404 220504 319410 220516
rect 339678 220504 339684 220516
rect 319404 220476 339684 220504
rect 319404 220464 319410 220476
rect 339678 220464 339684 220476
rect 339736 220464 339742 220516
rect 342898 220464 342904 220516
rect 342956 220504 342962 220516
rect 386782 220504 386788 220516
rect 342956 220476 386788 220504
rect 342956 220464 342962 220476
rect 386782 220464 386788 220476
rect 386840 220464 386846 220516
rect 222562 220396 222568 220448
rect 222620 220436 222626 220448
rect 264330 220436 264336 220448
rect 222620 220408 264336 220436
rect 222620 220396 222626 220408
rect 264330 220396 264336 220408
rect 264388 220396 264394 220448
rect 306098 220396 306104 220448
rect 306156 220436 306162 220448
rect 319530 220436 319536 220448
rect 306156 220408 319536 220436
rect 306156 220396 306162 220408
rect 319530 220396 319536 220408
rect 319588 220396 319594 220448
rect 331030 220396 331036 220448
rect 331088 220436 331094 220448
rect 375374 220436 375380 220448
rect 331088 220408 375380 220436
rect 331088 220396 331094 220408
rect 375374 220396 375380 220408
rect 375432 220396 375438 220448
rect 376018 220396 376024 220448
rect 376076 220436 376082 220448
rect 389146 220436 389174 220544
rect 394694 220532 394700 220544
rect 394752 220532 394758 220584
rect 395338 220532 395344 220584
rect 395396 220572 395402 220584
rect 519998 220572 520004 220584
rect 395396 220544 520004 220572
rect 395396 220532 395402 220544
rect 519998 220532 520004 220544
rect 520056 220572 520062 220584
rect 574922 220572 574928 220584
rect 520056 220544 574928 220572
rect 520056 220532 520062 220544
rect 574922 220532 574928 220544
rect 574980 220532 574986 220584
rect 391474 220464 391480 220516
rect 391532 220504 391538 220516
rect 522574 220504 522580 220516
rect 391532 220476 522580 220504
rect 391532 220464 391538 220476
rect 522574 220464 522580 220476
rect 522632 220464 522638 220516
rect 525058 220464 525064 220516
rect 525116 220504 525122 220516
rect 577130 220504 577136 220516
rect 525116 220476 577136 220504
rect 525116 220464 525122 220476
rect 577130 220464 577136 220476
rect 577188 220464 577194 220516
rect 376076 220408 389174 220436
rect 376076 220396 376082 220408
rect 394602 220396 394608 220448
rect 394660 220436 394666 220448
rect 527266 220436 527272 220448
rect 394660 220408 527272 220436
rect 394660 220396 394666 220408
rect 527266 220396 527272 220408
rect 527324 220436 527330 220448
rect 576302 220436 576308 220448
rect 527324 220408 576308 220436
rect 527324 220396 527330 220408
rect 576302 220396 576308 220408
rect 576360 220396 576366 220448
rect 192352 220340 219434 220368
rect 192352 220328 192358 220340
rect 224310 220328 224316 220380
rect 224368 220368 224374 220380
rect 265434 220368 265440 220380
rect 224368 220340 265440 220368
rect 224368 220328 224374 220340
rect 265434 220328 265440 220340
rect 265492 220328 265498 220380
rect 268010 220328 268016 220380
rect 268068 220368 268074 220380
rect 275370 220368 275376 220380
rect 268068 220340 275376 220368
rect 268068 220328 268074 220340
rect 275370 220328 275376 220340
rect 275428 220328 275434 220380
rect 307570 220328 307576 220380
rect 307628 220368 307634 220380
rect 321554 220368 321560 220380
rect 307628 220340 321560 220368
rect 307628 220328 307634 220340
rect 321554 220328 321560 220340
rect 321612 220328 321618 220380
rect 330478 220328 330484 220380
rect 330536 220368 330542 220380
rect 376938 220368 376944 220380
rect 330536 220340 376944 220368
rect 330536 220328 330542 220340
rect 376938 220328 376944 220340
rect 376996 220328 377002 220380
rect 378042 220328 378048 220380
rect 378100 220368 378106 220380
rect 387794 220368 387800 220380
rect 378100 220340 387800 220368
rect 378100 220328 378106 220340
rect 387794 220328 387800 220340
rect 387852 220328 387858 220380
rect 394510 220328 394516 220380
rect 394568 220368 394574 220380
rect 530118 220368 530124 220380
rect 394568 220340 530124 220368
rect 394568 220328 394574 220340
rect 530118 220328 530124 220340
rect 530176 220368 530182 220380
rect 574830 220368 574836 220380
rect 530176 220340 574836 220368
rect 530176 220328 530182 220340
rect 574830 220328 574836 220340
rect 574888 220328 574894 220380
rect 79594 220260 79600 220312
rect 79652 220300 79658 220312
rect 100754 220300 100760 220312
rect 79652 220272 100760 220300
rect 79652 220260 79658 220272
rect 100754 220260 100760 220272
rect 100812 220260 100818 220312
rect 104710 220260 104716 220312
rect 104768 220300 104774 220312
rect 204162 220300 204168 220312
rect 104768 220272 204168 220300
rect 104768 220260 104774 220272
rect 204162 220260 204168 220272
rect 204220 220260 204226 220312
rect 207474 220260 207480 220312
rect 207532 220300 207538 220312
rect 213822 220300 213828 220312
rect 207532 220272 213828 220300
rect 207532 220260 207538 220272
rect 213822 220260 213828 220272
rect 213880 220260 213886 220312
rect 217594 220260 217600 220312
rect 217652 220300 217658 220312
rect 260098 220300 260104 220312
rect 217652 220272 260104 220300
rect 217652 220260 217658 220272
rect 260098 220260 260104 220272
rect 260156 220260 260162 220312
rect 264698 220260 264704 220312
rect 264756 220300 264762 220312
rect 273806 220300 273812 220312
rect 264756 220272 273812 220300
rect 264756 220260 264762 220272
rect 273806 220260 273812 220272
rect 273864 220260 273870 220312
rect 307386 220260 307392 220312
rect 307444 220300 307450 220312
rect 322934 220300 322940 220312
rect 307444 220272 322940 220300
rect 307444 220260 307450 220272
rect 322934 220260 322940 220272
rect 322992 220260 322998 220312
rect 332226 220260 332232 220312
rect 332284 220300 332290 220312
rect 378410 220300 378416 220312
rect 332284 220272 378416 220300
rect 332284 220260 332290 220272
rect 378410 220260 378416 220272
rect 378468 220260 378474 220312
rect 378778 220260 378784 220312
rect 378836 220300 378842 220312
rect 391934 220300 391940 220312
rect 378836 220272 391940 220300
rect 378836 220260 378842 220272
rect 391934 220260 391940 220272
rect 391992 220260 391998 220312
rect 396718 220260 396724 220312
rect 396776 220300 396782 220312
rect 532694 220300 532700 220312
rect 396776 220272 532700 220300
rect 396776 220260 396782 220272
rect 532694 220260 532700 220272
rect 532752 220260 532758 220312
rect 66070 220192 66076 220244
rect 66128 220232 66134 220244
rect 69014 220232 69020 220244
rect 66128 220204 69020 220232
rect 66128 220192 66134 220204
rect 69014 220192 69020 220204
rect 69072 220192 69078 220244
rect 94774 220192 94780 220244
rect 94832 220232 94838 220244
rect 202414 220232 202420 220244
rect 94832 220204 202420 220232
rect 94832 220192 94838 220204
rect 202414 220192 202420 220204
rect 202472 220192 202478 220244
rect 206186 220192 206192 220244
rect 206244 220232 206250 220244
rect 213914 220232 213920 220244
rect 206244 220204 213920 220232
rect 206244 220192 206250 220204
rect 213914 220192 213920 220204
rect 213972 220192 213978 220244
rect 215846 220192 215852 220244
rect 215904 220232 215910 220244
rect 261478 220232 261484 220244
rect 215904 220204 261484 220232
rect 215904 220192 215910 220204
rect 261478 220192 261484 220204
rect 261536 220192 261542 220244
rect 262582 220192 262588 220244
rect 262640 220232 262646 220244
rect 267182 220232 267188 220244
rect 262640 220204 267188 220232
rect 262640 220192 262646 220204
rect 267182 220192 267188 220204
rect 267240 220192 267246 220244
rect 271414 220192 271420 220244
rect 271472 220232 271478 220244
rect 275278 220232 275284 220244
rect 271472 220204 275284 220232
rect 271472 220192 271478 220204
rect 275278 220192 275284 220204
rect 275336 220192 275342 220244
rect 308766 220192 308772 220244
rect 308824 220232 308830 220244
rect 326246 220232 326252 220244
rect 308824 220204 326252 220232
rect 308824 220192 308830 220204
rect 326246 220192 326252 220204
rect 326304 220192 326310 220244
rect 332410 220192 332416 220244
rect 332468 220232 332474 220244
rect 380066 220232 380072 220244
rect 332468 220204 380072 220232
rect 332468 220192 332474 220204
rect 380066 220192 380072 220204
rect 380124 220192 380130 220244
rect 380710 220192 380716 220244
rect 380768 220232 380774 220244
rect 395246 220232 395252 220244
rect 380768 220204 395252 220232
rect 380768 220192 380774 220204
rect 395246 220192 395252 220204
rect 395304 220192 395310 220244
rect 396810 220192 396816 220244
rect 396868 220232 396874 220244
rect 535362 220232 535368 220244
rect 396868 220204 535368 220232
rect 396868 220192 396874 220204
rect 535362 220192 535368 220204
rect 535420 220192 535426 220244
rect 672626 220192 672632 220244
rect 672684 220232 672690 220244
rect 676030 220232 676036 220244
rect 672684 220204 676036 220232
rect 672684 220192 672690 220204
rect 676030 220192 676036 220204
rect 676088 220192 676094 220244
rect 81250 220124 81256 220176
rect 81308 220164 81314 220176
rect 203518 220164 203524 220176
rect 81308 220136 203524 220164
rect 81308 220124 81314 220136
rect 203518 220124 203524 220136
rect 203576 220124 203582 220176
rect 204070 220124 204076 220176
rect 204128 220164 204134 220176
rect 209866 220164 209872 220176
rect 204128 220136 209872 220164
rect 204128 220124 204134 220136
rect 209866 220124 209872 220136
rect 209924 220124 209930 220176
rect 210786 220124 210792 220176
rect 210844 220164 210850 220176
rect 210844 220136 252232 220164
rect 210844 220124 210850 220136
rect 64506 220056 64512 220108
rect 64564 220096 64570 220108
rect 192846 220096 192852 220108
rect 64564 220068 192852 220096
rect 64564 220056 64570 220068
rect 192846 220056 192852 220068
rect 192904 220056 192910 220108
rect 209130 220056 209136 220108
rect 209188 220096 209194 220108
rect 252094 220096 252100 220108
rect 209188 220068 252100 220096
rect 209188 220056 209194 220068
rect 252094 220056 252100 220068
rect 252152 220056 252158 220108
rect 252204 220096 252232 220136
rect 254578 220124 254584 220176
rect 254636 220164 254642 220176
rect 255222 220164 255228 220176
rect 254636 220136 255228 220164
rect 254636 220124 254642 220136
rect 255222 220124 255228 220136
rect 255280 220124 255286 220176
rect 257890 220124 257896 220176
rect 257948 220164 257954 220176
rect 271230 220164 271236 220176
rect 257948 220136 271236 220164
rect 257948 220124 257954 220136
rect 271230 220124 271236 220136
rect 271288 220124 271294 220176
rect 279418 220164 279424 220176
rect 277366 220136 279424 220164
rect 255958 220096 255964 220108
rect 252204 220068 255964 220096
rect 255958 220056 255964 220068
rect 256016 220056 256022 220108
rect 266170 220056 266176 220108
rect 266228 220096 266234 220108
rect 277366 220096 277394 220136
rect 279418 220124 279424 220136
rect 279476 220124 279482 220176
rect 280614 220124 280620 220176
rect 280672 220164 280678 220176
rect 281442 220164 281448 220176
rect 280672 220136 281448 220164
rect 280672 220124 280678 220136
rect 281442 220124 281448 220136
rect 281500 220124 281506 220176
rect 287514 220164 287520 220176
rect 287026 220136 287520 220164
rect 266228 220068 277394 220096
rect 266228 220056 266234 220068
rect 278590 220056 278596 220108
rect 278648 220096 278654 220108
rect 287026 220096 287054 220136
rect 287514 220124 287520 220136
rect 287572 220124 287578 220176
rect 304442 220124 304448 220176
rect 304500 220164 304506 220176
rect 314654 220164 314660 220176
rect 304500 220136 314660 220164
rect 304500 220124 304506 220136
rect 314654 220124 314660 220136
rect 314712 220124 314718 220176
rect 315390 220124 315396 220176
rect 315448 220164 315454 220176
rect 332962 220164 332968 220176
rect 315448 220136 332968 220164
rect 315448 220124 315454 220136
rect 332962 220124 332968 220136
rect 333020 220124 333026 220176
rect 333790 220124 333796 220176
rect 333848 220164 333854 220176
rect 381814 220164 381820 220176
rect 333848 220136 381820 220164
rect 333848 220124 333854 220136
rect 381814 220124 381820 220136
rect 381872 220124 381878 220176
rect 382274 220124 382280 220176
rect 382332 220164 382338 220176
rect 396902 220164 396908 220176
rect 382332 220136 396908 220164
rect 382332 220124 382338 220136
rect 396902 220124 396908 220136
rect 396960 220124 396966 220176
rect 398558 220124 398564 220176
rect 398616 220164 398622 220176
rect 537386 220164 537392 220176
rect 398616 220136 537392 220164
rect 398616 220124 398622 220136
rect 537386 220124 537392 220136
rect 537444 220124 537450 220176
rect 548150 220124 548156 220176
rect 548208 220164 548214 220176
rect 548208 220136 552796 220164
rect 548208 220124 548214 220136
rect 278648 220068 287054 220096
rect 278648 220056 278654 220068
rect 301958 220056 301964 220108
rect 302016 220096 302022 220108
rect 309410 220096 309416 220108
rect 302016 220068 309416 220096
rect 302016 220056 302022 220068
rect 309410 220056 309416 220068
rect 309468 220056 309474 220108
rect 310238 220056 310244 220108
rect 310296 220096 310302 220108
rect 329834 220096 329840 220108
rect 310296 220068 329840 220096
rect 310296 220056 310302 220068
rect 329834 220056 329840 220068
rect 329892 220056 329898 220108
rect 333882 220056 333888 220108
rect 333940 220096 333946 220108
rect 383654 220096 383660 220108
rect 333940 220068 383660 220096
rect 333940 220056 333946 220068
rect 383654 220056 383660 220068
rect 383712 220056 383718 220108
rect 385494 220056 385500 220108
rect 385552 220096 385558 220108
rect 400306 220096 400312 220108
rect 385552 220068 400312 220096
rect 385552 220056 385558 220068
rect 400306 220056 400312 220068
rect 400364 220056 400370 220108
rect 404262 220056 404268 220108
rect 404320 220096 404326 220108
rect 404320 220068 528554 220096
rect 404320 220056 404326 220068
rect 148594 219988 148600 220040
rect 148652 220028 148658 220040
rect 223114 220028 223120 220040
rect 148652 220000 223120 220028
rect 148652 219988 148658 220000
rect 223114 219988 223120 220000
rect 223172 219988 223178 220040
rect 247862 219988 247868 220040
rect 247920 220028 247926 220040
rect 248322 220028 248328 220040
rect 247920 220000 248328 220028
rect 247920 219988 247926 220000
rect 248322 219988 248328 220000
rect 248380 219988 248386 220040
rect 272886 220028 272892 220040
rect 249536 220000 272892 220028
rect 151722 219920 151728 219972
rect 151780 219960 151786 219972
rect 224034 219960 224040 219972
rect 151780 219932 224040 219960
rect 151780 219920 151786 219932
rect 224034 219920 224040 219932
rect 224092 219920 224098 219972
rect 246114 219920 246120 219972
rect 246172 219960 246178 219972
rect 246942 219960 246948 219972
rect 246172 219932 246948 219960
rect 246172 219920 246178 219932
rect 246942 219920 246948 219932
rect 247000 219920 247006 219972
rect 249536 219960 249564 220000
rect 272886 219988 272892 220000
rect 272944 219988 272950 220040
rect 289630 219988 289636 220040
rect 289688 220028 289694 220040
rect 292850 220028 292856 220040
rect 289688 220000 292856 220028
rect 289688 219988 289694 220000
rect 292850 219988 292856 220000
rect 292908 219988 292914 220040
rect 318058 219988 318064 220040
rect 318116 220028 318122 220040
rect 336734 220028 336740 220040
rect 318116 220000 336740 220028
rect 318116 219988 318122 220000
rect 336734 219988 336740 220000
rect 336792 219988 336798 220040
rect 341518 219988 341524 220040
rect 341576 220028 341582 220040
rect 370038 220028 370044 220040
rect 341576 220000 370044 220028
rect 341576 219988 341582 220000
rect 370038 219988 370044 220000
rect 370096 219988 370102 220040
rect 370222 219988 370228 220040
rect 370280 220028 370286 220040
rect 382642 220028 382648 220040
rect 370280 220000 382648 220028
rect 370280 219988 370286 220000
rect 382642 219988 382648 220000
rect 382700 219988 382706 220040
rect 383378 219988 383384 220040
rect 383436 220028 383442 220040
rect 502426 220028 502432 220040
rect 383436 220000 502432 220028
rect 383436 219988 383442 220000
rect 502426 219988 502432 220000
rect 502484 219988 502490 220040
rect 528526 220028 528554 220068
rect 542998 220056 543004 220108
rect 543056 220096 543062 220108
rect 543056 220068 552704 220096
rect 543056 220056 543062 220068
rect 549622 220028 549628 220040
rect 528526 220000 549628 220028
rect 549622 219988 549628 220000
rect 549680 219988 549686 220040
rect 276198 219960 276204 219972
rect 248386 219932 249564 219960
rect 249628 219932 276204 219960
rect 158622 219852 158628 219904
rect 158680 219892 158686 219904
rect 227346 219892 227352 219904
rect 158680 219864 227352 219892
rect 158680 219852 158686 219864
rect 227346 219852 227352 219864
rect 227404 219852 227410 219904
rect 242802 219852 242808 219904
rect 242860 219892 242866 219904
rect 248386 219892 248414 219932
rect 242860 219864 248414 219892
rect 242860 219852 242866 219864
rect 249518 219852 249524 219904
rect 249576 219892 249582 219904
rect 249628 219892 249656 219932
rect 276198 219920 276204 219932
rect 276256 219920 276262 219972
rect 284846 219920 284852 219972
rect 284904 219960 284910 219972
rect 285582 219960 285588 219972
rect 284904 219932 285588 219960
rect 284904 219920 284910 219932
rect 285582 219920 285588 219932
rect 285640 219920 285646 219972
rect 340138 219920 340144 219972
rect 340196 219960 340202 219972
rect 360194 219960 360200 219972
rect 340196 219932 360200 219960
rect 340196 219920 340202 219932
rect 360194 219920 360200 219932
rect 360252 219920 360258 219972
rect 365254 219920 365260 219972
rect 365312 219960 365318 219972
rect 377582 219960 377588 219972
rect 365312 219932 377588 219960
rect 365312 219920 365318 219932
rect 377582 219920 377588 219932
rect 377640 219920 377646 219972
rect 384942 219920 384948 219972
rect 385000 219960 385006 219972
rect 504910 219960 504916 219972
rect 385000 219932 504916 219960
rect 385000 219920 385006 219932
rect 504910 219920 504916 219932
rect 504968 219920 504974 219972
rect 552676 219960 552704 220068
rect 552768 220028 552796 220136
rect 560754 220124 560760 220176
rect 560812 220164 560818 220176
rect 617150 220164 617156 220176
rect 560812 220136 617156 220164
rect 560812 220124 560818 220136
rect 617150 220124 617156 220136
rect 617208 220124 617214 220176
rect 552842 220056 552848 220108
rect 552900 220096 552906 220108
rect 609606 220096 609612 220108
rect 552900 220068 609612 220096
rect 552900 220056 552906 220068
rect 609606 220056 609612 220068
rect 609664 220056 609670 220108
rect 614114 220028 614120 220040
rect 552768 220000 614120 220028
rect 614114 219988 614120 220000
rect 614172 219988 614178 220040
rect 611722 219960 611728 219972
rect 552676 219932 611728 219960
rect 611722 219920 611728 219932
rect 611780 219920 611786 219972
rect 249576 219864 249656 219892
rect 249576 219852 249582 219864
rect 252922 219852 252928 219904
rect 252980 219892 252986 219904
rect 277578 219892 277584 219904
rect 252980 219864 277584 219892
rect 252980 219852 252986 219864
rect 277578 219852 277584 219864
rect 277636 219852 277642 219904
rect 322198 219852 322204 219904
rect 322256 219892 322262 219904
rect 343082 219892 343088 219904
rect 322256 219864 343088 219892
rect 322256 219852 322262 219864
rect 343082 219852 343088 219864
rect 343140 219852 343146 219904
rect 363138 219852 363144 219904
rect 363196 219892 363202 219904
rect 391014 219892 391020 219904
rect 363196 219864 391020 219892
rect 363196 219852 363202 219864
rect 391014 219852 391020 219864
rect 391072 219852 391078 219904
rect 399478 219852 399484 219904
rect 399536 219892 399542 219904
rect 513834 219892 513840 219904
rect 399536 219864 513840 219892
rect 399536 219852 399542 219864
rect 513834 219852 513840 219864
rect 513892 219852 513898 219904
rect 540422 219852 540428 219904
rect 540480 219892 540486 219904
rect 613010 219892 613016 219904
rect 540480 219864 613016 219892
rect 540480 219852 540486 219864
rect 613010 219852 613016 219864
rect 613068 219852 613074 219904
rect 673270 219852 673276 219904
rect 673328 219892 673334 219904
rect 676030 219892 676036 219904
rect 673328 219864 676036 219892
rect 673328 219852 673334 219864
rect 676030 219852 676036 219864
rect 676088 219852 676094 219904
rect 165430 219784 165436 219836
rect 165488 219824 165494 219836
rect 227714 219824 227720 219836
rect 165488 219796 227720 219824
rect 165488 219784 165494 219796
rect 227714 219784 227720 219796
rect 227772 219784 227778 219836
rect 256234 219784 256240 219836
rect 256292 219824 256298 219836
rect 278958 219824 278964 219836
rect 256292 219796 278964 219824
rect 256292 219784 256298 219796
rect 278958 219784 278964 219796
rect 279016 219784 279022 219836
rect 293218 219784 293224 219836
rect 293276 219824 293282 219836
rect 293954 219824 293960 219836
rect 293276 219796 293960 219824
rect 293276 219784 293282 219796
rect 293954 219784 293960 219796
rect 294012 219784 294018 219836
rect 338758 219784 338764 219836
rect 338816 219824 338822 219836
rect 356514 219824 356520 219836
rect 338816 219796 356520 219824
rect 338816 219784 338822 219796
rect 356514 219784 356520 219796
rect 356572 219784 356578 219836
rect 362954 219784 362960 219836
rect 363012 219824 363018 219836
rect 368474 219824 368480 219836
rect 363012 219796 368480 219824
rect 363012 219784 363018 219796
rect 368474 219784 368480 219796
rect 368532 219784 368538 219836
rect 375282 219784 375288 219836
rect 375340 219824 375346 219836
rect 379514 219824 379520 219836
rect 375340 219796 379520 219824
rect 375340 219784 375346 219796
rect 379514 219784 379520 219796
rect 379572 219784 379578 219836
rect 380986 219784 380992 219836
rect 381044 219824 381050 219836
rect 484394 219824 484400 219836
rect 381044 219796 484400 219824
rect 381044 219784 381050 219796
rect 484394 219784 484400 219796
rect 484452 219784 484458 219836
rect 535362 219784 535368 219836
rect 535420 219824 535426 219836
rect 609882 219824 609888 219836
rect 535420 219796 609888 219824
rect 535420 219784 535426 219796
rect 609882 219784 609888 219796
rect 609940 219784 609946 219836
rect 172146 219716 172152 219768
rect 172204 219756 172210 219768
rect 232406 219756 232412 219768
rect 172204 219728 232412 219756
rect 172204 219716 172210 219728
rect 232406 219716 232412 219728
rect 232464 219716 232470 219768
rect 250990 219716 250996 219768
rect 251048 219756 251054 219768
rect 271138 219756 271144 219768
rect 251048 219728 271144 219756
rect 251048 219716 251054 219728
rect 271138 219716 271144 219728
rect 271196 219716 271202 219768
rect 337378 219716 337384 219768
rect 337436 219756 337442 219768
rect 353294 219756 353300 219768
rect 337436 219728 353300 219756
rect 337436 219716 337442 219728
rect 353294 219716 353300 219728
rect 353352 219716 353358 219768
rect 372614 219716 372620 219768
rect 372672 219756 372678 219768
rect 384298 219756 384304 219768
rect 372672 219728 384304 219756
rect 372672 219716 372678 219728
rect 384298 219716 384304 219728
rect 384356 219716 384362 219768
rect 387150 219716 387156 219768
rect 387208 219756 387214 219768
rect 409874 219756 409880 219768
rect 387208 219728 409880 219756
rect 387208 219716 387214 219728
rect 409874 219716 409880 219728
rect 409932 219716 409938 219768
rect 409966 219716 409972 219768
rect 410024 219756 410030 219768
rect 416222 219756 416228 219768
rect 410024 219728 416228 219756
rect 410024 219716 410030 219728
rect 416222 219716 416228 219728
rect 416280 219716 416286 219768
rect 515398 219716 515404 219768
rect 515456 219756 515462 219768
rect 625338 219756 625344 219768
rect 515456 219728 625344 219756
rect 515456 219716 515462 219728
rect 625338 219716 625344 219728
rect 625396 219716 625402 219768
rect 185578 219648 185584 219700
rect 185636 219688 185642 219700
rect 186958 219688 186964 219700
rect 185636 219660 186964 219688
rect 185636 219648 185642 219660
rect 186958 219648 186964 219660
rect 187016 219648 187022 219700
rect 232774 219688 232780 219700
rect 187068 219660 232780 219688
rect 181990 219580 181996 219632
rect 182048 219620 182054 219632
rect 187068 219620 187096 219660
rect 232774 219648 232780 219660
rect 232832 219648 232838 219700
rect 252094 219648 252100 219700
rect 252152 219688 252158 219700
rect 257338 219688 257344 219700
rect 252152 219660 257344 219688
rect 252152 219648 252158 219660
rect 257338 219648 257344 219660
rect 257396 219648 257402 219700
rect 261294 219648 261300 219700
rect 261352 219688 261358 219700
rect 272978 219688 272984 219700
rect 261352 219660 272984 219688
rect 261352 219648 261358 219660
rect 272978 219648 272984 219660
rect 273036 219648 273042 219700
rect 334710 219648 334716 219700
rect 334768 219688 334774 219700
rect 349798 219688 349804 219700
rect 334768 219660 349804 219688
rect 334768 219648 334774 219660
rect 349798 219648 349804 219660
rect 349856 219648 349862 219700
rect 386414 219648 386420 219700
rect 386472 219688 386478 219700
rect 398834 219688 398840 219700
rect 386472 219660 398840 219688
rect 386472 219648 386478 219660
rect 398834 219648 398840 219660
rect 398892 219648 398898 219700
rect 415302 219648 415308 219700
rect 415360 219688 415366 219700
rect 418154 219688 418160 219700
rect 415360 219660 418160 219688
rect 415360 219648 415366 219660
rect 418154 219648 418160 219660
rect 418212 219648 418218 219700
rect 512822 219648 512828 219700
rect 512880 219688 512886 219700
rect 625246 219688 625252 219700
rect 512880 219660 625252 219688
rect 512880 219648 512886 219660
rect 625246 219648 625252 219660
rect 625304 219648 625310 219700
rect 182048 219592 187096 219620
rect 182048 219580 182054 219592
rect 188890 219580 188896 219632
rect 188948 219620 188954 219632
rect 234614 219620 234620 219632
rect 188948 219592 234620 219620
rect 188948 219580 188954 219592
rect 234614 219580 234620 219592
rect 234672 219580 234678 219632
rect 300486 219580 300492 219632
rect 300544 219620 300550 219632
rect 306926 219620 306932 219632
rect 300544 219592 306932 219620
rect 300544 219580 300550 219592
rect 306926 219580 306932 219592
rect 306984 219580 306990 219632
rect 334618 219580 334624 219632
rect 334676 219620 334682 219632
rect 346486 219620 346492 219632
rect 334676 219592 346492 219620
rect 334676 219580 334682 219592
rect 346486 219580 346492 219592
rect 346544 219580 346550 219632
rect 377306 219580 377312 219632
rect 377364 219620 377370 219632
rect 388530 219620 388536 219632
rect 377364 219592 388536 219620
rect 377364 219580 377370 219592
rect 388530 219580 388536 219592
rect 388588 219580 388594 219632
rect 498654 219580 498660 219632
rect 498712 219620 498718 219632
rect 505002 219620 505008 219632
rect 498712 219592 505008 219620
rect 498712 219580 498718 219592
rect 505002 219580 505008 219592
rect 505060 219580 505066 219632
rect 509878 219580 509884 219632
rect 509936 219620 509942 219632
rect 623866 219620 623872 219632
rect 509936 219592 623872 219620
rect 509936 219580 509942 219592
rect 623866 219580 623872 219592
rect 623924 219580 623930 219632
rect 97810 219512 97816 219564
rect 97868 219552 97874 219564
rect 97868 219524 103514 219552
rect 97868 219512 97874 219524
rect 54386 219444 54392 219496
rect 54444 219484 54450 219496
rect 56318 219484 56324 219496
rect 54444 219456 56324 219484
rect 54444 219444 54450 219456
rect 56318 219444 56324 219456
rect 56376 219444 56382 219496
rect 56594 219444 56600 219496
rect 56652 219444 56658 219496
rect 103486 219484 103514 219524
rect 195698 219512 195704 219564
rect 195756 219552 195762 219564
rect 234706 219552 234712 219564
rect 195756 219524 234712 219552
rect 195756 219512 195762 219524
rect 234706 219512 234712 219524
rect 234764 219512 234770 219564
rect 301590 219512 301596 219564
rect 301648 219552 301654 219564
rect 307754 219552 307760 219564
rect 301648 219524 307760 219552
rect 301648 219512 301654 219524
rect 307754 219512 307760 219524
rect 307812 219512 307818 219564
rect 406378 219512 406384 219564
rect 406436 219552 406442 219564
rect 412910 219552 412916 219564
rect 406436 219524 412916 219552
rect 406436 219512 406442 219524
rect 412910 219512 412916 219524
rect 412968 219512 412974 219564
rect 502426 219512 502432 219564
rect 502484 219552 502490 219564
rect 623038 219552 623044 219564
rect 502484 219524 623044 219552
rect 502484 219512 502490 219524
rect 623038 219512 623044 219524
rect 623096 219512 623102 219564
rect 195146 219484 195152 219496
rect 103486 219456 195152 219484
rect 195146 219444 195152 219456
rect 195204 219444 195210 219496
rect 202414 219444 202420 219496
rect 202472 219484 202478 219496
rect 237374 219484 237380 219496
rect 202472 219456 237380 219484
rect 202472 219444 202478 219456
rect 237374 219444 237380 219456
rect 237432 219444 237438 219496
rect 267182 219444 267188 219496
rect 267240 219484 267246 219496
rect 268378 219484 268384 219496
rect 267240 219456 268384 219484
rect 267240 219444 267246 219456
rect 268378 219444 268384 219456
rect 268436 219444 268442 219496
rect 276474 219444 276480 219496
rect 276532 219484 276538 219496
rect 278038 219484 278044 219496
rect 276532 219456 278044 219484
rect 276532 219444 276538 219456
rect 278038 219444 278044 219456
rect 278096 219444 278102 219496
rect 300578 219444 300584 219496
rect 300636 219484 300642 219496
rect 306374 219484 306380 219496
rect 300636 219456 306380 219484
rect 300636 219444 300642 219456
rect 306374 219444 306380 219456
rect 306432 219444 306438 219496
rect 360286 219444 360292 219496
rect 360344 219484 360350 219496
rect 364978 219484 364984 219496
rect 360344 219456 364984 219484
rect 360344 219444 360350 219456
rect 364978 219444 364984 219456
rect 365036 219444 365042 219496
rect 371326 219444 371332 219496
rect 371384 219484 371390 219496
rect 375926 219484 375932 219496
rect 371384 219456 375932 219484
rect 371384 219444 371390 219456
rect 375926 219444 375932 219456
rect 375984 219444 375990 219496
rect 378502 219444 378508 219496
rect 378560 219484 378566 219496
rect 385126 219484 385132 219496
rect 378560 219456 385132 219484
rect 378560 219444 378566 219456
rect 385126 219444 385132 219456
rect 385184 219444 385190 219496
rect 390646 219444 390652 219496
rect 390704 219484 390710 219496
rect 393590 219484 393596 219496
rect 390704 219456 393596 219484
rect 390704 219444 390710 219456
rect 393590 219444 393596 219456
rect 393648 219444 393654 219496
rect 408494 219444 408500 219496
rect 408552 219484 408558 219496
rect 414566 219484 414572 219496
rect 408552 219456 414572 219484
rect 408552 219444 408558 219456
rect 414566 219444 414572 219456
rect 414624 219444 414630 219496
rect 422220 219456 423168 219484
rect 52270 219376 52276 219428
rect 52328 219416 52334 219428
rect 56612 219416 56640 219444
rect 52328 219388 56640 219416
rect 52328 219376 52334 219388
rect 350166 219376 350172 219428
rect 350224 219416 350230 219428
rect 422220 219416 422248 219456
rect 350224 219388 422248 219416
rect 423140 219416 423168 219456
rect 504910 219444 504916 219496
rect 504968 219484 504974 219496
rect 623774 219484 623780 219496
rect 504968 219456 623780 219484
rect 504968 219444 504974 219456
rect 623774 219444 623780 219456
rect 623832 219444 623838 219496
rect 673362 219444 673368 219496
rect 673420 219484 673426 219496
rect 676030 219484 676036 219496
rect 673420 219456 676036 219484
rect 673420 219444 673426 219456
rect 676030 219444 676036 219456
rect 676088 219444 676094 219496
rect 423858 219416 423864 219428
rect 423140 219388 423864 219416
rect 350224 219376 350230 219388
rect 423858 219376 423864 219388
rect 423916 219376 423922 219428
rect 354398 219308 354404 219360
rect 354456 219348 354462 219360
rect 432230 219348 432236 219360
rect 354456 219320 432236 219348
rect 354456 219308 354462 219320
rect 432230 219308 432236 219320
rect 432288 219308 432294 219360
rect 353202 219240 353208 219292
rect 353260 219280 353266 219292
rect 430574 219280 430580 219292
rect 353260 219252 430580 219280
rect 353260 219240 353266 219252
rect 430574 219240 430580 219252
rect 430632 219240 430638 219292
rect 379422 219172 379428 219224
rect 379480 219212 379486 219224
rect 494514 219212 494520 219224
rect 379480 219184 494520 219212
rect 379480 219172 379486 219184
rect 494514 219172 494520 219184
rect 494572 219172 494578 219224
rect 570598 219172 570604 219224
rect 570656 219212 570662 219224
rect 635918 219212 635924 219224
rect 570656 219184 635924 219212
rect 570656 219172 570662 219184
rect 635918 219172 635924 219184
rect 635976 219172 635982 219224
rect 380802 219104 380808 219156
rect 380860 219144 380866 219156
rect 498194 219144 498200 219156
rect 380860 219116 498200 219144
rect 380860 219104 380866 219116
rect 498194 219104 498200 219116
rect 498252 219104 498258 219156
rect 555418 219104 555424 219156
rect 555476 219144 555482 219156
rect 577498 219144 577504 219156
rect 555476 219116 577504 219144
rect 555476 219104 555482 219116
rect 577498 219104 577504 219116
rect 577556 219104 577562 219156
rect 383470 219036 383476 219088
rect 383528 219076 383534 219088
rect 501230 219076 501236 219088
rect 383528 219048 501236 219076
rect 383528 219036 383534 219048
rect 501230 219036 501236 219048
rect 501288 219036 501294 219088
rect 548518 219036 548524 219088
rect 548576 219076 548582 219088
rect 576210 219076 576216 219088
rect 548576 219048 576216 219076
rect 548576 219036 548582 219048
rect 576210 219036 576216 219048
rect 576268 219036 576274 219088
rect 383562 218968 383568 219020
rect 383620 219008 383626 219020
rect 503714 219008 503720 219020
rect 383620 218980 503720 219008
rect 383620 218968 383626 218980
rect 503714 218968 503720 218980
rect 503772 218968 503778 219020
rect 505002 218968 505008 219020
rect 505060 219008 505066 219020
rect 622946 219008 622952 219020
rect 505060 218980 622952 219008
rect 505060 218968 505066 218980
rect 622946 218968 622952 218980
rect 623004 218968 623010 219020
rect 386322 218900 386328 218952
rect 386380 218940 386386 218952
rect 508774 218940 508780 218952
rect 386380 218912 508780 218940
rect 386380 218900 386386 218912
rect 508774 218900 508780 218912
rect 508832 218900 508838 218952
rect 557810 218900 557816 218952
rect 557868 218940 557874 218952
rect 607674 218940 607680 218952
rect 557868 218912 607680 218940
rect 557868 218900 557874 218912
rect 607674 218900 607680 218912
rect 607732 218900 607738 218952
rect 387702 218832 387708 218884
rect 387760 218872 387766 218884
rect 511350 218872 511356 218884
rect 387760 218844 511356 218872
rect 387760 218832 387766 218844
rect 511350 218832 511356 218844
rect 511408 218832 511414 218884
rect 561766 218832 561772 218884
rect 561824 218872 561830 218884
rect 562870 218872 562876 218884
rect 561824 218844 562876 218872
rect 561824 218832 561830 218844
rect 562870 218832 562876 218844
rect 562928 218872 562934 218884
rect 616782 218872 616788 218884
rect 562928 218844 616788 218872
rect 562928 218832 562934 218844
rect 616782 218832 616788 218844
rect 616840 218832 616846 218884
rect 391842 218764 391848 218816
rect 391900 218804 391906 218816
rect 521654 218804 521660 218816
rect 391900 218776 521660 218804
rect 391900 218764 391906 218776
rect 521654 218764 521660 218776
rect 521712 218764 521718 218816
rect 565446 218764 565452 218816
rect 565504 218804 565510 218816
rect 619542 218804 619548 218816
rect 565504 218776 619548 218804
rect 565504 218764 565510 218776
rect 619542 218764 619548 218776
rect 619600 218764 619606 218816
rect 44818 218696 44824 218748
rect 44876 218736 44882 218748
rect 659746 218736 659752 218748
rect 44876 218708 659752 218736
rect 44876 218696 44882 218708
rect 659746 218696 659752 218708
rect 659804 218696 659810 218748
rect 567930 218628 567936 218680
rect 567988 218668 567994 218680
rect 627454 218668 627460 218680
rect 567988 218640 627460 218668
rect 567988 218628 567994 218640
rect 627454 218628 627460 218640
rect 627512 218628 627518 218680
rect 515490 218560 515496 218612
rect 515548 218600 515554 218612
rect 576026 218600 576032 218612
rect 515548 218572 576032 218600
rect 515548 218560 515554 218572
rect 576026 218560 576032 218572
rect 576084 218560 576090 218612
rect 543182 218492 543188 218544
rect 543240 218532 543246 218544
rect 543642 218532 543648 218544
rect 543240 218504 543648 218532
rect 543240 218492 543246 218504
rect 543642 218492 543648 218504
rect 543700 218532 543706 218544
rect 576118 218532 576124 218544
rect 543700 218504 576124 218532
rect 543700 218492 543706 218504
rect 576118 218492 576124 218504
rect 576176 218492 576182 218544
rect 487798 218424 487804 218476
rect 487856 218464 487862 218476
rect 575934 218464 575940 218476
rect 487856 218436 575940 218464
rect 487856 218424 487862 218436
rect 575934 218424 575940 218436
rect 575992 218424 575998 218476
rect 495618 218356 495624 218408
rect 495676 218396 495682 218408
rect 495986 218396 495992 218408
rect 495676 218368 495992 218396
rect 495676 218356 495682 218368
rect 495986 218356 495992 218368
rect 496044 218396 496050 218408
rect 619726 218396 619732 218408
rect 496044 218368 619732 218396
rect 496044 218356 496050 218368
rect 619726 218356 619732 218368
rect 619784 218356 619790 218408
rect 500218 218288 500224 218340
rect 500276 218328 500282 218340
rect 637850 218328 637856 218340
rect 500276 218300 637856 218328
rect 500276 218288 500282 218300
rect 637850 218288 637856 218300
rect 637908 218288 637914 218340
rect 496078 218220 496084 218272
rect 496136 218260 496142 218272
rect 637390 218260 637396 218272
rect 496136 218232 637396 218260
rect 496136 218220 496142 218232
rect 637390 218220 637396 218232
rect 637448 218220 637454 218272
rect 493410 218152 493416 218204
rect 493468 218192 493474 218204
rect 636930 218192 636936 218204
rect 493468 218164 636936 218192
rect 493468 218152 493474 218164
rect 636930 218152 636936 218164
rect 636988 218152 636994 218204
rect 486418 218084 486424 218136
rect 486476 218124 486482 218136
rect 486476 218096 487936 218124
rect 486476 218084 486482 218096
rect 118694 218016 118700 218068
rect 118752 218056 118758 218068
rect 124858 218056 124864 218068
rect 118752 218028 124864 218056
rect 118752 218016 118758 218028
rect 124858 218016 124864 218028
rect 124916 218016 124922 218068
rect 487522 218016 487528 218068
rect 487580 218056 487586 218068
rect 487798 218056 487804 218068
rect 487580 218028 487804 218056
rect 487580 218016 487586 218028
rect 487798 218016 487804 218028
rect 487856 218016 487862 218068
rect 487908 218056 487936 218096
rect 489454 218084 489460 218136
rect 489512 218124 489518 218136
rect 633710 218124 633716 218136
rect 489512 218096 633716 218124
rect 489512 218084 489518 218096
rect 633710 218084 633716 218096
rect 633768 218084 633774 218136
rect 638310 218056 638316 218068
rect 487908 218028 638316 218056
rect 638310 218016 638316 218028
rect 638368 218016 638374 218068
rect 523034 217880 523040 217932
rect 523092 217920 523098 217932
rect 523954 217920 523960 217932
rect 523092 217892 523960 217920
rect 523092 217880 523098 217892
rect 523954 217880 523960 217892
rect 524012 217880 524018 217932
rect 538214 217880 538220 217932
rect 538272 217920 538278 217932
rect 539042 217920 539048 217932
rect 538272 217892 539048 217920
rect 538272 217880 538278 217892
rect 539042 217880 539048 217892
rect 539100 217880 539106 217932
rect 296806 217812 296812 217864
rect 296864 217852 296870 217864
rect 297634 217852 297640 217864
rect 296864 217824 297640 217852
rect 296864 217812 296870 217824
rect 297634 217812 297640 217824
rect 297692 217812 297698 217864
rect 331214 217812 331220 217864
rect 331272 217852 331278 217864
rect 332134 217852 332140 217864
rect 331272 217824 332140 217852
rect 331272 217812 331278 217824
rect 332134 217812 332140 217824
rect 332192 217812 332198 217864
rect 333974 217812 333980 217864
rect 334032 217852 334038 217864
rect 334710 217852 334716 217864
rect 334032 217824 334716 217852
rect 334032 217812 334038 217824
rect 334710 217812 334716 217824
rect 334768 217812 334774 217864
rect 350626 217812 350632 217864
rect 350684 217852 350690 217864
rect 351454 217852 351460 217864
rect 350684 217824 351460 217852
rect 350684 217812 350690 217824
rect 351454 217812 351460 217824
rect 351512 217812 351518 217864
rect 422294 217812 422300 217864
rect 422352 217852 422358 217864
rect 423030 217852 423036 217864
rect 422352 217824 423036 217852
rect 422352 217812 422358 217824
rect 423030 217812 423036 217824
rect 423088 217812 423094 217864
rect 434714 217812 434720 217864
rect 434772 217852 434778 217864
rect 435634 217852 435640 217864
rect 434772 217824 435640 217852
rect 434772 217812 434778 217824
rect 435634 217812 435640 217824
rect 435692 217812 435698 217864
rect 441614 217812 441620 217864
rect 441672 217852 441678 217864
rect 442350 217852 442356 217864
rect 441672 217824 442356 217852
rect 441672 217812 441678 217824
rect 442350 217812 442356 217824
rect 442408 217812 442414 217864
rect 454034 217812 454040 217864
rect 454092 217852 454098 217864
rect 454954 217852 454960 217864
rect 454092 217824 454960 217852
rect 454092 217812 454098 217824
rect 454954 217812 454960 217824
rect 455012 217812 455018 217864
rect 460934 217812 460940 217864
rect 460992 217852 460998 217864
rect 461670 217852 461676 217864
rect 460992 217824 461676 217852
rect 460992 217812 460998 217824
rect 461670 217812 461676 217824
rect 461728 217812 461734 217864
rect 465074 217812 465080 217864
rect 465132 217852 465138 217864
rect 465902 217852 465908 217864
rect 465132 217824 465908 217852
rect 465132 217812 465138 217824
rect 465902 217812 465908 217824
rect 465960 217812 465966 217864
rect 471974 217812 471980 217864
rect 472032 217852 472038 217864
rect 472618 217852 472624 217864
rect 472032 217824 472624 217852
rect 472032 217812 472038 217824
rect 472618 217812 472624 217824
rect 472676 217812 472682 217864
rect 476114 217812 476120 217864
rect 476172 217852 476178 217864
rect 476850 217852 476856 217864
rect 476172 217824 476856 217852
rect 476172 217812 476178 217824
rect 476850 217812 476856 217824
rect 476908 217812 476914 217864
rect 499574 217812 499580 217864
rect 499632 217852 499638 217864
rect 500862 217852 500868 217864
rect 499632 217824 500868 217852
rect 499632 217812 499638 217824
rect 500862 217812 500868 217824
rect 500920 217852 500926 217864
rect 608502 217852 608508 217864
rect 500920 217824 608508 217852
rect 500920 217812 500926 217824
rect 608502 217812 608508 217824
rect 608560 217812 608566 217864
rect 497642 217744 497648 217796
rect 497700 217784 497706 217796
rect 608042 217784 608048 217796
rect 497700 217756 608048 217784
rect 497700 217744 497706 217756
rect 608042 217744 608048 217756
rect 608100 217744 608106 217796
rect 490926 217676 490932 217728
rect 490984 217716 490990 217728
rect 607122 217716 607128 217728
rect 490984 217688 607128 217716
rect 490984 217676 490990 217688
rect 607122 217676 607128 217688
rect 607180 217676 607186 217728
rect 553716 217608 553722 217660
rect 553774 217648 553780 217660
rect 575842 217648 575848 217660
rect 553774 217620 575848 217648
rect 553774 217608 553780 217620
rect 575842 217608 575848 217620
rect 575900 217608 575906 217660
rect 609882 217608 609888 217660
rect 609940 217648 609946 217660
rect 629478 217648 629484 217660
rect 609940 217620 629484 217648
rect 609940 217608 609946 217620
rect 629478 217608 629484 217620
rect 629536 217608 629542 217660
rect 568804 217540 568810 217592
rect 568862 217580 568868 217592
rect 618346 217580 618352 217592
rect 568862 217552 618352 217580
rect 568862 217540 568868 217552
rect 618346 217540 618352 217552
rect 618404 217540 618410 217592
rect 556154 217472 556160 217524
rect 556212 217512 556218 217524
rect 618714 217512 618720 217524
rect 556212 217484 618720 217512
rect 556212 217472 556218 217484
rect 618714 217472 618720 217484
rect 618772 217472 618778 217524
rect 549622 217404 549628 217456
rect 549680 217444 549686 217456
rect 550542 217444 550548 217456
rect 549680 217416 550548 217444
rect 549680 217404 549686 217416
rect 550542 217404 550548 217416
rect 550600 217444 550606 217456
rect 632238 217444 632244 217456
rect 550600 217416 632244 217444
rect 550600 217404 550606 217416
rect 632238 217404 632244 217416
rect 632296 217404 632302 217456
rect 494330 217336 494336 217388
rect 494388 217376 494394 217388
rect 578142 217376 578148 217388
rect 494388 217348 578148 217376
rect 494388 217336 494394 217348
rect 578142 217336 578148 217348
rect 578200 217336 578206 217388
rect 609606 217336 609612 217388
rect 609664 217376 609670 217388
rect 632698 217376 632704 217388
rect 609664 217348 632704 217376
rect 609664 217336 609670 217348
rect 632698 217336 632704 217348
rect 632756 217336 632762 217388
rect 35802 217268 35808 217320
rect 35860 217308 35866 217320
rect 43806 217308 43812 217320
rect 35860 217280 43812 217308
rect 35860 217268 35866 217280
rect 43806 217268 43812 217280
rect 43864 217268 43870 217320
rect 545574 217268 545580 217320
rect 545632 217308 545638 217320
rect 631318 217308 631324 217320
rect 545632 217280 631324 217308
rect 545632 217268 545638 217280
rect 631318 217268 631324 217280
rect 631376 217268 631382 217320
rect 537938 217200 537944 217252
rect 537996 217240 538002 217252
rect 629938 217240 629944 217252
rect 537996 217212 629944 217240
rect 537996 217200 538002 217212
rect 629938 217200 629944 217212
rect 629996 217200 630002 217252
rect 513650 217132 513656 217184
rect 513708 217172 513714 217184
rect 610802 217172 610808 217184
rect 513708 217144 610808 217172
rect 513708 217132 513714 217144
rect 610802 217132 610808 217144
rect 610860 217132 610866 217184
rect 511074 217064 511080 217116
rect 511132 217104 511138 217116
rect 610342 217104 610348 217116
rect 511132 217076 610348 217104
rect 511132 217064 511138 217076
rect 610342 217064 610348 217076
rect 610400 217064 610406 217116
rect 508498 216996 508504 217048
rect 508556 217036 508562 217048
rect 609882 217036 609888 217048
rect 508556 217008 609888 217036
rect 508556 216996 508562 217008
rect 609882 216996 609888 217008
rect 609940 216996 609946 217048
rect 506106 216928 506112 216980
rect 506164 216968 506170 216980
rect 609422 216968 609428 216980
rect 506164 216940 609428 216968
rect 506164 216928 506170 216940
rect 609422 216928 609428 216940
rect 609480 216928 609486 216980
rect 502518 216860 502524 216912
rect 502576 216900 502582 216912
rect 503530 216900 503536 216912
rect 502576 216872 503536 216900
rect 502576 216860 502582 216872
rect 503530 216860 503536 216872
rect 503588 216900 503594 216912
rect 608962 216900 608968 216912
rect 503588 216872 608968 216900
rect 503588 216860 503594 216872
rect 608962 216860 608968 216872
rect 609020 216860 609026 216912
rect 564066 216792 564072 216844
rect 564124 216832 564130 216844
rect 577038 216832 577044 216844
rect 564124 216804 577044 216832
rect 564124 216792 564130 216804
rect 577038 216792 577044 216804
rect 577096 216792 577102 216844
rect 561398 216724 561404 216776
rect 561456 216764 561462 216776
rect 575750 216764 575756 216776
rect 561456 216736 575756 216764
rect 561456 216724 561462 216736
rect 575750 216724 575756 216736
rect 575808 216724 575814 216776
rect 558914 216656 558920 216708
rect 558972 216696 558978 216708
rect 575658 216696 575664 216708
rect 558972 216668 575664 216696
rect 558972 216656 558978 216668
rect 575658 216656 575664 216668
rect 575716 216656 575722 216708
rect 550606 216464 569954 216492
rect 118694 216424 118700 216436
rect 103486 216396 118700 216424
rect 52178 215908 52184 215960
rect 52236 215948 52242 215960
rect 103486 215948 103514 216396
rect 118694 216384 118700 216396
rect 118752 216384 118758 216436
rect 518710 216384 518716 216436
rect 518768 216424 518774 216436
rect 518768 216396 518894 216424
rect 518768 216384 518774 216396
rect 52236 215920 103514 215948
rect 52236 215908 52242 215920
rect 518866 215336 518894 216396
rect 521194 216384 521200 216436
rect 521252 216424 521258 216436
rect 521252 216396 523356 216424
rect 521252 216384 521258 216396
rect 523328 215404 523356 216396
rect 523770 216384 523776 216436
rect 523828 216424 523834 216436
rect 523828 216396 525104 216424
rect 523828 216384 523834 216396
rect 525076 215472 525104 216396
rect 526254 216384 526260 216436
rect 526312 216424 526318 216436
rect 526312 216396 526806 216424
rect 526312 216384 526318 216396
rect 526778 215540 526806 216396
rect 528554 216384 528560 216436
rect 528612 216424 528618 216436
rect 528612 216396 528692 216424
rect 528612 216384 528618 216396
rect 528664 215608 528692 216396
rect 531222 216384 531228 216436
rect 531280 216424 531286 216436
rect 531280 216396 533292 216424
rect 531280 216384 531286 216396
rect 533264 215676 533292 216396
rect 533798 216384 533804 216436
rect 533856 216424 533862 216436
rect 533856 216396 534856 216424
rect 533856 216384 533862 216396
rect 534828 215744 534856 216396
rect 536374 216384 536380 216436
rect 536432 216424 536438 216436
rect 536432 216396 538214 216424
rect 536432 216384 536438 216396
rect 538186 215812 538214 216396
rect 538858 216384 538864 216436
rect 538916 216384 538922 216436
rect 541434 216384 541440 216436
rect 541492 216424 541498 216436
rect 541492 216396 548012 216424
rect 541492 216384 541498 216396
rect 538876 216356 538904 216384
rect 538876 216328 547874 216356
rect 547846 215880 547874 216328
rect 547984 216084 548012 216396
rect 550606 216084 550634 216464
rect 551462 216384 551468 216436
rect 551520 216424 551526 216436
rect 551520 216396 560294 216424
rect 551520 216384 551526 216396
rect 547984 216056 550634 216084
rect 560266 216016 560294 216396
rect 566458 216384 566464 216436
rect 566516 216384 566522 216436
rect 566476 216016 566504 216384
rect 569926 216152 569954 216464
rect 574830 216384 574836 216436
rect 574888 216384 574894 216436
rect 574922 216384 574928 216436
rect 574980 216424 574986 216436
rect 574980 216396 576854 216424
rect 574980 216384 574986 216396
rect 574848 216152 574876 216384
rect 576826 216220 576854 216396
rect 613010 216316 613016 216368
rect 613068 216356 613074 216368
rect 630398 216356 630404 216368
rect 613068 216328 630404 216356
rect 613068 216316 613074 216328
rect 630398 216316 630404 216328
rect 630456 216316 630462 216368
rect 614114 216248 614120 216300
rect 614172 216288 614178 216300
rect 631778 216288 631784 216300
rect 614172 216260 631784 216288
rect 614172 216248 614178 216260
rect 631778 216248 631784 216260
rect 631836 216248 631842 216300
rect 626626 216220 626632 216232
rect 576826 216192 626632 216220
rect 626626 216180 626632 216192
rect 626684 216180 626690 216232
rect 628466 216152 628472 216164
rect 569926 216124 572714 216152
rect 574848 216124 628472 216152
rect 572686 216084 572714 216124
rect 628466 216112 628472 216124
rect 628524 216112 628530 216164
rect 672994 216112 673000 216164
rect 673052 216152 673058 216164
rect 676030 216152 676036 216164
rect 673052 216124 676036 216152
rect 673052 216112 673058 216124
rect 676030 216112 676036 216124
rect 676088 216112 676094 216164
rect 577866 216084 577872 216096
rect 572686 216056 577872 216084
rect 577866 216044 577872 216056
rect 577924 216044 577930 216096
rect 611722 216044 611728 216096
rect 611780 216084 611786 216096
rect 630858 216084 630864 216096
rect 611780 216056 630864 216084
rect 611780 216044 611786 216056
rect 630858 216044 630864 216056
rect 630916 216044 630922 216096
rect 620554 216016 620560 216028
rect 560266 215988 563054 216016
rect 566476 215988 620560 216016
rect 563026 215948 563054 215988
rect 620554 215976 620560 215988
rect 620612 215976 620618 216028
rect 563026 215920 617104 215948
rect 615494 215880 615500 215892
rect 547846 215852 615500 215880
rect 615494 215840 615500 215852
rect 615552 215840 615558 215892
rect 617076 215880 617104 215920
rect 617150 215908 617156 215960
rect 617208 215948 617214 215960
rect 634078 215948 634084 215960
rect 617208 215920 634084 215948
rect 617208 215908 617214 215920
rect 634078 215908 634084 215920
rect 634136 215908 634142 215960
rect 617794 215880 617800 215892
rect 617076 215852 617800 215880
rect 617794 215840 617800 215852
rect 617852 215840 617858 215892
rect 615034 215812 615040 215824
rect 538186 215784 615040 215812
rect 615034 215772 615040 215784
rect 615092 215772 615098 215824
rect 614574 215744 614580 215756
rect 534828 215716 614580 215744
rect 614574 215704 614580 215716
rect 614632 215704 614638 215756
rect 674558 215704 674564 215756
rect 674616 215744 674622 215756
rect 676030 215744 676036 215756
rect 674616 215716 676036 215744
rect 674616 215704 674622 215716
rect 676030 215704 676036 215716
rect 676088 215704 676094 215756
rect 614022 215676 614028 215688
rect 533264 215648 614028 215676
rect 614022 215636 614028 215648
rect 614080 215636 614086 215688
rect 613562 215608 613568 215620
rect 528664 215580 613568 215608
rect 613562 215568 613568 215580
rect 613620 215568 613626 215620
rect 613102 215540 613108 215552
rect 526778 215512 613108 215540
rect 613102 215500 613108 215512
rect 613160 215500 613166 215552
rect 676214 215500 676220 215552
rect 676272 215540 676278 215552
rect 676858 215540 676864 215552
rect 676272 215512 676864 215540
rect 676272 215500 676278 215512
rect 676858 215500 676864 215512
rect 676916 215500 676922 215552
rect 612642 215472 612648 215484
rect 525076 215444 612648 215472
rect 612642 215432 612648 215444
rect 612700 215432 612706 215484
rect 612182 215404 612188 215416
rect 523328 215376 612188 215404
rect 612182 215364 612188 215376
rect 612240 215364 612246 215416
rect 611722 215336 611728 215348
rect 518866 215308 611728 215336
rect 611722 215296 611728 215308
rect 611780 215296 611786 215348
rect 51356 215022 576186 215050
rect 35802 214548 35808 214600
rect 35860 214588 35866 214600
rect 46198 214588 46204 214600
rect 35860 214560 46204 214588
rect 35860 214548 35866 214560
rect 46198 214548 46204 214560
rect 46256 214548 46262 214600
rect 50338 214344 50344 214396
rect 50396 214384 50402 214396
rect 51356 214384 51384 215022
rect 50396 214356 51384 214384
rect 51424 214954 576118 214982
rect 50396 214344 50402 214356
rect 50062 214276 50068 214328
rect 50120 214316 50126 214328
rect 51424 214316 51452 214954
rect 50120 214288 51452 214316
rect 51492 214886 576050 214914
rect 50120 214276 50126 214288
rect 47210 214208 47216 214260
rect 47268 214248 47274 214260
rect 51492 214248 51520 214886
rect 47268 214220 51520 214248
rect 51560 214818 575982 214846
rect 47268 214208 47274 214220
rect 41322 214140 41328 214192
rect 41380 214180 41386 214192
rect 51560 214180 51588 214818
rect 41380 214152 51588 214180
rect 51628 214750 575914 214778
rect 41380 214140 41386 214152
rect 31110 214072 31116 214124
rect 31168 214112 31174 214124
rect 51628 214112 51656 214750
rect 31168 214084 51656 214112
rect 51696 214682 575846 214710
rect 31168 214072 31174 214084
rect 31294 214004 31300 214056
rect 31352 214044 31358 214056
rect 51696 214044 51724 214682
rect 31352 214016 51724 214044
rect 51764 214614 575778 214642
rect 31352 214004 31358 214016
rect 41506 213936 41512 213988
rect 41564 213976 41570 213988
rect 51764 213976 51792 214614
rect 41564 213948 51792 213976
rect 575750 213976 575778 214614
rect 575818 214044 575846 214682
rect 575886 214112 575914 214750
rect 575954 214180 575982 214818
rect 576022 214248 576050 214886
rect 576090 214316 576118 214954
rect 576158 214384 576186 215022
rect 576394 214752 576400 214804
rect 576452 214792 576458 214804
rect 626166 214792 626172 214804
rect 576452 214764 626172 214792
rect 576452 214752 576458 214764
rect 626166 214752 626172 214764
rect 626224 214752 626230 214804
rect 577130 214684 577136 214736
rect 577188 214724 577194 214736
rect 627546 214724 627552 214736
rect 577188 214696 627552 214724
rect 577188 214684 577194 214696
rect 627546 214684 627552 214696
rect 627604 214684 627610 214736
rect 577314 214616 577320 214668
rect 577372 214656 577378 214668
rect 627086 214656 627092 214668
rect 577372 214628 627092 214656
rect 577372 214616 577378 214628
rect 627086 214616 627092 214628
rect 627144 214616 627150 214668
rect 576302 214548 576308 214600
rect 576360 214588 576366 214600
rect 628006 214588 628012 214600
rect 576360 214560 628012 214588
rect 576360 214548 576366 214560
rect 628006 214548 628012 214560
rect 628064 214548 628070 214600
rect 662506 214548 662512 214600
rect 662564 214588 662570 214600
rect 663058 214588 663064 214600
rect 662564 214560 663064 214588
rect 662564 214548 662570 214560
rect 663058 214548 663064 214560
rect 663116 214548 663122 214600
rect 663794 214548 663800 214600
rect 663852 214588 663858 214600
rect 664438 214588 664444 214600
rect 663852 214560 664444 214588
rect 663852 214548 663858 214560
rect 664438 214548 664444 214560
rect 664496 214548 664502 214600
rect 623866 214480 623872 214532
rect 623924 214520 623930 214532
rect 624418 214520 624424 214532
rect 623924 214492 624424 214520
rect 623924 214480 623930 214492
rect 624418 214480 624424 214492
rect 624476 214480 624482 214532
rect 665266 214384 665272 214396
rect 576158 214356 665272 214384
rect 665266 214344 665272 214356
rect 665324 214344 665330 214396
rect 668854 214316 668860 214328
rect 576090 214288 668860 214316
rect 668854 214276 668860 214288
rect 668912 214276 668918 214328
rect 668118 214248 668124 214260
rect 576022 214220 668124 214248
rect 668118 214208 668124 214220
rect 668176 214208 668182 214260
rect 668946 214180 668952 214192
rect 575954 214152 668952 214180
rect 668946 214140 668952 214152
rect 669004 214140 669010 214192
rect 665726 214112 665732 214124
rect 575886 214084 665732 214112
rect 665726 214072 665732 214084
rect 665784 214072 665790 214124
rect 673178 214072 673184 214124
rect 673236 214112 673242 214124
rect 676030 214112 676036 214124
rect 673236 214084 676036 214112
rect 673236 214072 673242 214084
rect 676030 214072 676036 214084
rect 676088 214072 676094 214124
rect 666186 214044 666192 214056
rect 575818 214016 666192 214044
rect 666186 214004 666192 214016
rect 666244 214004 666250 214056
rect 669038 213976 669044 213988
rect 575750 213948 669044 213976
rect 41564 213936 41570 213948
rect 669038 213936 669044 213948
rect 669096 213936 669102 213988
rect 575934 213868 575940 213920
rect 575992 213908 575998 213920
rect 606662 213908 606668 213920
rect 575992 213880 606668 213908
rect 575992 213868 575998 213880
rect 606662 213868 606668 213880
rect 606720 213868 606726 213920
rect 607674 213868 607680 213920
rect 607732 213908 607738 213920
rect 633618 213908 633624 213920
rect 607732 213880 633624 213908
rect 607732 213868 607738 213880
rect 633618 213868 633624 213880
rect 633676 213868 633682 213920
rect 633710 213868 633716 213920
rect 633768 213908 633774 213920
rect 636378 213908 636384 213920
rect 633768 213880 636384 213908
rect 633768 213868 633774 213880
rect 636378 213868 636384 213880
rect 636436 213868 636442 213920
rect 636838 213868 636844 213920
rect 636896 213908 636902 213920
rect 639230 213908 639236 213920
rect 636896 213880 639236 213908
rect 636896 213868 636902 213880
rect 639230 213868 639236 213880
rect 639288 213868 639294 213920
rect 639598 213868 639604 213920
rect 639656 213908 639662 213920
rect 640610 213908 640616 213920
rect 639656 213880 640616 213908
rect 639656 213868 639662 213880
rect 640610 213868 640616 213880
rect 640668 213868 640674 213920
rect 576026 213800 576032 213852
rect 576084 213840 576090 213852
rect 611262 213840 611268 213852
rect 576084 213812 611268 213840
rect 576084 213800 576090 213812
rect 611262 213800 611268 213812
rect 611320 213800 611326 213852
rect 619726 213800 619732 213852
rect 619784 213840 619790 213852
rect 622486 213840 622492 213852
rect 619784 213812 622492 213840
rect 619784 213800 619790 213812
rect 622486 213800 622492 213812
rect 622544 213800 622550 213852
rect 577866 213732 577872 213784
rect 577924 213772 577930 213784
rect 615954 213772 615960 213784
rect 577924 213744 615960 213772
rect 577924 213732 577930 213744
rect 615954 213732 615960 213744
rect 616012 213732 616018 213784
rect 576118 213664 576124 213716
rect 576176 213704 576182 213716
rect 616414 213704 616420 213716
rect 576176 213676 616420 213704
rect 576176 213664 576182 213676
rect 616414 213664 616420 213676
rect 616472 213664 616478 213716
rect 616782 213664 616788 213716
rect 616840 213704 616846 213716
rect 634538 213704 634544 213716
rect 616840 213676 634544 213704
rect 616840 213664 616846 213676
rect 634538 213664 634544 213676
rect 634596 213664 634602 213716
rect 673086 213664 673092 213716
rect 673144 213704 673150 213716
rect 676030 213704 676036 213716
rect 673144 213676 676036 213704
rect 673144 213664 673150 213676
rect 676030 213664 676036 213676
rect 676088 213664 676094 213716
rect 576210 213596 576216 213648
rect 576268 213636 576274 213648
rect 617334 213636 617340 213648
rect 576268 213608 617340 213636
rect 576268 213596 576274 213608
rect 617334 213596 617340 213608
rect 617392 213596 617398 213648
rect 576486 213528 576492 213580
rect 576544 213568 576550 213580
rect 616874 213568 616880 213580
rect 576544 213540 616880 213568
rect 576544 213528 576550 213540
rect 616874 213528 616880 213540
rect 616932 213528 616938 213580
rect 575842 213460 575848 213512
rect 575900 213500 575906 213512
rect 618254 213500 618260 213512
rect 575900 213472 618260 213500
rect 575900 213460 575906 213472
rect 618254 213460 618260 213472
rect 618312 213460 618318 213512
rect 577038 213392 577044 213444
rect 577096 213432 577102 213444
rect 620094 213432 620100 213444
rect 577096 213404 620100 213432
rect 577096 213392 577102 213404
rect 620094 213392 620100 213404
rect 620152 213392 620158 213444
rect 627454 213392 627460 213444
rect 627512 213432 627518 213444
rect 635458 213432 635464 213444
rect 627512 213404 635464 213432
rect 627512 213392 627518 213404
rect 635458 213392 635464 213404
rect 635516 213392 635522 213444
rect 575658 213324 575664 213376
rect 575716 213364 575722 213376
rect 619174 213364 619180 213376
rect 575716 213336 619180 213364
rect 575716 213324 575722 213336
rect 619174 213324 619180 213336
rect 619232 213324 619238 213376
rect 619542 213324 619548 213376
rect 619600 213364 619606 213376
rect 634998 213364 635004 213376
rect 619600 213336 635004 213364
rect 619600 213324 619606 213336
rect 634998 213324 635004 213336
rect 635056 213324 635062 213376
rect 575750 213256 575756 213308
rect 575808 213296 575814 213308
rect 619634 213296 619640 213308
rect 575808 213268 619640 213296
rect 575808 213256 575814 213268
rect 619634 213256 619640 213268
rect 619692 213256 619698 213308
rect 621658 213256 621664 213308
rect 621716 213296 621722 213308
rect 641070 213296 641076 213308
rect 621716 213268 641076 213296
rect 621716 213256 621722 213268
rect 641070 213256 641076 213268
rect 641128 213256 641134 213308
rect 643830 213256 643836 213308
rect 643888 213296 643894 213308
rect 651466 213296 651472 213308
rect 643888 213268 651472 213296
rect 643888 213256 643894 213268
rect 651466 213256 651472 213268
rect 651524 213256 651530 213308
rect 577498 213188 577504 213240
rect 577556 213228 577562 213240
rect 633158 213228 633164 213240
rect 577556 213200 633164 213228
rect 577556 213188 577562 213200
rect 633158 213188 633164 213200
rect 633216 213188 633222 213240
rect 642726 213188 642732 213240
rect 642784 213228 642790 213240
rect 650086 213228 650092 213240
rect 642784 213200 650092 213228
rect 642784 213188 642790 213200
rect 650086 213188 650092 213200
rect 650144 213188 650150 213240
rect 578142 213120 578148 213172
rect 578200 213160 578206 213172
rect 607582 213160 607588 213172
rect 578200 213132 607588 213160
rect 578200 213120 578206 213132
rect 607582 213120 607588 213132
rect 607640 213120 607646 213172
rect 645578 213120 645584 213172
rect 645636 213160 645642 213172
rect 649994 213160 650000 213172
rect 645636 213132 650000 213160
rect 645636 213120 645642 213132
rect 649994 213120 650000 213132
rect 650052 213120 650058 213172
rect 646958 212984 646964 213036
rect 647016 213024 647022 213036
rect 651374 213024 651380 213036
rect 647016 212996 651380 213024
rect 647016 212984 647022 212996
rect 651374 212984 651380 212996
rect 651432 212984 651438 213036
rect 618346 212508 618352 212560
rect 618404 212548 618410 212560
rect 621014 212548 621020 212560
rect 618404 212520 621020 212548
rect 618404 212508 618410 212520
rect 621014 212508 621020 212520
rect 621072 212508 621078 212560
rect 583018 211148 583024 211200
rect 583076 211188 583082 211200
rect 638770 211188 638776 211200
rect 583076 211160 638776 211188
rect 583076 211148 583082 211160
rect 638770 211148 638776 211160
rect 638828 211148 638834 211200
rect 670326 211148 670332 211200
rect 670384 211188 670390 211200
rect 676030 211188 676036 211200
rect 670384 211160 676036 211188
rect 670384 211148 670390 211160
rect 676030 211148 676036 211160
rect 676088 211148 676094 211200
rect 652018 210400 652024 210452
rect 652076 210440 652082 210452
rect 667198 210440 667204 210452
rect 652076 210412 667204 210440
rect 652076 210400 652082 210412
rect 667198 210400 667204 210412
rect 667256 210400 667262 210452
rect 639046 210060 639052 210112
rect 639104 210100 639110 210112
rect 639782 210100 639788 210112
rect 639104 210072 639788 210100
rect 639104 210060 639110 210072
rect 639782 210060 639788 210072
rect 639840 210060 639846 210112
rect 578878 209720 578884 209772
rect 578936 209760 578942 209772
rect 603074 209760 603080 209772
rect 578936 209732 603080 209760
rect 578936 209720 578942 209732
rect 603074 209720 603080 209732
rect 603132 209720 603138 209772
rect 579246 209652 579252 209704
rect 579304 209692 579310 209704
rect 603166 209692 603172 209704
rect 579304 209664 603172 209692
rect 579304 209652 579310 209664
rect 603166 209652 603172 209664
rect 603224 209652 603230 209704
rect 578970 208292 578976 208344
rect 579028 208332 579034 208344
rect 603074 208332 603080 208344
rect 579028 208304 603080 208332
rect 579028 208292 579034 208304
rect 603074 208292 603080 208304
rect 603132 208292 603138 208344
rect 578418 206932 578424 206984
rect 578476 206972 578482 206984
rect 603074 206972 603080 206984
rect 578476 206944 603080 206972
rect 578476 206932 578482 206944
rect 603074 206932 603080 206944
rect 603132 206932 603138 206984
rect 578510 205572 578516 205624
rect 578568 205612 578574 205624
rect 603074 205612 603080 205624
rect 578568 205584 603080 205612
rect 578568 205572 578574 205584
rect 603074 205572 603080 205584
rect 603132 205572 603138 205624
rect 579522 205504 579528 205556
rect 579580 205544 579586 205556
rect 603166 205544 603172 205556
rect 579580 205516 603172 205544
rect 579580 205504 579586 205516
rect 603166 205504 603172 205516
rect 603224 205504 603230 205556
rect 578786 204212 578792 204264
rect 578844 204252 578850 204264
rect 603074 204252 603080 204264
rect 578844 204224 603080 204252
rect 578844 204212 578850 204224
rect 603074 204212 603080 204224
rect 603132 204212 603138 204264
rect 35802 202852 35808 202904
rect 35860 202892 35866 202904
rect 50338 202892 50344 202904
rect 35860 202864 50344 202892
rect 35860 202852 35866 202864
rect 50338 202852 50344 202864
rect 50396 202852 50402 202904
rect 579430 202784 579436 202836
rect 579488 202824 579494 202836
rect 603074 202824 603080 202836
rect 579488 202796 603080 202824
rect 579488 202784 579494 202796
rect 603074 202784 603080 202796
rect 603132 202784 603138 202836
rect 672994 201832 673000 201884
rect 673052 201872 673058 201884
rect 675386 201872 675392 201884
rect 673052 201844 675392 201872
rect 673052 201832 673058 201844
rect 675386 201832 675392 201844
rect 675444 201832 675450 201884
rect 578878 201424 578884 201476
rect 578936 201464 578942 201476
rect 603074 201464 603080 201476
rect 578936 201436 603080 201464
rect 578936 201424 578942 201436
rect 603074 201424 603080 201436
rect 603132 201424 603138 201476
rect 674558 201424 674564 201476
rect 674616 201464 674622 201476
rect 675386 201464 675392 201476
rect 674616 201436 675392 201464
rect 674616 201424 674622 201436
rect 675386 201424 675392 201436
rect 675444 201424 675450 201476
rect 579246 201356 579252 201408
rect 579304 201396 579310 201408
rect 603166 201396 603172 201408
rect 579304 201368 603172 201396
rect 579304 201356 579310 201368
rect 603166 201356 603172 201368
rect 603224 201356 603230 201408
rect 675110 200676 675116 200728
rect 675168 200716 675174 200728
rect 675386 200716 675392 200728
rect 675168 200688 675392 200716
rect 675168 200676 675174 200688
rect 675386 200676 675392 200688
rect 675444 200676 675450 200728
rect 578234 200064 578240 200116
rect 578292 200104 578298 200116
rect 603074 200104 603080 200116
rect 578292 200076 603080 200104
rect 578292 200064 578298 200076
rect 603074 200064 603080 200076
rect 603132 200064 603138 200116
rect 578418 198636 578424 198688
rect 578476 198676 578482 198688
rect 603074 198676 603080 198688
rect 578476 198648 603080 198676
rect 578476 198636 578482 198648
rect 603074 198636 603080 198648
rect 603132 198636 603138 198688
rect 673178 197412 673184 197464
rect 673236 197452 673242 197464
rect 675478 197452 675484 197464
rect 673236 197424 675484 197452
rect 673236 197412 673242 197424
rect 675478 197412 675484 197424
rect 675536 197412 675542 197464
rect 579062 197276 579068 197328
rect 579120 197316 579126 197328
rect 603166 197316 603172 197328
rect 579120 197288 603172 197316
rect 579120 197276 579126 197288
rect 603166 197276 603172 197288
rect 603224 197276 603230 197328
rect 674834 197004 674840 197056
rect 674892 197044 674898 197056
rect 675386 197044 675392 197056
rect 674892 197016 675392 197044
rect 674892 197004 674898 197016
rect 675386 197004 675392 197016
rect 675444 197004 675450 197056
rect 579522 196596 579528 196648
rect 579580 196636 579586 196648
rect 603074 196636 603080 196648
rect 579580 196608 603080 196636
rect 579580 196596 579586 196608
rect 603074 196596 603080 196608
rect 603132 196596 603138 196648
rect 673086 196528 673092 196580
rect 673144 196568 673150 196580
rect 675386 196568 675392 196580
rect 673144 196540 675392 196568
rect 673144 196528 673150 196540
rect 675386 196528 675392 196540
rect 675444 196528 675450 196580
rect 579522 195236 579528 195288
rect 579580 195276 579586 195288
rect 603074 195276 603080 195288
rect 579580 195248 603080 195276
rect 579580 195236 579586 195248
rect 603074 195236 603080 195248
rect 603132 195236 603138 195288
rect 579522 193808 579528 193860
rect 579580 193848 579586 193860
rect 603074 193848 603080 193860
rect 579580 193820 603080 193848
rect 579580 193808 579586 193820
rect 603074 193808 603080 193820
rect 603132 193808 603138 193860
rect 42058 193128 42064 193180
rect 42116 193168 42122 193180
rect 43346 193168 43352 193180
rect 42116 193140 43352 193168
rect 42116 193128 42122 193140
rect 43346 193128 43352 193140
rect 43404 193128 43410 193180
rect 579522 192448 579528 192500
rect 579580 192488 579586 192500
rect 603074 192488 603080 192500
rect 579580 192460 603080 192488
rect 579580 192448 579586 192460
rect 603074 192448 603080 192460
rect 603132 192448 603138 192500
rect 674834 192448 674840 192500
rect 674892 192488 674898 192500
rect 675386 192488 675392 192500
rect 674892 192460 675392 192488
rect 674892 192448 674898 192460
rect 675386 192448 675392 192460
rect 675444 192448 675450 192500
rect 579246 191836 579252 191888
rect 579304 191876 579310 191888
rect 603074 191876 603080 191888
rect 579304 191848 603080 191876
rect 579304 191836 579310 191848
rect 603074 191836 603080 191848
rect 603132 191836 603138 191888
rect 42150 191632 42156 191684
rect 42208 191672 42214 191684
rect 43254 191672 43260 191684
rect 42208 191644 43260 191672
rect 42208 191632 42214 191644
rect 43254 191632 43260 191644
rect 43312 191632 43318 191684
rect 42058 191428 42064 191480
rect 42116 191468 42122 191480
rect 43162 191468 43168 191480
rect 42116 191440 43168 191468
rect 42116 191428 42122 191440
rect 43162 191428 43168 191440
rect 43220 191428 43226 191480
rect 42150 190816 42156 190868
rect 42208 190856 42214 190868
rect 43438 190856 43444 190868
rect 42208 190828 43444 190856
rect 42208 190816 42214 190828
rect 43438 190816 43444 190828
rect 43496 190816 43502 190868
rect 675754 190612 675760 190664
rect 675812 190612 675818 190664
rect 578234 190476 578240 190528
rect 578292 190516 578298 190528
rect 603074 190516 603080 190528
rect 578292 190488 603080 190516
rect 578292 190476 578298 190488
rect 603074 190476 603080 190488
rect 603132 190476 603138 190528
rect 675772 190392 675800 190612
rect 675754 190340 675760 190392
rect 675812 190340 675818 190392
rect 579522 189116 579528 189168
rect 579580 189156 579586 189168
rect 603074 189156 603080 189168
rect 579580 189128 603080 189156
rect 579580 189116 579586 189128
rect 603074 189116 603080 189128
rect 603132 189116 603138 189168
rect 579246 189048 579252 189100
rect 579304 189088 579310 189100
rect 603166 189088 603172 189100
rect 579304 189060 603172 189088
rect 579304 189048 579310 189060
rect 603166 189048 603172 189060
rect 603224 189048 603230 189100
rect 578878 187688 578884 187740
rect 578936 187728 578942 187740
rect 603074 187728 603080 187740
rect 578936 187700 603080 187728
rect 578936 187688 578942 187700
rect 603074 187688 603080 187700
rect 603132 187688 603138 187740
rect 42150 187620 42156 187672
rect 42208 187660 42214 187672
rect 42978 187660 42984 187672
rect 42208 187632 42984 187660
rect 42208 187620 42214 187632
rect 42978 187620 42984 187632
rect 43036 187620 43042 187672
rect 579430 186328 579436 186380
rect 579488 186368 579494 186380
rect 603074 186368 603080 186380
rect 579488 186340 603080 186368
rect 579488 186328 579494 186340
rect 603074 186328 603080 186340
rect 603132 186328 603138 186380
rect 42058 186260 42064 186312
rect 42116 186300 42122 186312
rect 42886 186300 42892 186312
rect 42116 186272 42892 186300
rect 42116 186260 42122 186272
rect 42886 186260 42892 186272
rect 42944 186260 42950 186312
rect 42150 185852 42156 185904
rect 42208 185892 42214 185904
rect 42794 185892 42800 185904
rect 42208 185864 42800 185892
rect 42208 185852 42214 185864
rect 42794 185852 42800 185864
rect 42852 185852 42858 185904
rect 579522 184968 579528 185020
rect 579580 185008 579586 185020
rect 603166 185008 603172 185020
rect 579580 184980 603172 185008
rect 579580 184968 579586 184980
rect 603166 184968 603172 184980
rect 603224 184968 603230 185020
rect 578970 184900 578976 184952
rect 579028 184940 579034 184952
rect 603074 184940 603080 184952
rect 579028 184912 603080 184940
rect 579028 184900 579034 184912
rect 603074 184900 603080 184912
rect 603132 184900 603138 184952
rect 667934 183880 667940 183932
rect 667992 183920 667998 183932
rect 669958 183920 669964 183932
rect 667992 183892 669964 183920
rect 667992 183880 667998 183892
rect 669958 183880 669964 183892
rect 670016 183880 670022 183932
rect 579338 183540 579344 183592
rect 579396 183580 579402 183592
rect 603074 183580 603080 183592
rect 579396 183552 603080 183580
rect 579396 183540 579402 183552
rect 603074 183540 603080 183552
rect 603132 183540 603138 183592
rect 42150 183404 42156 183456
rect 42208 183444 42214 183456
rect 44174 183444 44180 183456
rect 42208 183416 44180 183444
rect 42208 183404 42214 183416
rect 44174 183404 44180 183416
rect 44232 183404 44238 183456
rect 578234 182180 578240 182232
rect 578292 182220 578298 182232
rect 603074 182220 603080 182232
rect 578292 182192 603080 182220
rect 578292 182180 578298 182192
rect 603074 182180 603080 182192
rect 603132 182180 603138 182232
rect 578326 180888 578332 180940
rect 578384 180928 578390 180940
rect 603166 180928 603172 180940
rect 578384 180900 603172 180928
rect 578384 180888 578390 180900
rect 603166 180888 603172 180900
rect 603224 180888 603230 180940
rect 578418 180820 578424 180872
rect 578476 180860 578482 180872
rect 603074 180860 603080 180872
rect 578476 180832 603080 180860
rect 578476 180820 578482 180832
rect 603074 180820 603080 180832
rect 603132 180820 603138 180872
rect 578786 179392 578792 179444
rect 578844 179432 578850 179444
rect 603074 179432 603080 179444
rect 578844 179404 603080 179432
rect 578844 179392 578850 179404
rect 603074 179392 603080 179404
rect 603132 179392 603138 179444
rect 667934 178780 667940 178832
rect 667992 178820 667998 178832
rect 670050 178820 670056 178832
rect 667992 178792 670056 178820
rect 667992 178780 667998 178792
rect 670050 178780 670056 178792
rect 670108 178780 670114 178832
rect 671522 178304 671528 178356
rect 671580 178344 671586 178356
rect 676030 178344 676036 178356
rect 671580 178316 676036 178344
rect 671580 178304 671586 178316
rect 676030 178304 676036 178316
rect 676088 178304 676094 178356
rect 668762 178168 668768 178220
rect 668820 178208 668826 178220
rect 675938 178208 675944 178220
rect 668820 178180 675944 178208
rect 668820 178168 668826 178180
rect 675938 178168 675944 178180
rect 675996 178168 676002 178220
rect 578694 178032 578700 178084
rect 578752 178072 578758 178084
rect 603074 178072 603080 178084
rect 578752 178044 603080 178072
rect 578752 178032 578758 178044
rect 603074 178032 603080 178044
rect 603132 178032 603138 178084
rect 674650 177284 674656 177336
rect 674708 177324 674714 177336
rect 676030 177324 676036 177336
rect 674708 177296 676036 177324
rect 674708 177284 674714 177296
rect 676030 177284 676036 177296
rect 676088 177284 676094 177336
rect 670234 176808 670240 176860
rect 670292 176848 670298 176860
rect 675938 176848 675944 176860
rect 670292 176820 675944 176848
rect 670292 176808 670298 176820
rect 675938 176808 675944 176820
rect 675996 176808 676002 176860
rect 579430 176740 579436 176792
rect 579488 176780 579494 176792
rect 603166 176780 603172 176792
rect 579488 176752 603172 176780
rect 579488 176740 579494 176752
rect 603166 176740 603172 176752
rect 603224 176740 603230 176792
rect 579338 176672 579344 176724
rect 579396 176712 579402 176724
rect 603074 176712 603080 176724
rect 579396 176684 603080 176712
rect 579396 176672 579402 176684
rect 603074 176672 603080 176684
rect 603132 176672 603138 176724
rect 672902 176672 672908 176724
rect 672960 176712 672966 176724
rect 676030 176712 676036 176724
rect 672960 176684 676036 176712
rect 672960 176672 672966 176684
rect 676030 176672 676036 176684
rect 676088 176672 676094 176724
rect 673178 175992 673184 176044
rect 673236 176032 673242 176044
rect 676030 176032 676036 176044
rect 673236 176004 676036 176032
rect 673236 175992 673242 176004
rect 676030 175992 676036 176004
rect 676088 175992 676094 176044
rect 672626 175652 672632 175704
rect 672684 175692 672690 175704
rect 676030 175692 676036 175704
rect 672684 175664 676036 175692
rect 672684 175652 672690 175664
rect 676030 175652 676036 175664
rect 676088 175652 676094 175704
rect 580258 175244 580264 175296
rect 580316 175284 580322 175296
rect 603074 175284 603080 175296
rect 580316 175256 603080 175284
rect 580316 175244 580322 175256
rect 603074 175244 603080 175256
rect 603132 175244 603138 175296
rect 673270 175176 673276 175228
rect 673328 175216 673334 175228
rect 676030 175216 676036 175228
rect 673328 175188 676036 175216
rect 673328 175176 673334 175188
rect 676030 175176 676036 175188
rect 676088 175176 676094 175228
rect 673362 174836 673368 174888
rect 673420 174876 673426 174888
rect 676030 174876 676036 174888
rect 673420 174848 676036 174876
rect 673420 174836 673426 174848
rect 676030 174836 676036 174848
rect 676088 174836 676094 174888
rect 580350 173884 580356 173936
rect 580408 173924 580414 173936
rect 603074 173924 603080 173936
rect 580408 173896 603080 173924
rect 580408 173884 580414 173896
rect 603074 173884 603080 173896
rect 603132 173884 603138 173936
rect 668302 173748 668308 173800
rect 668360 173788 668366 173800
rect 672718 173788 672724 173800
rect 668360 173760 672724 173788
rect 668360 173748 668366 173760
rect 672718 173748 672724 173760
rect 672776 173748 672782 173800
rect 579154 172524 579160 172576
rect 579212 172564 579218 172576
rect 603074 172564 603080 172576
rect 579212 172536 603080 172564
rect 579212 172524 579218 172536
rect 603074 172524 603080 172536
rect 603132 172524 603138 172576
rect 676214 171232 676220 171284
rect 676272 171272 676278 171284
rect 677042 171272 677048 171284
rect 676272 171244 677048 171272
rect 676272 171232 676278 171244
rect 677042 171232 677048 171244
rect 677100 171232 677106 171284
rect 579246 171096 579252 171148
rect 579304 171136 579310 171148
rect 603074 171136 603080 171148
rect 579304 171108 603080 171136
rect 579304 171096 579310 171108
rect 603074 171096 603080 171108
rect 603132 171096 603138 171148
rect 676214 171096 676220 171148
rect 676272 171136 676278 171148
rect 676858 171136 676864 171148
rect 676272 171108 676864 171136
rect 676272 171096 676278 171108
rect 676858 171096 676864 171108
rect 676916 171096 676922 171148
rect 674650 170280 674656 170332
rect 674708 170320 674714 170332
rect 676030 170320 676036 170332
rect 674708 170292 676036 170320
rect 674708 170280 674714 170292
rect 676030 170280 676036 170292
rect 676088 170280 676094 170332
rect 579062 169804 579068 169856
rect 579120 169844 579126 169856
rect 603166 169844 603172 169856
rect 579120 169816 603172 169844
rect 579120 169804 579126 169816
rect 603166 169804 603172 169816
rect 603224 169804 603230 169856
rect 578878 169736 578884 169788
rect 578936 169776 578942 169788
rect 603074 169776 603080 169788
rect 578936 169748 603080 169776
rect 578936 169736 578942 169748
rect 603074 169736 603080 169748
rect 603132 169736 603138 169788
rect 672994 169464 673000 169516
rect 673052 169504 673058 169516
rect 676030 169504 676036 169516
rect 673052 169476 676036 169504
rect 673052 169464 673058 169476
rect 676030 169464 676036 169476
rect 676088 169464 676094 169516
rect 674558 169056 674564 169108
rect 674616 169096 674622 169108
rect 676030 169096 676036 169108
rect 674616 169068 676036 169096
rect 674616 169056 674622 169068
rect 676030 169056 676036 169068
rect 676088 169056 676094 169108
rect 668302 168648 668308 168700
rect 668360 168688 668366 168700
rect 674190 168688 674196 168700
rect 668360 168660 674196 168688
rect 668360 168648 668366 168660
rect 674190 168648 674196 168660
rect 674248 168648 674254 168700
rect 673086 168580 673092 168632
rect 673144 168620 673150 168632
rect 676030 168620 676036 168632
rect 673144 168592 676036 168620
rect 673144 168580 673150 168592
rect 676030 168580 676036 168592
rect 676088 168580 676094 168632
rect 578970 168376 578976 168428
rect 579028 168416 579034 168428
rect 603074 168416 603080 168428
rect 579028 168388 603080 168416
rect 579028 168376 579034 168388
rect 603074 168376 603080 168388
rect 603132 168376 603138 168428
rect 669958 168240 669964 168292
rect 670016 168280 670022 168292
rect 676030 168280 676036 168292
rect 670016 168252 676036 168280
rect 670016 168240 670022 168252
rect 676030 168240 676036 168252
rect 676088 168240 676094 168292
rect 671522 167832 671528 167884
rect 671580 167872 671586 167884
rect 676030 167872 676036 167884
rect 671580 167844 676036 167872
rect 671580 167832 671586 167844
rect 676030 167832 676036 167844
rect 676088 167832 676094 167884
rect 583110 167016 583116 167068
rect 583168 167056 583174 167068
rect 603074 167056 603080 167068
rect 583168 167028 603080 167056
rect 583168 167016 583174 167028
rect 603074 167016 603080 167028
rect 603132 167016 603138 167068
rect 674190 167016 674196 167068
rect 674248 167056 674254 167068
rect 676030 167056 676036 167068
rect 674248 167028 676036 167056
rect 674248 167016 674254 167028
rect 676030 167016 676036 167028
rect 676088 167016 676094 167068
rect 578602 166948 578608 167000
rect 578660 166988 578666 167000
rect 580258 166988 580264 167000
rect 578660 166960 580264 166988
rect 578660 166948 578666 166960
rect 580258 166948 580264 166960
rect 580316 166948 580322 167000
rect 581638 165588 581644 165640
rect 581696 165628 581702 165640
rect 603074 165628 603080 165640
rect 581696 165600 603080 165628
rect 581696 165588 581702 165600
rect 603074 165588 603080 165600
rect 603132 165588 603138 165640
rect 578234 164432 578240 164484
rect 578292 164472 578298 164484
rect 580350 164472 580356 164484
rect 578292 164444 580356 164472
rect 578292 164432 578298 164444
rect 580350 164432 580356 164444
rect 580408 164432 580414 164484
rect 581730 164228 581736 164280
rect 581788 164268 581794 164280
rect 603074 164268 603080 164280
rect 581788 164240 603080 164268
rect 581788 164228 581794 164240
rect 603074 164228 603080 164240
rect 603132 164228 603138 164280
rect 579522 164160 579528 164212
rect 579580 164200 579586 164212
rect 603718 164200 603724 164212
rect 579580 164172 603724 164200
rect 579580 164160 579586 164172
rect 603718 164160 603724 164172
rect 603776 164160 603782 164212
rect 667934 163820 667940 163872
rect 667992 163860 667998 163872
rect 671338 163860 671344 163872
rect 667992 163832 671344 163860
rect 667992 163820 667998 163832
rect 671338 163820 671344 163832
rect 671396 163820 671402 163872
rect 580258 162868 580264 162920
rect 580316 162908 580322 162920
rect 603074 162908 603080 162920
rect 580316 162880 603080 162908
rect 580316 162868 580322 162880
rect 603074 162868 603080 162880
rect 603132 162868 603138 162920
rect 675754 162800 675760 162852
rect 675812 162840 675818 162852
rect 678238 162840 678244 162852
rect 675812 162812 678244 162840
rect 675812 162800 675818 162812
rect 678238 162800 678244 162812
rect 678296 162800 678302 162852
rect 584490 161440 584496 161492
rect 584548 161480 584554 161492
rect 603074 161480 603080 161492
rect 584548 161452 603080 161480
rect 584548 161440 584554 161452
rect 603074 161440 603080 161452
rect 603132 161440 603138 161492
rect 675754 160964 675760 161016
rect 675812 160964 675818 161016
rect 675772 160812 675800 160964
rect 675754 160760 675760 160812
rect 675812 160760 675818 160812
rect 579154 160080 579160 160132
rect 579212 160120 579218 160132
rect 603074 160120 603080 160132
rect 579212 160092 603080 160120
rect 579212 160080 579218 160092
rect 603074 160080 603080 160092
rect 603132 160080 603138 160132
rect 579338 158720 579344 158772
rect 579396 158760 579402 158772
rect 603074 158760 603080 158772
rect 579396 158732 603080 158760
rect 579396 158720 579402 158732
rect 603074 158720 603080 158732
rect 603132 158720 603138 158772
rect 592678 157428 592684 157480
rect 592736 157468 592742 157480
rect 603166 157468 603172 157480
rect 592736 157440 603172 157468
rect 592736 157428 592742 157440
rect 603166 157428 603172 157440
rect 603224 157428 603230 157480
rect 584398 157360 584404 157412
rect 584456 157400 584462 157412
rect 603074 157400 603080 157412
rect 584456 157372 603080 157400
rect 584456 157360 584462 157372
rect 603074 157360 603080 157372
rect 603132 157360 603138 157412
rect 585778 155932 585784 155984
rect 585836 155972 585842 155984
rect 603074 155972 603080 155984
rect 585836 155944 603080 155972
rect 585836 155932 585842 155944
rect 603074 155932 603080 155944
rect 603132 155932 603138 155984
rect 672994 155456 673000 155508
rect 673052 155496 673058 155508
rect 675478 155496 675484 155508
rect 673052 155468 675484 155496
rect 673052 155456 673058 155468
rect 675478 155456 675484 155468
rect 675536 155456 675542 155508
rect 578326 154844 578332 154896
rect 578384 154884 578390 154896
rect 583110 154884 583116 154896
rect 578384 154856 583116 154884
rect 578384 154844 578390 154856
rect 583110 154844 583116 154856
rect 583168 154844 583174 154896
rect 579246 154572 579252 154624
rect 579304 154612 579310 154624
rect 603074 154612 603080 154624
rect 579304 154584 603080 154612
rect 579304 154572 579310 154584
rect 603074 154572 603080 154584
rect 603132 154572 603138 154624
rect 579062 153280 579068 153332
rect 579120 153320 579126 153332
rect 603166 153320 603172 153332
rect 579120 153292 603172 153320
rect 579120 153280 579126 153292
rect 603166 153280 603172 153292
rect 603224 153280 603230 153332
rect 578878 153212 578884 153264
rect 578936 153252 578942 153264
rect 603074 153252 603080 153264
rect 578936 153224 603080 153252
rect 578936 153212 578942 153224
rect 603074 153212 603080 153224
rect 603132 153212 603138 153264
rect 579522 153144 579528 153196
rect 579580 153184 579586 153196
rect 603810 153184 603816 153196
rect 579580 153156 603816 153184
rect 579580 153144 579586 153156
rect 603810 153144 603816 153156
rect 603868 153144 603874 153196
rect 674558 152532 674564 152584
rect 674616 152572 674622 152584
rect 675386 152572 675392 152584
rect 674616 152544 675392 152572
rect 674616 152532 674622 152544
rect 675386 152532 675392 152544
rect 675444 152532 675450 152584
rect 580350 151784 580356 151836
rect 580408 151824 580414 151836
rect 603074 151824 603080 151836
rect 580408 151796 603080 151824
rect 580408 151784 580414 151796
rect 603074 151784 603080 151796
rect 603132 151784 603138 151836
rect 579430 151580 579436 151632
rect 579488 151620 579494 151632
rect 581638 151620 581644 151632
rect 579488 151592 581644 151620
rect 579488 151580 579494 151592
rect 581638 151580 581644 151592
rect 581696 151580 581702 151632
rect 673086 151376 673092 151428
rect 673144 151416 673150 151428
rect 675386 151416 675392 151428
rect 673144 151388 675392 151416
rect 673144 151376 673150 151388
rect 675386 151376 675392 151388
rect 675444 151376 675450 151428
rect 578970 150424 578976 150476
rect 579028 150464 579034 150476
rect 603074 150464 603080 150476
rect 579028 150436 603080 150464
rect 579028 150424 579034 150436
rect 603074 150424 603080 150436
rect 603132 150424 603138 150476
rect 674650 150356 674656 150408
rect 674708 150396 674714 150408
rect 675386 150396 675392 150408
rect 674708 150368 675392 150396
rect 674708 150356 674714 150368
rect 675386 150356 675392 150368
rect 675444 150356 675450 150408
rect 579430 150220 579436 150272
rect 579488 150260 579494 150272
rect 581730 150260 581736 150272
rect 579488 150232 581736 150260
rect 579488 150220 579494 150232
rect 581730 150220 581736 150232
rect 581788 150220 581794 150272
rect 589918 149064 589924 149116
rect 589976 149104 589982 149116
rect 603074 149104 603080 149116
rect 589976 149076 603080 149104
rect 589976 149064 589982 149076
rect 603074 149064 603080 149076
rect 603132 149064 603138 149116
rect 578510 148588 578516 148640
rect 578568 148628 578574 148640
rect 580258 148628 580264 148640
rect 578568 148600 580264 148628
rect 578568 148588 578574 148600
rect 580258 148588 580264 148600
rect 580316 148588 580322 148640
rect 668302 148384 668308 148436
rect 668360 148424 668366 148436
rect 674282 148424 674288 148436
rect 668360 148396 674288 148424
rect 668360 148384 668366 148396
rect 674282 148384 674288 148396
rect 674340 148384 674346 148436
rect 587250 147636 587256 147688
rect 587308 147676 587314 147688
rect 603074 147676 603080 147688
rect 587308 147648 603080 147676
rect 587308 147636 587314 147648
rect 603074 147636 603080 147648
rect 603132 147636 603138 147688
rect 579522 146956 579528 147008
rect 579580 146996 579586 147008
rect 583018 146996 583024 147008
rect 579580 146968 583024 146996
rect 579580 146956 579586 146968
rect 583018 146956 583024 146968
rect 583076 146956 583082 147008
rect 579614 146888 579620 146940
rect 579672 146928 579678 146940
rect 603718 146928 603724 146940
rect 579672 146900 603724 146928
rect 579672 146888 579678 146900
rect 603718 146888 603724 146900
rect 603776 146888 603782 146940
rect 591298 146276 591304 146328
rect 591356 146316 591362 146328
rect 603074 146316 603080 146328
rect 591356 146288 603080 146316
rect 591356 146276 591362 146288
rect 603074 146276 603080 146288
rect 603132 146276 603138 146328
rect 578694 146140 578700 146192
rect 578752 146180 578758 146192
rect 584490 146180 584496 146192
rect 578752 146152 584496 146180
rect 578752 146140 578758 146152
rect 584490 146140 584496 146152
rect 584548 146140 584554 146192
rect 583018 144916 583024 144968
rect 583076 144956 583082 144968
rect 603166 144956 603172 144968
rect 583076 144928 603172 144956
rect 583076 144916 583082 144928
rect 603166 144916 603172 144928
rect 603224 144916 603230 144968
rect 580258 143556 580264 143608
rect 580316 143596 580322 143608
rect 603074 143596 603080 143608
rect 580316 143568 603080 143596
rect 580316 143556 580322 143568
rect 603074 143556 603080 143568
rect 603132 143556 603138 143608
rect 578694 143488 578700 143540
rect 578752 143528 578758 143540
rect 592678 143528 592684 143540
rect 578752 143500 592684 143528
rect 578752 143488 578758 143500
rect 592678 143488 592684 143500
rect 592736 143488 592742 143540
rect 667934 143420 667940 143472
rect 667992 143460 667998 143472
rect 670142 143460 670148 143472
rect 667992 143432 670148 143460
rect 667992 143420 667998 143432
rect 670142 143420 670148 143432
rect 670200 143420 670206 143472
rect 591482 142128 591488 142180
rect 591540 142168 591546 142180
rect 603074 142168 603080 142180
rect 591540 142140 603080 142168
rect 591540 142128 591546 142140
rect 603074 142128 603080 142140
rect 603132 142128 603138 142180
rect 588630 140768 588636 140820
rect 588688 140808 588694 140820
rect 603074 140808 603080 140820
rect 588688 140780 603080 140808
rect 588688 140768 588694 140780
rect 603074 140768 603080 140780
rect 603132 140768 603138 140820
rect 584674 140020 584680 140072
rect 584732 140060 584738 140072
rect 603902 140060 603908 140072
rect 584732 140032 603908 140060
rect 584732 140020 584738 140032
rect 603902 140020 603908 140032
rect 603960 140020 603966 140072
rect 594150 139408 594156 139460
rect 594208 139448 594214 139460
rect 603074 139448 603080 139460
rect 594208 139420 603080 139448
rect 594208 139408 594214 139420
rect 603074 139408 603080 139420
rect 603132 139408 603138 139460
rect 667934 138184 667940 138236
rect 667992 138224 667998 138236
rect 671430 138224 671436 138236
rect 667992 138196 671436 138224
rect 667992 138184 667998 138196
rect 671430 138184 671436 138196
rect 671488 138184 671494 138236
rect 590102 138048 590108 138100
rect 590160 138088 590166 138100
rect 603074 138088 603080 138100
rect 590160 138060 603080 138088
rect 590160 138048 590166 138060
rect 603074 138048 603080 138060
rect 603132 138048 603138 138100
rect 587158 137980 587164 138032
rect 587216 138020 587222 138032
rect 603166 138020 603172 138032
rect 587216 137992 603172 138020
rect 587216 137980 587222 137992
rect 603166 137980 603172 137992
rect 603224 137980 603230 138032
rect 579522 137912 579528 137964
rect 579580 137952 579586 137964
rect 585778 137952 585784 137964
rect 579580 137924 585784 137952
rect 579580 137912 579586 137924
rect 585778 137912 585784 137924
rect 585836 137912 585842 137964
rect 588538 136620 588544 136672
rect 588596 136660 588602 136672
rect 603074 136660 603080 136672
rect 588596 136632 603080 136660
rect 588596 136620 588602 136632
rect 603074 136620 603080 136632
rect 603132 136620 603138 136672
rect 579522 136484 579528 136536
rect 579580 136524 579586 136536
rect 584398 136524 584404 136536
rect 579580 136496 584404 136524
rect 579580 136484 579586 136496
rect 584398 136484 584404 136496
rect 584456 136484 584462 136536
rect 585778 135260 585784 135312
rect 585836 135300 585842 135312
rect 603074 135300 603080 135312
rect 585836 135272 603080 135300
rect 585836 135260 585842 135272
rect 603074 135260 603080 135272
rect 603132 135260 603138 135312
rect 585962 133968 585968 134020
rect 586020 134008 586026 134020
rect 603166 134008 603172 134020
rect 586020 133980 603172 134008
rect 586020 133968 586026 133980
rect 603166 133968 603172 133980
rect 603224 133968 603230 134020
rect 581822 133900 581828 133952
rect 581880 133940 581886 133952
rect 603074 133940 603080 133952
rect 581880 133912 603080 133940
rect 581880 133900 581886 133912
rect 603074 133900 603080 133912
rect 603132 133900 603138 133952
rect 581638 133152 581644 133204
rect 581696 133192 581702 133204
rect 603718 133192 603724 133204
rect 581696 133164 603724 133192
rect 581696 133152 581702 133164
rect 603718 133152 603724 133164
rect 603776 133152 603782 133204
rect 674098 133016 674104 133068
rect 674156 133056 674162 133068
rect 676030 133056 676036 133068
rect 674156 133028 676036 133056
rect 674156 133016 674162 133028
rect 676030 133016 676036 133028
rect 676088 133016 676094 133068
rect 668578 132948 668584 133000
rect 668636 132988 668642 133000
rect 674374 132988 674380 133000
rect 668636 132960 674380 132988
rect 668636 132948 668642 132960
rect 674374 132948 674380 132960
rect 674432 132948 674438 133000
rect 672810 132744 672816 132796
rect 672868 132784 672874 132796
rect 676214 132784 676220 132796
rect 672868 132756 676220 132784
rect 672868 132744 672874 132756
rect 676214 132744 676220 132756
rect 676272 132744 676278 132796
rect 667198 132608 667204 132660
rect 667256 132648 667262 132660
rect 676122 132648 676128 132660
rect 667256 132620 676128 132648
rect 667256 132608 667262 132620
rect 676122 132608 676128 132620
rect 676180 132608 676186 132660
rect 592770 132472 592776 132524
rect 592828 132512 592834 132524
rect 603074 132512 603080 132524
rect 592828 132484 603080 132512
rect 592828 132472 592834 132484
rect 603074 132472 603080 132484
rect 603132 132472 603138 132524
rect 672902 131384 672908 131436
rect 672960 131424 672966 131436
rect 676214 131424 676220 131436
rect 672960 131396 676220 131424
rect 672960 131384 672966 131396
rect 676214 131384 676220 131396
rect 676272 131384 676278 131436
rect 673178 131248 673184 131300
rect 673236 131288 673242 131300
rect 676030 131288 676036 131300
rect 673236 131260 676036 131288
rect 673236 131248 673242 131260
rect 676030 131248 676036 131260
rect 676088 131248 676094 131300
rect 584582 131112 584588 131164
rect 584640 131152 584646 131164
rect 603074 131152 603080 131164
rect 584640 131124 603080 131152
rect 584640 131112 584646 131124
rect 603074 131112 603080 131124
rect 603132 131112 603138 131164
rect 668670 131112 668676 131164
rect 668728 131152 668734 131164
rect 669038 131152 669044 131164
rect 668728 131124 669044 131152
rect 668728 131112 668734 131124
rect 669038 131112 669044 131124
rect 669096 131152 669102 131164
rect 676122 131152 676128 131164
rect 669096 131124 676128 131152
rect 669096 131112 669102 131124
rect 676122 131112 676128 131124
rect 676180 131112 676186 131164
rect 578326 130500 578332 130552
rect 578384 130540 578390 130552
rect 580350 130540 580356 130552
rect 578384 130512 580356 130540
rect 578384 130500 578390 130512
rect 580350 130500 580356 130512
rect 580408 130500 580414 130552
rect 673270 129956 673276 130008
rect 673328 129996 673334 130008
rect 676214 129996 676220 130008
rect 673328 129968 676220 129996
rect 673328 129956 673334 129968
rect 676214 129956 676220 129968
rect 676272 129956 676278 130008
rect 583110 129820 583116 129872
rect 583168 129860 583174 129872
rect 603166 129860 603172 129872
rect 583168 129832 603172 129860
rect 583168 129820 583174 129832
rect 603166 129820 603172 129832
rect 603224 129820 603230 129872
rect 672718 129820 672724 129872
rect 672776 129860 672782 129872
rect 676122 129860 676128 129872
rect 672776 129832 676128 129860
rect 672776 129820 672782 129832
rect 676122 129820 676128 129832
rect 676180 129820 676186 129872
rect 581730 129752 581736 129804
rect 581788 129792 581794 129804
rect 603074 129792 603080 129804
rect 581788 129764 603080 129792
rect 581788 129752 581794 129764
rect 603074 129752 603080 129764
rect 603132 129752 603138 129804
rect 668578 129752 668584 129804
rect 668636 129792 668642 129804
rect 668946 129792 668952 129804
rect 668636 129764 668952 129792
rect 668636 129752 668642 129764
rect 668946 129752 668952 129764
rect 669004 129792 669010 129804
rect 676214 129792 676220 129804
rect 669004 129764 676220 129792
rect 669004 129752 669010 129764
rect 676214 129752 676220 129764
rect 676272 129752 676278 129804
rect 584490 128324 584496 128376
rect 584548 128364 584554 128376
rect 603074 128364 603080 128376
rect 584548 128336 603080 128364
rect 584548 128324 584554 128336
rect 603074 128324 603080 128336
rect 603132 128324 603138 128376
rect 668762 128324 668768 128376
rect 668820 128364 668826 128376
rect 676214 128364 676220 128376
rect 668820 128336 676220 128364
rect 668820 128324 668826 128336
rect 676214 128324 676220 128336
rect 676272 128324 676278 128376
rect 579522 128256 579528 128308
rect 579580 128296 579586 128308
rect 587250 128296 587256 128308
rect 579580 128268 587256 128296
rect 579580 128256 579586 128268
rect 587250 128256 587256 128268
rect 587308 128256 587314 128308
rect 667934 127916 667940 127968
rect 667992 127956 667998 127968
rect 671614 127956 671620 127968
rect 667992 127928 671620 127956
rect 667992 127916 667998 127928
rect 671614 127916 671620 127928
rect 671672 127916 671678 127968
rect 580350 126964 580356 127016
rect 580408 127004 580414 127016
rect 603074 127004 603080 127016
rect 580408 126976 603080 127004
rect 580408 126964 580414 126976
rect 603074 126964 603080 126976
rect 603132 126964 603138 127016
rect 675110 126964 675116 127016
rect 675168 127004 675174 127016
rect 676030 127004 676036 127016
rect 675168 126976 676036 127004
rect 675168 126964 675174 126976
rect 676030 126964 676036 126976
rect 676088 126964 676094 127016
rect 578694 126012 578700 126064
rect 578752 126052 578758 126064
rect 584674 126052 584680 126064
rect 578752 126024 584680 126052
rect 578752 126012 578758 126024
rect 584674 126012 584680 126024
rect 584732 126012 584738 126064
rect 594058 125672 594064 125724
rect 594116 125712 594122 125724
rect 603074 125712 603080 125724
rect 594116 125684 603080 125712
rect 594116 125672 594122 125684
rect 603074 125672 603080 125684
rect 603132 125672 603138 125724
rect 587250 125604 587256 125656
rect 587308 125644 587314 125656
rect 603166 125644 603172 125656
rect 587308 125616 603172 125644
rect 587308 125604 587314 125616
rect 603166 125604 603172 125616
rect 603224 125604 603230 125656
rect 578418 125536 578424 125588
rect 578476 125576 578482 125588
rect 589918 125576 589924 125588
rect 578476 125548 589924 125576
rect 578476 125536 578482 125548
rect 589918 125536 589924 125548
rect 589976 125536 589982 125588
rect 591390 124176 591396 124228
rect 591448 124216 591454 124228
rect 603074 124216 603080 124228
rect 591448 124188 603080 124216
rect 591448 124176 591454 124188
rect 603074 124176 603080 124188
rect 603132 124176 603138 124228
rect 579246 124108 579252 124160
rect 579304 124148 579310 124160
rect 591298 124148 591304 124160
rect 579304 124120 591304 124148
rect 579304 124108 579310 124120
rect 591298 124108 591304 124120
rect 591356 124108 591362 124160
rect 667934 124040 667940 124092
rect 667992 124080 667998 124092
rect 670326 124080 670332 124092
rect 667992 124052 670332 124080
rect 667992 124040 667998 124052
rect 670326 124040 670332 124052
rect 670384 124040 670390 124092
rect 674650 123904 674656 123956
rect 674708 123944 674714 123956
rect 676030 123944 676036 123956
rect 674708 123916 676036 123944
rect 674708 123904 674714 123916
rect 676030 123904 676036 123916
rect 676088 123904 676094 123956
rect 598198 122884 598204 122936
rect 598256 122924 598262 122936
rect 603166 122924 603172 122936
rect 598256 122896 603172 122924
rect 598256 122884 598262 122896
rect 603166 122884 603172 122896
rect 603224 122884 603230 122936
rect 592678 122816 592684 122868
rect 592736 122856 592742 122868
rect 603074 122856 603080 122868
rect 592736 122828 603080 122856
rect 592736 122816 592742 122828
rect 603074 122816 603080 122828
rect 603132 122816 603138 122868
rect 668854 122816 668860 122868
rect 668912 122856 668918 122868
rect 676214 122856 676220 122868
rect 668912 122828 676220 122856
rect 668912 122816 668918 122828
rect 676214 122816 676220 122828
rect 676272 122816 676278 122868
rect 579430 122068 579436 122120
rect 579488 122108 579494 122120
rect 591482 122108 591488 122120
rect 579488 122080 591488 122108
rect 579488 122068 579494 122080
rect 591482 122068 591488 122080
rect 591540 122068 591546 122120
rect 591298 121456 591304 121508
rect 591356 121496 591362 121508
rect 603074 121496 603080 121508
rect 591356 121468 603080 121496
rect 591356 121456 591362 121468
rect 603074 121456 603080 121468
rect 603132 121456 603138 121508
rect 671338 121456 671344 121508
rect 671396 121496 671402 121508
rect 676122 121496 676128 121508
rect 671396 121468 676128 121496
rect 671396 121456 671402 121468
rect 676122 121456 676128 121468
rect 676180 121456 676186 121508
rect 579522 121388 579528 121440
rect 579580 121428 579586 121440
rect 583018 121428 583024 121440
rect 579580 121400 583024 121428
rect 579580 121388 579586 121400
rect 583018 121388 583024 121400
rect 583076 121388 583082 121440
rect 670050 120708 670056 120760
rect 670108 120748 670114 120760
rect 676214 120748 676220 120760
rect 670108 120720 676220 120748
rect 670108 120708 670114 120720
rect 676214 120708 676220 120720
rect 676272 120708 676278 120760
rect 590010 120096 590016 120148
rect 590068 120136 590074 120148
rect 603074 120136 603080 120148
rect 590068 120108 603080 120136
rect 590068 120096 590074 120108
rect 603074 120096 603080 120108
rect 603132 120096 603138 120148
rect 579246 120028 579252 120080
rect 579304 120068 579310 120080
rect 581638 120068 581644 120080
rect 579304 120040 581644 120068
rect 579304 120028 579310 120040
rect 581638 120028 581644 120040
rect 581696 120028 581702 120080
rect 579154 118668 579160 118720
rect 579212 118708 579218 118720
rect 603074 118708 603080 118720
rect 579212 118680 603080 118708
rect 579212 118668 579218 118680
rect 603074 118668 603080 118680
rect 603132 118668 603138 118720
rect 578510 118532 578516 118584
rect 578568 118572 578574 118584
rect 580258 118572 580264 118584
rect 578568 118544 580264 118572
rect 578568 118532 578574 118544
rect 580258 118532 580264 118544
rect 580316 118532 580322 118584
rect 667934 117716 667940 117768
rect 667992 117756 667998 117768
rect 669958 117756 669964 117768
rect 667992 117728 669964 117756
rect 667992 117716 667998 117728
rect 669958 117716 669964 117728
rect 670016 117716 670022 117768
rect 579062 117308 579068 117360
rect 579120 117348 579126 117360
rect 603074 117348 603080 117360
rect 579120 117320 603080 117348
rect 579120 117308 579126 117320
rect 603074 117308 603080 117320
rect 603132 117308 603138 117360
rect 579522 117240 579528 117292
rect 579580 117280 579586 117292
rect 603810 117280 603816 117292
rect 579580 117252 603816 117280
rect 579580 117240 579586 117252
rect 603810 117240 603816 117252
rect 603868 117240 603874 117292
rect 668394 116968 668400 117020
rect 668452 117008 668458 117020
rect 671522 117008 671528 117020
rect 668452 116980 671528 117008
rect 668452 116968 668458 116980
rect 671522 116968 671528 116980
rect 671580 116968 671586 117020
rect 675478 116696 675484 116748
rect 675536 116736 675542 116748
rect 677594 116736 677600 116748
rect 675536 116708 677600 116736
rect 675536 116696 675542 116708
rect 677594 116696 677600 116708
rect 677652 116696 677658 116748
rect 675202 116560 675208 116612
rect 675260 116600 675266 116612
rect 683298 116600 683304 116612
rect 675260 116572 683304 116600
rect 675260 116560 675266 116572
rect 683298 116560 683304 116572
rect 683356 116560 683362 116612
rect 678238 116192 678244 116204
rect 675036 116164 678244 116192
rect 675036 115444 675064 116164
rect 678238 116152 678244 116164
rect 678296 116152 678302 116204
rect 675478 115744 675484 115796
rect 675536 115744 675542 115796
rect 675110 115540 675116 115592
rect 675168 115580 675174 115592
rect 675386 115580 675392 115592
rect 675168 115552 675392 115580
rect 675168 115540 675174 115552
rect 675386 115540 675392 115552
rect 675444 115540 675450 115592
rect 675110 115444 675116 115456
rect 675036 115416 675116 115444
rect 675110 115404 675116 115416
rect 675168 115404 675174 115456
rect 675202 114792 675208 114844
rect 675260 114832 675266 114844
rect 675386 114832 675392 114844
rect 675260 114804 675392 114832
rect 675260 114792 675266 114804
rect 675386 114792 675392 114804
rect 675444 114792 675450 114844
rect 596818 114588 596824 114640
rect 596876 114628 596882 114640
rect 603166 114628 603172 114640
rect 596876 114600 603172 114628
rect 596876 114588 596882 114600
rect 603166 114588 603172 114600
rect 603224 114588 603230 114640
rect 675110 114588 675116 114640
rect 675168 114628 675174 114640
rect 675496 114628 675524 115744
rect 675168 114600 675524 114628
rect 675168 114588 675174 114600
rect 578970 114520 578976 114572
rect 579028 114560 579034 114572
rect 603074 114560 603080 114572
rect 579028 114532 603080 114560
rect 579028 114520 579034 114532
rect 603074 114520 603080 114532
rect 603132 114520 603138 114572
rect 579246 114452 579252 114504
rect 579304 114492 579310 114504
rect 588630 114492 588636 114504
rect 579304 114464 588636 114492
rect 579304 114452 579310 114464
rect 588630 114452 588636 114464
rect 588688 114452 588694 114504
rect 669222 114316 669228 114368
rect 669280 114356 669286 114368
rect 674190 114356 674196 114368
rect 669280 114328 674196 114356
rect 669280 114316 669286 114328
rect 674190 114316 674196 114328
rect 674248 114316 674254 114368
rect 578878 113160 578884 113212
rect 578936 113200 578942 113212
rect 603074 113200 603080 113212
rect 578936 113172 603080 113200
rect 578936 113160 578942 113172
rect 603074 113160 603080 113172
rect 603132 113160 603138 113212
rect 579522 113092 579528 113144
rect 579580 113132 579586 113144
rect 594150 113132 594156 113144
rect 579580 113104 594156 113132
rect 579580 113092 579586 113104
rect 594150 113092 594156 113104
rect 594208 113092 594214 113144
rect 595438 111800 595444 111852
rect 595496 111840 595502 111852
rect 603074 111840 603080 111852
rect 595496 111812 603080 111840
rect 595496 111800 595502 111812
rect 603074 111800 603080 111812
rect 603132 111800 603138 111852
rect 578694 111732 578700 111784
rect 578752 111772 578758 111784
rect 587158 111772 587164 111784
rect 578752 111744 587164 111772
rect 578752 111732 578758 111744
rect 587158 111732 587164 111744
rect 587216 111732 587222 111784
rect 668302 111732 668308 111784
rect 668360 111772 668366 111784
rect 671338 111772 671344 111784
rect 668360 111744 671344 111772
rect 668360 111732 668366 111744
rect 671338 111732 671344 111744
rect 671396 111732 671402 111784
rect 675202 111120 675208 111172
rect 675260 111160 675266 111172
rect 675386 111160 675392 111172
rect 675260 111132 675392 111160
rect 675260 111120 675266 111132
rect 675386 111120 675392 111132
rect 675444 111120 675450 111172
rect 675110 110644 675116 110696
rect 675168 110684 675174 110696
rect 675386 110684 675392 110696
rect 675168 110656 675392 110684
rect 675168 110644 675174 110656
rect 675386 110644 675392 110656
rect 675444 110644 675450 110696
rect 589918 110440 589924 110492
rect 589976 110480 589982 110492
rect 603074 110480 603080 110492
rect 589976 110452 603080 110480
rect 589976 110440 589982 110452
rect 603074 110440 603080 110452
rect 603132 110440 603138 110492
rect 579522 110372 579528 110424
rect 579580 110412 579586 110424
rect 590102 110412 590108 110424
rect 579580 110384 590108 110412
rect 579580 110372 579586 110384
rect 590102 110372 590108 110384
rect 590160 110372 590166 110424
rect 667934 109284 667940 109336
rect 667992 109324 667998 109336
rect 670050 109324 670056 109336
rect 667992 109296 670056 109324
rect 667992 109284 667998 109296
rect 670050 109284 670056 109296
rect 670108 109284 670114 109336
rect 588630 109012 588636 109064
rect 588688 109052 588694 109064
rect 603074 109052 603080 109064
rect 588688 109024 603080 109052
rect 588688 109012 588694 109024
rect 603074 109012 603080 109024
rect 603132 109012 603138 109064
rect 578786 108944 578792 108996
rect 578844 108984 578850 108996
rect 588538 108984 588544 108996
rect 578844 108956 588544 108984
rect 578844 108944 578850 108956
rect 588538 108944 588544 108956
rect 588596 108944 588602 108996
rect 585870 107652 585876 107704
rect 585928 107692 585934 107704
rect 603074 107692 603080 107704
rect 585928 107664 603080 107692
rect 585928 107652 585934 107664
rect 603074 107652 603080 107664
rect 603132 107652 603138 107704
rect 674650 107516 674656 107568
rect 674708 107556 674714 107568
rect 675386 107556 675392 107568
rect 674708 107528 675392 107556
rect 674708 107516 674714 107528
rect 675386 107516 675392 107528
rect 675444 107516 675450 107568
rect 579430 107040 579436 107092
rect 579488 107080 579494 107092
rect 585778 107080 585784 107092
rect 579488 107052 585784 107080
rect 579488 107040 579494 107052
rect 585778 107040 585784 107052
rect 585836 107040 585842 107092
rect 675110 106700 675116 106752
rect 675168 106740 675174 106752
rect 675386 106740 675392 106752
rect 675168 106712 675392 106740
rect 675168 106700 675174 106712
rect 675386 106700 675392 106712
rect 675444 106700 675450 106752
rect 588538 106360 588544 106412
rect 588596 106400 588602 106412
rect 603166 106400 603172 106412
rect 588596 106372 603172 106400
rect 588596 106360 588602 106372
rect 603166 106360 603172 106372
rect 603224 106360 603230 106412
rect 587158 106292 587164 106344
rect 587216 106332 587222 106344
rect 603074 106332 603080 106344
rect 587216 106304 603080 106332
rect 587216 106292 587222 106304
rect 603074 106292 603080 106304
rect 603132 106292 603138 106344
rect 674742 106224 674748 106276
rect 674800 106264 674806 106276
rect 675386 106264 675392 106276
rect 674800 106236 675392 106264
rect 674800 106224 674806 106236
rect 675386 106224 675392 106236
rect 675444 106224 675450 106276
rect 669222 106088 669228 106140
rect 669280 106128 669286 106140
rect 672718 106128 672724 106140
rect 669280 106100 672724 106128
rect 669280 106088 669286 106100
rect 672718 106088 672724 106100
rect 672776 106088 672782 106140
rect 578234 105136 578240 105188
rect 578292 105176 578298 105188
rect 585962 105176 585968 105188
rect 578292 105148 585968 105176
rect 578292 105136 578298 105148
rect 585962 105136 585968 105148
rect 586020 105136 586026 105188
rect 585778 104864 585784 104916
rect 585836 104904 585842 104916
rect 603074 104904 603080 104916
rect 585836 104876 603080 104904
rect 585836 104864 585842 104876
rect 603074 104864 603080 104876
rect 603132 104864 603138 104916
rect 584398 103504 584404 103556
rect 584456 103544 584462 103556
rect 603074 103544 603080 103556
rect 584456 103516 603080 103544
rect 584456 103504 584462 103516
rect 603074 103504 603080 103516
rect 603132 103504 603138 103556
rect 579338 103436 579344 103488
rect 579396 103476 579402 103488
rect 581822 103476 581828 103488
rect 579396 103448 581828 103476
rect 579396 103436 579402 103448
rect 581822 103436 581828 103448
rect 581880 103436 581886 103488
rect 583018 102212 583024 102264
rect 583076 102252 583082 102264
rect 603166 102252 603172 102264
rect 583076 102224 603172 102252
rect 583076 102212 583082 102224
rect 603166 102212 603172 102224
rect 603224 102212 603230 102264
rect 581638 102144 581644 102196
rect 581696 102184 581702 102196
rect 603074 102184 603080 102196
rect 581696 102156 603080 102184
rect 581696 102144 581702 102156
rect 603074 102144 603080 102156
rect 603132 102144 603138 102196
rect 578326 102076 578332 102128
rect 578384 102116 578390 102128
rect 592770 102116 592776 102128
rect 578384 102088 592776 102116
rect 578384 102076 578390 102088
rect 592770 102076 592776 102088
rect 592828 102076 592834 102128
rect 580258 100716 580264 100768
rect 580316 100756 580322 100768
rect 603074 100756 603080 100768
rect 580316 100728 603080 100756
rect 580316 100716 580322 100728
rect 603074 100716 603080 100728
rect 603132 100716 603138 100768
rect 578694 100308 578700 100360
rect 578752 100348 578758 100360
rect 584582 100348 584588 100360
rect 578752 100320 584588 100348
rect 578752 100308 578758 100320
rect 584582 100308 584588 100320
rect 584640 100308 584646 100360
rect 600958 99356 600964 99408
rect 601016 99396 601022 99408
rect 603442 99396 603448 99408
rect 601016 99368 603448 99396
rect 601016 99356 601022 99368
rect 603442 99356 603448 99368
rect 603500 99356 603506 99408
rect 579522 99084 579528 99136
rect 579580 99124 579586 99136
rect 583110 99124 583116 99136
rect 579580 99096 583116 99124
rect 579580 99084 579586 99096
rect 583110 99084 583116 99096
rect 583168 99084 583174 99136
rect 624602 97928 624608 97980
rect 624660 97968 624666 97980
rect 625798 97968 625804 97980
rect 624660 97940 625804 97968
rect 624660 97928 624666 97940
rect 625798 97928 625804 97940
rect 625856 97928 625862 97980
rect 633802 97928 633808 97980
rect 633860 97968 633866 97980
rect 636378 97968 636384 97980
rect 633860 97940 636384 97968
rect 633860 97928 633866 97940
rect 636378 97928 636384 97940
rect 636436 97928 636442 97980
rect 663058 97928 663064 97980
rect 663116 97968 663122 97980
rect 665358 97968 665364 97980
rect 663116 97940 665364 97968
rect 663116 97928 663122 97940
rect 665358 97928 665364 97940
rect 665416 97928 665422 97980
rect 633066 97860 633072 97912
rect 633124 97900 633130 97912
rect 635274 97900 635280 97912
rect 633124 97872 635280 97900
rect 633124 97860 633130 97872
rect 635274 97860 635280 97872
rect 635332 97860 635338 97912
rect 637482 97860 637488 97912
rect 637540 97900 637546 97912
rect 644658 97900 644664 97912
rect 637540 97872 644664 97900
rect 637540 97860 637546 97872
rect 644658 97860 644664 97872
rect 644716 97860 644722 97912
rect 649442 97860 649448 97912
rect 649500 97900 649506 97912
rect 658826 97900 658832 97912
rect 649500 97872 658832 97900
rect 649500 97860 649506 97872
rect 658826 97860 658832 97872
rect 658884 97860 658890 97912
rect 638310 97792 638316 97844
rect 638368 97832 638374 97844
rect 644750 97832 644756 97844
rect 638368 97804 644756 97832
rect 638368 97792 638374 97804
rect 644750 97792 644756 97804
rect 644808 97792 644814 97844
rect 647510 97792 647516 97844
rect 647568 97832 647574 97844
rect 654778 97832 654784 97844
rect 647568 97804 654784 97832
rect 647568 97792 647574 97804
rect 654778 97792 654784 97804
rect 654836 97792 654842 97844
rect 635090 97724 635096 97776
rect 635148 97764 635154 97776
rect 639046 97764 639052 97776
rect 635148 97736 639052 97764
rect 635148 97724 635154 97736
rect 639046 97724 639052 97736
rect 639104 97724 639110 97776
rect 634446 97656 634452 97708
rect 634504 97696 634510 97708
rect 637574 97696 637580 97708
rect 634504 97668 637580 97696
rect 634504 97656 634510 97668
rect 637574 97656 637580 97668
rect 637632 97656 637638 97708
rect 578694 97588 578700 97640
rect 578752 97628 578758 97640
rect 581730 97628 581736 97640
rect 578752 97600 581736 97628
rect 578752 97588 578758 97600
rect 581730 97588 581736 97600
rect 581788 97588 581794 97640
rect 631134 97588 631140 97640
rect 631192 97628 631198 97640
rect 632146 97628 632152 97640
rect 631192 97600 632152 97628
rect 631192 97588 631198 97600
rect 632146 97588 632152 97600
rect 632204 97588 632210 97640
rect 635734 97588 635740 97640
rect 635792 97628 635798 97640
rect 639874 97628 639880 97640
rect 635792 97600 639880 97628
rect 635792 97588 635798 97600
rect 639874 97588 639880 97600
rect 639932 97588 639938 97640
rect 637022 97520 637028 97572
rect 637080 97560 637086 97572
rect 642174 97560 642180 97572
rect 637080 97532 642180 97560
rect 637080 97520 637086 97532
rect 642174 97520 642180 97532
rect 642232 97520 642238 97572
rect 614850 97452 614856 97504
rect 614908 97492 614914 97504
rect 621658 97492 621664 97504
rect 614908 97464 621664 97492
rect 614908 97452 614914 97464
rect 621658 97452 621664 97464
rect 621716 97452 621722 97504
rect 643554 97452 643560 97504
rect 643612 97492 643618 97504
rect 660390 97492 660396 97504
rect 643612 97464 660396 97492
rect 643612 97452 643618 97464
rect 660390 97452 660396 97464
rect 660448 97452 660454 97504
rect 620738 97384 620744 97436
rect 620796 97424 620802 97436
rect 646038 97424 646044 97436
rect 620796 97396 646044 97424
rect 620796 97384 620802 97396
rect 646038 97384 646044 97396
rect 646096 97384 646102 97436
rect 648154 97384 648160 97436
rect 648212 97424 648218 97436
rect 660114 97424 660120 97436
rect 648212 97396 660120 97424
rect 648212 97384 648218 97396
rect 660114 97384 660120 97396
rect 660172 97384 660178 97436
rect 652018 97316 652024 97368
rect 652076 97356 652082 97368
rect 652076 97328 654640 97356
rect 652076 97316 652082 97328
rect 622026 97248 622032 97300
rect 622084 97288 622090 97300
rect 648614 97288 648620 97300
rect 622084 97260 648620 97288
rect 622084 97248 622090 97260
rect 648614 97248 648620 97260
rect 648672 97248 648678 97300
rect 621382 97180 621388 97232
rect 621440 97220 621446 97232
rect 647418 97220 647424 97232
rect 621440 97192 647424 97220
rect 621440 97180 621446 97192
rect 647418 97180 647424 97192
rect 647476 97180 647482 97232
rect 631778 97112 631784 97164
rect 631836 97152 631842 97164
rect 632974 97152 632980 97164
rect 631836 97124 632980 97152
rect 631836 97112 631842 97124
rect 632974 97112 632980 97124
rect 633032 97112 633038 97164
rect 654612 97152 654640 97328
rect 655974 97316 655980 97368
rect 656032 97356 656038 97368
rect 659562 97356 659568 97368
rect 656032 97328 659568 97356
rect 656032 97316 656038 97328
rect 659562 97316 659568 97328
rect 659620 97316 659626 97368
rect 657722 97248 657728 97300
rect 657780 97288 657786 97300
rect 660666 97288 660672 97300
rect 657780 97260 660672 97288
rect 657780 97248 657786 97260
rect 660666 97248 660672 97260
rect 660724 97248 660730 97300
rect 654686 97180 654692 97232
rect 654744 97220 654750 97232
rect 658366 97220 658372 97232
rect 654744 97192 658372 97220
rect 654744 97180 654750 97192
rect 658366 97180 658372 97192
rect 658424 97180 658430 97232
rect 660574 97180 660580 97232
rect 660632 97220 660638 97232
rect 661402 97220 661408 97232
rect 660632 97192 661408 97220
rect 660632 97180 660638 97192
rect 661402 97180 661408 97192
rect 661460 97180 661466 97232
rect 661954 97152 661960 97164
rect 654612 97124 661960 97152
rect 661954 97112 661960 97124
rect 662012 97112 662018 97164
rect 662322 97112 662328 97164
rect 662380 97152 662386 97164
rect 663978 97152 663984 97164
rect 662380 97124 663984 97152
rect 662380 97112 662386 97124
rect 663978 97112 663984 97124
rect 664036 97112 664042 97164
rect 610066 96908 610072 96960
rect 610124 96948 610130 96960
rect 610894 96948 610900 96960
rect 610124 96920 610900 96948
rect 610124 96908 610130 96920
rect 610894 96908 610900 96920
rect 610952 96908 610958 96960
rect 611354 96908 611360 96960
rect 611412 96948 611418 96960
rect 612182 96948 612188 96960
rect 611412 96920 612188 96948
rect 611412 96908 611418 96920
rect 612182 96908 612188 96920
rect 612240 96908 612246 96960
rect 616138 96908 616144 96960
rect 616196 96948 616202 96960
rect 616782 96948 616788 96960
rect 616196 96920 616788 96948
rect 616196 96908 616202 96920
rect 616782 96908 616788 96920
rect 616840 96908 616846 96960
rect 617426 96908 617432 96960
rect 617484 96948 617490 96960
rect 618162 96948 618168 96960
rect 617484 96920 618168 96948
rect 617484 96908 617490 96920
rect 618162 96908 618168 96920
rect 618220 96908 618226 96960
rect 623682 96908 623688 96960
rect 623740 96948 623746 96960
rect 624418 96948 624424 96960
rect 623740 96920 624424 96948
rect 623740 96908 623746 96920
rect 624418 96908 624424 96920
rect 624476 96908 624482 96960
rect 625890 96908 625896 96960
rect 625948 96948 625954 96960
rect 626442 96948 626448 96960
rect 625948 96920 626448 96948
rect 625948 96908 625954 96920
rect 626442 96908 626448 96920
rect 626500 96908 626506 96960
rect 645486 96908 645492 96960
rect 645544 96948 645550 96960
rect 646498 96948 646504 96960
rect 645544 96920 646504 96948
rect 645544 96908 645550 96920
rect 646498 96908 646504 96920
rect 646556 96908 646562 96960
rect 655422 96908 655428 96960
rect 655480 96948 655486 96960
rect 659286 96948 659292 96960
rect 655480 96920 659292 96948
rect 655480 96908 655486 96920
rect 659286 96908 659292 96920
rect 659344 96908 659350 96960
rect 618714 96840 618720 96892
rect 618772 96880 618778 96892
rect 619542 96880 619548 96892
rect 618772 96852 619548 96880
rect 618772 96840 618778 96852
rect 619542 96840 619548 96852
rect 619600 96840 619606 96892
rect 620002 96840 620008 96892
rect 620060 96880 620066 96892
rect 620922 96880 620928 96892
rect 620060 96852 620928 96880
rect 620060 96840 620066 96852
rect 620922 96840 620928 96852
rect 620980 96840 620986 96892
rect 632422 96840 632428 96892
rect 632480 96880 632486 96892
rect 634078 96880 634084 96892
rect 632480 96852 634084 96880
rect 632480 96840 632486 96852
rect 634078 96840 634084 96852
rect 634136 96840 634142 96892
rect 640978 96840 640984 96892
rect 641036 96880 641042 96892
rect 643278 96880 643284 96892
rect 641036 96852 643284 96880
rect 641036 96840 641042 96852
rect 643278 96840 643284 96852
rect 643336 96840 643342 96892
rect 650730 96840 650736 96892
rect 650788 96880 650794 96892
rect 651282 96880 651288 96892
rect 650788 96852 651288 96880
rect 650788 96840 650794 96852
rect 651282 96840 651288 96852
rect 651340 96840 651346 96892
rect 661862 96840 661868 96892
rect 661920 96880 661926 96892
rect 663058 96880 663064 96892
rect 661920 96852 663064 96880
rect 661920 96840 661926 96852
rect 663058 96840 663064 96852
rect 663116 96840 663122 96892
rect 622670 96772 622676 96824
rect 622728 96812 622734 96824
rect 623682 96812 623688 96824
rect 622728 96784 623688 96812
rect 622728 96772 622734 96784
rect 623682 96772 623688 96784
rect 623740 96772 623746 96824
rect 659194 96772 659200 96824
rect 659252 96812 659258 96824
rect 662506 96812 662512 96824
rect 659252 96784 662512 96812
rect 659252 96772 659258 96784
rect 662506 96772 662512 96784
rect 662564 96772 662570 96824
rect 636102 96704 636108 96756
rect 636160 96744 636166 96756
rect 640978 96744 640984 96756
rect 636160 96716 640984 96744
rect 636160 96704 636166 96716
rect 640978 96704 640984 96716
rect 641036 96704 641042 96756
rect 639598 96568 639604 96620
rect 639656 96608 639662 96620
rect 643094 96608 643100 96620
rect 639656 96580 643100 96608
rect 639656 96568 639662 96580
rect 643094 96568 643100 96580
rect 643152 96568 643158 96620
rect 644842 96568 644848 96620
rect 644900 96608 644906 96620
rect 651926 96608 651932 96620
rect 644900 96580 651932 96608
rect 644900 96568 644906 96580
rect 651926 96568 651932 96580
rect 651984 96568 651990 96620
rect 656802 96568 656808 96620
rect 656860 96608 656866 96620
rect 658274 96608 658280 96620
rect 656860 96580 658280 96608
rect 656860 96568 656866 96580
rect 658274 96568 658280 96580
rect 658332 96568 658338 96620
rect 656618 96160 656624 96212
rect 656676 96200 656682 96212
rect 663886 96200 663892 96212
rect 656676 96172 663892 96200
rect 656676 96160 656682 96172
rect 663886 96160 663892 96172
rect 663944 96160 663950 96212
rect 646774 96024 646780 96076
rect 646832 96064 646838 96076
rect 663794 96064 663800 96076
rect 646832 96036 663800 96064
rect 646832 96024 646838 96036
rect 663794 96024 663800 96036
rect 663852 96024 663858 96076
rect 578510 95956 578516 96008
rect 578568 95996 578574 96008
rect 584490 95996 584496 96008
rect 578568 95968 584496 95996
rect 578568 95956 578574 95968
rect 584490 95956 584496 95968
rect 584548 95956 584554 96008
rect 653306 95956 653312 96008
rect 653364 95996 653370 96008
rect 665266 95996 665272 96008
rect 653364 95968 665272 95996
rect 653364 95956 653370 95968
rect 665266 95956 665272 95968
rect 665324 95956 665330 96008
rect 640058 95888 640064 95940
rect 640116 95928 640122 95940
rect 644566 95928 644572 95940
rect 640116 95900 644572 95928
rect 640116 95888 640122 95900
rect 644566 95888 644572 95900
rect 644624 95888 644630 95940
rect 646130 95888 646136 95940
rect 646188 95928 646194 95940
rect 665174 95928 665180 95940
rect 646188 95900 665180 95928
rect 646188 95888 646194 95900
rect 665174 95888 665180 95900
rect 665232 95888 665238 95940
rect 641622 95616 641628 95668
rect 641680 95656 641686 95668
rect 645946 95656 645952 95668
rect 641680 95628 645952 95656
rect 641680 95616 641686 95628
rect 645946 95616 645952 95628
rect 646004 95616 646010 95668
rect 638862 95548 638868 95600
rect 638920 95588 638926 95600
rect 644474 95588 644480 95600
rect 638920 95560 644480 95588
rect 638920 95548 638926 95560
rect 644474 95548 644480 95560
rect 644532 95548 644538 95600
rect 607214 95480 607220 95532
rect 607272 95520 607278 95532
rect 607674 95520 607680 95532
rect 607272 95492 607680 95520
rect 607272 95480 607278 95492
rect 607674 95480 607680 95492
rect 607732 95480 607738 95532
rect 657262 95208 657268 95260
rect 657320 95248 657326 95260
rect 664070 95248 664076 95260
rect 657320 95220 664076 95248
rect 657320 95208 657326 95220
rect 664070 95208 664076 95220
rect 664128 95208 664134 95260
rect 578602 95140 578608 95192
rect 578660 95180 578666 95192
rect 580350 95180 580356 95192
rect 578660 95152 580356 95180
rect 578660 95140 578666 95152
rect 580350 95140 580356 95152
rect 580408 95140 580414 95192
rect 579522 93780 579528 93832
rect 579580 93820 579586 93832
rect 587250 93820 587256 93832
rect 579580 93792 587256 93820
rect 579580 93780 579586 93792
rect 587250 93780 587256 93792
rect 587308 93780 587314 93832
rect 579522 92420 579528 92472
rect 579580 92460 579586 92472
rect 594058 92460 594064 92472
rect 579580 92432 594064 92460
rect 579580 92420 579586 92432
rect 594058 92420 594064 92432
rect 594116 92420 594122 92472
rect 644382 92420 644388 92472
rect 644440 92460 644446 92472
rect 654318 92460 654324 92472
rect 644440 92432 654324 92460
rect 644440 92420 644446 92432
rect 654318 92420 654324 92432
rect 654376 92420 654382 92472
rect 579522 90992 579528 91044
rect 579580 91032 579586 91044
rect 591390 91032 591396 91044
rect 579580 91004 591396 91032
rect 579580 90992 579586 91004
rect 591390 90992 591396 91004
rect 591448 90992 591454 91044
rect 651926 90924 651932 90976
rect 651984 90964 651990 90976
rect 654318 90964 654324 90976
rect 651984 90936 654324 90964
rect 651984 90924 651990 90936
rect 654318 90924 654324 90936
rect 654376 90924 654382 90976
rect 579522 89632 579528 89684
rect 579580 89672 579586 89684
rect 592678 89672 592684 89684
rect 579580 89644 592684 89672
rect 579580 89632 579586 89644
rect 592678 89632 592684 89644
rect 592736 89632 592742 89684
rect 616690 89632 616696 89684
rect 616748 89672 616754 89684
rect 626442 89672 626448 89684
rect 616748 89644 626448 89672
rect 616748 89632 616754 89644
rect 626442 89632 626448 89644
rect 626500 89632 626506 89684
rect 656802 88816 656808 88868
rect 656860 88856 656866 88868
rect 658090 88856 658096 88868
rect 656860 88828 658096 88856
rect 656860 88816 656866 88828
rect 658090 88816 658096 88828
rect 658148 88816 658154 88868
rect 662322 88816 662328 88868
rect 662380 88856 662386 88868
rect 663978 88856 663984 88868
rect 662380 88828 663984 88856
rect 662380 88816 662386 88828
rect 663978 88816 663984 88828
rect 664036 88816 664042 88868
rect 616782 88272 616788 88324
rect 616840 88312 616846 88324
rect 626442 88312 626448 88324
rect 616840 88284 626448 88312
rect 616840 88272 616846 88284
rect 626442 88272 626448 88284
rect 626500 88272 626506 88324
rect 659470 88272 659476 88324
rect 659528 88312 659534 88324
rect 663150 88312 663156 88324
rect 659528 88284 663156 88312
rect 659528 88272 659534 88284
rect 663150 88272 663156 88284
rect 663208 88272 663214 88324
rect 620922 88204 620928 88256
rect 620980 88244 620986 88256
rect 626350 88244 626356 88256
rect 620980 88216 626356 88244
rect 620980 88204 620986 88216
rect 626350 88204 626356 88216
rect 626408 88204 626414 88256
rect 584490 87592 584496 87644
rect 584548 87632 584554 87644
rect 603718 87632 603724 87644
rect 584548 87604 603724 87632
rect 584548 87592 584554 87604
rect 603718 87592 603724 87604
rect 603776 87592 603782 87644
rect 646498 86980 646504 87032
rect 646556 87020 646562 87032
rect 660114 87020 660120 87032
rect 646556 86992 660120 87020
rect 646556 86980 646562 86992
rect 660114 86980 660120 86992
rect 660172 86980 660178 87032
rect 579522 86912 579528 86964
rect 579580 86952 579586 86964
rect 598198 86952 598204 86964
rect 579580 86924 598204 86952
rect 579580 86912 579586 86924
rect 598198 86912 598204 86924
rect 598256 86912 598262 86964
rect 651190 86912 651196 86964
rect 651248 86952 651254 86964
rect 657170 86952 657176 86964
rect 651248 86924 657176 86952
rect 651248 86912 651254 86924
rect 657170 86912 657176 86924
rect 657228 86912 657234 86964
rect 651282 86844 651288 86896
rect 651340 86884 651346 86896
rect 657722 86884 657728 86896
rect 651340 86856 657728 86884
rect 651340 86844 651346 86856
rect 657722 86844 657728 86856
rect 657780 86844 657786 86896
rect 649902 86776 649908 86828
rect 649960 86816 649966 86828
rect 660666 86816 660672 86828
rect 649960 86788 660672 86816
rect 649960 86776 649966 86788
rect 660666 86776 660672 86788
rect 660724 86776 660730 86828
rect 648522 86708 648528 86760
rect 648580 86748 648586 86760
rect 661402 86748 661408 86760
rect 648580 86720 661408 86748
rect 648580 86708 648586 86720
rect 661402 86708 661408 86720
rect 661460 86708 661466 86760
rect 653950 86640 653956 86692
rect 654008 86680 654014 86692
rect 658826 86680 658832 86692
rect 654008 86652 658832 86680
rect 654008 86640 654014 86652
rect 658826 86640 658832 86652
rect 658884 86640 658890 86692
rect 652662 86572 652668 86624
rect 652720 86612 652726 86624
rect 662506 86612 662512 86624
rect 652720 86584 662512 86612
rect 652720 86572 652726 86584
rect 662506 86572 662512 86584
rect 662564 86572 662570 86624
rect 619450 86232 619456 86284
rect 619508 86272 619514 86284
rect 626442 86272 626448 86284
rect 619508 86244 626448 86272
rect 619508 86232 619514 86244
rect 626442 86232 626448 86244
rect 626500 86232 626506 86284
rect 579522 85484 579528 85536
rect 579580 85524 579586 85536
rect 591298 85524 591304 85536
rect 579580 85496 591304 85524
rect 579580 85484 579586 85496
rect 591298 85484 591304 85496
rect 591356 85484 591362 85536
rect 619542 85484 619548 85536
rect 619600 85524 619606 85536
rect 626442 85524 626448 85536
rect 619600 85496 626448 85524
rect 619600 85484 619606 85496
rect 626442 85484 626448 85496
rect 626500 85484 626506 85536
rect 579522 84124 579528 84176
rect 579580 84164 579586 84176
rect 590010 84164 590016 84176
rect 579580 84136 590016 84164
rect 579580 84124 579586 84136
rect 590010 84124 590016 84136
rect 590068 84124 590074 84176
rect 618162 84124 618168 84176
rect 618220 84164 618226 84176
rect 626074 84164 626080 84176
rect 618220 84136 626080 84164
rect 618220 84124 618226 84136
rect 626074 84124 626080 84136
rect 626132 84124 626138 84176
rect 618070 84056 618076 84108
rect 618128 84096 618134 84108
rect 625614 84096 625620 84108
rect 618128 84068 625620 84096
rect 618128 84056 618134 84068
rect 625614 84056 625620 84068
rect 625672 84056 625678 84108
rect 581730 82084 581736 82136
rect 581788 82124 581794 82136
rect 603810 82124 603816 82136
rect 581788 82096 603816 82124
rect 581788 82084 581794 82096
rect 603810 82084 603816 82096
rect 603868 82084 603874 82136
rect 579522 80860 579528 80912
rect 579580 80900 579586 80912
rect 584490 80900 584496 80912
rect 579580 80872 584496 80900
rect 579580 80860 579586 80872
rect 584490 80860 584496 80872
rect 584548 80860 584554 80912
rect 624418 80656 624424 80708
rect 624476 80696 624482 80708
rect 648706 80696 648712 80708
rect 624476 80668 648712 80696
rect 624476 80656 624482 80668
rect 648706 80656 648712 80668
rect 648764 80656 648770 80708
rect 623590 79296 623596 79348
rect 623648 79336 623654 79348
rect 647326 79336 647332 79348
rect 623648 79308 647332 79336
rect 623648 79296 623654 79308
rect 647326 79296 647332 79308
rect 647384 79296 647390 79348
rect 579522 78616 579528 78668
rect 579580 78656 579586 78668
rect 602338 78656 602344 78668
rect 579580 78628 602344 78656
rect 579580 78616 579586 78628
rect 602338 78616 602344 78628
rect 602396 78616 602402 78668
rect 626442 78140 626448 78192
rect 626500 78180 626506 78192
rect 642450 78180 642456 78192
rect 626500 78152 642456 78180
rect 626500 78140 626506 78152
rect 642450 78140 642456 78152
rect 642508 78140 642514 78192
rect 631042 78072 631048 78124
rect 631100 78112 631106 78124
rect 638954 78112 638960 78124
rect 631100 78084 638960 78112
rect 631100 78072 631106 78084
rect 638954 78072 638960 78084
rect 639012 78072 639018 78124
rect 629202 78004 629208 78056
rect 629260 78044 629266 78056
rect 645302 78044 645308 78056
rect 629260 78016 645308 78044
rect 629260 78004 629266 78016
rect 645302 78004 645308 78016
rect 645360 78004 645366 78056
rect 605742 77936 605748 77988
rect 605800 77976 605806 77988
rect 636746 77976 636752 77988
rect 605800 77948 636752 77976
rect 605800 77936 605806 77948
rect 636746 77936 636752 77948
rect 636804 77936 636810 77988
rect 628374 77596 628380 77648
rect 628432 77636 628438 77648
rect 631502 77636 631508 77648
rect 628432 77608 631508 77636
rect 628432 77596 628438 77608
rect 631502 77596 631508 77608
rect 631560 77596 631566 77648
rect 579062 77324 579068 77376
rect 579120 77364 579126 77376
rect 628374 77364 628380 77376
rect 579120 77336 628380 77364
rect 579120 77324 579126 77336
rect 628374 77324 628380 77336
rect 628432 77324 628438 77376
rect 576118 77256 576124 77308
rect 576176 77296 576182 77308
rect 631042 77296 631048 77308
rect 576176 77268 631048 77296
rect 576176 77256 576182 77268
rect 631042 77256 631048 77268
rect 631100 77256 631106 77308
rect 623682 76508 623688 76560
rect 623740 76548 623746 76560
rect 646130 76548 646136 76560
rect 623740 76520 646136 76548
rect 623740 76508 623746 76520
rect 646130 76508 646136 76520
rect 646188 76508 646194 76560
rect 579522 75828 579528 75880
rect 579580 75868 579586 75880
rect 596818 75868 596824 75880
rect 579580 75840 596824 75868
rect 579580 75828 579586 75840
rect 596818 75828 596824 75840
rect 596876 75828 596882 75880
rect 617518 75216 617524 75268
rect 617576 75256 617582 75268
rect 631134 75256 631140 75268
rect 617576 75228 631140 75256
rect 617576 75216 617582 75228
rect 631134 75216 631140 75228
rect 631192 75216 631198 75268
rect 615402 75148 615408 75200
rect 615460 75188 615466 75200
rect 646866 75188 646872 75200
rect 615460 75160 646872 75188
rect 615460 75148 615466 75160
rect 646866 75148 646872 75160
rect 646924 75148 646930 75200
rect 579522 71680 579528 71732
rect 579580 71720 579586 71732
rect 595438 71720 595444 71732
rect 579580 71692 595444 71720
rect 579580 71680 579586 71692
rect 595438 71680 595444 71692
rect 595496 71680 595502 71732
rect 579246 70252 579252 70304
rect 579304 70292 579310 70304
rect 581730 70292 581736 70304
rect 579304 70264 581736 70292
rect 579304 70252 579310 70264
rect 581730 70252 581736 70264
rect 581788 70252 581794 70304
rect 578694 68960 578700 69012
rect 578752 69000 578758 69012
rect 589918 69000 589924 69012
rect 578752 68972 589924 69000
rect 578752 68960 578758 68972
rect 589918 68960 589924 68972
rect 589976 68960 589982 69012
rect 579522 67532 579528 67584
rect 579580 67572 579586 67584
rect 588630 67572 588636 67584
rect 579580 67544 588636 67572
rect 579580 67532 579586 67544
rect 588630 67532 588636 67544
rect 588688 67532 588694 67584
rect 579522 65900 579528 65952
rect 579580 65940 579586 65952
rect 585870 65940 585876 65952
rect 579580 65912 585876 65940
rect 579580 65900 579586 65912
rect 585870 65900 585876 65912
rect 585928 65900 585934 65952
rect 578694 64812 578700 64864
rect 578752 64852 578758 64864
rect 588538 64852 588544 64864
rect 578752 64824 588544 64852
rect 578752 64812 578758 64824
rect 588538 64812 588544 64824
rect 588596 64812 588602 64864
rect 579522 63452 579528 63504
rect 579580 63492 579586 63504
rect 587158 63492 587164 63504
rect 579580 63464 587164 63492
rect 579580 63452 579586 63464
rect 587158 63452 587164 63464
rect 587216 63452 587222 63504
rect 617518 62132 617524 62144
rect 615466 62104 617524 62132
rect 578694 62024 578700 62076
rect 578752 62064 578758 62076
rect 585778 62064 585784 62076
rect 578752 62036 585784 62064
rect 578752 62024 578758 62036
rect 585778 62024 585784 62036
rect 585836 62024 585842 62076
rect 614758 62024 614764 62076
rect 614816 62064 614822 62076
rect 615466 62064 615494 62104
rect 617518 62092 617524 62104
rect 617576 62092 617582 62144
rect 614816 62036 615494 62064
rect 614816 62024 614822 62036
rect 578878 60664 578884 60716
rect 578936 60704 578942 60716
rect 584398 60704 584404 60716
rect 578936 60676 584404 60704
rect 578936 60664 578942 60676
rect 584398 60664 584404 60676
rect 584456 60664 584462 60716
rect 578878 58760 578884 58812
rect 578936 58800 578942 58812
rect 583018 58800 583024 58812
rect 578936 58772 583024 58800
rect 578936 58760 578942 58772
rect 583018 58760 583024 58772
rect 583076 58760 583082 58812
rect 578878 57876 578884 57928
rect 578936 57916 578942 57928
rect 581638 57916 581644 57928
rect 578936 57888 581644 57916
rect 578936 57876 578942 57888
rect 581638 57876 581644 57888
rect 581696 57876 581702 57928
rect 578326 57196 578332 57248
rect 578384 57236 578390 57248
rect 600958 57236 600964 57248
rect 578384 57208 600964 57236
rect 578384 57196 578390 57208
rect 600958 57196 600964 57208
rect 601016 57196 601022 57248
rect 621658 57196 621664 57248
rect 621716 57236 621722 57248
rect 662414 57236 662420 57248
rect 621716 57208 662420 57236
rect 621716 57196 621722 57208
rect 662414 57196 662420 57208
rect 662472 57196 662478 57248
rect 578234 55632 578240 55684
rect 578292 55672 578298 55684
rect 580258 55672 580264 55684
rect 578292 55644 580264 55672
rect 578292 55632 578298 55644
rect 580258 55632 580264 55644
rect 580316 55632 580322 55684
rect 405090 53116 405096 53168
rect 405148 53156 405154 53168
rect 608778 53156 608784 53168
rect 405148 53128 608784 53156
rect 405148 53116 405154 53128
rect 608778 53116 608784 53128
rect 608836 53116 608842 53168
rect 145374 53048 145380 53100
rect 145432 53088 145438 53100
rect 579062 53088 579068 53100
rect 145432 53060 579068 53088
rect 145432 53048 145438 53060
rect 579062 53048 579068 53060
rect 579120 53048 579126 53100
rect 52270 52436 52276 52488
rect 52328 52476 52334 52488
rect 346808 52476 346814 52488
rect 52328 52448 346814 52476
rect 52328 52436 52334 52448
rect 346808 52436 346814 52448
rect 346866 52476 346872 52488
rect 614758 52476 614764 52488
rect 346866 52448 614764 52476
rect 346866 52436 346872 52448
rect 614758 52436 614764 52448
rect 614816 52436 614822 52488
rect 478138 49716 478144 49768
rect 478196 49756 478202 49768
rect 478782 49756 478788 49768
rect 478196 49728 478788 49756
rect 478196 49716 478202 49728
rect 478782 49716 478788 49728
rect 478840 49716 478846 49768
rect 664254 49512 664260 49564
rect 664312 49552 664318 49564
rect 672074 49552 672080 49564
rect 664312 49524 672080 49552
rect 664312 49512 664318 49524
rect 672074 49512 672080 49524
rect 672132 49512 672138 49564
rect 194042 46180 194048 46232
rect 194100 46220 194106 46232
rect 661466 46220 661472 46232
rect 194100 46192 661472 46220
rect 194100 46180 194106 46192
rect 661466 46180 661472 46192
rect 661524 46180 661530 46232
rect 473170 42476 473176 42528
rect 473228 42476 473234 42528
rect 415118 42340 415124 42392
rect 415176 42340 415182 42392
<< via1 >>
rect 195336 1007088 195388 1007140
rect 203892 1007088 203944 1007140
rect 92612 1006544 92664 1006596
rect 99932 1006544 99984 1006596
rect 95976 1006476 96028 1006528
rect 104808 1006476 104860 1006528
rect 249064 1006476 249116 1006528
rect 258172 1006476 258224 1006528
rect 302884 1006476 302936 1006528
rect 308128 1006476 308180 1006528
rect 428372 1006476 428424 1006528
rect 93216 1006408 93268 1006460
rect 104348 1006408 104400 1006460
rect 253296 1006408 253348 1006460
rect 99104 1006340 99156 1006392
rect 126244 1006340 126296 1006392
rect 149704 1006340 149756 1006392
rect 150900 1006340 150952 1006392
rect 93124 1006272 93176 1006324
rect 100668 1006272 100720 1006324
rect 146944 1006272 146996 1006324
rect 154120 1006272 154172 1006324
rect 145564 1006204 145616 1006256
rect 151728 1006204 151780 1006256
rect 201868 1006340 201920 1006392
rect 228364 1006340 228416 1006392
rect 248328 1006340 248380 1006392
rect 254860 1006340 254912 1006392
rect 177304 1006272 177356 1006324
rect 195152 1006272 195204 1006324
rect 202696 1006272 202748 1006324
rect 207664 1006272 207716 1006324
rect 210056 1006272 210108 1006324
rect 301504 1006408 301556 1006460
rect 307300 1006408 307352 1006460
rect 358176 1006408 358228 1006460
rect 369124 1006408 369176 1006460
rect 427544 1006408 427596 1006460
rect 356060 1006340 356112 1006392
rect 380164 1006340 380216 1006392
rect 280804 1006272 280856 1006324
rect 298744 1006272 298796 1006324
rect 310612 1006272 310664 1006324
rect 357716 1006272 357768 1006324
rect 374644 1006272 374696 1006324
rect 504548 1006340 504600 1006392
rect 514208 1006340 514260 1006392
rect 196624 1006204 196676 1006256
rect 204352 1006204 204404 1006256
rect 249156 1006204 249208 1006256
rect 257344 1006204 257396 1006256
rect 300308 1006204 300360 1006256
rect 306472 1006204 306524 1006256
rect 358912 1006204 358964 1006256
rect 376024 1006204 376076 1006256
rect 445760 1006272 445812 1006324
rect 555976 1006272 556028 1006324
rect 456064 1006204 456116 1006256
rect 505376 1006204 505428 1006256
rect 514116 1006204 514168 1006256
rect 94688 1006136 94740 1006188
rect 103612 1006136 103664 1006188
rect 147036 1006136 147088 1006188
rect 152096 1006136 152148 1006188
rect 197360 1006136 197412 1006188
rect 98276 1006068 98328 1006120
rect 99104 1006068 99156 1006120
rect 102784 1006068 102836 1006120
rect 108856 1006068 108908 1006120
rect 154488 1006068 154540 1006120
rect 160652 1006068 160704 1006120
rect 198004 1006068 198056 1006120
rect 94504 1006000 94556 1006052
rect 103152 1006000 103204 1006052
rect 144184 1006000 144236 1006052
rect 150900 1006000 150952 1006052
rect 159088 1006000 159140 1006052
rect 162124 1006000 162176 1006052
rect 201040 1006068 201092 1006120
rect 201868 1006068 201920 1006120
rect 204996 1006136 205048 1006188
rect 210424 1006136 210476 1006188
rect 247684 1006136 247736 1006188
rect 255320 1006136 255372 1006188
rect 425152 1006136 425204 1006188
rect 449256 1006136 449308 1006188
rect 505008 1006136 505060 1006188
rect 516784 1006136 516836 1006188
rect 557172 1006136 557224 1006188
rect 565176 1006136 565228 1006188
rect 207204 1006068 207256 1006120
rect 209596 1006068 209648 1006120
rect 228456 1006068 228508 1006120
rect 248420 1006068 248472 1006120
rect 207572 1006000 207624 1006052
rect 252468 1006000 252520 1006052
rect 253296 1006000 253348 1006052
rect 254676 1006068 254728 1006120
rect 258540 1006068 258592 1006120
rect 303528 1006068 303580 1006120
rect 304080 1006068 304132 1006120
rect 304908 1006068 304960 1006120
rect 356888 1006068 356940 1006120
rect 360844 1006068 360896 1006120
rect 361396 1006068 361448 1006120
rect 368480 1006068 368532 1006120
rect 369124 1006068 369176 1006120
rect 380900 1006068 380952 1006120
rect 420828 1006068 420880 1006120
rect 422668 1006068 422720 1006120
rect 428004 1006068 428056 1006120
rect 465724 1006068 465776 1006120
rect 502524 1006068 502576 1006120
rect 256976 1006000 257028 1006052
rect 257344 1006000 257396 1006052
rect 259000 1006000 259052 1006052
rect 261024 1006000 261076 1006052
rect 269764 1006000 269816 1006052
rect 298836 1006000 298888 1006052
rect 305276 1006000 305328 1006052
rect 315120 1006000 315172 1006052
rect 319444 1006000 319496 1006052
rect 353116 1006000 353168 1006052
rect 354496 1006000 354548 1006052
rect 358544 1006000 358596 1006052
rect 362224 1006000 362276 1006052
rect 423496 1006000 423548 1006052
rect 426348 1006000 426400 1006052
rect 430028 1006000 430080 1006052
rect 468484 1006000 468536 1006052
rect 498108 1006000 498160 1006052
rect 499672 1006000 499724 1006052
rect 500500 1006000 500552 1006052
rect 504364 1006000 504416 1006052
rect 518900 1006000 518952 1006052
rect 549168 1006000 549220 1006052
rect 550272 1006000 550324 1006052
rect 551100 1006000 551152 1006052
rect 552296 1006000 552348 1006052
rect 556712 1006000 556764 1006052
rect 556804 1006000 556856 1006052
rect 570604 1006000 570656 1006052
rect 573364 1006000 573416 1006052
rect 143724 1005388 143776 1005440
rect 169024 1005388 169076 1005440
rect 361028 1005388 361080 1005440
rect 371884 1005388 371936 1005440
rect 360568 1005320 360620 1005372
rect 378784 1005320 378836 1005372
rect 360200 1005252 360252 1005304
rect 381544 1005252 381596 1005304
rect 426348 1005252 426400 1005304
rect 462964 1005252 463016 1005304
rect 503352 1005252 503404 1005304
rect 518992 1005252 519044 1005304
rect 508688 1005048 508740 1005100
rect 511264 1005048 511316 1005100
rect 507032 1004980 507084 1005032
rect 509792 1004980 509844 1005032
rect 508228 1004912 508280 1004964
rect 510620 1004912 510672 1004964
rect 159824 1004844 159876 1004896
rect 162308 1004844 162360 1004896
rect 363420 1004844 363472 1004896
rect 366364 1004844 366416 1004896
rect 159456 1004776 159508 1004828
rect 161480 1004776 161532 1004828
rect 208768 1004776 208820 1004828
rect 211804 1004776 211856 1004828
rect 304264 1004776 304316 1004828
rect 306932 1004776 306984 1004828
rect 313832 1004776 313884 1004828
rect 316040 1004776 316092 1004828
rect 364248 1004776 364300 1004828
rect 366548 1004776 366600 1004828
rect 499488 1004776 499540 1004828
rect 501328 1004776 501380 1004828
rect 507860 1004776 507912 1004828
rect 510068 1004776 510120 1004828
rect 160284 1004708 160336 1004760
rect 163504 1004708 163556 1004760
rect 209228 1004708 209280 1004760
rect 211160 1004708 211212 1004760
rect 305828 1004708 305880 1004760
rect 308588 1004708 308640 1004760
rect 314660 1004708 314712 1004760
rect 316684 1004708 316736 1004760
rect 354312 1004708 354364 1004760
rect 356888 1004708 356940 1004760
rect 361856 1004708 361908 1004760
rect 364984 1004708 365036 1004760
rect 499028 1004708 499080 1004760
rect 500868 1004708 500920 1004760
rect 509056 1004708 509108 1004760
rect 510712 1004708 510764 1004760
rect 556344 1004708 556396 1004760
rect 559748 1004708 559800 1004760
rect 94596 1004640 94648 1004692
rect 103152 1004640 103204 1004692
rect 160652 1004640 160704 1004692
rect 162952 1004640 163004 1004692
rect 199384 1004640 199436 1004692
rect 202236 1004640 202288 1004692
rect 208400 1004640 208452 1004692
rect 209780 1004640 209832 1004692
rect 305644 1004640 305696 1004692
rect 307760 1004640 307812 1004692
rect 315488 1004640 315540 1004692
rect 318064 1004640 318116 1004692
rect 354588 1004640 354640 1004692
rect 356060 1004640 356112 1004692
rect 362592 1004640 362644 1004692
rect 365168 1004640 365220 1004692
rect 499212 1004640 499264 1004692
rect 500500 1004640 500552 1004692
rect 507400 1004640 507452 1004692
rect 509240 1004640 509292 1004692
rect 557632 1004640 557684 1004692
rect 559564 1004640 559616 1004692
rect 298928 1004572 298980 1004624
rect 308956 1004572 309008 1004624
rect 422024 1004572 422076 1004624
rect 423864 1004572 423916 1004624
rect 424692 1004028 424744 1004080
rect 451280 1004028 451332 1004080
rect 423496 1003892 423548 1003944
rect 454316 1003892 454368 1003944
rect 503720 1003892 503772 1003944
rect 519268 1003892 519320 1003944
rect 92520 1003280 92572 1003332
rect 99472 1003280 99524 1003332
rect 380900 1003280 380952 1003332
rect 383568 1003280 383620 1003332
rect 553400 1003280 553452 1003332
rect 554688 1003280 554740 1003332
rect 445760 1003212 445812 1003264
rect 449808 1003212 449860 1003264
rect 553952 1002600 554004 1002652
rect 564992 1002600 565044 1002652
rect 144092 1002532 144144 1002584
rect 154580 1002532 154632 1002584
rect 354588 1002532 354640 1002584
rect 359188 1002532 359240 1002584
rect 425980 1002532 426032 1002584
rect 469312 1002532 469364 1002584
rect 554320 1002532 554372 1002584
rect 567292 1002532 567344 1002584
rect 559196 1002396 559248 1002448
rect 562508 1002396 562560 1002448
rect 106832 1002328 106884 1002380
rect 109868 1002328 109920 1002380
rect 560852 1002328 560904 1002380
rect 565084 1002328 565136 1002380
rect 106188 1002260 106240 1002312
rect 108488 1002260 108540 1002312
rect 261852 1002260 261904 1002312
rect 264244 1002260 264296 1002312
rect 558460 1002260 558512 1002312
rect 560944 1002260 560996 1002312
rect 95884 1002192 95936 1002244
rect 101496 1002192 101548 1002244
rect 106004 1002192 106056 1002244
rect 108304 1002192 108356 1002244
rect 158260 1002192 158312 1002244
rect 160744 1002192 160796 1002244
rect 202144 1002192 202196 1002244
rect 205180 1002192 205232 1002244
rect 211620 1002192 211672 1002244
rect 215944 1002192 215996 1002244
rect 252468 1002192 252520 1002244
rect 254492 1002192 254544 1002244
rect 261484 1002192 261536 1002244
rect 263600 1002192 263652 1002244
rect 559656 1002192 559708 1002244
rect 561772 1002192 561824 1002244
rect 97356 1002124 97408 1002176
rect 102324 1002124 102376 1002176
rect 105636 1002124 105688 1002176
rect 107936 1002124 107988 1002176
rect 108028 1002124 108080 1002176
rect 110512 1002124 110564 1002176
rect 157800 1002124 157852 1002176
rect 160192 1002124 160244 1002176
rect 200948 1002124 201000 1002176
rect 203524 1002124 203576 1002176
rect 210424 1002124 210476 1002176
rect 213184 1002124 213236 1002176
rect 253756 1002124 253808 1002176
rect 256148 1002124 256200 1002176
rect 260840 1002124 260892 1002176
rect 261852 1002124 261904 1002176
rect 262680 1002124 262732 1002176
rect 265808 1002124 265860 1002176
rect 550272 1002124 550324 1002176
rect 553124 1002124 553176 1002176
rect 560484 1002124 560536 1002176
rect 563060 1002124 563112 1002176
rect 97264 1002056 97316 1002108
rect 100300 1002056 100352 1002108
rect 107660 1002056 107712 1002108
rect 109592 1002056 109644 1002108
rect 157432 1002056 157484 1002108
rect 159364 1002056 159416 1002108
rect 203708 1002056 203760 1002108
rect 205916 1002056 205968 1002108
rect 211252 1002056 211304 1002108
rect 213368 1002056 213420 1002108
rect 253848 1002056 253900 1002108
rect 255688 1002056 255740 1002108
rect 259828 1002056 259880 1002108
rect 261484 1002056 261536 1002108
rect 263508 1002056 263560 1002108
rect 267004 1002056 267056 1002108
rect 310152 1002056 310204 1002108
rect 311900 1002056 311952 1002108
rect 365076 1002056 365128 1002108
rect 367928 1002056 367980 1002108
rect 423312 1002056 423364 1002108
rect 425980 1002056 426032 1002108
rect 502156 1002056 502208 1002108
rect 503720 1002056 503772 1002108
rect 509516 1002056 509568 1002108
rect 514024 1002056 514076 1002108
rect 550364 1002056 550416 1002108
rect 552296 1002056 552348 1002108
rect 560024 1002056 560076 1002108
rect 562324 1002056 562376 1002108
rect 92336 1001988 92388 1002040
rect 92612 1001988 92664 1002040
rect 98644 1001988 98696 1002040
rect 101128 1001988 101180 1002040
rect 104348 1001988 104400 1002040
rect 106648 1001988 106700 1002040
rect 107200 1001988 107252 1002040
rect 109040 1001988 109092 1002040
rect 109684 1001988 109736 1002040
rect 111800 1001988 111852 1002040
rect 158628 1001988 158680 1002040
rect 160100 1001988 160152 1002040
rect 200304 1001988 200356 1002040
rect 203064 1001988 203116 1002040
rect 203524 1001988 203576 1002040
rect 205548 1001988 205600 1002040
rect 212540 1001988 212592 1002040
rect 214564 1001988 214616 1002040
rect 260196 1001988 260248 1002040
rect 262864 1001988 262916 1002040
rect 263048 1001988 263100 1002040
rect 265624 1001988 265676 1002040
rect 300124 1001988 300176 1002040
rect 306104 1001988 306156 1002040
rect 307024 1001988 307076 1002040
rect 309324 1001988 309376 1002040
rect 312268 1001988 312320 1002040
rect 314660 1001988 314712 1002040
rect 357164 1001988 357216 1002040
rect 359372 1001988 359424 1002040
rect 365904 1001988 365956 1002040
rect 369124 1001988 369176 1002040
rect 424968 1001988 425020 1002040
rect 426348 1001988 426400 1002040
rect 505836 1001988 505888 1002040
rect 508688 1001988 508740 1002040
rect 509884 1001988 509936 1002040
rect 512828 1001988 512880 1002040
rect 550456 1001988 550508 1002040
rect 552664 1001988 552716 1002040
rect 553124 1001988 553176 1002040
rect 555148 1001988 555200 1002040
rect 558000 1001988 558052 1002040
rect 560576 1001988 560628 1002040
rect 561680 1001988 561732 1002040
rect 563704 1001988 563756 1002040
rect 100024 1001920 100076 1001972
rect 101956 1001920 102008 1001972
rect 106464 1001920 106516 1001972
rect 107752 1001920 107804 1001972
rect 108488 1001920 108540 1001972
rect 111064 1001920 111116 1001972
rect 156972 1001920 157024 1001972
rect 158720 1001920 158772 1001972
rect 195152 1001920 195204 1001972
rect 197360 1001920 197412 1001972
rect 202328 1001920 202380 1001972
rect 204720 1001920 204772 1001972
rect 204904 1001920 204956 1001972
rect 206744 1001920 206796 1001972
rect 212080 1001920 212132 1001972
rect 213920 1001920 213972 1001972
rect 251824 1001920 251876 1001972
rect 254124 1001920 254176 1001972
rect 254584 1001920 254636 1001972
rect 256516 1001920 256568 1001972
rect 260656 1001920 260708 1001972
rect 262220 1001920 262272 1001972
rect 263876 1001920 263928 1001972
rect 267096 1001920 267148 1001972
rect 300216 1001920 300268 1001972
rect 305736 1001920 305788 1001972
rect 311440 1001920 311492 1001972
rect 313556 1001920 313608 1001972
rect 357348 1001920 357400 1001972
rect 358912 1001920 358964 1001972
rect 365444 1001920 365496 1001972
rect 367744 1001920 367796 1001972
rect 420828 1001920 420880 1001972
rect 421472 1001920 421524 1001972
rect 423404 1001920 423456 1001972
rect 425152 1001920 425204 1001972
rect 425704 1001920 425756 1001972
rect 426808 1001920 426860 1001972
rect 506204 1001920 506256 1001972
rect 508504 1001920 508556 1001972
rect 510344 1001920 510396 1001972
rect 512644 1001920 512696 1001972
rect 549076 1001920 549128 1001972
rect 551468 1001920 551520 1001972
rect 551928 1001920 551980 1001972
rect 553492 1001920 553544 1001972
rect 558828 1001920 558880 1001972
rect 560300 1001920 560352 1001972
rect 561312 1001920 561364 1001972
rect 563888 1001920 563940 1001972
rect 298376 1001852 298428 1001904
rect 310152 1001852 310204 1001904
rect 518900 1001852 518952 1001904
rect 523868 1001852 523920 1001904
rect 449256 1001784 449308 1001836
rect 452568 1001784 452620 1001836
rect 424968 1001240 425020 1001292
rect 447140 1001240 447192 1001292
rect 92428 1001172 92480 1001224
rect 98644 1001172 98696 1001224
rect 195428 1001172 195480 1001224
rect 200948 1001172 201000 1001224
rect 423312 1001172 423364 1001224
rect 469220 1001172 469272 1001224
rect 299388 1000560 299440 1000612
rect 302884 1000560 302936 1000612
rect 92704 1000492 92756 1000544
rect 94688 1000492 94740 1000544
rect 152740 1000492 152792 1000544
rect 154948 1000492 155000 1000544
rect 298560 1000492 298612 1000544
rect 300308 1000492 300360 1000544
rect 611360 1000492 611412 1000544
rect 625712 1000492 625764 1000544
rect 514208 1000424 514260 1000476
rect 520188 1000424 520240 1000476
rect 451280 1000220 451332 1000272
rect 459560 1000220 459612 1000272
rect 247040 999948 247092 1000000
rect 252468 999948 252520 1000000
rect 551928 999812 551980 999864
rect 568212 999812 568264 999864
rect 143816 999744 143868 999796
rect 155776 999744 155828 999796
rect 428832 999744 428884 999796
rect 469404 999744 469456 999796
rect 499488 999744 499540 999796
rect 504272 999744 504324 999796
rect 508688 999744 508740 999796
rect 513932 999744 513984 999796
rect 550272 999744 550324 999796
rect 567936 999744 567988 999796
rect 247132 999472 247184 999524
rect 253756 999472 253808 999524
rect 249708 999132 249760 999184
rect 254676 999132 254728 999184
rect 469312 999132 469364 999184
rect 472072 999132 472124 999184
rect 92336 999064 92388 999116
rect 94596 999064 94648 999116
rect 250720 999064 250772 999116
rect 253848 999064 253900 999116
rect 514116 999064 514168 999116
rect 520096 999064 520148 999116
rect 357164 998996 357216 999048
rect 361580 998996 361632 999048
rect 469220 998860 469272 998912
rect 472256 998860 472308 998912
rect 516784 998656 516836 998708
rect 524052 998656 524104 998708
rect 452568 998588 452620 998640
rect 459652 998588 459704 998640
rect 499028 998588 499080 998640
rect 516876 998588 516928 998640
rect 423404 998520 423456 998572
rect 472164 998520 472216 998572
rect 499212 998520 499264 998572
rect 516968 998520 517020 998572
rect 368480 998452 368532 998504
rect 383384 998452 383436 998504
rect 425704 998452 425756 998504
rect 472624 998452 472676 998504
rect 504364 998452 504416 998504
rect 522396 998452 522448 998504
rect 360844 998384 360896 998436
rect 380900 998384 380952 998436
rect 422024 998384 422076 998436
rect 465724 998384 465776 998436
rect 472532 998384 472584 998436
rect 502156 998384 502208 998436
rect 524052 998384 524104 998436
rect 549076 998384 549128 998436
rect 572720 998384 572772 998436
rect 472348 998180 472400 998232
rect 430856 998112 430908 998164
rect 433984 998112 434036 998164
rect 149060 998044 149112 998096
rect 152924 998044 152976 998096
rect 431684 998044 431736 998096
rect 434168 998044 434220 998096
rect 148324 997976 148376 998028
rect 151268 997976 151320 998028
rect 429660 997976 429712 998028
rect 431960 997976 432012 998028
rect 151084 997908 151136 997960
rect 153752 997908 153804 997960
rect 246672 997908 246724 997960
rect 248420 997908 248472 997960
rect 428464 997908 428516 997960
rect 430856 997908 430908 997960
rect 432880 997908 432932 997960
rect 436744 997908 436796 997960
rect 518992 997908 519044 997960
rect 523960 997908 524012 997960
rect 92612 997840 92664 997892
rect 94504 997840 94556 997892
rect 150348 997840 150400 997892
rect 152556 997840 152608 997892
rect 298284 997840 298336 997892
rect 151268 997772 151320 997824
rect 153384 997772 153436 997824
rect 246764 997772 246816 997824
rect 253664 997772 253716 997824
rect 303252 997772 303304 997824
rect 305828 997772 305880 997824
rect 430396 997840 430448 997892
rect 432144 997840 432196 997892
rect 432420 997840 432472 997892
rect 435548 997840 435600 997892
rect 328368 997772 328420 997824
rect 378784 997772 378836 997824
rect 383476 997772 383528 997824
rect 429200 997772 429252 997824
rect 431224 997772 431276 997824
rect 432052 997772 432104 997824
rect 433340 997772 433392 997824
rect 109868 997704 109920 997756
rect 117228 997704 117280 997756
rect 160744 997704 160796 997756
rect 167552 997704 167604 997756
rect 195244 997704 195296 997756
rect 211160 997704 211212 997756
rect 213368 997704 213420 997756
rect 218888 997704 218940 997756
rect 246580 997704 246632 997756
rect 260840 997704 260892 997756
rect 265808 997704 265860 997756
rect 270408 997704 270460 997756
rect 298744 997704 298796 997756
rect 316040 997704 316092 997756
rect 362224 997704 362276 997756
rect 372344 997704 372396 997756
rect 399944 997704 399996 997756
rect 433432 997704 433484 997756
rect 434168 997704 434220 997756
rect 439688 997704 439740 997756
rect 488908 997704 488960 997756
rect 510712 997704 510764 997756
rect 513932 997704 513984 997756
rect 516692 997704 516744 997756
rect 540888 997704 540940 997756
rect 563060 997704 563112 997756
rect 567292 997704 567344 997756
rect 625804 997772 625856 997824
rect 111064 997636 111116 997688
rect 116308 997636 116360 997688
rect 144828 997636 144880 997688
rect 160192 997636 160244 997688
rect 162308 997636 162360 997688
rect 167644 997636 167696 997688
rect 201408 997636 201460 997688
rect 203708 997636 203760 997688
rect 366548 997636 366600 997688
rect 372436 997636 372488 997688
rect 400036 997636 400088 997688
rect 432144 997636 432196 997688
rect 511264 997636 511316 997688
rect 516784 997636 516836 997688
rect 568212 997636 568264 997688
rect 611360 997636 611412 997688
rect 144736 997568 144788 997620
rect 161480 997568 161532 997620
rect 365168 997568 365220 997620
rect 372528 997568 372580 997620
rect 550364 997568 550416 997620
rect 564992 997500 565044 997552
rect 565176 997432 565228 997484
rect 590476 997480 590528 997532
rect 590568 997392 590620 997444
rect 144000 997296 144052 997348
rect 147036 997296 147088 997348
rect 202052 997296 202104 997348
rect 204904 997296 204956 997348
rect 590384 997284 590436 997336
rect 200212 997228 200264 997280
rect 204996 997228 205048 997280
rect 573364 997160 573416 997212
rect 620284 997160 620336 997212
rect 559748 997092 559800 997144
rect 618168 997092 618220 997144
rect 328368 997024 328420 997076
rect 381176 997024 381228 997076
rect 550456 997024 550508 997076
rect 622400 997024 622452 997076
rect 195244 996820 195296 996872
rect 199384 996820 199436 996872
rect 195980 996752 196032 996804
rect 202328 996752 202380 996804
rect 303252 996412 303304 996464
rect 304264 996412 304316 996464
rect 299296 996344 299348 996396
rect 305644 996344 305696 996396
rect 159364 996140 159416 996192
rect 209780 996140 209832 996192
rect 262864 996140 262916 996192
rect 313556 996140 313608 996192
rect 364984 996140 365036 996192
rect 431960 996140 432012 996192
rect 433984 996140 434036 996192
rect 510620 996140 510672 996192
rect 556712 996140 556764 996192
rect 108304 996072 108356 996124
rect 158720 996072 158772 996124
rect 162124 996072 162176 996124
rect 207664 996072 207716 996124
rect 211804 996072 211856 996124
rect 261484 996072 261536 996124
rect 264244 996072 264296 996124
rect 313372 996072 313424 996124
rect 366364 996072 366416 996124
rect 428464 996072 428516 996124
rect 431224 996072 431276 996124
rect 506572 996072 506624 996124
rect 508504 996072 508556 996124
rect 560576 996072 560628 996124
rect 109592 996004 109644 996056
rect 160100 996004 160152 996056
rect 228456 996004 228508 996056
rect 262220 996004 262272 996056
rect 269764 996004 269816 996056
rect 314660 996004 314712 996056
rect 361580 996004 361632 996056
rect 150348 995868 150400 995920
rect 213184 995868 213236 995920
rect 263600 995868 263652 995920
rect 298928 995936 298980 995988
rect 298468 995868 298520 995920
rect 468484 996004 468536 996056
rect 509240 996004 509292 996056
rect 510068 996004 510120 996056
rect 561772 996004 561824 996056
rect 504272 995936 504324 995988
rect 472348 995868 472400 995920
rect 509792 995868 509844 995920
rect 85304 995800 85356 995852
rect 92244 995800 92296 995852
rect 139216 995800 139268 995852
rect 140504 995800 140556 995852
rect 143724 995800 143776 995852
rect 192484 995800 192536 995852
rect 195152 995800 195204 995852
rect 242072 995800 242124 995852
rect 247684 995800 247736 995852
rect 290648 995800 290700 995852
rect 291108 995800 291160 995852
rect 292488 995800 292540 995852
rect 298836 995800 298888 995852
rect 383384 995800 383436 995852
rect 385684 995800 385736 995852
rect 391756 995800 391808 995852
rect 472532 995800 472584 995852
rect 473360 995800 473412 995852
rect 478236 995800 478288 995852
rect 523960 995800 524012 995852
rect 525340 995800 525392 995852
rect 91560 995732 91612 995784
rect 92336 995732 92388 995784
rect 141056 995732 141108 995784
rect 143816 995732 143868 995784
rect 190460 995732 190512 995784
rect 195336 995732 195388 995784
rect 245568 995732 245620 995784
rect 246672 995732 246724 995784
rect 297272 995732 297324 995784
rect 298048 995732 298100 995784
rect 383640 995732 383692 995784
rect 384396 995732 384448 995784
rect 432052 995732 432104 995784
rect 439780 995732 439832 995784
rect 472440 995732 472492 995784
rect 474740 995732 474792 995784
rect 524144 995732 524196 995784
rect 524788 995732 524840 995784
rect 533436 995800 533488 995852
rect 560300 995868 560352 995920
rect 557540 995800 557592 995852
rect 568212 995800 568264 995852
rect 634728 995800 634780 995852
rect 625804 995732 625856 995784
rect 627184 995732 627236 995784
rect 87880 995664 87932 995716
rect 92428 995664 92480 995716
rect 136272 995664 136324 995716
rect 144092 995664 144144 995716
rect 235264 995664 235316 995716
rect 247132 995664 247184 995716
rect 294880 995664 294932 995716
rect 298284 995664 298336 995716
rect 383732 995664 383784 995716
rect 388628 995664 388680 995716
rect 472256 995664 472308 995716
rect 474004 995664 474056 995716
rect 523868 995664 523920 995716
rect 529020 995664 529072 995716
rect 625712 995664 625764 995716
rect 630864 995664 630916 995716
rect 169024 995596 169076 995648
rect 184296 995596 184348 995648
rect 240876 995596 240928 995648
rect 246764 995596 246816 995648
rect 295432 995596 295484 995648
rect 298376 995596 298428 995648
rect 472164 995596 472216 995648
rect 477684 995596 477736 995648
rect 472072 995528 472124 995580
rect 476948 995528 477000 995580
rect 288072 995460 288124 995512
rect 300124 995460 300176 995512
rect 286784 995392 286836 995444
rect 299296 995392 299348 995444
rect 81256 995324 81308 995376
rect 95884 995324 95936 995376
rect 287520 995324 287572 995376
rect 301504 995324 301556 995376
rect 78312 995256 78364 995308
rect 95976 995256 96028 995308
rect 133420 995256 133472 995308
rect 145564 995256 145616 995308
rect 239266 995256 239318 995308
rect 251824 995256 251876 995308
rect 359188 995256 359240 995308
rect 392676 995256 392728 995308
rect 572720 995256 572772 995308
rect 636154 995256 636206 995308
rect 80704 995188 80756 995240
rect 100024 995188 100076 995240
rect 184158 995188 184210 995240
rect 196624 995188 196676 995240
rect 235586 995188 235638 995240
rect 250720 995188 250772 995240
rect 284116 995188 284168 995240
rect 298652 995188 298704 995240
rect 567936 995188 567988 995240
rect 637350 995188 637402 995240
rect 77668 995120 77720 995172
rect 97356 995120 97408 995172
rect 129096 995120 129148 995172
rect 151084 995120 151136 995172
rect 187608 995120 187660 995172
rect 201408 995120 201460 995172
rect 231584 995120 231636 995172
rect 249064 995120 249116 995172
rect 283472 995120 283524 995172
rect 299388 995120 299440 995172
rect 354312 995120 354364 995172
rect 393228 995120 393280 995172
rect 520096 995120 520148 995172
rect 537392 995120 537444 995172
rect 570604 995120 570656 995172
rect 638960 995120 639012 995172
rect 77024 995052 77076 995104
rect 106648 995052 106700 995104
rect 129740 995052 129792 995104
rect 155224 995052 155276 995104
rect 181444 995052 181496 995104
rect 198004 995052 198056 995104
rect 232228 995052 232280 995104
rect 254584 995052 254636 995104
rect 282828 995052 282880 995104
rect 311900 995052 311952 995104
rect 371884 995052 371936 995104
rect 397000 995052 397052 995104
rect 501972 995052 502024 995104
rect 528744 995052 528796 995104
rect 553124 995052 553176 995104
rect 633992 995052 634044 995104
rect 88708 994984 88760 995036
rect 121736 994984 121788 995036
rect 180708 994984 180760 995036
rect 202144 994984 202196 995036
rect 243268 994984 243320 995036
rect 316408 994984 316460 995036
rect 357348 994984 357400 995036
rect 398840 994984 398892 995036
rect 447140 994984 447192 995036
rect 487804 994984 487856 995036
rect 501696 994984 501748 995036
rect 535552 994984 535604 995036
rect 553400 994984 553452 995036
rect 640708 995052 640760 995104
rect 638868 994984 638920 995036
rect 640800 994984 640852 995036
rect 319444 992944 319496 992996
rect 332600 992944 332652 992996
rect 367928 992944 367980 992996
rect 429936 992944 429988 992996
rect 562508 992944 562560 992996
rect 661684 992944 661736 992996
rect 48964 992876 49016 992928
rect 110512 992876 110564 992928
rect 215300 992876 215352 992928
rect 251456 992876 251508 992928
rect 265624 992876 265676 992928
rect 300032 992876 300084 992928
rect 316684 992876 316736 992928
rect 364984 992876 365036 992928
rect 420828 992876 420880 992928
rect 666744 992876 666796 992928
rect 47584 991516 47636 991568
rect 107752 991516 107804 991568
rect 512828 991516 512880 991568
rect 527640 991516 527692 991568
rect 559564 991516 559616 991568
rect 660304 991516 660356 991568
rect 44824 991448 44876 991500
rect 109040 991448 109092 991500
rect 138296 991448 138348 991500
rect 162952 991448 163004 991500
rect 203156 991448 203208 991500
rect 213920 991448 213972 991500
rect 367744 991448 367796 991500
rect 397828 991448 397880 991500
rect 435548 991448 435600 991500
rect 495164 991448 495216 991500
rect 498108 991448 498160 991500
rect 666560 991448 666612 991500
rect 214564 991176 214616 991228
rect 219440 991176 219492 991228
rect 184296 990836 184348 990888
rect 186964 990836 187016 990888
rect 267096 990836 267148 990888
rect 268752 990836 268804 990888
rect 560944 990224 560996 990276
rect 658924 990224 658976 990276
rect 562324 990156 562376 990208
rect 669964 990156 670016 990208
rect 50344 990088 50396 990140
rect 107936 990088 107988 990140
rect 353116 990088 353168 990140
rect 666836 990088 666888 990140
rect 512644 988728 512696 988780
rect 543832 988728 543884 988780
rect 563888 988728 563940 988780
rect 592500 988728 592552 988780
rect 435364 987368 435416 987420
rect 478972 987368 479024 987420
rect 563704 987368 563756 987420
rect 608784 987368 608836 987420
rect 267004 986620 267056 986672
rect 268108 986620 268160 986672
rect 89628 986008 89680 986060
rect 111800 986008 111852 986060
rect 73436 985940 73488 985992
rect 102784 985940 102836 985992
rect 215944 985940 215996 985992
rect 235632 985940 235684 985992
rect 268752 985940 268804 985992
rect 284300 985940 284352 985992
rect 318064 985940 318116 985992
rect 349160 985940 349212 985992
rect 369124 985940 369176 985992
rect 414112 985940 414164 985992
rect 436744 985940 436796 985992
rect 462780 985940 462832 985992
rect 514024 985940 514076 985992
rect 560116 985940 560168 985992
rect 565084 985940 565136 985992
rect 624976 985940 625028 985992
rect 163504 985872 163556 985924
rect 170772 985872 170824 985924
rect 549168 984920 549220 984972
rect 666652 984920 666704 984972
rect 303528 984852 303580 984904
rect 665456 984852 665508 984904
rect 280804 984784 280856 984836
rect 650092 984784 650144 984836
rect 228364 984716 228416 984768
rect 651472 984716 651524 984768
rect 177304 984648 177356 984700
rect 650000 984648 650052 984700
rect 126244 984580 126296 984632
rect 651380 984580 651432 984632
rect 42708 975672 42760 975724
rect 62120 975672 62172 975724
rect 651656 975672 651708 975724
rect 671344 975672 671396 975724
rect 42156 967240 42208 967292
rect 42708 967240 42760 967292
rect 42156 963976 42208 964028
rect 42800 963976 42852 964028
rect 42156 962820 42208 962872
rect 42892 962820 42944 962872
rect 674840 962684 674892 962736
rect 675484 962684 675536 962736
rect 675024 962004 675076 962056
rect 675392 962004 675444 962056
rect 47676 961868 47728 961920
rect 62120 961868 62172 961920
rect 42064 959692 42116 959744
rect 44180 959692 44232 959744
rect 42156 959080 42208 959132
rect 42984 959080 43036 959132
rect 673276 958332 673328 958384
rect 675392 958332 675444 958384
rect 659016 957788 659068 957840
rect 674840 957788 674892 957840
rect 674748 956972 674800 957024
rect 675392 956972 675444 957024
rect 672356 956496 672408 956548
rect 675024 956496 675076 956548
rect 674564 955680 674616 955732
rect 675484 955680 675536 955732
rect 42340 955544 42392 955596
rect 42708 955544 42760 955596
rect 674840 955476 674892 955528
rect 675484 955476 675536 955528
rect 42248 954252 42300 954304
rect 42708 954252 42760 954304
rect 36544 952212 36596 952264
rect 42340 952212 42392 952264
rect 675760 952008 675812 952060
rect 675760 951736 675812 951788
rect 31024 951464 31076 951516
rect 41880 951464 41932 951516
rect 675760 949424 675812 949476
rect 678244 949424 678296 949476
rect 651564 948064 651616 948116
rect 674196 948064 674248 948116
rect 34520 945956 34572 946008
rect 62120 945956 62172 946008
rect 35808 943236 35860 943288
rect 48412 943236 48464 943288
rect 35716 943168 35768 943220
rect 47676 943168 47728 943220
rect 41788 941808 41840 941860
rect 42064 941808 42116 941860
rect 652024 939768 652076 939820
rect 676036 939768 676088 939820
rect 674196 939156 674248 939208
rect 676036 939156 676088 939208
rect 671344 938680 671396 938732
rect 676220 938680 676272 938732
rect 669964 938544 670016 938596
rect 676036 938544 676088 938596
rect 661684 937320 661736 937372
rect 676220 937320 676272 937372
rect 658924 937184 658976 937236
rect 676220 937184 676272 937236
rect 672632 937116 672684 937168
rect 676128 937116 676180 937168
rect 673184 937048 673236 937100
rect 676036 937048 676088 937100
rect 48412 936980 48464 937032
rect 62120 936980 62172 937032
rect 651564 936980 651616 937032
rect 659016 936980 659068 937032
rect 673644 936640 673696 936692
rect 676036 936640 676088 936692
rect 674656 935824 674708 935876
rect 676036 935824 676088 935876
rect 660304 935620 660356 935672
rect 676220 935620 676272 935672
rect 39948 932084 40000 932136
rect 41880 932084 41932 932136
rect 674564 931948 674616 932000
rect 676220 931948 676272 932000
rect 673276 930248 673328 930300
rect 676220 930248 676272 930300
rect 669964 927392 670016 927444
rect 683120 927392 683172 927444
rect 51724 923244 51776 923296
rect 62120 923244 62172 923296
rect 651564 921816 651616 921868
rect 664444 921816 664496 921868
rect 40684 909440 40736 909492
rect 62120 909440 62172 909492
rect 651564 909440 651616 909492
rect 661684 909440 661736 909492
rect 53104 896996 53156 897048
rect 62120 896996 62172 897048
rect 651564 895636 651616 895688
rect 660304 895636 660356 895688
rect 44824 884620 44876 884672
rect 62120 884620 62172 884672
rect 671988 879044 672040 879096
rect 675300 879044 675352 879096
rect 673092 873536 673144 873588
rect 675392 873536 675444 873588
rect 55956 870816 56008 870868
rect 62120 870816 62172 870868
rect 674380 869796 674432 869848
rect 675392 869796 675444 869848
rect 673000 869592 673052 869644
rect 675392 869592 675444 869644
rect 651564 869388 651616 869440
rect 671344 869388 671396 869440
rect 672908 868980 672960 869032
rect 675392 868980 675444 869032
rect 652024 868640 652076 868692
rect 674932 868640 674984 868692
rect 674564 868028 674616 868080
rect 675392 868028 675444 868080
rect 674472 866804 674524 866856
rect 675392 866804 675444 866856
rect 674932 866192 674984 866244
rect 675392 866192 675444 866244
rect 672816 862792 672868 862844
rect 675484 862792 675536 862844
rect 43628 858372 43680 858424
rect 62120 858372 62172 858424
rect 652576 855584 652628 855636
rect 672724 855584 672776 855636
rect 54484 844568 54536 844620
rect 62120 844568 62172 844620
rect 651564 841780 651616 841832
rect 663064 841780 663116 841832
rect 50436 832124 50488 832176
rect 62120 832124 62172 832176
rect 651564 829404 651616 829456
rect 659016 829404 659068 829456
rect 47584 818320 47636 818372
rect 62120 818320 62172 818372
rect 41328 817504 41380 817556
rect 44824 817504 44876 817556
rect 41236 817368 41288 817420
rect 53104 817368 53156 817420
rect 651564 815600 651616 815652
rect 665824 815600 665876 815652
rect 41512 814852 41564 814904
rect 41788 814852 41840 814904
rect 35808 806420 35860 806472
rect 41880 806420 41932 806472
rect 50344 805944 50396 805996
rect 62120 805944 62172 805996
rect 42156 803836 42208 803888
rect 42616 803836 42668 803888
rect 42064 803768 42116 803820
rect 42708 803768 42760 803820
rect 651564 803156 651616 803208
rect 658924 803156 658976 803208
rect 35256 801116 35308 801168
rect 43076 801116 43128 801168
rect 32404 801048 32456 801100
rect 42892 801048 42944 801100
rect 40684 800504 40736 800556
rect 42984 800504 43036 800556
rect 42156 799960 42208 800012
rect 42340 799960 42392 800012
rect 51724 799688 51776 799740
rect 42708 799076 42760 799128
rect 42156 798124 42208 798176
rect 42616 798124 42668 798176
rect 42156 797240 42208 797292
rect 42708 797240 42760 797292
rect 42156 796288 42208 796340
rect 42708 796288 42760 796340
rect 42156 794996 42208 795048
rect 42432 794996 42484 795048
rect 42432 794860 42484 794912
rect 42984 794860 43036 794912
rect 43168 794860 43220 794912
rect 44456 794860 44508 794912
rect 42156 794248 42208 794300
rect 42708 794248 42760 794300
rect 42156 793772 42208 793824
rect 43168 793772 43220 793824
rect 44824 793500 44876 793552
rect 62120 793500 62172 793552
rect 42156 793160 42208 793212
rect 42432 793160 42484 793212
rect 42432 793024 42484 793076
rect 44364 793024 44416 793076
rect 42156 790644 42208 790696
rect 42708 790644 42760 790696
rect 42156 790100 42208 790152
rect 42432 790100 42484 790152
rect 42156 789420 42208 789472
rect 42340 789420 42392 789472
rect 651656 789352 651708 789404
rect 661776 789352 661828 789404
rect 674288 787312 674340 787364
rect 675392 787312 675444 787364
rect 42064 786428 42116 786480
rect 42432 786428 42484 786480
rect 42156 785612 42208 785664
rect 42708 785612 42760 785664
rect 674196 784252 674248 784304
rect 675392 784252 675444 784304
rect 674012 782892 674064 782944
rect 675484 782892 675536 782944
rect 671896 780716 671948 780768
rect 675484 780716 675536 780768
rect 673276 779968 673328 780020
rect 675484 779968 675536 780020
rect 51724 779696 51776 779748
rect 62120 779696 62172 779748
rect 672540 779288 672592 779340
rect 675392 779288 675444 779340
rect 659016 778948 659068 779000
rect 674748 778948 674800 779000
rect 673736 778608 673788 778660
rect 675484 778608 675536 778660
rect 673920 777316 673972 777368
rect 675392 777316 675444 777368
rect 674748 777044 674800 777096
rect 675392 777044 675444 777096
rect 651564 775548 651616 775600
rect 659016 775548 659068 775600
rect 670516 775548 670568 775600
rect 675392 775548 675444 775600
rect 35808 774188 35860 774240
rect 54484 774188 54536 774240
rect 672448 773576 672500 773628
rect 675484 773576 675536 773628
rect 48964 767320 49016 767372
rect 62120 767320 62172 767372
rect 675208 766572 675260 766624
rect 675668 766572 675720 766624
rect 651564 763172 651616 763224
rect 664536 763172 664588 763224
rect 41512 761744 41564 761796
rect 55864 761744 55916 761796
rect 664444 760792 664496 760844
rect 676220 760792 676272 760844
rect 661684 760656 661736 760708
rect 676128 760656 676180 760708
rect 660304 760520 660356 760572
rect 676036 760520 676088 760572
rect 31024 759636 31076 759688
rect 41880 759636 41932 759688
rect 672632 759296 672684 759348
rect 676220 759296 676272 759348
rect 673184 759160 673236 759212
rect 676220 759160 676272 759212
rect 673828 759024 673880 759076
rect 676036 759024 676088 759076
rect 673644 758820 673696 758872
rect 676220 758820 676272 758872
rect 33784 758480 33836 758532
rect 41788 758480 41840 758532
rect 32496 758344 32548 758396
rect 42708 758344 42760 758396
rect 32404 758276 32456 758328
rect 42432 758276 42484 758328
rect 673552 758208 673604 758260
rect 676036 758208 676088 758260
rect 41880 756984 41932 757036
rect 42432 756848 42484 756900
rect 55956 756848 56008 756900
rect 41880 756712 41932 756764
rect 42708 756508 42760 756560
rect 42984 756508 43036 756560
rect 673368 756236 673420 756288
rect 676220 756236 676272 756288
rect 674380 755556 674432 755608
rect 676220 755556 676272 755608
rect 42432 755488 42484 755540
rect 42616 755216 42668 755268
rect 672816 755080 672868 755132
rect 676220 755080 676272 755132
rect 671988 754944 672040 754996
rect 676128 754944 676180 754996
rect 42064 754264 42116 754316
rect 42616 754264 42668 754316
rect 673092 753584 673144 753636
rect 676220 753584 676272 753636
rect 43628 753516 43680 753568
rect 62120 753516 62172 753568
rect 674472 753380 674524 753432
rect 676036 753380 676088 753432
rect 673000 752360 673052 752412
rect 676220 752360 676272 752412
rect 672908 752224 672960 752276
rect 676128 752224 676180 752276
rect 674564 751884 674616 751936
rect 676220 751884 676272 751936
rect 42156 751748 42208 751800
rect 42616 751748 42668 751800
rect 42616 751612 42668 751664
rect 42984 751612 43036 751664
rect 42156 751068 42208 751120
rect 43260 751068 43312 751120
rect 42156 749776 42208 749828
rect 43168 749776 43220 749828
rect 42984 749368 43036 749420
rect 44456 749368 44508 749420
rect 651564 749368 651616 749420
rect 668584 749368 668636 749420
rect 670056 749368 670108 749420
rect 683120 749368 683172 749420
rect 43076 747940 43128 747992
rect 44364 747940 44416 747992
rect 42984 746988 43036 747040
rect 42064 746920 42116 746972
rect 42156 746920 42208 746972
rect 42616 746920 42668 746972
rect 42156 746036 42208 746088
rect 43076 746036 43128 746088
rect 42156 745628 42208 745680
rect 42708 745628 42760 745680
rect 42708 745492 42760 745544
rect 42892 745492 42944 745544
rect 670608 743792 670660 743844
rect 42156 743724 42208 743776
rect 42708 743724 42760 743776
rect 675392 743724 675444 743776
rect 42156 743248 42208 743300
rect 42616 743248 42668 743300
rect 673184 742500 673236 742552
rect 675392 742500 675444 742552
rect 54484 741072 54536 741124
rect 62120 741072 62172 741124
rect 674840 739916 674892 739968
rect 675392 739916 675444 739968
rect 673000 739100 673052 739152
rect 675392 739100 675444 739152
rect 673092 738624 673144 738676
rect 675392 738624 675444 738676
rect 673644 738216 673696 738268
rect 675392 738216 675444 738268
rect 674380 735632 674432 735684
rect 675392 735632 675444 735684
rect 651564 735564 651616 735616
rect 660304 735564 660356 735616
rect 672908 734952 672960 735004
rect 675392 734952 675444 735004
rect 659016 734816 659068 734868
rect 674656 734816 674708 734868
rect 672632 733864 672684 733916
rect 675392 733864 675444 733916
rect 674656 732028 674708 732080
rect 675392 732028 675444 732080
rect 31392 731348 31444 731400
rect 44548 731348 44600 731400
rect 31484 731212 31536 731264
rect 44824 731212 44876 731264
rect 31576 731076 31628 731128
rect 50344 731076 50396 731128
rect 31668 730940 31720 730992
rect 51724 730940 51776 730992
rect 671804 730464 671856 730516
rect 675392 730464 675444 730516
rect 674656 728628 674708 728680
rect 675484 728628 675536 728680
rect 51724 727268 51776 727320
rect 62120 727268 62172 727320
rect 652024 723120 652076 723172
rect 668676 723120 668728 723172
rect 41512 719652 41564 719704
rect 50344 719652 50396 719704
rect 35808 716864 35860 716916
rect 42432 716864 42484 716916
rect 672724 716524 672776 716576
rect 676036 716524 676088 716576
rect 40776 716184 40828 716236
rect 41880 716184 41932 716236
rect 671344 716116 671396 716168
rect 676036 716116 676088 716168
rect 35716 715504 35768 715556
rect 42524 715504 42576 715556
rect 663064 714960 663116 715012
rect 676036 714960 676088 715012
rect 50436 714824 50488 714876
rect 62120 714824 62172 714876
rect 673828 714484 673880 714536
rect 676036 714484 676088 714536
rect 40684 714212 40736 714264
rect 42800 714212 42852 714264
rect 40868 714144 40920 714196
rect 42892 714144 42944 714196
rect 673828 714008 673880 714060
rect 676036 714008 676088 714060
rect 41880 713804 41932 713856
rect 673552 713668 673604 713720
rect 676036 713668 676088 713720
rect 41880 713532 41932 713584
rect 674564 713192 674616 713244
rect 676036 713192 676088 713244
rect 673368 712852 673420 712904
rect 676036 712852 676088 712904
rect 672172 712376 672224 712428
rect 676036 712376 676088 712428
rect 43076 712104 43128 712156
rect 47584 712104 47636 712156
rect 42156 711628 42208 711680
rect 42800 711628 42852 711680
rect 670516 711628 670568 711680
rect 676036 711628 676088 711680
rect 42524 710948 42576 711000
rect 42800 710948 42852 711000
rect 42156 710880 42208 710932
rect 43076 710880 43128 710932
rect 671896 710404 671948 710456
rect 676036 710404 676088 710456
rect 672448 709996 672500 710048
rect 676036 709996 676088 710048
rect 42156 709860 42208 709912
rect 42892 709860 42944 709912
rect 674288 709588 674340 709640
rect 676036 709588 676088 709640
rect 42892 709316 42944 709368
rect 44180 709316 44232 709368
rect 651564 709316 651616 709368
rect 671436 709316 671488 709368
rect 674196 709180 674248 709232
rect 676036 709180 676088 709232
rect 676036 709044 676088 709096
rect 676956 709044 677008 709096
rect 42156 708568 42208 708620
rect 42524 708568 42576 708620
rect 673920 708364 673972 708416
rect 676036 708364 676088 708416
rect 42156 708024 42208 708076
rect 42984 708024 43036 708076
rect 672540 707956 672592 708008
rect 676036 707956 676088 708008
rect 674012 707548 674064 707600
rect 676036 707548 676088 707600
rect 42156 707208 42208 707260
rect 42892 707208 42944 707260
rect 673736 706732 673788 706784
rect 675944 706732 675996 706784
rect 673276 706664 673328 706716
rect 676036 706664 676088 706716
rect 42432 706052 42484 706104
rect 44456 706596 44508 706648
rect 42064 704216 42116 704268
rect 42432 704216 42484 704268
rect 672724 703808 672776 703860
rect 676036 703808 676088 703860
rect 42156 703672 42208 703724
rect 42800 703672 42852 703724
rect 42800 701020 42852 701072
rect 44364 701020 44416 701072
rect 42156 700408 42208 700460
rect 42432 700408 42484 700460
rect 42156 699864 42208 699916
rect 42708 699864 42760 699916
rect 671988 698164 672040 698216
rect 675392 698164 675444 698216
rect 672264 697348 672316 697400
rect 675392 697348 675444 697400
rect 30288 696192 30340 696244
rect 43628 696192 43680 696244
rect 674472 694288 674524 694340
rect 675484 694288 675536 694340
rect 673552 692996 673604 693048
rect 675484 692996 675536 693048
rect 673368 690412 673420 690464
rect 675392 690412 675444 690464
rect 674012 690004 674064 690056
rect 675392 690004 675444 690056
rect 672816 689324 672868 689376
rect 675484 689324 675536 689376
rect 674196 688712 674248 688764
rect 675392 688712 675444 688764
rect 43720 688644 43772 688696
rect 62120 688644 62172 688696
rect 668676 688644 668728 688696
rect 674288 688644 674340 688696
rect 35808 687896 35860 687948
rect 51724 687896 51776 687948
rect 35624 687760 35676 687812
rect 54484 687760 54536 687812
rect 674288 687012 674340 687064
rect 675484 687012 675536 687064
rect 673920 684224 673972 684276
rect 675392 684224 675444 684276
rect 651840 683136 651892 683188
rect 659016 683136 659068 683188
rect 40684 683000 40736 683052
rect 41696 683000 41748 683052
rect 40776 681776 40828 681828
rect 41696 681776 41748 681828
rect 30472 676812 30524 676864
rect 51724 676812 51776 676864
rect 55956 674840 56008 674892
rect 62120 674840 62172 674892
rect 35164 672800 35216 672852
rect 42432 672800 42484 672852
rect 31024 672732 31076 672784
rect 41880 672732 41932 672784
rect 40776 670964 40828 671016
rect 42064 670964 42116 671016
rect 40684 670896 40736 670948
rect 41788 670896 41840 670948
rect 665824 670896 665876 670948
rect 676036 670896 676088 670948
rect 658924 670760 658976 670812
rect 676220 670760 676272 670812
rect 41880 670556 41932 670608
rect 41972 670556 42024 670608
rect 42892 670556 42944 670608
rect 41880 670352 41932 670404
rect 42708 670012 42760 670064
rect 48964 670012 49016 670064
rect 673828 669468 673880 669520
rect 676036 669468 676088 669520
rect 661776 669400 661828 669452
rect 676128 669400 676180 669452
rect 651564 669332 651616 669384
rect 658924 669332 658976 669384
rect 672448 669332 672500 669384
rect 676220 669332 676272 669384
rect 674564 668516 674616 668568
rect 676036 668516 676088 668568
rect 672540 667904 672592 667956
rect 676220 667904 676272 667956
rect 42156 667836 42208 667888
rect 42708 667836 42760 667888
rect 42800 667768 42852 667820
rect 42800 667564 42852 667616
rect 673828 667224 673880 667276
rect 676036 667224 676088 667276
rect 42156 666680 42208 666732
rect 44180 666680 44232 666732
rect 672172 666680 672224 666732
rect 676220 666680 676272 666732
rect 671804 665456 671856 665508
rect 676128 665456 676180 665508
rect 670608 665320 670660 665372
rect 676220 665320 676272 665372
rect 674380 665252 674432 665304
rect 676036 665252 676088 665304
rect 42892 665184 42944 665236
rect 44456 665184 44508 665236
rect 674656 664980 674708 665032
rect 676220 664980 676272 665032
rect 42156 663960 42208 664012
rect 42892 663960 42944 664012
rect 673184 663960 673236 664012
rect 676220 663960 676272 664012
rect 42708 663756 42760 663808
rect 42892 663756 42944 663808
rect 673000 663756 673052 663808
rect 676220 663756 676272 663808
rect 42800 662600 42852 662652
rect 43076 662600 43128 662652
rect 42708 662396 42760 662448
rect 42984 662396 43036 662448
rect 47584 662396 47636 662448
rect 62120 662396 62172 662448
rect 673092 662396 673144 662448
rect 676220 662396 676272 662448
rect 673644 662328 673696 662380
rect 676036 662328 676088 662380
rect 672908 661240 672960 661292
rect 676220 661240 676272 661292
rect 672632 661104 672684 661156
rect 676128 661104 676180 661156
rect 42156 661036 42208 661088
rect 42800 661036 42852 661088
rect 42156 659676 42208 659728
rect 42892 659676 42944 659728
rect 674196 659676 674248 659728
rect 683120 659676 683172 659728
rect 42156 658996 42208 659048
rect 42708 658996 42760 659048
rect 42156 657228 42208 657280
rect 42524 657228 42576 657280
rect 651564 656888 651616 656940
rect 663064 656888 663116 656940
rect 42156 656820 42208 656872
rect 43076 656820 43128 656872
rect 42156 656140 42208 656192
rect 42340 656140 42392 656192
rect 675208 653760 675260 653812
rect 675484 653760 675536 653812
rect 671896 652740 671948 652792
rect 675392 652740 675444 652792
rect 674656 652128 674708 652180
rect 675484 652128 675536 652180
rect 671804 651516 671856 651568
rect 675392 651516 675444 651568
rect 674380 649068 674432 649120
rect 675392 649068 675444 649120
rect 43628 647844 43680 647896
rect 62120 647844 62172 647896
rect 673184 647708 673236 647760
rect 675484 647708 675536 647760
rect 673736 645396 673788 645448
rect 675392 645396 675444 645448
rect 673000 644988 673052 645040
rect 675392 644988 675444 645040
rect 35624 644580 35676 644632
rect 43720 644580 43772 644632
rect 35808 644512 35860 644564
rect 55956 644512 56008 644564
rect 658924 643696 658976 643748
rect 674564 643696 674616 643748
rect 673092 643356 673144 643408
rect 675392 643356 675444 643408
rect 651564 643084 651616 643136
rect 668676 643084 668728 643136
rect 674564 641860 674616 641912
rect 675392 641860 675444 641912
rect 670516 640296 670568 640348
rect 675392 640296 675444 640348
rect 673276 639072 673328 639124
rect 675392 639072 675444 639124
rect 55956 636216 56008 636268
rect 62120 636216 62172 636268
rect 675484 633768 675536 633820
rect 681096 633768 681148 633820
rect 32404 629892 32456 629944
rect 41788 629892 41840 629944
rect 651564 629280 651616 629332
rect 661684 629280 661736 629332
rect 39304 629212 39356 629264
rect 42524 629212 42576 629264
rect 41788 627376 41840 627428
rect 42892 627172 42944 627224
rect 50436 627172 50488 627224
rect 41788 627036 41840 627088
rect 668584 625472 668636 625524
rect 676128 625472 676180 625524
rect 664536 625336 664588 625388
rect 676220 625336 676272 625388
rect 42156 625268 42208 625320
rect 42524 625268 42576 625320
rect 660304 625132 660356 625184
rect 676220 625132 676272 625184
rect 42156 624656 42208 624708
rect 42892 624656 42944 624708
rect 672448 624112 672500 624164
rect 676220 624112 676272 624164
rect 672540 623908 672592 623960
rect 676220 623908 676272 623960
rect 42524 623840 42576 623892
rect 672448 623840 672500 623892
rect 676128 623840 676180 623892
rect 42156 623432 42208 623484
rect 51816 623772 51868 623824
rect 62120 623772 62172 623824
rect 672540 623772 672592 623824
rect 676036 623772 676088 623824
rect 674748 623636 674800 623688
rect 676220 623636 676272 623688
rect 673460 623024 673512 623076
rect 676036 623024 676088 623076
rect 673828 622820 673880 622872
rect 676220 622820 676272 622872
rect 42064 622140 42116 622192
rect 42524 622140 42576 622192
rect 42524 622004 42576 622056
rect 44548 622412 44600 622464
rect 673828 622208 673880 622260
rect 676036 622208 676088 622260
rect 671988 621120 672040 621172
rect 676220 621120 676272 621172
rect 42524 621052 42576 621104
rect 42524 620916 42576 620968
rect 42800 620916 42852 620968
rect 42064 620780 42116 620832
rect 42064 620304 42116 620356
rect 42984 620304 43036 620356
rect 673920 619828 673972 619880
rect 676036 619828 676088 619880
rect 673368 619760 673420 619812
rect 676220 619760 676272 619812
rect 674472 619012 674524 619064
rect 676036 619012 676088 619064
rect 672264 618400 672316 618452
rect 676220 618400 676272 618452
rect 42156 617856 42208 617908
rect 42524 617856 42576 617908
rect 42524 617720 42576 617772
rect 44456 618264 44508 618316
rect 673552 617380 673604 617432
rect 676036 617380 676088 617432
rect 42064 617108 42116 617160
rect 42524 617108 42576 617160
rect 674012 616972 674064 617024
rect 676036 616972 676088 617024
rect 652392 616836 652444 616888
rect 658924 616836 658976 616888
rect 672816 616836 672868 616888
rect 676220 616836 676272 616888
rect 674288 616700 674340 616752
rect 676220 616700 676272 616752
rect 42156 614184 42208 614236
rect 42524 614184 42576 614236
rect 671344 614116 671396 614168
rect 683120 614116 683172 614168
rect 42156 612756 42208 612808
rect 42524 612756 42576 612808
rect 48964 609968 49016 610020
rect 62120 609968 62172 610020
rect 670608 607996 670660 608048
rect 675392 607996 675444 608048
rect 673368 607588 673420 607640
rect 675392 607588 675444 607640
rect 675208 604528 675260 604580
rect 675392 604528 675444 604580
rect 674472 604324 674524 604376
rect 675392 604324 675444 604376
rect 674564 603236 674616 603288
rect 675484 603236 675536 603288
rect 651564 603100 651616 603152
rect 660304 603100 660356 603152
rect 673552 603032 673604 603084
rect 675392 603032 675444 603084
rect 35808 601672 35860 601724
rect 55956 601672 56008 601724
rect 35716 601604 35768 601656
rect 43628 601604 43680 601656
rect 35624 601468 35676 601520
rect 44180 601468 44232 601520
rect 35808 601332 35860 601384
rect 51816 601332 51868 601384
rect 672816 600380 672868 600432
rect 675484 600380 675536 600432
rect 674288 599768 674340 599820
rect 675484 599768 675536 599820
rect 658924 599564 658976 599616
rect 674748 599564 674800 599616
rect 674012 598408 674064 598460
rect 675484 598408 675536 598460
rect 672908 597728 672960 597780
rect 675484 597728 675536 597780
rect 50436 597524 50488 597576
rect 62120 597524 62172 597576
rect 674748 596844 674800 596896
rect 675392 596844 675444 596896
rect 672632 593376 672684 593428
rect 675484 593376 675536 593428
rect 651564 590656 651616 590708
rect 664444 590656 664496 590708
rect 41512 589908 41564 589960
rect 53104 589908 53156 589960
rect 33784 585896 33836 585948
rect 41880 585896 41932 585948
rect 32404 585760 32456 585812
rect 41604 585760 41656 585812
rect 41880 584196 41932 584248
rect 42064 584196 42116 584248
rect 42708 584196 42760 584248
rect 41880 583924 41932 583976
rect 51816 583720 51868 583772
rect 62120 583720 62172 583772
rect 42156 581272 42208 581324
rect 47584 581272 47636 581324
rect 652024 581000 652076 581052
rect 676036 581000 676088 581052
rect 672448 580048 672500 580100
rect 676220 580048 676272 580100
rect 671436 579912 671488 579964
rect 676128 579912 676180 579964
rect 659016 579776 659068 579828
rect 676036 579776 676088 579828
rect 42984 579640 43036 579692
rect 44640 579640 44692 579692
rect 42156 578416 42208 578468
rect 42984 578416 43036 578468
rect 672540 578416 672592 578468
rect 676220 578416 676272 578468
rect 672448 578280 672500 578332
rect 676312 578280 676364 578332
rect 42984 578212 43036 578264
rect 44364 578212 44416 578264
rect 672540 578212 672592 578264
rect 676128 578212 676180 578264
rect 673460 578144 673512 578196
rect 676036 578144 676088 578196
rect 673920 577600 673972 577652
rect 676220 577600 676272 577652
rect 673828 577396 673880 577448
rect 676036 577396 676088 577448
rect 42156 576920 42208 576972
rect 42984 576920 43036 576972
rect 673644 576920 673696 576972
rect 676036 576920 676088 576972
rect 44456 576852 44508 576904
rect 651564 576852 651616 576904
rect 659016 576852 659068 576904
rect 42156 576580 42208 576632
rect 42708 576376 42760 576428
rect 42432 576308 42484 576360
rect 42156 576172 42208 576224
rect 42340 575968 42392 576020
rect 671896 575832 671948 575884
rect 676036 575832 676088 575884
rect 671804 575696 671856 575748
rect 676128 575696 676180 575748
rect 670516 575560 670568 575612
rect 676220 575560 676272 575612
rect 673736 574948 673788 575000
rect 676036 574948 676088 575000
rect 42156 574676 42208 574728
rect 42340 574676 42392 574728
rect 673276 574200 673328 574252
rect 676220 574200 676272 574252
rect 42340 574132 42392 574184
rect 42708 574132 42760 574184
rect 674656 574132 674708 574184
rect 676036 574132 676088 574184
rect 674380 573724 674432 573776
rect 676036 573724 676088 573776
rect 42156 573452 42208 573504
rect 42892 573452 42944 573504
rect 41972 572704 42024 572756
rect 42708 572704 42760 572756
rect 673184 571616 673236 571668
rect 676220 571616 676272 571668
rect 42340 571480 42392 571532
rect 673000 571480 673052 571532
rect 676220 571480 676272 571532
rect 42064 570868 42116 570920
rect 43720 571344 43772 571396
rect 62120 571344 62172 571396
rect 673092 569916 673144 569968
rect 676220 569916 676272 569968
rect 42064 569576 42116 569628
rect 42708 569576 42760 569628
rect 671436 568556 671488 568608
rect 683120 568556 683172 568608
rect 35624 566448 35676 566500
rect 43720 566448 43772 566500
rect 652116 563048 652168 563100
rect 658924 563048 658976 563100
rect 671988 561892 672040 561944
rect 675392 561892 675444 561944
rect 673276 559104 673328 559156
rect 675392 559104 675444 559156
rect 35716 558288 35768 558340
rect 50436 558288 50488 558340
rect 35808 558152 35860 558204
rect 51816 558152 51868 558204
rect 47584 557540 47636 557592
rect 62120 557540 62172 557592
rect 673184 557540 673236 557592
rect 675484 557540 675536 557592
rect 674748 555228 674800 555280
rect 675392 555228 675444 555280
rect 673092 554752 673144 554804
rect 675300 554752 675352 554804
rect 658924 554004 658976 554056
rect 675300 554004 675352 554056
rect 674380 553392 674432 553444
rect 675392 553392 675444 553444
rect 651564 550604 651616 550656
rect 661776 550604 661828 550656
rect 674656 549312 674708 549364
rect 674932 549312 674984 549364
rect 674932 549176 674984 549228
rect 675300 549176 675352 549228
rect 674748 548428 674800 548480
rect 674748 548292 674800 548344
rect 675300 548292 675352 548344
rect 674656 547952 674708 548004
rect 675760 547952 675812 548004
rect 674380 547884 674432 547936
rect 31668 547136 31720 547188
rect 35808 547136 35860 547188
rect 53196 547136 53248 547188
rect 43628 545096 43680 545148
rect 62120 545096 62172 545148
rect 31024 542988 31076 543040
rect 41788 542988 41840 543040
rect 40684 542308 40736 542360
rect 42708 542308 42760 542360
rect 41788 541016 41840 541068
rect 41788 540744 41840 540796
rect 42984 540200 43036 540252
rect 48964 540200 49016 540252
rect 42064 538908 42116 538960
rect 42708 538908 42760 538960
rect 42984 538364 43036 538416
rect 42156 538228 42208 538280
rect 42984 538228 43036 538280
rect 44180 538228 44232 538280
rect 42064 537072 42116 537124
rect 42984 537072 43036 537124
rect 42616 536800 42668 536852
rect 44548 536800 44600 536852
rect 651564 536800 651616 536852
rect 660396 536800 660448 536852
rect 42616 535984 42668 536036
rect 42156 535780 42208 535832
rect 668676 535712 668728 535764
rect 676220 535712 676272 535764
rect 663064 535576 663116 535628
rect 676036 535576 676088 535628
rect 42064 535236 42116 535288
rect 43076 535236 43128 535288
rect 672448 534488 672500 534540
rect 676220 534488 676272 534540
rect 672540 534352 672592 534404
rect 676220 534352 676272 534404
rect 661684 534216 661736 534268
rect 676128 534216 676180 534268
rect 42156 533944 42208 533996
rect 42616 533944 42668 533996
rect 673920 533264 673972 533316
rect 676036 533264 676088 533316
rect 55956 532720 56008 532772
rect 62120 532720 62172 532772
rect 673644 532652 673696 532704
rect 676220 532652 676272 532704
rect 42156 530884 42208 530936
rect 42616 530884 42668 530936
rect 42616 530748 42668 530800
rect 44456 531292 44508 531344
rect 672816 530136 672868 530188
rect 676220 530136 676272 530188
rect 42156 530068 42208 530120
rect 42616 530068 42668 530120
rect 670608 530000 670660 530052
rect 676128 530000 676180 530052
rect 42156 529456 42208 529508
rect 42340 529592 42392 529644
rect 674472 528980 674524 529032
rect 676404 528980 676456 529032
rect 673368 528776 673420 528828
rect 676220 528776 676272 528828
rect 672632 528640 672684 528692
rect 676128 528640 676180 528692
rect 674564 528368 674616 528420
rect 675852 528368 675904 528420
rect 672908 527416 672960 527468
rect 676220 527416 676272 527468
rect 42064 527212 42116 527264
rect 42340 527212 42392 527264
rect 42156 527144 42208 527196
rect 42892 527144 42944 527196
rect 673552 527076 673604 527128
rect 675852 527076 675904 527128
rect 674288 526940 674340 526992
rect 676220 526940 676272 526992
rect 42156 526600 42208 526652
rect 42616 526600 42668 526652
rect 674012 526532 674064 526584
rect 676220 526532 676272 526584
rect 674472 524424 674524 524476
rect 683120 524424 683172 524476
rect 651564 522996 651616 523048
rect 663248 522996 663300 523048
rect 677324 520276 677376 520328
rect 683856 520276 683908 520328
rect 40684 518916 40736 518968
rect 62120 518916 62172 518968
rect 651564 510620 651616 510672
rect 661684 510620 661736 510672
rect 48964 506472 49016 506524
rect 62120 506472 62172 506524
rect 675024 500896 675076 500948
rect 681004 500896 681056 500948
rect 674932 498244 674984 498296
rect 679716 498244 679768 498296
rect 675760 498176 675812 498228
rect 679624 498176 679676 498228
rect 651564 496816 651616 496868
rect 658924 496816 658976 496868
rect 46204 491920 46256 491972
rect 62120 491920 62172 491972
rect 664444 491648 664496 491700
rect 675852 491648 675904 491700
rect 660304 491512 660356 491564
rect 675944 491512 675996 491564
rect 659016 491376 659068 491428
rect 675944 491376 675996 491428
rect 675944 490152 675996 490204
rect 676128 490152 676180 490204
rect 676036 488792 676088 488844
rect 677324 488792 677376 488844
rect 676036 488452 676088 488504
rect 677232 488452 677284 488504
rect 676036 487976 676088 488028
rect 677232 487976 677284 488028
rect 676036 486820 676088 486872
rect 677508 486820 677560 486872
rect 674380 486004 674432 486056
rect 676036 486004 676088 486056
rect 671988 485188 672040 485240
rect 675944 485188 675996 485240
rect 673276 484780 673328 484832
rect 675944 484780 675996 484832
rect 651564 484372 651616 484424
rect 660488 484372 660540 484424
rect 673184 483148 673236 483200
rect 675944 483148 675996 483200
rect 673092 482740 673144 482792
rect 675944 482740 675996 482792
rect 44824 480224 44876 480276
rect 62120 480224 62172 480276
rect 674288 480224 674340 480276
rect 678980 480224 679032 480276
rect 668584 475804 668636 475856
rect 674472 475804 674524 475856
rect 668676 474512 668728 474564
rect 671436 474512 671488 474564
rect 651656 470568 651708 470620
rect 664536 470568 664588 470620
rect 51816 466420 51868 466472
rect 62120 466420 62172 466472
rect 651564 456764 651616 456816
rect 663156 456764 663208 456816
rect 50436 454044 50488 454096
rect 62120 454044 62172 454096
rect 651564 444388 651616 444440
rect 659016 444388 659068 444440
rect 43720 440240 43772 440292
rect 62120 440240 62172 440292
rect 40684 432556 40736 432608
rect 41788 432556 41840 432608
rect 43168 430584 43220 430636
rect 55956 430584 56008 430636
rect 651564 430584 651616 430636
rect 660304 430584 660356 430636
rect 46296 427796 46348 427848
rect 62120 427796 62172 427848
rect 41788 419432 41840 419484
rect 43628 419432 43680 419484
rect 651564 416780 651616 416832
rect 663064 416780 663116 416832
rect 55956 415420 56008 415472
rect 62120 415420 62172 415472
rect 32496 414808 32548 414860
rect 41880 414808 41932 414860
rect 31024 414672 31076 414724
rect 42524 414672 42576 414724
rect 41880 413380 41932 413432
rect 41880 413108 41932 413160
rect 42156 410660 42208 410712
rect 47584 410660 47636 410712
rect 42064 408144 42116 408196
rect 44640 408144 44692 408196
rect 42156 407600 42208 407652
rect 42524 407600 42576 407652
rect 42064 406784 42116 406836
rect 42984 406784 43036 406836
rect 652024 404336 652076 404388
rect 661868 404336 661920 404388
rect 42156 403860 42208 403912
rect 44456 403860 44508 403912
rect 663248 403384 663300 403436
rect 676404 403384 676456 403436
rect 661776 403248 661828 403300
rect 676220 403248 676272 403300
rect 660396 403112 660448 403164
rect 676312 403112 676364 403164
rect 42156 402908 42208 402960
rect 42892 402908 42944 402960
rect 47584 401616 47636 401668
rect 62120 401616 62172 401668
rect 673276 401616 673328 401668
rect 676220 401616 676272 401668
rect 673368 400188 673420 400240
rect 676220 400188 676272 400240
rect 674656 399576 674708 399628
rect 676220 399576 676272 399628
rect 675024 398216 675076 398268
rect 676036 398216 676088 398268
rect 674932 397468 674984 397520
rect 676036 397468 676088 397520
rect 674564 394272 674616 394324
rect 676220 394272 676272 394324
rect 673184 393320 673236 393372
rect 676220 393320 676272 393372
rect 670148 391960 670200 392012
rect 683120 391960 683172 392012
rect 651564 390532 651616 390584
rect 664444 390532 664496 390584
rect 45008 389172 45060 389224
rect 62120 389172 62172 389224
rect 675208 389104 675260 389156
rect 676956 389104 677008 389156
rect 35716 387744 35768 387796
rect 44180 387744 44232 387796
rect 35808 387608 35860 387660
rect 44824 387608 44876 387660
rect 675116 387540 675168 387592
rect 676496 387540 676548 387592
rect 35624 387472 35676 387524
rect 46204 387472 46256 387524
rect 35808 387336 35860 387388
rect 51816 387336 51868 387388
rect 675300 387064 675352 387116
rect 678244 387064 678296 387116
rect 675024 386112 675076 386164
rect 675392 386112 675444 386164
rect 675024 385976 675076 386028
rect 675300 385976 675352 386028
rect 675024 383868 675076 383920
rect 675300 383868 675352 383920
rect 674932 383052 674984 383104
rect 675392 383052 675444 383104
rect 675116 381080 675168 381132
rect 675392 381080 675444 381132
rect 651564 378156 651616 378208
rect 665824 378156 665876 378208
rect 674564 377952 674616 378004
rect 675484 377952 675536 378004
rect 673184 376592 673236 376644
rect 675484 376592 675536 376644
rect 35808 376048 35860 376100
rect 41512 376048 41564 376100
rect 44824 376048 44876 376100
rect 49056 375368 49108 375420
rect 62120 375368 62172 375420
rect 31024 371832 31076 371884
rect 42340 371832 42392 371884
rect 40868 371220 40920 371272
rect 42708 371220 42760 371272
rect 40684 370540 40736 370592
rect 41788 370540 41840 370592
rect 42156 369656 42208 369708
rect 42340 369656 42392 369708
rect 42156 368092 42208 368144
rect 42708 368092 42760 368144
rect 42156 366800 42208 366852
rect 42708 366800 42760 366852
rect 42156 364964 42208 365016
rect 44548 364964 44600 365016
rect 652024 364352 652076 364404
rect 660396 364352 660448 364404
rect 42156 364284 42208 364336
rect 44456 364284 44508 364336
rect 42708 364216 42760 364268
rect 48964 364216 49016 364268
rect 56048 362924 56100 362976
rect 62120 362924 62172 362976
rect 42064 360680 42116 360732
rect 43076 360680 43128 360732
rect 42156 359456 42208 359508
rect 42984 359456 43036 359508
rect 661684 357824 661736 357876
rect 675944 357824 675996 357876
rect 660488 357688 660540 357740
rect 676036 357688 676088 357740
rect 658924 357552 658976 357604
rect 675852 357552 675904 357604
rect 673276 357484 673328 357536
rect 676036 357484 676088 357536
rect 673276 357008 673328 357060
rect 676036 357008 676088 357060
rect 673368 356668 673420 356720
rect 676036 356668 676088 356720
rect 673000 356192 673052 356244
rect 676036 356192 676088 356244
rect 42156 355988 42208 356040
rect 43168 355988 43220 356040
rect 674656 355036 674708 355088
rect 676036 355036 676088 355088
rect 674656 354560 674708 354612
rect 676036 354560 676088 354612
rect 27620 351160 27672 351212
rect 46296 351160 46348 351212
rect 676220 351092 676272 351144
rect 676864 351092 676916 351144
rect 674472 350888 674524 350940
rect 676036 350888 676088 350940
rect 651564 350548 651616 350600
rect 671528 350548 671580 350600
rect 673184 350548 673236 350600
rect 676036 350548 676088 350600
rect 674564 349256 674616 349308
rect 676036 349256 676088 349308
rect 673092 348848 673144 348900
rect 676036 348848 676088 348900
rect 44916 347012 44968 347064
rect 62120 347012 62172 347064
rect 671436 346400 671488 346452
rect 676036 346400 676088 346452
rect 35716 344292 35768 344344
rect 43720 344292 43772 344344
rect 35808 344156 35860 344208
rect 55956 344156 56008 344208
rect 651656 338104 651708 338156
rect 668768 338104 668820 338156
rect 46296 336744 46348 336796
rect 62120 336744 62172 336796
rect 674472 336540 674524 336592
rect 675484 336540 675536 336592
rect 674840 336268 674892 336320
rect 675392 336268 675444 336320
rect 30380 333208 30432 333260
rect 64144 333208 64196 333260
rect 674564 332596 674616 332648
rect 675392 332596 675444 332648
rect 673092 331576 673144 331628
rect 675392 331576 675444 331628
rect 674840 329468 674892 329520
rect 675392 329468 675444 329520
rect 673184 328380 673236 328432
rect 674840 328380 674892 328432
rect 675116 327632 675168 327684
rect 675484 327632 675536 327684
rect 42064 326748 42116 326800
rect 44180 326748 44232 326800
rect 675760 325796 675812 325848
rect 675760 325592 675812 325644
rect 651564 324300 651616 324352
rect 670240 324300 670292 324352
rect 42156 323280 42208 323332
rect 42616 323280 42668 323332
rect 47676 322940 47728 322992
rect 62120 322940 62172 322992
rect 42064 322872 42116 322924
rect 44364 322872 44416 322924
rect 42616 321512 42668 321564
rect 50436 321512 50488 321564
rect 42156 321444 42208 321496
rect 44456 321444 44508 321496
rect 42156 319948 42208 320000
rect 43076 319948 43128 320000
rect 42156 316684 42208 316736
rect 42984 316684 43036 316736
rect 664536 313488 664588 313540
rect 676220 313488 676272 313540
rect 663156 313352 663208 313404
rect 676036 313352 676088 313404
rect 673276 312128 673328 312180
rect 676220 312128 676272 312180
rect 659016 311992 659068 312044
rect 676128 311992 676180 312044
rect 673368 311856 673420 311908
rect 676220 311856 676272 311908
rect 673000 310632 673052 310684
rect 676220 310632 676272 310684
rect 651564 310564 651616 310616
rect 674104 310564 674156 310616
rect 46204 310496 46256 310548
rect 62120 310496 62172 310548
rect 673276 310496 673328 310548
rect 676128 310496 676180 310548
rect 674748 310224 674800 310276
rect 676220 310224 676272 310276
rect 674656 310020 674708 310072
rect 676036 310020 676088 310072
rect 674748 309408 674800 309460
rect 676220 309408 676272 309460
rect 673184 303764 673236 303816
rect 676220 303764 676272 303816
rect 673092 303696 673144 303748
rect 676128 303696 676180 303748
rect 673000 303628 673052 303680
rect 676312 303628 676364 303680
rect 674380 302200 674432 302252
rect 683120 302200 683172 302252
rect 35808 301044 35860 301096
rect 49056 300976 49108 301028
rect 35808 300908 35860 300960
rect 56048 300908 56100 300960
rect 43720 298120 43772 298172
rect 62120 298120 62172 298172
rect 675208 298052 675260 298104
rect 676864 298052 676916 298104
rect 675760 297984 675812 298036
rect 678244 297984 678296 298036
rect 675116 297372 675168 297424
rect 676496 297372 676548 297424
rect 675760 296148 675812 296200
rect 675760 295944 675812 295996
rect 675208 295400 675260 295452
rect 675392 295400 675444 295452
rect 675116 294040 675168 294092
rect 675024 293972 675076 294024
rect 675024 291728 675076 291780
rect 675392 291728 675444 291780
rect 673000 291048 673052 291100
rect 675392 291048 675444 291100
rect 673092 287920 673144 287972
rect 675392 287920 675444 287972
rect 673184 286560 673236 286612
rect 675392 286560 675444 286612
rect 32404 284928 32456 284980
rect 41880 284928 41932 284980
rect 43812 284316 43864 284368
rect 62120 284316 62172 284368
rect 651564 284316 651616 284368
rect 672816 284316 672868 284368
rect 41880 283772 41932 283824
rect 41880 283568 41932 283620
rect 42156 280168 42208 280220
rect 47584 280168 47636 280220
rect 42064 278604 42116 278656
rect 44548 278604 44600 278656
rect 43444 278196 43496 278248
rect 646044 278196 646096 278248
rect 53196 278128 53248 278180
rect 656900 278128 656952 278180
rect 51816 278060 51868 278112
rect 662420 278060 662472 278112
rect 43628 277992 43680 278044
rect 658280 277992 658332 278044
rect 332508 277924 332560 277976
rect 436652 277924 436704 277976
rect 333888 277856 333940 277908
rect 440332 277856 440384 277908
rect 335084 277788 335136 277840
rect 443828 277788 443880 277840
rect 336372 277720 336424 277772
rect 447324 277720 447376 277772
rect 338028 277652 338080 277704
rect 452476 277652 452528 277704
rect 339224 277584 339276 277636
rect 454776 277584 454828 277636
rect 360108 277516 360160 277568
rect 507952 277516 508004 277568
rect 391664 277448 391716 277500
rect 594340 277448 594392 277500
rect 398748 277380 398800 277432
rect 612004 277380 612056 277432
rect 353208 277312 353260 277364
rect 492588 277312 492640 277364
rect 355968 277244 356020 277296
rect 499764 277244 499816 277296
rect 358728 277176 358780 277228
rect 506848 277176 506900 277228
rect 42156 277108 42208 277160
rect 43168 277108 43220 277160
rect 380808 277108 380860 277160
rect 563520 277108 563572 277160
rect 383476 277040 383528 277092
rect 570696 277040 570748 277092
rect 383568 276972 383620 277024
rect 571800 276972 571852 277024
rect 387248 276904 387300 276956
rect 582472 276904 582524 276956
rect 389916 276836 389968 276888
rect 589556 276836 589608 276888
rect 403900 276768 403952 276820
rect 627368 276768 627420 276820
rect 42064 276700 42116 276752
rect 42892 276700 42944 276752
rect 406660 276700 406712 276752
rect 634452 276700 634504 276752
rect 409788 276632 409840 276684
rect 641628 276632 641680 276684
rect 350448 276564 350500 276616
rect 485504 276564 485556 276616
rect 349068 276496 349120 276548
rect 478420 276496 478472 276548
rect 332416 276428 332468 276480
rect 435916 276428 435968 276480
rect 329748 276360 329800 276412
rect 428832 276360 428884 276412
rect 326712 276292 326764 276344
rect 421656 276292 421708 276344
rect 324044 276224 324096 276276
rect 414572 276224 414624 276276
rect 146208 275952 146260 276004
rect 195980 275952 196032 276004
rect 348976 275952 349028 276004
rect 480812 275952 480864 276004
rect 487160 275952 487212 276004
rect 163964 275884 164016 275936
rect 216680 275884 216732 275936
rect 351828 275884 351880 275936
rect 487896 275884 487948 275936
rect 583760 275952 583812 276004
rect 600228 275952 600280 276004
rect 581276 275884 581328 275936
rect 171048 275816 171100 275868
rect 226984 275816 227036 275868
rect 354404 275816 354456 275868
rect 494980 275816 495032 275868
rect 496728 275816 496780 275868
rect 513932 275816 513984 275868
rect 581644 275816 581696 275868
rect 599032 275816 599084 275868
rect 149796 275748 149848 275800
rect 220636 275748 220688 275800
rect 258540 275748 258592 275800
rect 264612 275748 264664 275800
rect 357348 275748 357400 275800
rect 502064 275748 502116 275800
rect 502248 275748 502300 275800
rect 584864 275748 584916 275800
rect 107200 275680 107252 275732
rect 208308 275680 208360 275732
rect 214840 275680 214892 275732
rect 227720 275680 227772 275732
rect 251456 275680 251508 275732
rect 252376 275680 252428 275732
rect 362224 275680 362276 275732
rect 509148 275680 509200 275732
rect 513472 275680 513524 275732
rect 593144 275680 593196 275732
rect 100116 275612 100168 275664
rect 205824 275612 205876 275664
rect 207756 275612 207808 275664
rect 213460 275612 213512 275664
rect 223120 275612 223172 275664
rect 241428 275612 241480 275664
rect 363512 275612 363564 275664
rect 516232 275612 516284 275664
rect 521568 275612 521620 275664
rect 596640 275612 596692 275664
rect 597836 275612 597888 275664
rect 610808 275612 610860 275664
rect 90640 275544 90692 275596
rect 201684 275544 201736 275596
rect 212448 275544 212500 275596
rect 222476 275544 222528 275596
rect 224224 275544 224276 275596
rect 243544 275544 243596 275596
rect 367008 275544 367060 275596
rect 523408 275544 523460 275596
rect 523684 275544 523736 275596
rect 591948 275544 592000 275596
rect 593420 275544 593472 275596
rect 607312 275544 607364 275596
rect 83556 275476 83608 275528
rect 199108 275476 199160 275528
rect 210056 275476 210108 275528
rect 224960 275476 225012 275528
rect 227812 275476 227864 275528
rect 249616 275476 249668 275528
rect 368388 275476 368440 275528
rect 530492 275476 530544 275528
rect 543740 275476 543792 275528
rect 595444 275476 595496 275528
rect 600044 275476 600096 275528
rect 614396 275476 614448 275528
rect 81256 275408 81308 275460
rect 197820 275408 197872 275460
rect 213644 275408 213696 275460
rect 234620 275408 234672 275460
rect 239588 275408 239640 275460
rect 249708 275408 249760 275460
rect 340604 275408 340656 275460
rect 459560 275408 459612 275460
rect 459652 275408 459704 275460
rect 626172 275408 626224 275460
rect 66996 275340 67048 275392
rect 187700 275340 187752 275392
rect 208860 275340 208912 275392
rect 233884 275340 233936 275392
rect 249064 275340 249116 275392
rect 260748 275340 260800 275392
rect 336648 275340 336700 275392
rect 448888 275340 448940 275392
rect 448980 275340 449032 275392
rect 633348 275340 633400 275392
rect 71780 275272 71832 275324
rect 194876 275272 194928 275324
rect 206560 275272 206612 275324
rect 237380 275272 237432 275324
rect 240784 275272 240836 275324
rect 258264 275272 258316 275324
rect 263232 275272 263284 275324
rect 266544 275272 266596 275324
rect 388168 275272 388220 275324
rect 402796 275272 402848 275324
rect 412548 275272 412600 275324
rect 647516 275272 647568 275324
rect 128544 275204 128596 275256
rect 131120 275204 131172 275256
rect 156880 275204 156932 275256
rect 204904 275204 204956 275256
rect 234896 275204 234948 275256
rect 235908 275204 235960 275256
rect 259736 275204 259788 275256
rect 264980 275204 265032 275256
rect 346124 275204 346176 275256
rect 473728 275204 473780 275256
rect 474188 275204 474240 275256
rect 577780 275204 577832 275256
rect 139124 275136 139176 275188
rect 185032 275136 185084 275188
rect 188804 275136 188856 275188
rect 210424 275136 210476 275188
rect 343364 275136 343416 275188
rect 466644 275136 466696 275188
rect 466736 275136 466788 275188
rect 510344 275136 510396 275188
rect 178132 275068 178184 275120
rect 221464 275068 221516 275120
rect 335176 275068 335228 275120
rect 441804 275068 441856 275120
rect 185216 275000 185268 275052
rect 214564 275000 214616 275052
rect 329656 275000 329708 275052
rect 427636 275000 427688 275052
rect 427728 275000 427780 275052
rect 458364 275000 458416 275052
rect 260932 274932 260984 274984
rect 265072 274932 265124 274984
rect 375196 274932 375248 274984
rect 434720 274932 434772 274984
rect 401784 274864 401836 274916
rect 407488 274864 407540 274916
rect 409972 274864 410024 274916
rect 419356 274864 419408 274916
rect 243176 274796 243228 274848
rect 245844 274796 245896 274848
rect 250260 274796 250312 274848
rect 254216 274796 254268 274848
rect 407028 274796 407080 274848
rect 411076 274796 411128 274848
rect 458180 274796 458232 274848
rect 461860 274796 461912 274848
rect 262128 274728 262180 274780
rect 265900 274728 265952 274780
rect 401600 274728 401652 274780
rect 406292 274728 406344 274780
rect 408592 274728 408644 274780
rect 412272 274728 412324 274780
rect 516140 274728 516192 274780
rect 74080 274660 74132 274712
rect 76012 274660 76064 274712
rect 88340 274660 88392 274712
rect 93124 274660 93176 274712
rect 160468 274660 160520 274712
rect 161388 274660 161440 274712
rect 220728 274660 220780 274712
rect 223580 274660 223632 274712
rect 225420 274660 225472 274712
rect 229836 274660 229888 274712
rect 264428 274660 264480 274712
rect 266728 274660 266780 274712
rect 266820 274660 266872 274712
rect 267740 274660 267792 274712
rect 398840 274660 398892 274712
rect 403992 274660 404044 274712
rect 404268 274660 404320 274712
rect 409880 274660 409932 274712
rect 510528 274660 510580 274712
rect 517428 274660 517480 274712
rect 521016 274660 521068 274712
rect 136824 274592 136876 274644
rect 218244 274592 218296 274644
rect 297364 274592 297416 274644
rect 319996 274592 320048 274644
rect 320088 274592 320140 274644
rect 338948 274592 339000 274644
rect 348516 274592 348568 274644
rect 479616 274592 479668 274644
rect 145012 274524 145064 274576
rect 222200 274524 222252 274576
rect 309784 274524 309836 274576
rect 333060 274524 333112 274576
rect 350356 274524 350408 274576
rect 483204 274524 483256 274576
rect 137928 274456 137980 274508
rect 219624 274456 219676 274508
rect 289636 274456 289688 274508
rect 321192 274456 321244 274508
rect 351736 274456 351788 274508
rect 486700 274456 486752 274508
rect 123760 274388 123812 274440
rect 214104 274388 214156 274440
rect 291844 274388 291896 274440
rect 311716 274388 311768 274440
rect 317788 274388 317840 274440
rect 349620 274388 349672 274440
rect 353024 274388 353076 274440
rect 490288 274388 490340 274440
rect 121368 274320 121420 274372
rect 213092 274320 213144 274372
rect 295984 274320 296036 274372
rect 329472 274320 329524 274372
rect 357256 274320 357308 274372
rect 500868 274320 500920 274372
rect 42156 274252 42208 274304
rect 42984 274252 43036 274304
rect 116676 274252 116728 274304
rect 211344 274252 211396 274304
rect 237288 274252 237340 274304
rect 256884 274252 256936 274304
rect 288348 274252 288400 274304
rect 318800 274252 318852 274304
rect 319444 274252 319496 274304
rect 353116 274252 353168 274304
rect 362592 274252 362644 274304
rect 518624 274252 518676 274304
rect 111984 274184 112036 274236
rect 208952 274184 209004 274236
rect 229008 274184 229060 274236
rect 253480 274184 253532 274236
rect 293684 274184 293736 274236
rect 335360 274184 335412 274236
rect 365628 274184 365680 274236
rect 525708 274184 525760 274236
rect 97724 274116 97776 274168
rect 203616 274116 203668 274168
rect 205364 274116 205416 274168
rect 244556 274116 244608 274168
rect 298008 274116 298060 274168
rect 346032 274116 346084 274168
rect 372528 274116 372580 274168
rect 543464 274116 543516 274168
rect 94228 274048 94280 274100
rect 201592 274048 201644 274100
rect 202972 274048 203024 274100
rect 242900 274048 242952 274100
rect 279424 274048 279476 274100
rect 288072 274048 288124 274100
rect 289728 274048 289780 274100
rect 322388 274048 322440 274100
rect 323676 274048 323728 274100
rect 374368 274048 374420 274100
rect 376668 274048 376720 274100
rect 551744 274048 551796 274100
rect 84752 273980 84804 274032
rect 198832 273980 198884 274032
rect 201776 273980 201828 274032
rect 242992 273980 243044 274032
rect 243544 273980 243596 274032
rect 251640 273980 251692 274032
rect 253848 273980 253900 274032
rect 262772 273980 262824 274032
rect 275928 273980 275980 274032
rect 285772 273980 285824 274032
rect 287704 273980 287756 274032
rect 297548 273980 297600 274032
rect 303344 273980 303396 274032
rect 360200 273980 360252 274032
rect 378048 273980 378100 274032
rect 558828 273980 558880 274032
rect 72976 273912 73028 273964
rect 194600 273912 194652 273964
rect 195888 273912 195940 273964
rect 240232 273912 240284 273964
rect 277308 273912 277360 273964
rect 289268 273912 289320 273964
rect 291108 273912 291160 273964
rect 324780 273912 324832 273964
rect 326344 273912 326396 273964
rect 385040 273912 385092 273964
rect 390376 273912 390428 273964
rect 590752 273912 590804 273964
rect 155684 273844 155736 273896
rect 225880 273844 225932 273896
rect 245568 273844 245620 273896
rect 259644 273844 259696 273896
rect 307024 273844 307076 273896
rect 325976 273844 326028 273896
rect 347688 273844 347740 273896
rect 476120 273844 476172 273896
rect 132040 273776 132092 273828
rect 196624 273776 196676 273828
rect 197084 273776 197136 273828
rect 236644 273776 236696 273828
rect 305644 273776 305696 273828
rect 315304 273776 315356 273828
rect 315396 273776 315448 273828
rect 328276 273776 328328 273828
rect 346216 273776 346268 273828
rect 472532 273776 472584 273828
rect 182916 273708 182968 273760
rect 231124 273708 231176 273760
rect 311164 273708 311216 273760
rect 323584 273708 323636 273760
rect 344560 273708 344612 273760
rect 468944 273708 468996 273760
rect 194692 273640 194744 273692
rect 240140 273640 240192 273692
rect 343456 273640 343508 273692
rect 465448 273640 465500 273692
rect 204168 273572 204220 273624
rect 239404 273572 239456 273624
rect 273168 273572 273220 273624
rect 279792 273572 279844 273624
rect 341892 273572 341944 273624
rect 458180 273572 458232 273624
rect 187700 273504 187752 273556
rect 192392 273504 192444 273556
rect 327724 273504 327776 273556
rect 416964 273504 417016 273556
rect 340696 273436 340748 273488
rect 427728 273436 427780 273488
rect 322204 273368 322256 273420
rect 367284 273368 367336 273420
rect 319536 273232 319588 273284
rect 320088 273232 320140 273284
rect 148600 273164 148652 273216
rect 222292 273164 222344 273216
rect 303528 273164 303580 273216
rect 357900 273164 357952 273216
rect 368296 273164 368348 273216
rect 532792 273164 532844 273216
rect 141516 273096 141568 273148
rect 220820 273096 220872 273148
rect 306288 273096 306340 273148
rect 364984 273096 365036 273148
rect 394424 273096 394476 273148
rect 583760 273096 583812 273148
rect 42156 273028 42208 273080
rect 44456 273028 44508 273080
rect 131120 273028 131172 273080
rect 216036 273028 216088 273080
rect 313096 273028 313148 273080
rect 383844 273028 383896 273080
rect 397276 273028 397328 273080
rect 593420 273028 593472 273080
rect 127348 272960 127400 273012
rect 215392 272960 215444 273012
rect 314476 272960 314528 273012
rect 387432 272960 387484 273012
rect 398932 272960 398984 273012
rect 600044 272960 600096 273012
rect 120264 272892 120316 272944
rect 212632 272892 212684 272944
rect 315856 272892 315908 272944
rect 390928 272892 390980 272944
rect 398656 272892 398708 272944
rect 597836 272892 597888 272944
rect 113180 272824 113232 272876
rect 209964 272824 210016 272876
rect 288440 272824 288492 272876
rect 304632 272824 304684 272876
rect 317236 272824 317288 272876
rect 394516 272824 394568 272876
rect 400312 272824 400364 272876
rect 617984 272824 618036 272876
rect 108396 272756 108448 272808
rect 207572 272756 207624 272808
rect 233700 272756 233752 272808
rect 255504 272756 255556 272808
rect 282736 272756 282788 272808
rect 305828 272756 305880 272808
rect 318616 272756 318668 272808
rect 398012 272756 398064 272808
rect 401968 272756 402020 272808
rect 621480 272756 621532 272808
rect 101312 272688 101364 272740
rect 204812 272688 204864 272740
rect 222476 272688 222528 272740
rect 247224 272688 247276 272740
rect 285588 272688 285640 272740
rect 308220 272688 308272 272740
rect 321284 272688 321336 272740
rect 401600 272688 401652 272740
rect 402980 272688 403032 272740
rect 625068 272688 625120 272740
rect 89536 272620 89588 272672
rect 200488 272620 200540 272672
rect 200580 272620 200632 272672
rect 243084 272620 243136 272672
rect 285404 272620 285456 272672
rect 312912 272620 312964 272672
rect 319904 272620 319956 272672
rect 401692 272620 401744 272672
rect 405648 272620 405700 272672
rect 632152 272620 632204 272672
rect 76012 272552 76064 272604
rect 194784 272552 194836 272604
rect 198280 272552 198332 272604
rect 241888 272552 241940 272604
rect 246764 272552 246816 272604
rect 260104 272552 260156 272604
rect 285864 272552 285916 272604
rect 314108 272552 314160 272604
rect 321376 272552 321428 272604
rect 405188 272552 405240 272604
rect 408316 272552 408368 272604
rect 639236 272552 639288 272604
rect 68192 272484 68244 272536
rect 193220 272484 193272 272536
rect 193496 272484 193548 272536
rect 240324 272484 240376 272536
rect 241980 272484 242032 272536
rect 258356 272484 258408 272536
rect 274732 272484 274784 272536
rect 284576 272484 284628 272536
rect 286784 272484 286836 272536
rect 316500 272484 316552 272536
rect 321192 272484 321244 272536
rect 408408 272484 408460 272536
rect 409604 272484 409656 272536
rect 642732 272484 642784 272536
rect 159272 272416 159324 272468
rect 226892 272416 226944 272468
rect 301504 272416 301556 272468
rect 317696 272416 317748 272468
rect 358636 272416 358688 272468
rect 504456 272416 504508 272468
rect 179328 272348 179380 272400
rect 233792 272348 233844 272400
rect 363604 272348 363656 272400
rect 392124 272348 392176 272400
rect 393136 272348 393188 272400
rect 521568 272348 521620 272400
rect 191196 272280 191248 272332
rect 239220 272280 239272 272332
rect 391756 272280 391808 272332
rect 513472 272280 513524 272332
rect 153292 272212 153344 272264
rect 192484 272212 192536 272264
rect 192576 272212 192628 272264
rect 238852 272212 238904 272264
rect 322664 272212 322716 272264
rect 408592 272212 408644 272264
rect 410432 272212 410484 272264
rect 199476 272144 199528 272196
rect 241612 272144 241664 272196
rect 325608 272144 325660 272196
rect 409972 272144 410024 272196
rect 422944 272212 422996 272264
rect 431132 272212 431184 272264
rect 431224 272212 431276 272264
rect 438216 272212 438268 272264
rect 424048 272144 424100 272196
rect 322756 272076 322808 272128
rect 404268 272076 404320 272128
rect 404360 272076 404412 272128
rect 459652 272076 459704 272128
rect 349804 272008 349856 272060
rect 422852 272008 422904 272060
rect 347044 271940 347096 271992
rect 415768 271940 415820 271992
rect 273812 271872 273864 271924
rect 282184 271872 282236 271924
rect 360844 271872 360896 271924
rect 399208 271872 399260 271924
rect 403440 271872 403492 271924
rect 404360 271872 404412 271924
rect 161572 271804 161624 271856
rect 227812 271804 227864 271856
rect 295248 271804 295300 271856
rect 336556 271804 336608 271856
rect 366916 271804 366968 271856
rect 529296 271804 529348 271856
rect 142712 271736 142764 271788
rect 162124 271736 162176 271788
rect 162768 271736 162820 271788
rect 228272 271736 228324 271788
rect 296444 271736 296496 271788
rect 340144 271736 340196 271788
rect 368112 271736 368164 271788
rect 531596 271736 531648 271788
rect 93032 271668 93084 271720
rect 153844 271668 153896 271720
rect 158076 271668 158128 271720
rect 226432 271668 226484 271720
rect 300768 271668 300820 271720
rect 350724 271668 350776 271720
rect 360016 271668 360068 271720
rect 362224 271668 362276 271720
rect 369492 271668 369544 271720
rect 535184 271668 535236 271720
rect 152188 271600 152240 271652
rect 224500 271600 224552 271652
rect 303160 271600 303212 271652
rect 359004 271600 359056 271652
rect 365536 271600 365588 271652
rect 367008 271600 367060 271652
rect 370780 271600 370832 271652
rect 538772 271600 538824 271652
rect 150992 271532 151044 271584
rect 223672 271532 223724 271584
rect 241428 271532 241480 271584
rect 251272 271532 251324 271584
rect 304448 271532 304500 271584
rect 362316 271532 362368 271584
rect 362684 271532 362736 271584
rect 363512 271532 363564 271584
rect 372160 271532 372212 271584
rect 542268 271532 542320 271584
rect 78864 271464 78916 271516
rect 152464 271464 152516 271516
rect 154488 271464 154540 271516
rect 225052 271464 225104 271516
rect 233884 271464 233936 271516
rect 246028 271464 246080 271516
rect 306196 271464 306248 271516
rect 366088 271464 366140 271516
rect 373816 271464 373868 271516
rect 547052 271464 547104 271516
rect 143908 271396 143960 271448
rect 96620 271328 96672 271380
rect 144184 271328 144236 271380
rect 147404 271396 147456 271448
rect 222476 271396 222528 271448
rect 224960 271396 225012 271448
rect 245936 271396 245988 271448
rect 281540 271396 281592 271448
rect 294052 271396 294104 271448
rect 307484 271396 307536 271448
rect 369676 271396 369728 271448
rect 375288 271396 375340 271448
rect 550548 271396 550600 271448
rect 220912 271328 220964 271380
rect 231400 271328 231452 271380
rect 254308 271328 254360 271380
rect 275652 271328 275704 271380
rect 286508 271328 286560 271380
rect 124956 271260 125008 271312
rect 214012 271260 214064 271312
rect 230204 271260 230256 271312
rect 254032 271260 254084 271312
rect 254216 271260 254268 271312
rect 261484 271260 261536 271312
rect 273352 271260 273404 271312
rect 280988 271260 281040 271312
rect 114284 271192 114336 271244
rect 209872 271192 209924 271244
rect 226616 271192 226668 271244
rect 252652 271192 252704 271244
rect 256148 271192 256200 271244
rect 263692 271192 263744 271244
rect 279148 271192 279200 271244
rect 296352 271328 296404 271380
rect 307576 271328 307628 271380
rect 370872 271328 370924 271380
rect 376576 271328 376628 271380
rect 554136 271328 554188 271380
rect 287796 271260 287848 271312
rect 303436 271260 303488 271312
rect 308956 271260 309008 271312
rect 373264 271260 373316 271312
rect 377956 271260 378008 271312
rect 557632 271260 557684 271312
rect 104900 271124 104952 271176
rect 206284 271124 206336 271176
rect 223580 271124 223632 271176
rect 250352 271124 250404 271176
rect 252928 271124 252980 271176
rect 262312 271124 262364 271176
rect 280528 271124 280580 271176
rect 299940 271192 299992 271244
rect 310336 271192 310388 271244
rect 376760 271192 376812 271244
rect 379428 271192 379480 271244
rect 561220 271192 561272 271244
rect 165160 271056 165212 271108
rect 229284 271056 229336 271108
rect 168656 270988 168708 271040
rect 230664 270988 230716 271040
rect 280988 270988 281040 271040
rect 301136 271124 301188 271176
rect 311808 271124 311860 271176
rect 380348 271124 380400 271176
rect 385960 271124 386012 271176
rect 578884 271124 578936 271176
rect 312452 271056 312504 271108
rect 343640 271056 343692 271108
rect 367008 271056 367060 271108
rect 528100 271056 528152 271108
rect 333244 270988 333296 271040
rect 354312 270988 354364 271040
rect 365444 270988 365496 271040
rect 524512 270988 524564 271040
rect 172244 270920 172296 270972
rect 232044 270920 232096 270972
rect 286968 270920 287020 270972
rect 287796 270920 287848 270972
rect 327816 270920 327868 270972
rect 347228 270920 347280 270972
rect 364156 270920 364208 270972
rect 516140 270920 516192 270972
rect 175832 270852 175884 270904
rect 233424 270852 233476 270904
rect 362776 270852 362828 270904
rect 510528 270852 510580 270904
rect 190000 270784 190052 270836
rect 235356 270784 235408 270836
rect 361488 270784 361540 270836
rect 496728 270784 496780 270836
rect 221924 270716 221976 270768
rect 238116 270716 238168 270768
rect 359924 270716 359976 270768
rect 466736 270716 466788 270768
rect 329564 270648 329616 270700
rect 429936 270648 429988 270700
rect 332324 270580 332376 270632
rect 375196 270580 375248 270632
rect 70584 270444 70636 270496
rect 71780 270444 71832 270496
rect 169852 270444 169904 270496
rect 231492 270444 231544 270496
rect 296536 270444 296588 270496
rect 342260 270444 342312 270496
rect 346400 270444 346452 270496
rect 474740 270444 474792 270496
rect 166908 270376 166960 270428
rect 230204 270376 230256 270428
rect 297456 270376 297508 270428
rect 343824 270376 343876 270428
rect 354864 270376 354916 270428
rect 496820 270376 496872 270428
rect 140688 270308 140740 270360
rect 219992 270308 220044 270360
rect 220636 270308 220688 270360
rect 224408 270308 224460 270360
rect 298744 270308 298796 270360
rect 347780 270308 347832 270360
rect 360200 270308 360252 270360
rect 510620 270308 510672 270360
rect 133788 270240 133840 270292
rect 216956 270240 217008 270292
rect 300124 270240 300176 270292
rect 351920 270240 351972 270292
rect 364248 270240 364300 270292
rect 521660 270240 521712 270292
rect 129648 270172 129700 270224
rect 215944 270172 215996 270224
rect 301412 270172 301464 270224
rect 354680 270172 354732 270224
rect 369584 270172 369636 270224
rect 535460 270172 535512 270224
rect 103704 270104 103756 270156
rect 125968 270104 126020 270156
rect 126888 270104 126940 270156
rect 214656 270104 214708 270156
rect 119068 270036 119120 270088
rect 110788 269968 110840 270020
rect 119620 269968 119672 270020
rect 122748 270036 122800 270088
rect 212908 270036 212960 270088
rect 234620 270036 234672 270088
rect 248052 270104 248104 270156
rect 301872 270104 301924 270156
rect 356060 270104 356112 270156
rect 374000 270104 374052 270156
rect 547880 270104 547932 270156
rect 211896 269968 211948 270020
rect 237380 269968 237432 270020
rect 245292 270036 245344 270088
rect 248328 270036 248380 270088
rect 260932 270036 260984 270088
rect 293408 270036 293460 270088
rect 333980 270036 334032 270088
rect 339776 270036 339828 270088
rect 456800 270036 456852 270088
rect 457996 270036 458048 270088
rect 636200 270036 636252 270088
rect 244372 269968 244424 270020
rect 259552 269968 259604 270020
rect 303344 269968 303396 270020
rect 303528 269968 303580 270020
rect 304540 269968 304592 270020
rect 362960 269968 363012 270020
rect 381636 269968 381688 270020
rect 567200 269968 567252 270020
rect 85948 269900 86000 269952
rect 110512 269900 110564 269952
rect 118608 269900 118660 269952
rect 212356 269900 212408 269952
rect 236092 269900 236144 269952
rect 256424 269900 256476 269952
rect 274272 269900 274324 269952
rect 282920 269900 282972 269952
rect 283564 269900 283616 269952
rect 292580 269900 292632 269952
rect 314292 269900 314344 269952
rect 376944 269900 376996 269952
rect 380716 269900 380768 269952
rect 565912 269900 565964 269952
rect 77208 269832 77260 269884
rect 113180 269832 113232 269884
rect 115848 269832 115900 269884
rect 210608 269832 210660 269884
rect 227720 269832 227772 269884
rect 248420 269832 248472 269884
rect 276940 269832 276992 269884
rect 289820 269832 289872 269884
rect 294788 269832 294840 269884
rect 336740 269832 336792 269884
rect 337108 269832 337160 269884
rect 449900 269832 449952 269884
rect 451372 269832 451424 269884
rect 644480 269832 644532 269884
rect 110328 269764 110380 269816
rect 208860 269764 208912 269816
rect 216680 269764 216732 269816
rect 229468 269764 229520 269816
rect 229836 269764 229888 269816
rect 252468 269764 252520 269816
rect 278688 269764 278740 269816
rect 294144 269764 294196 269816
rect 319260 269764 319312 269816
rect 388168 269764 388220 269816
rect 388720 269764 388772 269816
rect 586520 269764 586572 269816
rect 173808 269696 173860 269748
rect 232872 269696 232924 269748
rect 296076 269696 296128 269748
rect 340880 269696 340932 269748
rect 345112 269696 345164 269748
rect 470600 269696 470652 269748
rect 470692 269696 470744 269748
rect 476304 269696 476356 269748
rect 176936 269628 176988 269680
rect 234160 269628 234212 269680
rect 292580 269628 292632 269680
rect 331220 269628 331272 269680
rect 343732 269628 343784 269680
rect 467840 269628 467892 269680
rect 180708 269560 180760 269612
rect 235540 269560 235592 269612
rect 292120 269560 292172 269612
rect 329840 269560 329892 269612
rect 342444 269560 342496 269612
rect 463700 269560 463752 269612
rect 135628 269492 135680 269544
rect 184756 269492 184808 269544
rect 184848 269492 184900 269544
rect 236920 269492 236972 269544
rect 290740 269492 290792 269544
rect 327080 269492 327132 269544
rect 341064 269492 341116 269544
rect 459744 269492 459796 269544
rect 187516 269424 187568 269476
rect 238208 269424 238260 269476
rect 338396 269424 338448 269476
rect 452660 269424 452712 269476
rect 335728 269356 335780 269408
rect 445760 269356 445812 269408
rect 334348 269288 334400 269340
rect 443000 269288 443052 269340
rect 353300 269220 353352 269272
rect 380900 269220 380952 269272
rect 102508 269016 102560 269068
rect 206192 269016 206244 269068
rect 249616 269016 249668 269068
rect 253388 269016 253440 269068
rect 303712 269016 303764 269068
rect 360384 269016 360436 269068
rect 361580 269016 361632 269068
rect 514760 269016 514812 269068
rect 99288 268948 99340 269000
rect 204444 268948 204496 269000
rect 249708 268948 249760 269000
rect 257804 268948 257856 269000
rect 308864 268948 308916 269000
rect 375380 268948 375432 269000
rect 391848 268948 391900 269000
rect 543740 268948 543792 269000
rect 95424 268880 95476 268932
rect 203524 268880 203576 268932
rect 306656 268880 306708 268932
rect 368480 268880 368532 268932
rect 370872 268880 370924 268932
rect 539600 268880 539652 268932
rect 92388 268812 92440 268864
rect 202144 268812 202196 268864
rect 321008 268812 321060 268864
rect 401784 268812 401836 268864
rect 404360 268812 404412 268864
rect 587900 268812 587952 268864
rect 87144 268744 87196 268796
rect 200396 268744 200448 268796
rect 204904 268744 204956 268796
rect 226708 268744 226760 268796
rect 310428 268744 310480 268796
rect 378140 268744 378192 268796
rect 393228 268744 393280 268796
rect 581644 268744 581696 268796
rect 82728 268676 82780 268728
rect 198556 268676 198608 268728
rect 218336 268676 218388 268728
rect 242808 268676 242860 268728
rect 277400 268676 277452 268728
rect 291200 268676 291252 268728
rect 313004 268676 313056 268728
rect 385224 268676 385276 268728
rect 394056 268676 394108 268728
rect 600320 268676 600372 268728
rect 80060 268608 80112 268660
rect 197268 268608 197320 268660
rect 219532 268608 219584 268660
rect 250260 268608 250312 268660
rect 280068 268608 280120 268660
rect 298100 268608 298152 268660
rect 314384 268608 314436 268660
rect 389180 268608 389232 268660
rect 394516 268608 394568 268660
rect 601700 268608 601752 268660
rect 77668 268540 77720 268592
rect 196808 268540 196860 268592
rect 217140 268540 217192 268592
rect 249340 268540 249392 268592
rect 289912 268540 289964 268592
rect 310520 268540 310572 268592
rect 315672 268540 315724 268592
rect 393320 268540 393372 268592
rect 395804 268540 395856 268592
rect 605840 268540 605892 268592
rect 75828 268472 75880 268524
rect 195428 268472 195480 268524
rect 216588 268472 216640 268524
rect 248880 268472 248932 268524
rect 283196 268472 283248 268524
rect 306380 268472 306432 268524
rect 317052 268472 317104 268524
rect 396080 268472 396132 268524
rect 397184 268472 397236 268524
rect 608600 268472 608652 268524
rect 69388 268404 69440 268456
rect 193680 268404 193732 268456
rect 213460 268404 213512 268456
rect 245752 268404 245804 268456
rect 245844 268404 245896 268456
rect 259184 268404 259236 268456
rect 281448 268404 281500 268456
rect 302240 268404 302292 268456
rect 319720 268404 319772 268456
rect 398840 268404 398892 268456
rect 399852 268404 399904 268456
rect 615684 268404 615736 268456
rect 66168 268336 66220 268388
rect 192116 268336 192168 268388
rect 211252 268336 211304 268388
rect 247132 268336 247184 268388
rect 257988 268336 258040 268388
rect 264520 268336 264572 268388
rect 284116 268336 284168 268388
rect 309140 268336 309192 268388
rect 318340 268336 318392 268388
rect 400220 268336 400272 268388
rect 401140 268336 401192 268388
rect 619640 268336 619692 268388
rect 106188 268268 106240 268320
rect 207480 268268 207532 268320
rect 307668 268268 307720 268320
rect 371332 268268 371384 268320
rect 372712 268268 372764 268320
rect 391940 268268 391992 268320
rect 131028 268200 131080 268252
rect 216864 268200 216916 268252
rect 339408 268200 339460 268252
rect 382280 268200 382332 268252
rect 388168 268200 388220 268252
rect 502248 268200 502300 268252
rect 135168 268132 135220 268184
rect 218152 268132 218204 268184
rect 386512 268132 386564 268184
rect 487160 268132 487212 268184
rect 186412 268064 186464 268116
rect 237288 268064 237340 268116
rect 331128 268064 331180 268116
rect 419540 268064 419592 268116
rect 663064 268064 663116 268116
rect 676220 268064 676272 268116
rect 185032 267996 185084 268048
rect 220360 267996 220412 268048
rect 385132 267996 385184 268048
rect 474188 267996 474240 268048
rect 195980 267928 196032 267980
rect 223028 267928 223080 267980
rect 322388 267928 322440 267980
rect 407028 267928 407080 267980
rect 661868 267928 661920 267980
rect 676220 267928 676272 267980
rect 343640 267860 343692 267912
rect 426440 267860 426492 267912
rect 371884 267792 371936 267844
rect 394700 267792 394752 267844
rect 409880 267792 409932 267844
rect 412640 267792 412692 267844
rect 365720 267724 365772 267776
rect 387800 267724 387852 267776
rect 390468 267724 390520 267776
rect 523684 267724 523736 267776
rect 660304 267724 660356 267776
rect 676128 267724 676180 267776
rect 175188 267656 175240 267708
rect 233792 267656 233844 267708
rect 276480 267656 276532 267708
rect 277308 267656 277360 267708
rect 287612 267656 287664 267708
rect 288348 267656 288400 267708
rect 289820 267656 289872 267708
rect 291108 267656 291160 267708
rect 299204 267656 299256 267708
rect 309324 267656 309376 267708
rect 311716 267656 311768 267708
rect 162124 267588 162176 267640
rect 221740 267588 221792 267640
rect 231124 267588 231176 267640
rect 236000 267588 236052 267640
rect 300584 267588 300636 267640
rect 319444 267588 319496 267640
rect 144184 267520 144236 267572
rect 204352 267520 204404 267572
rect 284944 267520 284996 267572
rect 291844 267520 291896 267572
rect 295156 267520 295208 267572
rect 319536 267520 319588 267572
rect 168288 267452 168340 267504
rect 231124 267452 231176 267504
rect 287152 267452 287204 267504
rect 301504 267452 301556 267504
rect 306380 267452 306432 267504
rect 311164 267452 311216 267504
rect 311256 267452 311308 267504
rect 316040 267452 316092 267504
rect 344652 267656 344704 267708
rect 469220 267656 469272 267708
rect 324136 267588 324188 267640
rect 347044 267588 347096 267640
rect 349988 267588 350040 267640
rect 483388 267588 483440 267640
rect 326804 267520 326856 267572
rect 349804 267520 349856 267572
rect 352656 267520 352708 267572
rect 491392 267520 491444 267572
rect 339408 267452 339460 267504
rect 355324 267452 355376 267504
rect 498200 267452 498252 267504
rect 161388 267384 161440 267436
rect 228456 267384 228508 267436
rect 236644 267384 236696 267436
rect 241796 267384 241848 267436
rect 278320 267384 278372 267436
rect 281540 267384 281592 267436
rect 283656 267384 283708 267436
rect 285588 267384 285640 267436
rect 298284 267384 298336 267436
rect 327816 267384 327868 267436
rect 357992 267384 358044 267436
rect 505100 267384 505152 267436
rect 125968 267316 126020 267368
rect 207020 267316 207072 267368
rect 276020 267316 276072 267368
rect 279424 267316 279476 267368
rect 288072 267316 288124 267368
rect 297364 267316 297416 267368
rect 300952 267316 301004 267368
rect 333244 267316 333296 267368
rect 360660 267316 360712 267368
rect 512000 267316 512052 267368
rect 113180 267248 113232 267300
rect 196348 267248 196400 267300
rect 196624 267248 196676 267300
rect 217692 267248 217744 267300
rect 238116 267248 238168 267300
rect 251088 267248 251140 267300
rect 281816 267248 281868 267300
rect 286968 267248 287020 267300
rect 288532 267248 288584 267300
rect 289636 267248 289688 267300
rect 292948 267248 293000 267300
rect 110512 267180 110564 267232
rect 199936 267180 199988 267232
rect 221464 267180 221516 267232
rect 235080 267180 235132 267232
rect 235908 267180 235960 267232
rect 256056 267180 256108 267232
rect 272524 267180 272576 267232
rect 277860 267180 277912 267232
rect 290280 267180 290332 267232
rect 307024 267180 307076 267232
rect 309324 267248 309376 267300
rect 317788 267248 317840 267300
rect 317880 267248 317932 267300
rect 360844 267248 360896 267300
rect 363328 267248 363380 267300
rect 518900 267248 518952 267300
rect 309784 267180 309836 267232
rect 313924 267180 313976 267232
rect 316040 267180 316092 267232
rect 316132 267180 316184 267232
rect 353300 267180 353352 267232
rect 119620 267112 119672 267164
rect 209688 267112 209740 267164
rect 226984 267112 227036 267164
rect 232412 267112 232464 267164
rect 233148 267112 233200 267164
rect 255136 267112 255188 267164
rect 255228 267112 255280 267164
rect 263600 267112 263652 267164
rect 286324 267112 286376 267164
rect 305644 267112 305696 267164
rect 93124 267044 93176 267096
rect 201224 267044 201276 267096
rect 214564 267044 214616 267096
rect 237748 267044 237800 267096
rect 238668 267044 238720 267096
rect 257344 267044 257396 267096
rect 289452 267044 289504 267096
rect 306380 267044 306432 267096
rect 71780 266976 71832 267028
rect 194140 266976 194192 267028
rect 210424 266976 210476 267028
rect 239128 266976 239180 267028
rect 252376 266976 252428 267028
rect 262220 266976 262272 267028
rect 272432 266976 272484 267028
rect 277768 266976 277820 267028
rect 279608 266976 279660 267028
rect 287704 266976 287756 267028
rect 291200 266976 291252 267028
rect 315212 267112 315264 267164
rect 363604 267180 363656 267232
rect 356244 267112 356296 267164
rect 357256 267112 357308 267164
rect 358912 267112 358964 267164
rect 360108 267112 360160 267164
rect 362040 267112 362092 267164
rect 362684 267112 362736 267164
rect 315396 267044 315448 267096
rect 316040 267044 316092 267096
rect 365720 267180 365772 267232
rect 365996 267180 366048 267232
rect 525800 267180 525852 267232
rect 368664 267112 368716 267164
rect 532884 267112 532936 267164
rect 371332 267044 371384 267096
rect 540980 267044 541032 267096
rect 182088 266908 182140 266960
rect 236460 266908 236512 266960
rect 153844 266840 153896 266892
rect 203064 266840 203116 266892
rect 152464 266772 152516 266824
rect 197728 266772 197780 266824
rect 296996 266772 297048 266824
rect 312452 266976 312504 267028
rect 316592 266976 316644 267028
rect 371884 266976 371936 267028
rect 375380 266976 375432 267028
rect 376668 266976 376720 267028
rect 382464 266976 382516 267028
rect 383476 266976 383528 267028
rect 397644 266976 397696 267028
rect 398656 266976 398708 267028
rect 399024 266976 399076 267028
rect 409880 266976 409932 267028
rect 417424 266976 417476 267028
rect 643100 266976 643152 267028
rect 673920 266976 673972 267028
rect 676036 266976 676088 267028
rect 184756 266704 184808 266756
rect 219072 266704 219124 266756
rect 282276 266704 282328 266756
rect 288440 266704 288492 266756
rect 192484 266636 192536 266688
rect 225788 266636 225840 266688
rect 305920 266636 305972 266688
rect 322204 266908 322256 266960
rect 324596 266908 324648 266960
rect 327724 266908 327776 266960
rect 328184 266908 328236 266960
rect 343640 266908 343692 266960
rect 347320 266908 347372 266960
rect 470692 266908 470744 266960
rect 271604 266568 271656 266620
rect 276296 266568 276348 266620
rect 277860 266568 277912 266620
rect 283564 266568 283616 266620
rect 308588 266568 308640 266620
rect 323676 266840 323728 266892
rect 341984 266840 342036 266892
rect 462320 266840 462372 266892
rect 339316 266772 339368 266824
rect 455420 266772 455472 266824
rect 312544 266704 312596 266756
rect 335268 266704 335320 266756
rect 444380 266704 444432 266756
rect 326344 266636 326396 266688
rect 329932 266636 329984 266688
rect 325976 266568 326028 266620
rect 331128 266568 331180 266620
rect 332600 266636 332652 266688
rect 431224 266636 431276 266688
rect 422944 266568 422996 266620
rect 673368 266568 673420 266620
rect 676220 266568 676272 266620
rect 271144 266500 271196 266552
rect 274640 266500 274692 266552
rect 323216 266500 323268 266552
rect 399024 266500 399076 266552
rect 239404 266432 239456 266484
rect 244464 266432 244516 266484
rect 270684 266432 270736 266484
rect 273260 266432 273312 266484
rect 291660 266432 291712 266484
rect 295984 266432 296036 266484
rect 305000 266432 305052 266484
rect 306288 266432 306340 266484
rect 309876 266432 309928 266484
rect 314292 266432 314344 266484
rect 320180 266432 320232 266484
rect 321376 266432 321428 266484
rect 328644 266432 328696 266484
rect 329656 266432 329708 266484
rect 233884 266364 233936 266416
rect 234620 266364 234672 266416
rect 235356 266364 235408 266416
rect 238668 266364 238720 266416
rect 242808 266364 242860 266416
rect 249800 266364 249852 266416
rect 270316 266364 270368 266416
rect 272064 266364 272116 266416
rect 284484 266364 284536 266416
rect 289912 266364 289964 266416
rect 294328 266364 294380 266416
rect 295248 266364 295300 266416
rect 295616 266364 295668 266416
rect 296444 266364 296496 266416
rect 299664 266364 299716 266416
rect 300768 266364 300820 266416
rect 302332 266364 302384 266416
rect 303436 266364 303488 266416
rect 305460 266364 305512 266416
rect 306196 266364 306248 266416
rect 306748 266364 306800 266416
rect 307484 266364 307536 266416
rect 308128 266364 308180 266416
rect 308956 266364 309008 266416
rect 309416 266364 309468 266416
rect 310336 266364 310388 266416
rect 310796 266364 310848 266416
rect 311808 266364 311860 266416
rect 312084 266364 312136 266416
rect 313096 266364 313148 266416
rect 313464 266364 313516 266416
rect 314476 266364 314528 266416
rect 314844 266364 314896 266416
rect 315856 266364 315908 266416
rect 316132 266364 316184 266416
rect 317236 266364 317288 266416
rect 317512 266364 317564 266416
rect 318616 266364 318668 266416
rect 318800 266364 318852 266416
rect 319904 266364 319956 266416
rect 320548 266364 320600 266416
rect 321284 266364 321336 266416
rect 321928 266364 321980 266416
rect 322756 266364 322808 266416
rect 327264 266364 327316 266416
rect 329012 266364 329064 266416
rect 329748 266364 329800 266416
rect 408776 266432 408828 266484
rect 409696 266432 409748 266484
rect 410064 266500 410116 266552
rect 417424 266500 417476 266552
rect 410432 266432 410484 266484
rect 411444 266432 411496 266484
rect 412548 266432 412600 266484
rect 673276 266432 673328 266484
rect 676220 266432 676272 266484
rect 331312 266364 331364 266416
rect 332324 266364 332376 266416
rect 333980 266364 334032 266416
rect 335176 266364 335228 266416
rect 340144 266364 340196 266416
rect 340696 266364 340748 266416
rect 342812 266364 342864 266416
rect 343456 266364 343508 266416
rect 345480 266364 345532 266416
rect 346216 266364 346268 266416
rect 346860 266364 346912 266416
rect 347688 266364 347740 266416
rect 347780 266364 347832 266416
rect 349068 266364 349120 266416
rect 349528 266364 349580 266416
rect 350356 266364 350408 266416
rect 350908 266364 350960 266416
rect 351736 266364 351788 266416
rect 352196 266364 352248 266416
rect 353024 266364 353076 266416
rect 356612 266364 356664 266416
rect 357348 266364 357400 266416
rect 357532 266364 357584 266416
rect 358636 266364 358688 266416
rect 359372 266364 359424 266416
rect 360016 266364 360068 266416
rect 362408 266364 362460 266416
rect 362776 266364 362828 266416
rect 364708 266364 364760 266416
rect 365536 266364 365588 266416
rect 366456 266364 366508 266416
rect 367008 266364 367060 266416
rect 367376 266364 367428 266416
rect 368388 266364 368440 266416
rect 370044 266364 370096 266416
rect 371056 266364 371108 266416
rect 376484 266364 376536 266416
rect 376668 266364 376720 266416
rect 378876 266364 378928 266416
rect 379428 266364 379480 266416
rect 379796 266364 379848 266416
rect 380808 266364 380860 266416
rect 382924 266364 382976 266416
rect 383568 266364 383620 266416
rect 390928 266364 390980 266416
rect 391756 266364 391808 266416
rect 392308 266364 392360 266416
rect 393136 266364 393188 266416
rect 393596 266364 393648 266416
rect 394424 266364 394476 266416
rect 396264 266364 396316 266416
rect 397276 266364 397328 266416
rect 398104 266364 398156 266416
rect 398748 266364 398800 266416
rect 409236 266364 409288 266416
rect 409788 266364 409840 266416
rect 410524 266364 410576 266416
rect 451372 266364 451424 266416
rect 354404 266296 354456 266348
rect 495440 266296 495492 266348
rect 357072 266228 357124 266280
rect 502340 266228 502392 266280
rect 373172 266160 373224 266212
rect 545120 266160 545172 266212
rect 374460 266092 374512 266144
rect 549260 266092 549312 266144
rect 375840 266024 375892 266076
rect 552020 266024 552072 266076
rect 674012 266024 674064 266076
rect 676220 266024 676272 266076
rect 377128 265956 377180 266008
rect 556160 265956 556212 266008
rect 378508 265888 378560 265940
rect 558920 265888 558972 265940
rect 380256 265820 380308 265872
rect 564440 265820 564492 265872
rect 674656 265820 674708 265872
rect 676036 265820 676088 265872
rect 381176 265752 381228 265804
rect 566004 265752 566056 265804
rect 384304 265684 384356 265736
rect 574284 265684 574336 265736
rect 28356 265616 28408 265668
rect 46296 265616 46348 265668
rect 383844 265616 383896 265668
rect 574100 265616 574152 265668
rect 194784 265548 194836 265600
rect 195612 265548 195664 265600
rect 201592 265548 201644 265600
rect 202236 265548 202288 265600
rect 209872 265548 209924 265600
rect 210700 265548 210752 265600
rect 214012 265548 214064 265600
rect 214748 265548 214800 265600
rect 222292 265548 222344 265600
rect 223212 265548 223264 265600
rect 238852 265548 238904 265600
rect 239680 265548 239732 265600
rect 240140 265548 240192 265600
rect 240508 265548 240560 265600
rect 241612 265548 241664 265600
rect 242348 265548 242400 265600
rect 242992 265548 243044 265600
rect 243268 265548 243320 265600
rect 266360 265548 266412 265600
rect 267280 265548 267332 265600
rect 351736 265548 351788 265600
rect 488540 265548 488592 265600
rect 194600 265480 194652 265532
rect 194968 265480 195020 265532
rect 240232 265480 240284 265532
rect 241060 265480 241112 265532
rect 242900 265480 242952 265532
rect 243636 265480 243688 265532
rect 349068 265480 349120 265532
rect 481640 265480 481692 265532
rect 333060 265412 333112 265464
rect 438860 265412 438912 265464
rect 330852 265344 330904 265396
rect 433340 265344 433392 265396
rect 330392 265276 330444 265328
rect 431960 265276 432012 265328
rect 327724 265208 327776 265260
rect 425060 265208 425112 265260
rect 325056 265140 325108 265192
rect 418160 265140 418212 265192
rect 245844 264936 245896 264988
rect 246396 264936 246448 264988
rect 673368 264936 673420 264988
rect 676220 264936 676272 264988
rect 337476 264528 337528 264580
rect 451280 264528 451332 264580
rect 353852 264460 353904 264512
rect 492680 264460 492732 264512
rect 384948 264392 385000 264444
rect 575480 264392 575532 264444
rect 387616 264324 387668 264376
rect 582564 264324 582616 264376
rect 393044 264256 393096 264308
rect 597560 264256 597612 264308
rect 45008 264188 45060 264240
rect 662512 264188 662564 264240
rect 399760 264120 399812 264172
rect 401232 264120 401284 264172
rect 607404 264120 607456 264172
rect 615500 264052 615552 264104
rect 673276 263576 673328 263628
rect 676220 263576 676272 263628
rect 675024 262624 675076 262676
rect 676036 262624 676088 262676
rect 415308 262216 415360 262268
rect 572720 262216 572772 262268
rect 675208 262216 675260 262268
rect 676036 262216 676088 262268
rect 674472 261944 674524 261996
rect 676220 261944 676272 261996
rect 674748 261536 674800 261588
rect 676220 261536 676272 261588
rect 673000 260856 673052 260908
rect 676220 260856 676272 260908
rect 674564 259904 674616 259956
rect 676220 259904 676272 259956
rect 675484 259360 675536 259412
rect 676312 259360 676364 259412
rect 185216 258340 185268 258392
rect 189080 258340 189132 258392
rect 673184 258136 673236 258188
rect 676220 258136 676272 258188
rect 414204 258068 414256 258120
rect 571524 258068 571576 258120
rect 673092 258068 673144 258120
rect 676128 258068 676180 258120
rect 31576 258000 31628 258052
rect 44364 258000 44416 258052
rect 31484 257864 31536 257916
rect 44916 257864 44968 257916
rect 31668 257728 31720 257780
rect 47676 257728 47728 257780
rect 671620 256708 671672 256760
rect 683120 256708 683172 256760
rect 415308 255280 415360 255332
rect 571432 255280 571484 255332
rect 414388 252560 414440 252612
rect 574744 252560 574796 252612
rect 674656 251676 674708 251728
rect 675024 251676 675076 251728
rect 675024 251540 675076 251592
rect 675484 251540 675536 251592
rect 675392 251200 675444 251252
rect 675392 250928 675444 250980
rect 674748 250180 674800 250232
rect 675484 250180 675536 250232
rect 675024 249704 675076 249756
rect 675392 249704 675444 249756
rect 674656 249568 674708 249620
rect 675024 249568 675076 249620
rect 675208 248480 675260 248532
rect 414204 248412 414256 248464
rect 438216 248412 438268 248464
rect 675208 248276 675260 248328
rect 675024 247868 675076 247920
rect 675484 247868 675536 247920
rect 673000 246984 673052 247036
rect 675392 246984 675444 247036
rect 35808 245624 35860 245676
rect 117964 245624 118016 245676
rect 415308 245624 415360 245676
rect 438124 245624 438176 245676
rect 674748 243856 674800 243908
rect 675116 243856 675168 243908
rect 675208 243856 675260 243908
rect 675300 243584 675352 243636
rect 414388 242904 414440 242956
rect 621664 242904 621716 242956
rect 32404 242292 32456 242344
rect 41972 242292 42024 242344
rect 31116 242224 31168 242276
rect 42432 242224 42484 242276
rect 31024 242156 31076 242208
rect 42708 242156 42760 242208
rect 674564 242156 674616 242208
rect 675392 242156 675444 242208
rect 673092 241612 673144 241664
rect 675300 241612 675352 241664
rect 175004 241544 175056 241596
rect 155868 240796 155920 240848
rect 673184 241068 673236 241120
rect 675300 241068 675352 241120
rect 42432 240048 42484 240100
rect 42800 240048 42852 240100
rect 42156 239980 42208 240032
rect 44180 239980 44232 240032
rect 414940 238756 414992 238808
rect 428464 238756 428516 238808
rect 674748 238756 674800 238808
rect 675392 238688 675444 238740
rect 438216 238008 438268 238060
rect 574100 238008 574152 238060
rect 184940 237396 184992 237448
rect 189080 237396 189132 237448
rect 153108 235968 153160 236020
rect 155868 235968 155920 236020
rect 42156 235356 42208 235408
rect 44640 235356 44692 235408
rect 42156 234540 42208 234592
rect 44548 234540 44600 234592
rect 42156 233996 42208 234048
rect 44916 233996 44968 234048
rect 130384 233860 130436 233912
rect 153108 233860 153160 233912
rect 438124 233860 438176 233912
rect 572812 233860 572864 233912
rect 42156 233248 42208 233300
rect 43168 233248 43220 233300
rect 415308 233248 415360 233300
rect 427084 233248 427136 233300
rect 177120 232500 177172 232552
rect 184848 232500 184900 232552
rect 414204 232500 414256 232552
rect 639604 232500 639656 232552
rect 427084 232432 427136 232484
rect 639144 232432 639196 232484
rect 428464 231752 428516 231804
rect 639052 231752 639104 231804
rect 190368 231684 190420 231736
rect 604460 231684 604512 231736
rect 191104 231616 191156 231668
rect 663800 231616 663852 231668
rect 65156 231548 65208 231600
rect 177120 231548 177172 231600
rect 189724 231548 189776 231600
rect 663892 231548 663944 231600
rect 55864 231480 55916 231532
rect 649356 231480 649408 231532
rect 64144 231412 64196 231464
rect 661040 231412 661092 231464
rect 54484 231344 54536 231396
rect 654140 231344 654192 231396
rect 50344 231276 50396 231328
rect 650644 231276 650696 231328
rect 51724 231208 51776 231260
rect 652760 231208 652812 231260
rect 53104 231140 53156 231192
rect 655520 231140 655572 231192
rect 42156 231072 42208 231124
rect 43260 231072 43312 231124
rect 43904 231072 43956 231124
rect 662604 231072 662656 231124
rect 42156 230528 42208 230580
rect 42432 230528 42484 230580
rect 179328 230392 179380 230444
rect 246120 230392 246172 230444
rect 262220 230392 262272 230444
rect 263232 230392 263284 230444
rect 263600 230392 263652 230444
rect 263784 230392 263836 230444
rect 175188 230324 175240 230376
rect 244648 230324 244700 230376
rect 246948 230324 247000 230376
rect 333612 230460 333664 230512
rect 274640 230392 274692 230444
rect 276756 230392 276808 230444
rect 277768 230392 277820 230444
rect 271328 230324 271380 230376
rect 272800 230324 272852 230376
rect 169668 230256 169720 230308
rect 241796 230256 241848 230308
rect 244188 230256 244240 230308
rect 274272 230256 274324 230308
rect 274548 230256 274600 230308
rect 285312 230392 285364 230444
rect 288348 230392 288400 230444
rect 292764 230392 292816 230444
rect 299940 230392 299992 230444
rect 303988 230392 304040 230444
rect 314936 230392 314988 230444
rect 315948 230392 316000 230444
rect 318800 230392 318852 230444
rect 326344 230392 326396 230444
rect 331312 230392 331364 230444
rect 332232 230392 332284 230444
rect 333060 230392 333112 230444
rect 333888 230392 333940 230444
rect 385132 230460 385184 230512
rect 507952 230460 508004 230512
rect 604460 230460 604512 230512
rect 605748 230460 605800 230512
rect 636844 230460 636896 230512
rect 371884 230392 371936 230444
rect 279424 230324 279476 230376
rect 283196 230324 283248 230376
rect 278044 230256 278096 230308
rect 287428 230324 287480 230376
rect 305644 230324 305696 230376
rect 306196 230324 306248 230376
rect 307024 230324 307076 230376
rect 307576 230324 307628 230376
rect 312084 230324 312136 230376
rect 313188 230324 313240 230376
rect 314568 230324 314620 230376
rect 286968 230256 287020 230308
rect 291752 230256 291804 230308
rect 316316 230324 316368 230376
rect 317328 230324 317380 230376
rect 317788 230324 317840 230376
rect 318708 230324 318760 230376
rect 319260 230324 319312 230376
rect 319904 230324 319956 230376
rect 320640 230324 320692 230376
rect 321376 230324 321428 230376
rect 321652 230324 321704 230376
rect 338764 230324 338816 230376
rect 341984 230324 342036 230376
rect 380716 230392 380768 230444
rect 393688 230392 393740 230444
rect 400680 230392 400732 230444
rect 401876 230392 401928 230444
rect 456156 230392 456208 230444
rect 374092 230324 374144 230376
rect 377404 230324 377456 230376
rect 390836 230324 390888 230376
rect 391848 230324 391900 230376
rect 393320 230324 393372 230376
rect 394608 230324 394660 230376
rect 397644 230324 397696 230376
rect 398564 230324 398616 230376
rect 399024 230324 399076 230376
rect 400128 230324 400180 230376
rect 403348 230324 403400 230376
rect 404176 230324 404228 230376
rect 404360 230324 404412 230376
rect 406660 230324 406712 230376
rect 406844 230324 406896 230376
rect 410984 230324 411036 230376
rect 411168 230324 411220 230376
rect 461584 230324 461636 230376
rect 319352 230256 319404 230308
rect 339132 230256 339184 230308
rect 378232 230256 378284 230308
rect 395436 230256 395488 230308
rect 396724 230256 396776 230308
rect 398656 230256 398708 230308
rect 400864 230256 400916 230308
rect 402980 230256 403032 230308
rect 404268 230256 404320 230308
rect 404728 230256 404780 230308
rect 409788 230256 409840 230308
rect 136364 230188 136416 230240
rect 213276 230188 213328 230240
rect 219256 230188 219308 230240
rect 262220 230188 262272 230240
rect 262772 230188 262824 230240
rect 269948 230188 270000 230240
rect 276664 230188 276716 230240
rect 287060 230188 287112 230240
rect 311716 230188 311768 230240
rect 315304 230188 315356 230240
rect 320272 230188 320324 230240
rect 337384 230188 337436 230240
rect 347688 230188 347740 230240
rect 386420 230188 386472 230240
rect 398104 230188 398156 230240
rect 403072 230188 403124 230240
rect 406200 230188 406252 230240
rect 467104 230256 467156 230308
rect 409972 230188 410024 230240
rect 469220 230188 469272 230240
rect 155868 230120 155920 230172
rect 236092 230120 236144 230172
rect 240048 230120 240100 230172
rect 271788 230120 271840 230172
rect 275284 230120 275336 230172
rect 277676 230120 277728 230172
rect 277768 230120 277820 230172
rect 286048 230120 286100 230172
rect 317420 230120 317472 230172
rect 334624 230120 334676 230172
rect 336648 230120 336700 230172
rect 376024 230120 376076 230172
rect 378324 230120 378376 230172
rect 443644 230120 443696 230172
rect 146208 230052 146260 230104
rect 231860 230052 231912 230104
rect 233148 230052 233200 230104
rect 139308 229984 139360 230036
rect 229008 229984 229060 230036
rect 234528 229984 234580 230036
rect 262772 229984 262824 230036
rect 271144 230052 271196 230104
rect 277124 230052 277176 230104
rect 277216 230052 277268 230104
rect 282460 230052 282512 230104
rect 315856 230052 315908 230104
rect 322204 230052 322256 230104
rect 323768 230052 323820 230104
rect 364524 230052 364576 230104
rect 387984 230052 388036 230104
rect 515404 230052 515456 230104
rect 268936 229984 268988 230036
rect 270408 229984 270460 230036
rect 283840 229984 283892 230036
rect 285496 229984 285548 230036
rect 290648 229984 290700 230036
rect 312360 229984 312412 230036
rect 337016 229984 337068 230036
rect 343732 229984 343784 230036
rect 385684 229984 385736 230036
rect 387616 229984 387668 230036
rect 399484 229984 399536 230036
rect 400864 229984 400916 230036
rect 407764 229984 407816 230036
rect 408316 229984 408368 230036
rect 132408 229916 132460 229968
rect 226156 229916 226208 229968
rect 226248 229916 226300 229968
rect 259920 229916 259972 229968
rect 260104 229916 260156 229968
rect 262864 229916 262916 229968
rect 270316 229916 270368 229968
rect 284576 229916 284628 229968
rect 285588 229916 285640 229968
rect 291384 229916 291436 229968
rect 313832 229916 313884 229968
rect 341248 229916 341300 229968
rect 345572 229916 345624 229968
rect 354772 229916 354824 229968
rect 356244 229916 356296 229968
rect 357072 229916 357124 229968
rect 359096 229916 359148 229968
rect 360108 229916 360160 229968
rect 360568 229916 360620 229968
rect 361304 229916 361356 229968
rect 361948 229916 362000 229968
rect 362684 229916 362736 229968
rect 364248 229916 364300 229968
rect 407028 229916 407080 229968
rect 409328 229916 409380 229968
rect 411996 229984 412048 230036
rect 539600 229984 539652 230036
rect 42156 229848 42208 229900
rect 43076 229848 43128 229900
rect 91744 229848 91796 229900
rect 206192 229848 206244 229900
rect 212448 229848 212500 229900
rect 260380 229848 260432 229900
rect 263508 229848 263560 229900
rect 281724 229848 281776 229900
rect 284116 229848 284168 229900
rect 290280 229848 290332 229900
rect 304908 229848 304960 229900
rect 311624 229848 311676 229900
rect 316684 229848 316736 229900
rect 346492 229848 346544 229900
rect 352012 229848 352064 229900
rect 398104 229848 398156 229900
rect 399760 229848 399812 229900
rect 407856 229848 407908 229900
rect 410432 229848 410484 229900
rect 547144 229916 547196 229968
rect 82820 229780 82872 229832
rect 203340 229780 203392 229832
rect 203524 229780 203576 229832
rect 204720 229780 204772 229832
rect 206744 229780 206796 229832
rect 257528 229780 257580 229832
rect 259368 229780 259420 229832
rect 280344 229780 280396 229832
rect 281356 229780 281408 229832
rect 289912 229780 289964 229832
rect 298836 229780 298888 229832
rect 302516 229780 302568 229832
rect 303528 229780 303580 229832
rect 312544 229780 312596 229832
rect 318064 229780 318116 229832
rect 350908 229780 350960 229832
rect 362316 229780 362368 229832
rect 364156 229780 364208 229832
rect 364248 229780 364300 229832
rect 407396 229780 407448 229832
rect 73804 229712 73856 229764
rect 200488 229712 200540 229764
rect 200672 229712 200724 229764
rect 254676 229712 254728 229764
rect 255228 229712 255280 229764
rect 278504 229712 278556 229764
rect 278688 229712 278740 229764
rect 288532 229712 288584 229764
rect 302056 229712 302108 229764
rect 311164 229712 311216 229764
rect 326344 229712 326396 229764
rect 334716 229712 334768 229764
rect 344836 229712 344888 229764
rect 406384 229712 406436 229764
rect 406660 229712 406712 229764
rect 409052 229780 409104 229832
rect 411076 229780 411128 229832
rect 551284 229848 551336 229900
rect 563704 229780 563756 229832
rect 411168 229712 411220 229764
rect 411536 229712 411588 229764
rect 570604 229712 570656 229764
rect 140044 229644 140096 229696
rect 205824 229644 205876 229696
rect 227536 229644 227588 229696
rect 151820 229576 151872 229628
rect 218980 229576 219032 229628
rect 248328 229576 248380 229628
rect 149704 229508 149756 229560
rect 216128 229508 216180 229560
rect 244924 229508 244976 229560
rect 254308 229508 254360 229560
rect 146392 229440 146444 229492
rect 209044 229440 209096 229492
rect 259920 229644 259972 229696
rect 266084 229644 266136 229696
rect 268384 229644 268436 229696
rect 277216 229644 277268 229696
rect 280068 229644 280120 229696
rect 288900 229644 288952 229696
rect 323124 229644 323176 229696
rect 340144 229644 340196 229696
rect 340880 229644 340932 229696
rect 380256 229644 380308 229696
rect 400772 229644 400824 229696
rect 453304 229644 453356 229696
rect 267096 229508 267148 229560
rect 275652 229576 275704 229628
rect 277308 229576 277360 229628
rect 277492 229576 277544 229628
rect 277676 229576 277728 229628
rect 285680 229576 285732 229628
rect 313464 229576 313516 229628
rect 314568 229576 314620 229628
rect 331680 229576 331732 229628
rect 332416 229576 332468 229628
rect 270132 229508 270184 229560
rect 271420 229508 271472 229560
rect 272984 229508 273036 229560
rect 281080 229508 281132 229560
rect 300676 229508 300728 229560
rect 305552 229508 305604 229560
rect 327356 229508 327408 229560
rect 341524 229576 341576 229628
rect 350540 229576 350592 229628
rect 387800 229576 387852 229628
rect 398104 229576 398156 229628
rect 404360 229576 404412 229628
rect 407856 229576 407908 229628
rect 449164 229576 449216 229628
rect 332692 229508 332744 229560
rect 333796 229508 333848 229560
rect 338028 229508 338080 229560
rect 352564 229508 352616 229560
rect 354864 229508 354916 229560
rect 364248 229508 364300 229560
rect 366548 229508 366600 229560
rect 409880 229508 409932 229560
rect 411904 229508 411956 229560
rect 422300 229508 422352 229560
rect 273904 229440 273956 229492
rect 282828 229440 282880 229492
rect 339500 229440 339552 229492
rect 353944 229440 353996 229492
rect 355508 229440 355560 229492
rect 379520 229440 379572 229492
rect 382096 229440 382148 229492
rect 393412 229440 393464 229492
rect 401508 229440 401560 229492
rect 405004 229440 405056 229492
rect 407764 229440 407816 229492
rect 438952 229440 439004 229492
rect 186964 229372 187016 229424
rect 248972 229372 249024 229424
rect 275376 229372 275428 229424
rect 284208 229372 284260 229424
rect 298468 229372 298520 229424
rect 301136 229372 301188 229424
rect 310612 229372 310664 229424
rect 314476 229372 314528 229424
rect 334532 229372 334584 229424
rect 342904 229372 342956 229424
rect 361212 229372 361264 229424
rect 382464 229372 382516 229424
rect 392216 229372 392268 229424
rect 431960 229372 432012 229424
rect 162860 229304 162912 229356
rect 223304 229304 223356 229356
rect 277492 229304 277544 229356
rect 286692 229304 286744 229356
rect 296720 229304 296772 229356
rect 300124 229304 300176 229356
rect 315212 229304 315264 229356
rect 180800 229236 180852 229288
rect 238944 229236 238996 229288
rect 271236 229236 271288 229288
rect 279976 229236 280028 229288
rect 281448 229236 281500 229288
rect 288164 229236 288216 229288
rect 296352 229236 296404 229288
rect 298468 229236 298520 229288
rect 313096 229236 313148 229288
rect 318064 229236 318116 229288
rect 342352 229304 342404 229356
rect 343272 229304 343324 229356
rect 363420 229304 363472 229356
rect 364156 229304 364208 229356
rect 371976 229304 372028 229356
rect 398104 229304 398156 229356
rect 407212 229304 407264 229356
rect 411996 229304 412048 229356
rect 343824 229236 343876 229288
rect 357716 229236 357768 229288
rect 376116 229236 376168 229288
rect 379704 229236 379756 229288
rect 255964 229168 256016 229220
rect 260012 229168 260064 229220
rect 282828 229168 282880 229220
rect 289268 229168 289320 229220
rect 295248 229168 295300 229220
rect 296904 229168 296956 229220
rect 297456 229168 297508 229220
rect 299480 229168 299532 229220
rect 324872 229168 324924 229220
rect 325516 229168 325568 229220
rect 328460 229168 328512 229220
rect 329564 229168 329616 229220
rect 369400 229168 369452 229220
rect 382096 229168 382148 229220
rect 382280 229168 382332 229220
rect 383476 229168 383528 229220
rect 384396 229236 384448 229288
rect 411260 229236 411312 229288
rect 386604 229168 386656 229220
rect 386880 229168 386932 229220
rect 388444 229168 388496 229220
rect 390100 229168 390152 229220
rect 395344 229168 395396 229220
rect 395436 229168 395488 229220
rect 407304 229168 407356 229220
rect 407396 229168 407448 229220
rect 407764 229168 407816 229220
rect 410064 229168 410116 229220
rect 416228 229168 416280 229220
rect 62120 229100 62172 229152
rect 65156 229100 65208 229152
rect 257344 229100 257396 229152
rect 258908 229100 258960 229152
rect 284208 229100 284260 229152
rect 289544 229100 289596 229152
rect 292580 229100 292632 229152
rect 293868 229100 293920 229152
rect 298100 229100 298152 229152
rect 299388 229100 299440 229152
rect 299572 229100 299624 229152
rect 300492 229100 300544 229152
rect 323492 229100 323544 229152
rect 324228 229100 324280 229152
rect 324504 229100 324556 229152
rect 325332 229100 325384 229152
rect 328828 229100 328880 229152
rect 329656 229100 329708 229152
rect 329840 229100 329892 229152
rect 331036 229100 331088 229152
rect 381176 229100 381228 229152
rect 382188 229100 382240 229152
rect 382648 229100 382700 229152
rect 383384 229100 383436 229152
rect 383660 229100 383712 229152
rect 384948 229100 385000 229152
rect 385500 229100 385552 229152
rect 386328 229100 386380 229152
rect 386512 229100 386564 229152
rect 387708 229100 387760 229152
rect 405096 229100 405148 229152
rect 409972 229100 410024 229152
rect 410892 229100 410944 229152
rect 421012 229100 421064 229152
rect 120816 229032 120868 229084
rect 220820 229032 220872 229084
rect 365168 229032 365220 229084
rect 460940 229032 460992 229084
rect 117228 228964 117280 229016
rect 219348 228964 219400 229016
rect 332048 228964 332100 229016
rect 370228 228964 370280 229016
rect 373356 228964 373408 229016
rect 480260 228964 480312 229016
rect 114192 228896 114244 228948
rect 217968 228896 218020 228948
rect 224040 228896 224092 228948
rect 234712 228896 234764 228948
rect 329196 228896 329248 228948
rect 371332 228896 371384 228948
rect 375104 228896 375156 228948
rect 483480 228896 483532 228948
rect 110696 228828 110748 228880
rect 216496 228828 216548 228880
rect 227720 228828 227772 228880
rect 240416 228828 240468 228880
rect 327724 228828 327776 228880
rect 372712 228828 372764 228880
rect 376576 228828 376628 228880
rect 487712 228828 487764 228880
rect 107476 228760 107528 228812
rect 215116 228760 215168 228812
rect 216680 228760 216732 228812
rect 224684 228760 224736 228812
rect 230296 228760 230348 228812
rect 103980 228692 104032 228744
rect 213644 228692 213696 228744
rect 222108 228692 222160 228744
rect 230388 228692 230440 228744
rect 233516 228760 233568 228812
rect 268200 228760 268252 228812
rect 330576 228760 330628 228812
rect 375288 228760 375340 228812
rect 377956 228760 378008 228812
rect 491300 228760 491352 228812
rect 266728 228692 266780 228744
rect 328092 228692 328144 228744
rect 374092 228692 374144 228744
rect 391940 228692 391992 228744
rect 523040 228692 523092 228744
rect 100668 228624 100720 228676
rect 212264 228624 212316 228676
rect 215116 228624 215168 228676
rect 260748 228624 260800 228676
rect 334900 228624 334952 228676
rect 389272 228624 389324 228676
rect 392952 228624 393004 228676
rect 526352 228624 526404 228676
rect 97264 228556 97316 228608
rect 210792 228556 210844 228608
rect 213828 228556 213880 228608
rect 258540 228556 258592 228608
rect 336280 228556 336332 228608
rect 392584 228556 392636 228608
rect 397276 228556 397328 228608
rect 536840 228556 536892 228608
rect 93768 228488 93820 228540
rect 209412 228488 209464 228540
rect 209872 228488 209924 228540
rect 257160 228488 257212 228540
rect 306656 228488 306708 228540
rect 323676 228488 323728 228540
rect 337752 228488 337804 228540
rect 396172 228488 396224 228540
rect 398288 228488 398340 228540
rect 538220 228488 538272 228540
rect 56324 228420 56376 228472
rect 193312 228420 193364 228472
rect 194968 228420 195020 228472
rect 252192 228420 252244 228472
rect 53656 228352 53708 228404
rect 192300 228352 192352 228404
rect 194140 228352 194192 228404
rect 252836 228352 252888 228404
rect 127532 228284 127584 228336
rect 223672 228284 223724 228336
rect 252008 228284 252060 228336
rect 276388 228420 276440 228472
rect 309876 228420 309928 228472
rect 327816 228420 327868 228472
rect 345204 228420 345256 228472
rect 408500 228420 408552 228472
rect 409788 228420 409840 228472
rect 553400 228420 553452 228472
rect 260564 228352 260616 228404
rect 279608 228352 279660 228404
rect 131028 228216 131080 228268
rect 225052 228216 225104 228268
rect 294236 228352 294288 228404
rect 308128 228352 308180 228404
rect 327080 228352 327132 228404
rect 346308 228352 346360 228404
rect 409972 228352 410024 228404
rect 410800 228352 410852 228404
rect 568580 228352 568632 228404
rect 353392 228284 353444 228336
rect 433340 228284 433392 228336
rect 349160 228216 349212 228268
rect 422208 228216 422260 228268
rect 422300 228216 422352 228268
rect 485136 228216 485188 228268
rect 137744 228148 137796 228200
rect 227904 228148 227956 228200
rect 294052 228148 294104 228200
rect 340604 228148 340656 228200
rect 402980 228148 403032 228200
rect 404360 228148 404412 228200
rect 476120 228148 476172 228200
rect 144368 228080 144420 228132
rect 230756 228080 230808 228132
rect 334164 228080 334216 228132
rect 378508 228080 378560 228132
rect 380716 228080 380768 228132
rect 406016 228080 406068 228132
rect 407028 228080 407080 228132
rect 454040 228080 454092 228132
rect 154488 228012 154540 228064
rect 235080 228012 235132 228064
rect 343456 228012 343508 228064
rect 387156 228012 387208 228064
rect 387800 228012 387852 228064
rect 426440 228012 426492 228064
rect 161296 227944 161348 227996
rect 237932 227944 237984 227996
rect 386420 227944 386472 227996
rect 419540 227944 419592 227996
rect 171048 227876 171100 227928
rect 242164 227876 242216 227928
rect 378232 227876 378284 227928
rect 399392 227876 399444 227928
rect 403072 227876 403124 227928
rect 429660 227876 429712 227928
rect 375472 227808 375524 227860
rect 380992 227808 381044 227860
rect 77944 227740 77996 227792
rect 82820 227740 82872 227792
rect 84660 227740 84712 227792
rect 91744 227740 91796 227792
rect 377312 227740 377364 227792
rect 380348 227740 380400 227792
rect 160376 227672 160428 227724
rect 238576 227672 238628 227724
rect 364432 227672 364484 227724
rect 457352 227672 457404 227724
rect 157064 227604 157116 227656
rect 237196 227604 237248 227656
rect 358728 227604 358780 227656
rect 444380 227604 444432 227656
rect 449164 227604 449216 227656
rect 543004 227604 543056 227656
rect 153660 227536 153712 227588
rect 235724 227536 235776 227588
rect 365904 227536 365956 227588
rect 461216 227536 461268 227588
rect 461584 227536 461636 227588
rect 552664 227536 552716 227588
rect 108212 227468 108264 227520
rect 149704 227468 149756 227520
rect 150348 227468 150400 227520
rect 234344 227468 234396 227520
rect 367284 227468 367336 227520
rect 464160 227468 464212 227520
rect 147588 227400 147640 227452
rect 232228 227400 232280 227452
rect 309508 227400 309560 227452
rect 330392 227400 330444 227452
rect 368756 227400 368808 227452
rect 467840 227400 467892 227452
rect 469220 227400 469272 227452
rect 555424 227400 555476 227452
rect 91376 227332 91428 227384
rect 146392 227332 146444 227384
rect 146944 227332 146996 227384
rect 232872 227332 232924 227384
rect 315580 227332 315632 227384
rect 341340 227332 341392 227384
rect 370136 227332 370188 227384
rect 470876 227332 470928 227384
rect 143448 227264 143500 227316
rect 231492 227264 231544 227316
rect 312728 227264 312780 227316
rect 333980 227264 334032 227316
rect 335176 227264 335228 227316
rect 363144 227264 363196 227316
rect 371608 227264 371660 227316
rect 474188 227264 474240 227316
rect 141056 227196 141108 227248
rect 229376 227196 229428 227248
rect 232780 227196 232832 227248
rect 247500 227196 247552 227248
rect 318432 227196 318484 227248
rect 348056 227196 348108 227248
rect 372988 227196 373040 227248
rect 477592 227196 477644 227248
rect 478144 227196 478196 227248
rect 500224 227196 500276 227248
rect 82728 227128 82780 227180
rect 140044 227128 140096 227180
rect 140136 227128 140188 227180
rect 230020 227128 230072 227180
rect 237380 227128 237432 227180
rect 256056 227128 256108 227180
rect 258816 227128 258868 227180
rect 279240 227128 279292 227180
rect 321284 227128 321336 227180
rect 354772 227128 354824 227180
rect 374460 227128 374512 227180
rect 480904 227128 480956 227180
rect 134248 227060 134300 227112
rect 226524 227060 226576 227112
rect 234712 227060 234764 227112
rect 253204 227060 253256 227112
rect 255136 227060 255188 227112
rect 277860 227060 277912 227112
rect 329472 227060 329524 227112
rect 365260 227060 365312 227112
rect 374828 227060 374880 227112
rect 483112 227060 483164 227112
rect 124128 226992 124180 227044
rect 222200 226992 222252 227044
rect 237012 226992 237064 227044
rect 269580 226992 269632 227044
rect 305276 226992 305328 227044
rect 320272 226992 320324 227044
rect 325608 226992 325660 227044
rect 360292 226992 360344 227044
rect 409696 226992 409748 227044
rect 565912 226992 565964 227044
rect 125048 226924 125100 226976
rect 162860 226924 162912 226976
rect 163688 226924 163740 226976
rect 239772 226924 239824 226976
rect 293960 226924 294012 226976
rect 294604 226924 294656 226976
rect 363052 226924 363104 226976
rect 454132 226924 454184 226976
rect 166908 226856 166960 226908
rect 241428 226856 241480 226908
rect 361580 226856 361632 226908
rect 450636 226856 450688 226908
rect 164608 226788 164660 226840
rect 239312 226788 239364 226840
rect 360200 226788 360252 226840
rect 447324 226788 447376 226840
rect 173808 226720 173860 226772
rect 244280 226720 244332 226772
rect 357348 226720 357400 226772
rect 440608 226720 440660 226772
rect 42156 226652 42208 226704
rect 44364 226652 44416 226704
rect 174636 226652 174688 226704
rect 243636 226652 243688 226704
rect 355876 226652 355928 226704
rect 437480 226652 437532 226704
rect 177212 226584 177264 226636
rect 245752 226584 245804 226636
rect 354496 226584 354548 226636
rect 433800 226584 433852 226636
rect 190276 226516 190328 226568
rect 251456 226516 251508 226568
rect 351644 226516 351696 226568
rect 427084 226516 427136 226568
rect 124864 226312 124916 226364
rect 130384 226312 130436 226364
rect 116584 226244 116636 226296
rect 220084 226244 220136 226296
rect 364064 226244 364116 226296
rect 455696 226244 455748 226296
rect 456156 226244 456208 226296
rect 548156 226244 548208 226296
rect 42156 226176 42208 226228
rect 42984 226176 43036 226228
rect 112996 226176 113048 226228
rect 218612 226176 218664 226228
rect 223120 226176 223172 226228
rect 233240 226176 233292 226228
rect 365536 226176 365588 226228
rect 459560 226176 459612 226228
rect 109868 226108 109920 226160
rect 217232 226108 217284 226160
rect 218060 226108 218112 226160
rect 227260 226108 227312 226160
rect 227352 226108 227404 226160
rect 237564 226108 237616 226160
rect 366916 226108 366968 226160
rect 462412 226108 462464 226160
rect 106556 226040 106608 226092
rect 215760 226040 215812 226092
rect 224960 226040 225012 226092
rect 251824 226040 251876 226092
rect 253848 226040 253900 226092
rect 276480 226040 276532 226092
rect 335912 226040 335964 226092
rect 367652 226040 367704 226092
rect 368388 226040 368440 226092
rect 465080 226040 465132 226092
rect 103244 225972 103296 226024
rect 214380 225972 214432 226024
rect 220636 225972 220688 226024
rect 264244 225972 264296 226024
rect 322756 225972 322808 226024
rect 358176 225972 358228 226024
rect 369768 225972 369820 226024
rect 469220 225972 469272 226024
rect 99840 225904 99892 225956
rect 212908 225904 212960 225956
rect 215300 225904 215352 225956
rect 261392 225904 261444 225956
rect 326988 225904 327040 225956
rect 362960 225904 363012 225956
rect 371240 225904 371292 225956
rect 471980 225904 472032 225956
rect 96528 225836 96580 225888
rect 211528 225836 211580 225888
rect 211712 225836 211764 225888
rect 259000 225836 259052 225888
rect 356980 225836 357032 225888
rect 438860 225836 438912 225888
rect 438952 225836 439004 225888
rect 540428 225836 540480 225888
rect 86316 225768 86368 225820
rect 207204 225768 207256 225820
rect 208308 225768 208360 225820
rect 257896 225768 257948 225820
rect 324136 225768 324188 225820
rect 361580 225768 361632 225820
rect 372620 225768 372672 225820
rect 476212 225768 476264 225820
rect 76288 225700 76340 225752
rect 202972 225700 203024 225752
rect 206836 225700 206888 225752
rect 256792 225700 256844 225752
rect 303804 225700 303856 225752
rect 317420 225700 317472 225752
rect 343088 225700 343140 225752
rect 407120 225700 407172 225752
rect 407304 225700 407356 225752
rect 531412 225700 531464 225752
rect 539600 225700 539652 225752
rect 560852 225700 560904 225752
rect 56048 225632 56100 225684
rect 194416 225632 194468 225684
rect 199016 225632 199068 225684
rect 200672 225632 200724 225684
rect 203248 225632 203300 225684
rect 255320 225632 255372 225684
rect 263416 225632 263468 225684
rect 280988 225632 281040 225684
rect 302424 225632 302476 225684
rect 313556 225632 313608 225684
rect 314476 225632 314528 225684
rect 331220 225632 331272 225684
rect 341616 225632 341668 225684
rect 403532 225632 403584 225684
rect 403624 225632 403676 225684
rect 552020 225632 552072 225684
rect 52736 225564 52788 225616
rect 192668 225564 192720 225616
rect 201408 225564 201460 225616
rect 255044 225564 255096 225616
rect 257068 225564 257120 225616
rect 278136 225564 278188 225616
rect 310980 225564 311032 225616
rect 334072 225564 334124 225616
rect 344468 225564 344520 225616
rect 410248 225564 410300 225616
rect 410984 225564 411036 225616
rect 559196 225564 559248 225616
rect 119896 225496 119948 225548
rect 221188 225496 221240 225548
rect 362868 225496 362920 225548
rect 452660 225496 452712 225548
rect 123392 225428 123444 225480
rect 222936 225428 222988 225480
rect 359832 225428 359884 225480
rect 445760 225428 445812 225480
rect 126796 225360 126848 225412
rect 224316 225360 224368 225412
rect 358360 225360 358412 225412
rect 441620 225360 441672 225412
rect 130108 225292 130160 225344
rect 225788 225292 225840 225344
rect 348792 225292 348844 225344
rect 420368 225292 420420 225344
rect 133512 225224 133564 225276
rect 227168 225224 227220 225276
rect 345940 225224 345992 225276
rect 414020 225224 414072 225276
rect 170496 225156 170548 225208
rect 242900 225156 242952 225208
rect 339040 225156 339092 225208
rect 382280 225156 382332 225208
rect 382464 225156 382516 225208
rect 448980 225156 449032 225208
rect 180616 225088 180668 225140
rect 247132 225088 247184 225140
rect 340236 225088 340288 225140
rect 385500 225088 385552 225140
rect 386604 225088 386656 225140
rect 434720 225088 434772 225140
rect 192852 224952 192904 225004
rect 197636 224952 197688 225004
rect 162768 224884 162820 224936
rect 238208 224884 238260 224936
rect 368020 224884 368072 224936
rect 468300 224884 468352 224936
rect 159548 224816 159600 224868
rect 236828 224816 236880 224868
rect 377404 224816 377456 224868
rect 479248 224816 479300 224868
rect 155776 224748 155828 224800
rect 235356 224748 235408 224800
rect 370872 224748 370924 224800
rect 475016 224748 475068 224800
rect 114928 224680 114980 224732
rect 151820 224680 151872 224732
rect 152924 224680 152976 224732
rect 233976 224680 234028 224732
rect 372252 224680 372304 224732
rect 478972 224680 479024 224732
rect 149428 224612 149480 224664
rect 232320 224612 232372 224664
rect 373724 224612 373776 224664
rect 481824 224612 481876 224664
rect 146116 224544 146168 224596
rect 231124 224544 231176 224596
rect 335544 224544 335596 224596
rect 377312 224544 377364 224596
rect 388720 224544 388772 224596
rect 516232 224544 516284 224596
rect 142712 224476 142764 224528
rect 229652 224476 229704 224528
rect 332324 224476 332376 224528
rect 372620 224476 372672 224528
rect 389732 224476 389784 224528
rect 518900 224476 518952 224528
rect 139216 224408 139268 224460
rect 228272 224408 228324 224460
rect 234620 224408 234672 224460
rect 250352 224408 250404 224460
rect 268936 224408 268988 224460
rect 283564 224408 283616 224460
rect 333704 224408 333756 224460
rect 378048 224408 378100 224460
rect 400036 224408 400088 224460
rect 543188 224408 543240 224460
rect 135996 224340 136048 224392
rect 226800 224340 226852 224392
rect 246856 224340 246908 224392
rect 273628 224340 273680 224392
rect 307760 224340 307812 224392
rect 325700 224340 325752 224392
rect 339868 224340 339920 224392
rect 386420 224340 386472 224392
rect 402244 224340 402296 224392
rect 548524 224340 548576 224392
rect 101496 224272 101548 224324
rect 136364 224272 136416 224324
rect 136548 224272 136600 224324
rect 228640 224272 228692 224324
rect 232412 224272 232464 224324
rect 243268 224272 243320 224324
rect 243636 224272 243688 224324
rect 272248 224272 272300 224324
rect 309232 224272 309284 224324
rect 328736 224272 328788 224324
rect 341432 224272 341484 224324
rect 401876 224272 401928 224324
rect 405464 224272 405516 224324
rect 556160 224272 556212 224324
rect 88156 224204 88208 224256
rect 207572 224204 207624 224256
rect 239956 224204 240008 224256
rect 271052 224204 271104 224256
rect 292580 224204 292632 224256
rect 293500 224204 293552 224256
rect 311348 224204 311400 224256
rect 331312 224204 331364 224256
rect 344100 224204 344152 224256
rect 408592 224204 408644 224256
rect 408684 224204 408736 224256
rect 563612 224204 563664 224256
rect 166264 224136 166316 224188
rect 239680 224136 239732 224188
rect 342720 224136 342772 224188
rect 405832 224136 405884 224188
rect 411260 224136 411312 224188
rect 506480 224136 506532 224188
rect 169576 224068 169628 224120
rect 241060 224068 241112 224120
rect 338396 224068 338448 224120
rect 380716 224068 380768 224120
rect 393412 224068 393464 224120
rect 472072 224068 472124 224120
rect 172980 224000 173032 224052
rect 242532 224000 242584 224052
rect 349804 224000 349856 224052
rect 422392 224000 422444 224052
rect 176476 223932 176528 223984
rect 243912 223932 243964 223984
rect 347320 223932 347372 223984
rect 417056 223932 417108 223984
rect 179696 223864 179748 223916
rect 245384 223864 245436 223916
rect 348424 223864 348476 223916
rect 418712 223864 418764 223916
rect 183192 223796 183244 223848
rect 246764 223796 246816 223848
rect 346952 223796 347004 223848
rect 415492 223796 415544 223848
rect 186228 223728 186280 223780
rect 248236 223728 248288 223780
rect 354864 223728 354916 223780
rect 411996 223728 412048 223780
rect 337292 223660 337344 223712
rect 378784 223660 378836 223712
rect 409880 223660 409932 223712
rect 465172 223660 465224 223712
rect 56600 223524 56652 223576
rect 62028 223592 62080 223644
rect 125876 223524 125928 223576
rect 222568 223524 222620 223576
rect 359464 223524 359516 223576
rect 448612 223524 448664 223576
rect 115756 223456 115808 223508
rect 108856 223388 108908 223440
rect 105728 223320 105780 223372
rect 209596 223320 209648 223372
rect 101956 223252 102008 223304
rect 95608 223184 95660 223236
rect 209688 223184 209740 223236
rect 213920 223456 213972 223508
rect 221832 223456 221884 223508
rect 361120 223456 361172 223508
rect 451464 223456 451516 223508
rect 352288 223388 352340 223440
rect 431316 223388 431368 223440
rect 431960 223388 432012 223440
rect 525064 223388 525116 223440
rect 218244 223320 218296 223372
rect 389088 223320 389140 223372
rect 395712 223320 395764 223372
rect 215392 223252 215444 223304
rect 212540 223184 212592 223236
rect 319260 223184 319312 223236
rect 350632 223184 350684 223236
rect 391572 223184 391624 223236
rect 82176 223116 82228 223168
rect 203984 223116 204036 223168
rect 209596 223116 209648 223168
rect 214012 223116 214064 223168
rect 250352 223116 250404 223168
rect 275100 223116 275152 223168
rect 311624 223116 311676 223168
rect 318892 223116 318944 223168
rect 330944 223116 330996 223168
rect 367008 223116 367060 223168
rect 385868 223116 385920 223168
rect 387800 223116 387852 223168
rect 523132 223320 523184 223372
rect 398288 223252 398340 223304
rect 530584 223252 530636 223304
rect 395988 223184 396040 223236
rect 533068 223184 533120 223236
rect 397920 223116 397972 223168
rect 538312 223116 538364 223168
rect 75368 223048 75420 223100
rect 201132 223048 201184 223100
rect 204904 223048 204956 223100
rect 256424 223048 256476 223100
rect 314200 223048 314252 223100
rect 338120 223048 338172 223100
rect 348148 223048 348200 223100
rect 421196 223048 421248 223100
rect 421288 223048 421340 223100
rect 569316 223048 569368 223100
rect 69020 222980 69072 223032
rect 68744 222912 68796 222964
rect 193956 222912 194008 222964
rect 198188 222980 198240 223032
rect 253572 222980 253624 223032
rect 306380 222980 306432 223032
rect 321928 222980 321980 223032
rect 326620 222980 326672 223032
rect 371240 222980 371292 223032
rect 379796 222980 379848 223032
rect 389180 222980 389232 223032
rect 394792 222980 394844 223032
rect 398288 222980 398340 223032
rect 404636 222980 404688 223032
rect 553676 222980 553728 223032
rect 198372 222912 198424 222964
rect 199936 222912 199988 222964
rect 253940 222912 253992 222964
rect 265532 222912 265584 222964
rect 282092 222912 282144 222964
rect 317052 222912 317104 222964
rect 345020 222912 345072 222964
rect 346676 222912 346728 222964
rect 415308 222912 415360 222964
rect 416228 222912 416280 222964
rect 567200 222912 567252 222964
rect 65340 222844 65392 222896
rect 196900 222844 196952 222896
rect 200764 222844 200816 222896
rect 255688 222844 255740 222896
rect 262128 222844 262180 222896
rect 280712 222844 280764 222896
rect 308496 222844 308548 222896
rect 324504 222844 324556 222896
rect 337660 222844 337712 222896
rect 390652 222844 390704 222896
rect 407580 222844 407632 222896
rect 560944 222844 560996 222896
rect 132316 222776 132368 222828
rect 225420 222776 225472 222828
rect 357992 222776 358044 222828
rect 444748 222776 444800 222828
rect 177856 222708 177908 222760
rect 245016 222708 245068 222760
rect 356612 222708 356664 222760
rect 441712 222708 441764 222760
rect 162032 222640 162084 222692
rect 180800 222640 180852 222692
rect 181352 222640 181404 222692
rect 246488 222640 246540 222692
rect 355140 222640 355192 222692
rect 438032 222640 438084 222692
rect 187332 222572 187384 222624
rect 249984 222572 250036 222624
rect 353760 222572 353812 222624
rect 434812 222572 434864 222624
rect 184756 222504 184808 222556
rect 247868 222504 247920 222556
rect 352656 222504 352708 222556
rect 429292 222504 429344 222556
rect 665824 222504 665876 222556
rect 675944 222504 675996 222556
rect 188160 222436 188212 222488
rect 249340 222436 249392 222488
rect 351184 222436 351236 222488
rect 427912 222436 427964 222488
rect 428648 222436 428700 222488
rect 488540 222436 488592 222488
rect 191564 222368 191616 222420
rect 250720 222368 250772 222420
rect 349436 222368 349488 222420
rect 425060 222368 425112 222420
rect 664444 222368 664496 222420
rect 676036 222368 676088 222420
rect 196532 222300 196584 222352
rect 252284 222300 252336 222352
rect 193956 222232 194008 222284
rect 198280 222232 198332 222284
rect 673920 222232 673972 222284
rect 676036 222232 676088 222284
rect 660396 222164 660448 222216
rect 675852 222164 675904 222216
rect 122472 222096 122524 222148
rect 221004 222096 221056 222148
rect 228456 222096 228508 222148
rect 266452 222096 266504 222148
rect 311164 222096 311216 222148
rect 311992 222096 312044 222148
rect 312544 222096 312596 222148
rect 315304 222096 315356 222148
rect 318708 222096 318760 222148
rect 349160 222096 349212 222148
rect 362684 222096 362736 222148
rect 453212 222096 453264 222148
rect 453304 222096 453356 222148
rect 545212 222096 545264 222148
rect 574744 222096 574796 222148
rect 575480 222096 575532 222148
rect 119160 222028 119212 222080
rect 219624 222028 219676 222080
rect 226800 222028 226852 222080
rect 265256 222028 265308 222080
rect 321376 222028 321428 222080
rect 356060 222028 356112 222080
rect 364156 222028 364208 222080
rect 456800 222028 456852 222080
rect 100760 221960 100812 222012
rect 204352 221960 204404 222012
rect 223488 221960 223540 222012
rect 263692 221960 263744 222012
rect 321192 221960 321244 222012
rect 357532 221960 357584 222012
rect 363972 221960 364024 222012
rect 458364 221960 458416 222012
rect 112444 221892 112496 221944
rect 216864 221892 216916 221944
rect 224868 221892 224920 221944
rect 265164 221892 265216 221944
rect 322296 221892 322348 221944
rect 359096 221892 359148 221944
rect 365076 221892 365128 221944
rect 460020 221892 460072 221944
rect 88892 221824 88944 221876
rect 85488 221756 85540 221808
rect 205180 221756 205232 221808
rect 83832 221688 83884 221740
rect 204812 221688 204864 221740
rect 205548 221824 205600 221876
rect 206744 221824 206796 221876
rect 220084 221824 220136 221876
rect 262312 221824 262364 221876
rect 322664 221824 322716 221876
rect 360752 221824 360804 221876
rect 366456 221824 366508 221876
rect 463700 221824 463752 221876
rect 674656 221824 674708 221876
rect 676036 221824 676088 221876
rect 206928 221756 206980 221808
rect 217324 221756 217376 221808
rect 218428 221756 218480 221808
rect 261852 221756 261904 221808
rect 324228 221756 324280 221808
rect 362408 221756 362460 221808
rect 367928 221756 367980 221808
rect 466736 221756 466788 221808
rect 467104 221756 467156 221808
rect 557816 221756 557868 221808
rect 206652 221688 206704 221740
rect 208216 221688 208268 221740
rect 220176 221688 220228 221740
rect 221740 221688 221792 221740
rect 263784 221688 263836 221740
rect 325516 221688 325568 221740
rect 365812 221688 365864 221740
rect 369308 221688 369360 221740
rect 470140 221688 470192 221740
rect 80428 221620 80480 221672
rect 203432 221620 203484 221672
rect 204168 221620 204220 221672
rect 214472 221620 214524 221672
rect 216588 221620 216640 221672
rect 261024 221620 261076 221672
rect 326528 221620 326580 221672
rect 369124 221620 369176 221672
rect 370780 221620 370832 221672
rect 473544 221620 473596 221672
rect 77024 221552 77076 221604
rect 201960 221552 202012 221604
rect 202420 221552 202472 221604
rect 210148 221552 210200 221604
rect 213368 221552 213420 221604
rect 259644 221552 259696 221604
rect 325424 221552 325476 221604
rect 367468 221552 367520 221604
rect 400128 221552 400180 221604
rect 541072 221552 541124 221604
rect 547144 221552 547196 221604
rect 561772 221552 561824 221604
rect 63408 221484 63460 221536
rect 196256 221484 196308 221536
rect 197268 221484 197320 221536
rect 244924 221484 244976 221536
rect 245292 221484 245344 221536
rect 273444 221484 273496 221536
rect 275560 221484 275612 221536
rect 286140 221484 286192 221536
rect 319444 221484 319496 221536
rect 352380 221484 352432 221536
rect 352564 221484 352616 221536
rect 397736 221484 397788 221536
rect 404176 221484 404228 221536
rect 550824 221484 550876 221536
rect 551284 221484 551336 221536
rect 565452 221484 565504 221536
rect 674012 221484 674064 221536
rect 676036 221484 676088 221536
rect 28724 221416 28776 221468
rect 43720 221416 43772 221468
rect 60280 221416 60332 221468
rect 194876 221416 194928 221468
rect 209688 221416 209740 221468
rect 258264 221416 258316 221468
rect 272248 221416 272300 221468
rect 284668 221416 284720 221468
rect 301228 221416 301280 221468
rect 310520 221416 310572 221468
rect 319812 221416 319864 221468
rect 354036 221416 354088 221468
rect 129280 221348 129332 221400
rect 223764 221348 223816 221400
rect 231676 221348 231728 221400
rect 267832 221348 267884 221400
rect 317328 221348 317380 221400
rect 345572 221348 345624 221400
rect 151084 221280 151136 221332
rect 233424 221280 233476 221332
rect 235264 221280 235316 221332
rect 269212 221280 269264 221332
rect 315948 221280 316000 221332
rect 342260 221280 342312 221332
rect 353944 221280 353996 221332
rect 401140 221416 401192 221468
rect 406752 221416 406804 221468
rect 558460 221416 558512 221468
rect 361304 221348 361356 221400
rect 449900 221348 449952 221400
rect 360108 221280 360160 221332
rect 446588 221280 446640 221332
rect 157800 221212 157852 221264
rect 236184 221212 236236 221264
rect 238576 221212 238628 221264
rect 270684 221212 270736 221264
rect 314568 221212 314620 221264
rect 338856 221212 338908 221264
rect 357072 221212 357124 221264
rect 439780 221212 439832 221264
rect 443644 221212 443696 221264
rect 491944 221212 491996 221264
rect 167920 221144 167972 221196
rect 240508 221144 240560 221196
rect 241980 221144 242032 221196
rect 271972 221144 272024 221196
rect 313188 221144 313240 221196
rect 335544 221144 335596 221196
rect 351552 221144 351604 221196
rect 425520 221144 425572 221196
rect 183928 221076 183980 221128
rect 248604 221076 248656 221128
rect 248696 221076 248748 221128
rect 274824 221076 274876 221128
rect 376116 221076 376168 221128
rect 443184 221076 443236 221128
rect 189816 221008 189868 221060
rect 249432 221008 249484 221060
rect 343272 221008 343324 221060
rect 407856 221008 407908 221060
rect 407948 221008 408000 221060
rect 436468 221008 436520 221060
rect 192944 220940 192996 220992
rect 250812 220940 250864 220992
rect 385684 220940 385736 220992
rect 411260 220940 411312 220992
rect 195152 220872 195204 220924
rect 211620 220872 211672 220924
rect 380256 220872 380308 220924
rect 404452 220872 404504 220924
rect 61108 220736 61160 220788
rect 64144 220736 64196 220788
rect 71228 220736 71280 220788
rect 73804 220736 73856 220788
rect 131764 220736 131816 220788
rect 132408 220736 132460 220788
rect 138480 220736 138532 220788
rect 139308 220736 139360 220788
rect 141884 220736 141936 220788
rect 222108 220736 222160 220788
rect 232688 220736 232740 220788
rect 233148 220736 233200 220788
rect 239404 220736 239456 220788
rect 240048 220736 240100 220788
rect 241152 220736 241204 220788
rect 269672 220736 269724 220788
rect 270316 220736 270368 220788
rect 305552 220804 305604 220856
rect 308588 220804 308640 220856
rect 563704 220804 563756 220856
rect 567936 220804 567988 220856
rect 271328 220736 271380 220788
rect 273904 220736 273956 220788
rect 274548 220736 274600 220788
rect 278136 220736 278188 220788
rect 278688 220736 278740 220788
rect 282368 220736 282420 220788
rect 282828 220736 282880 220788
rect 283196 220736 283248 220788
rect 284116 220736 284168 220788
rect 286508 220736 286560 220788
rect 286968 220736 287020 220788
rect 287336 220736 287388 220788
rect 290648 220736 290700 220788
rect 290740 220736 290792 220788
rect 292212 220736 292264 220788
rect 292488 220736 292540 220788
rect 293224 220736 293276 220788
rect 294972 220736 295024 220788
rect 295524 220736 295576 220788
rect 298008 220736 298060 220788
rect 302240 220736 302292 220788
rect 325332 220736 325384 220788
rect 363236 220736 363288 220788
rect 367008 220736 367060 220788
rect 380900 220736 380952 220788
rect 387800 220736 387852 220788
rect 509884 220736 509936 220788
rect 134984 220668 135036 220720
rect 128176 220600 128228 220652
rect 214196 220668 214248 220720
rect 215300 220668 215352 220720
rect 237748 220668 237800 220720
rect 270132 220668 270184 220720
rect 274456 220668 274508 220720
rect 276664 220668 276716 220720
rect 289084 220668 289136 220720
rect 291844 220668 291896 220720
rect 303068 220668 303120 220720
rect 311164 220668 311216 220720
rect 326252 220668 326304 220720
rect 366640 220668 366692 220720
rect 367652 220668 367704 220720
rect 390560 220668 390612 220720
rect 395712 220668 395764 220720
rect 517520 220668 517572 220720
rect 576400 220736 576452 220788
rect 522580 220668 522632 220720
rect 577320 220668 577372 220720
rect 673368 220668 673420 220720
rect 676036 220668 676088 220720
rect 118332 220532 118384 220584
rect 218060 220600 218112 220652
rect 235908 220600 235960 220652
rect 270040 220600 270092 220652
rect 273076 220600 273128 220652
rect 276756 220600 276808 220652
rect 291476 220600 291528 220652
rect 294052 220600 294104 220652
rect 303436 220600 303488 220652
rect 312820 220600 312872 220652
rect 329564 220600 329616 220652
rect 371700 220600 371752 220652
rect 371884 220600 371936 220652
rect 385960 220600 386012 220652
rect 388444 220600 388496 220652
rect 512828 220600 512880 220652
rect 545764 220600 545816 220652
rect 576492 220600 576544 220652
rect 121276 220464 121328 220516
rect 206192 220464 206244 220516
rect 216680 220532 216732 220584
rect 229376 220532 229428 220584
rect 262588 220532 262640 220584
rect 262956 220532 263008 220584
rect 263508 220532 263560 220584
rect 299388 220532 299440 220584
rect 303620 220532 303672 220584
rect 304816 220532 304868 220584
rect 316132 220532 316184 220584
rect 329656 220532 329708 220584
rect 373356 220532 373408 220584
rect 208216 220464 208268 220516
rect 111616 220396 111668 220448
rect 206928 220396 206980 220448
rect 145196 220328 145248 220380
rect 146208 220328 146260 220380
rect 155316 220328 155368 220380
rect 155868 220328 155920 220380
rect 168748 220328 168800 220380
rect 169668 220328 169720 220380
rect 178868 220328 178920 220380
rect 179328 220328 179380 220380
rect 192300 220328 192352 220380
rect 224960 220464 225012 220516
rect 231032 220464 231084 220516
rect 268292 220464 268344 220516
rect 299296 220464 299348 220516
rect 305276 220464 305328 220516
rect 306196 220464 306248 220516
rect 317880 220464 317932 220516
rect 319352 220464 319404 220516
rect 339684 220464 339736 220516
rect 342904 220464 342956 220516
rect 386788 220464 386840 220516
rect 222568 220396 222620 220448
rect 264336 220396 264388 220448
rect 306104 220396 306156 220448
rect 319536 220396 319588 220448
rect 331036 220396 331088 220448
rect 375380 220396 375432 220448
rect 376024 220396 376076 220448
rect 394700 220532 394752 220584
rect 395344 220532 395396 220584
rect 520004 220532 520056 220584
rect 574928 220532 574980 220584
rect 391480 220464 391532 220516
rect 522580 220464 522632 220516
rect 525064 220464 525116 220516
rect 577136 220464 577188 220516
rect 394608 220396 394660 220448
rect 527272 220396 527324 220448
rect 576308 220396 576360 220448
rect 224316 220328 224368 220380
rect 265440 220328 265492 220380
rect 268016 220328 268068 220380
rect 275376 220328 275428 220380
rect 307576 220328 307628 220380
rect 321560 220328 321612 220380
rect 330484 220328 330536 220380
rect 376944 220328 376996 220380
rect 378048 220328 378100 220380
rect 387800 220328 387852 220380
rect 394516 220328 394568 220380
rect 530124 220328 530176 220380
rect 574836 220328 574888 220380
rect 79600 220260 79652 220312
rect 100760 220260 100812 220312
rect 104716 220260 104768 220312
rect 204168 220260 204220 220312
rect 207480 220260 207532 220312
rect 213828 220260 213880 220312
rect 217600 220260 217652 220312
rect 260104 220260 260156 220312
rect 264704 220260 264756 220312
rect 273812 220260 273864 220312
rect 307392 220260 307444 220312
rect 322940 220260 322992 220312
rect 332232 220260 332284 220312
rect 378416 220260 378468 220312
rect 378784 220260 378836 220312
rect 391940 220260 391992 220312
rect 396724 220260 396776 220312
rect 532700 220260 532752 220312
rect 66076 220192 66128 220244
rect 69020 220192 69072 220244
rect 94780 220192 94832 220244
rect 202420 220192 202472 220244
rect 206192 220192 206244 220244
rect 213920 220192 213972 220244
rect 215852 220192 215904 220244
rect 261484 220192 261536 220244
rect 262588 220192 262640 220244
rect 267188 220192 267240 220244
rect 271420 220192 271472 220244
rect 275284 220192 275336 220244
rect 308772 220192 308824 220244
rect 326252 220192 326304 220244
rect 332416 220192 332468 220244
rect 380072 220192 380124 220244
rect 380716 220192 380768 220244
rect 395252 220192 395304 220244
rect 396816 220192 396868 220244
rect 535368 220192 535420 220244
rect 672632 220192 672684 220244
rect 676036 220192 676088 220244
rect 81256 220124 81308 220176
rect 203524 220124 203576 220176
rect 204076 220124 204128 220176
rect 209872 220124 209924 220176
rect 210792 220124 210844 220176
rect 64512 220056 64564 220108
rect 192852 220056 192904 220108
rect 209136 220056 209188 220108
rect 252100 220056 252152 220108
rect 254584 220124 254636 220176
rect 255228 220124 255280 220176
rect 257896 220124 257948 220176
rect 271236 220124 271288 220176
rect 255964 220056 256016 220108
rect 266176 220056 266228 220108
rect 279424 220124 279476 220176
rect 280620 220124 280672 220176
rect 281448 220124 281500 220176
rect 278596 220056 278648 220108
rect 287520 220124 287572 220176
rect 304448 220124 304500 220176
rect 314660 220124 314712 220176
rect 315396 220124 315448 220176
rect 332968 220124 333020 220176
rect 333796 220124 333848 220176
rect 381820 220124 381872 220176
rect 382280 220124 382332 220176
rect 396908 220124 396960 220176
rect 398564 220124 398616 220176
rect 537392 220124 537444 220176
rect 548156 220124 548208 220176
rect 301964 220056 302016 220108
rect 309416 220056 309468 220108
rect 310244 220056 310296 220108
rect 329840 220056 329892 220108
rect 333888 220056 333940 220108
rect 383660 220056 383712 220108
rect 385500 220056 385552 220108
rect 400312 220056 400364 220108
rect 404268 220056 404320 220108
rect 148600 219988 148652 220040
rect 223120 219988 223172 220040
rect 247868 219988 247920 220040
rect 248328 219988 248380 220040
rect 151728 219920 151780 219972
rect 224040 219920 224092 219972
rect 246120 219920 246172 219972
rect 246948 219920 247000 219972
rect 272892 219988 272944 220040
rect 289636 219988 289688 220040
rect 292856 219988 292908 220040
rect 318064 219988 318116 220040
rect 336740 219988 336792 220040
rect 341524 219988 341576 220040
rect 370044 219988 370096 220040
rect 370228 219988 370280 220040
rect 382648 219988 382700 220040
rect 383384 219988 383436 220040
rect 502432 219988 502484 220040
rect 543004 220056 543056 220108
rect 549628 219988 549680 220040
rect 158628 219852 158680 219904
rect 227352 219852 227404 219904
rect 242808 219852 242860 219904
rect 249524 219852 249576 219904
rect 276204 219920 276256 219972
rect 284852 219920 284904 219972
rect 285588 219920 285640 219972
rect 340144 219920 340196 219972
rect 360200 219920 360252 219972
rect 365260 219920 365312 219972
rect 377588 219920 377640 219972
rect 384948 219920 385000 219972
rect 504916 219920 504968 219972
rect 560760 220124 560812 220176
rect 617156 220124 617208 220176
rect 552848 220056 552900 220108
rect 609612 220056 609664 220108
rect 614120 219988 614172 220040
rect 611728 219920 611780 219972
rect 252928 219852 252980 219904
rect 277584 219852 277636 219904
rect 322204 219852 322256 219904
rect 343088 219852 343140 219904
rect 363144 219852 363196 219904
rect 391020 219852 391072 219904
rect 399484 219852 399536 219904
rect 513840 219852 513892 219904
rect 540428 219852 540480 219904
rect 613016 219852 613068 219904
rect 673276 219852 673328 219904
rect 676036 219852 676088 219904
rect 165436 219784 165488 219836
rect 227720 219784 227772 219836
rect 256240 219784 256292 219836
rect 278964 219784 279016 219836
rect 293224 219784 293276 219836
rect 293960 219784 294012 219836
rect 338764 219784 338816 219836
rect 356520 219784 356572 219836
rect 362960 219784 363012 219836
rect 368480 219784 368532 219836
rect 375288 219784 375340 219836
rect 379520 219784 379572 219836
rect 380992 219784 381044 219836
rect 484400 219784 484452 219836
rect 535368 219784 535420 219836
rect 609888 219784 609940 219836
rect 172152 219716 172204 219768
rect 232412 219716 232464 219768
rect 250996 219716 251048 219768
rect 271144 219716 271196 219768
rect 337384 219716 337436 219768
rect 353300 219716 353352 219768
rect 372620 219716 372672 219768
rect 384304 219716 384356 219768
rect 387156 219716 387208 219768
rect 409880 219716 409932 219768
rect 409972 219716 410024 219768
rect 416228 219716 416280 219768
rect 515404 219716 515456 219768
rect 625344 219716 625396 219768
rect 185584 219648 185636 219700
rect 186964 219648 187016 219700
rect 181996 219580 182048 219632
rect 232780 219648 232832 219700
rect 252100 219648 252152 219700
rect 257344 219648 257396 219700
rect 261300 219648 261352 219700
rect 272984 219648 273036 219700
rect 334716 219648 334768 219700
rect 349804 219648 349856 219700
rect 386420 219648 386472 219700
rect 398840 219648 398892 219700
rect 415308 219648 415360 219700
rect 418160 219648 418212 219700
rect 512828 219648 512880 219700
rect 625252 219648 625304 219700
rect 188896 219580 188948 219632
rect 234620 219580 234672 219632
rect 300492 219580 300544 219632
rect 306932 219580 306984 219632
rect 334624 219580 334676 219632
rect 346492 219580 346544 219632
rect 377312 219580 377364 219632
rect 388536 219580 388588 219632
rect 498660 219580 498712 219632
rect 505008 219580 505060 219632
rect 509884 219580 509936 219632
rect 623872 219580 623924 219632
rect 97816 219512 97868 219564
rect 54392 219444 54444 219496
rect 56324 219444 56376 219496
rect 56600 219444 56652 219496
rect 195704 219512 195756 219564
rect 234712 219512 234764 219564
rect 301596 219512 301648 219564
rect 307760 219512 307812 219564
rect 406384 219512 406436 219564
rect 412916 219512 412968 219564
rect 502432 219512 502484 219564
rect 623044 219512 623096 219564
rect 195152 219444 195204 219496
rect 202420 219444 202472 219496
rect 237380 219444 237432 219496
rect 267188 219444 267240 219496
rect 268384 219444 268436 219496
rect 276480 219444 276532 219496
rect 278044 219444 278096 219496
rect 300584 219444 300636 219496
rect 306380 219444 306432 219496
rect 360292 219444 360344 219496
rect 364984 219444 365036 219496
rect 371332 219444 371384 219496
rect 375932 219444 375984 219496
rect 378508 219444 378560 219496
rect 385132 219444 385184 219496
rect 390652 219444 390704 219496
rect 393596 219444 393648 219496
rect 408500 219444 408552 219496
rect 414572 219444 414624 219496
rect 52276 219376 52328 219428
rect 350172 219376 350224 219428
rect 504916 219444 504968 219496
rect 623780 219444 623832 219496
rect 673368 219444 673420 219496
rect 676036 219444 676088 219496
rect 423864 219376 423916 219428
rect 354404 219308 354456 219360
rect 432236 219308 432288 219360
rect 353208 219240 353260 219292
rect 430580 219240 430632 219292
rect 379428 219172 379480 219224
rect 494520 219172 494572 219224
rect 570604 219172 570656 219224
rect 635924 219172 635976 219224
rect 380808 219104 380860 219156
rect 498200 219104 498252 219156
rect 555424 219104 555476 219156
rect 577504 219104 577556 219156
rect 383476 219036 383528 219088
rect 501236 219036 501288 219088
rect 548524 219036 548576 219088
rect 576216 219036 576268 219088
rect 383568 218968 383620 219020
rect 503720 218968 503772 219020
rect 505008 218968 505060 219020
rect 622952 218968 623004 219020
rect 386328 218900 386380 218952
rect 508780 218900 508832 218952
rect 557816 218900 557868 218952
rect 607680 218900 607732 218952
rect 387708 218832 387760 218884
rect 511356 218832 511408 218884
rect 561772 218832 561824 218884
rect 562876 218832 562928 218884
rect 616788 218832 616840 218884
rect 391848 218764 391900 218816
rect 521660 218764 521712 218816
rect 565452 218764 565504 218816
rect 619548 218764 619600 218816
rect 44824 218696 44876 218748
rect 659752 218696 659804 218748
rect 567936 218628 567988 218680
rect 627460 218628 627512 218680
rect 515496 218560 515548 218612
rect 576032 218560 576084 218612
rect 543188 218492 543240 218544
rect 543648 218492 543700 218544
rect 576124 218492 576176 218544
rect 487804 218424 487856 218476
rect 575940 218424 575992 218476
rect 495624 218356 495676 218408
rect 495992 218356 496044 218408
rect 619732 218356 619784 218408
rect 500224 218288 500276 218340
rect 637856 218288 637908 218340
rect 496084 218220 496136 218272
rect 637396 218220 637448 218272
rect 493416 218152 493468 218204
rect 636936 218152 636988 218204
rect 486424 218084 486476 218136
rect 118700 218016 118752 218068
rect 124864 218016 124916 218068
rect 487528 218016 487580 218068
rect 487804 218016 487856 218068
rect 489460 218084 489512 218136
rect 633716 218084 633768 218136
rect 638316 218016 638368 218068
rect 523040 217880 523092 217932
rect 523960 217880 524012 217932
rect 538220 217880 538272 217932
rect 539048 217880 539100 217932
rect 296812 217812 296864 217864
rect 297640 217812 297692 217864
rect 331220 217812 331272 217864
rect 332140 217812 332192 217864
rect 333980 217812 334032 217864
rect 334716 217812 334768 217864
rect 350632 217812 350684 217864
rect 351460 217812 351512 217864
rect 422300 217812 422352 217864
rect 423036 217812 423088 217864
rect 434720 217812 434772 217864
rect 435640 217812 435692 217864
rect 441620 217812 441672 217864
rect 442356 217812 442408 217864
rect 454040 217812 454092 217864
rect 454960 217812 455012 217864
rect 460940 217812 460992 217864
rect 461676 217812 461728 217864
rect 465080 217812 465132 217864
rect 465908 217812 465960 217864
rect 471980 217812 472032 217864
rect 472624 217812 472676 217864
rect 476120 217812 476172 217864
rect 476856 217812 476908 217864
rect 499580 217812 499632 217864
rect 500868 217812 500920 217864
rect 608508 217812 608560 217864
rect 497648 217744 497700 217796
rect 608048 217744 608100 217796
rect 490932 217676 490984 217728
rect 607128 217676 607180 217728
rect 553722 217608 553774 217660
rect 575848 217608 575900 217660
rect 609888 217608 609940 217660
rect 629484 217608 629536 217660
rect 568810 217540 568862 217592
rect 618352 217540 618404 217592
rect 556160 217472 556212 217524
rect 618720 217472 618772 217524
rect 549628 217404 549680 217456
rect 550548 217404 550600 217456
rect 632244 217404 632296 217456
rect 494336 217336 494388 217388
rect 578148 217336 578200 217388
rect 609612 217336 609664 217388
rect 632704 217336 632756 217388
rect 35808 217268 35860 217320
rect 43812 217268 43864 217320
rect 545580 217268 545632 217320
rect 631324 217268 631376 217320
rect 537944 217200 537996 217252
rect 629944 217200 629996 217252
rect 513656 217132 513708 217184
rect 610808 217132 610860 217184
rect 511080 217064 511132 217116
rect 610348 217064 610400 217116
rect 508504 216996 508556 217048
rect 609888 216996 609940 217048
rect 506112 216928 506164 216980
rect 609428 216928 609480 216980
rect 502524 216860 502576 216912
rect 503536 216860 503588 216912
rect 608968 216860 609020 216912
rect 564072 216792 564124 216844
rect 577044 216792 577096 216844
rect 561404 216724 561456 216776
rect 575756 216724 575808 216776
rect 558920 216656 558972 216708
rect 575664 216656 575716 216708
rect 52184 215908 52236 215960
rect 118700 216384 118752 216436
rect 518716 216384 518768 216436
rect 521200 216384 521252 216436
rect 523776 216384 523828 216436
rect 526260 216384 526312 216436
rect 528560 216384 528612 216436
rect 531228 216384 531280 216436
rect 533804 216384 533856 216436
rect 536380 216384 536432 216436
rect 538864 216384 538916 216436
rect 541440 216384 541492 216436
rect 551468 216384 551520 216436
rect 566464 216384 566516 216436
rect 574836 216384 574888 216436
rect 574928 216384 574980 216436
rect 613016 216316 613068 216368
rect 630404 216316 630456 216368
rect 614120 216248 614172 216300
rect 631784 216248 631836 216300
rect 626632 216180 626684 216232
rect 628472 216112 628524 216164
rect 673000 216112 673052 216164
rect 676036 216112 676088 216164
rect 577872 216044 577924 216096
rect 611728 216044 611780 216096
rect 630864 216044 630916 216096
rect 620560 215976 620612 216028
rect 615500 215840 615552 215892
rect 617156 215908 617208 215960
rect 634084 215908 634136 215960
rect 617800 215840 617852 215892
rect 615040 215772 615092 215824
rect 614580 215704 614632 215756
rect 674564 215704 674616 215756
rect 676036 215704 676088 215756
rect 614028 215636 614080 215688
rect 613568 215568 613620 215620
rect 613108 215500 613160 215552
rect 676220 215500 676272 215552
rect 676864 215500 676916 215552
rect 612648 215432 612700 215484
rect 612188 215364 612240 215416
rect 611728 215296 611780 215348
rect 35808 214548 35860 214600
rect 46204 214548 46256 214600
rect 50344 214344 50396 214396
rect 50068 214276 50120 214328
rect 47216 214208 47268 214260
rect 41328 214140 41380 214192
rect 31116 214072 31168 214124
rect 31300 214004 31352 214056
rect 41512 213936 41564 213988
rect 576400 214752 576452 214804
rect 626172 214752 626224 214804
rect 577136 214684 577188 214736
rect 627552 214684 627604 214736
rect 577320 214616 577372 214668
rect 627092 214616 627144 214668
rect 576308 214548 576360 214600
rect 628012 214548 628064 214600
rect 662512 214548 662564 214600
rect 663064 214548 663116 214600
rect 663800 214548 663852 214600
rect 664444 214548 664496 214600
rect 623872 214480 623924 214532
rect 624424 214480 624476 214532
rect 665272 214344 665324 214396
rect 668860 214276 668912 214328
rect 668124 214208 668176 214260
rect 668952 214140 669004 214192
rect 665732 214072 665784 214124
rect 673184 214072 673236 214124
rect 676036 214072 676088 214124
rect 666192 214004 666244 214056
rect 669044 213936 669096 213988
rect 575940 213868 575992 213920
rect 606668 213868 606720 213920
rect 607680 213868 607732 213920
rect 633624 213868 633676 213920
rect 633716 213868 633768 213920
rect 636384 213868 636436 213920
rect 636844 213868 636896 213920
rect 639236 213868 639288 213920
rect 639604 213868 639656 213920
rect 640616 213868 640668 213920
rect 576032 213800 576084 213852
rect 611268 213800 611320 213852
rect 619732 213800 619784 213852
rect 622492 213800 622544 213852
rect 577872 213732 577924 213784
rect 615960 213732 616012 213784
rect 576124 213664 576176 213716
rect 616420 213664 616472 213716
rect 616788 213664 616840 213716
rect 634544 213664 634596 213716
rect 673092 213664 673144 213716
rect 676036 213664 676088 213716
rect 576216 213596 576268 213648
rect 617340 213596 617392 213648
rect 576492 213528 576544 213580
rect 616880 213528 616932 213580
rect 575848 213460 575900 213512
rect 618260 213460 618312 213512
rect 577044 213392 577096 213444
rect 620100 213392 620152 213444
rect 627460 213392 627512 213444
rect 635464 213392 635516 213444
rect 575664 213324 575716 213376
rect 619180 213324 619232 213376
rect 619548 213324 619600 213376
rect 635004 213324 635056 213376
rect 575756 213256 575808 213308
rect 619640 213256 619692 213308
rect 621664 213256 621716 213308
rect 641076 213256 641128 213308
rect 643836 213256 643888 213308
rect 651472 213256 651524 213308
rect 577504 213188 577556 213240
rect 633164 213188 633216 213240
rect 642732 213188 642784 213240
rect 650092 213188 650144 213240
rect 578148 213120 578200 213172
rect 607588 213120 607640 213172
rect 645584 213120 645636 213172
rect 650000 213120 650052 213172
rect 646964 212984 647016 213036
rect 651380 212984 651432 213036
rect 618352 212508 618404 212560
rect 621020 212508 621072 212560
rect 583024 211148 583076 211200
rect 638776 211148 638828 211200
rect 670332 211148 670384 211200
rect 676036 211148 676088 211200
rect 652024 210400 652076 210452
rect 667204 210400 667256 210452
rect 639052 210060 639104 210112
rect 639788 210060 639840 210112
rect 578884 209720 578936 209772
rect 603080 209720 603132 209772
rect 579252 209652 579304 209704
rect 603172 209652 603224 209704
rect 578976 208292 579028 208344
rect 603080 208292 603132 208344
rect 578424 206932 578476 206984
rect 603080 206932 603132 206984
rect 578516 205572 578568 205624
rect 603080 205572 603132 205624
rect 579528 205504 579580 205556
rect 603172 205504 603224 205556
rect 578792 204212 578844 204264
rect 603080 204212 603132 204264
rect 35808 202852 35860 202904
rect 50344 202852 50396 202904
rect 579436 202784 579488 202836
rect 603080 202784 603132 202836
rect 673000 201832 673052 201884
rect 675392 201832 675444 201884
rect 578884 201424 578936 201476
rect 603080 201424 603132 201476
rect 674564 201424 674616 201476
rect 675392 201424 675444 201476
rect 579252 201356 579304 201408
rect 603172 201356 603224 201408
rect 675116 200676 675168 200728
rect 675392 200676 675444 200728
rect 578240 200064 578292 200116
rect 603080 200064 603132 200116
rect 578424 198636 578476 198688
rect 603080 198636 603132 198688
rect 673184 197412 673236 197464
rect 675484 197412 675536 197464
rect 579068 197276 579120 197328
rect 603172 197276 603224 197328
rect 674840 197004 674892 197056
rect 675392 197004 675444 197056
rect 579528 196596 579580 196648
rect 603080 196596 603132 196648
rect 673092 196528 673144 196580
rect 675392 196528 675444 196580
rect 579528 195236 579580 195288
rect 603080 195236 603132 195288
rect 579528 193808 579580 193860
rect 603080 193808 603132 193860
rect 42064 193128 42116 193180
rect 43352 193128 43404 193180
rect 579528 192448 579580 192500
rect 603080 192448 603132 192500
rect 674840 192448 674892 192500
rect 675392 192448 675444 192500
rect 579252 191836 579304 191888
rect 603080 191836 603132 191888
rect 42156 191632 42208 191684
rect 43260 191632 43312 191684
rect 42064 191428 42116 191480
rect 43168 191428 43220 191480
rect 42156 190816 42208 190868
rect 43444 190816 43496 190868
rect 675760 190612 675812 190664
rect 578240 190476 578292 190528
rect 603080 190476 603132 190528
rect 675760 190340 675812 190392
rect 579528 189116 579580 189168
rect 603080 189116 603132 189168
rect 579252 189048 579304 189100
rect 603172 189048 603224 189100
rect 578884 187688 578936 187740
rect 603080 187688 603132 187740
rect 42156 187620 42208 187672
rect 42984 187620 43036 187672
rect 579436 186328 579488 186380
rect 603080 186328 603132 186380
rect 42064 186260 42116 186312
rect 42892 186260 42944 186312
rect 42156 185852 42208 185904
rect 42800 185852 42852 185904
rect 579528 184968 579580 185020
rect 603172 184968 603224 185020
rect 578976 184900 579028 184952
rect 603080 184900 603132 184952
rect 667940 183880 667992 183932
rect 669964 183880 670016 183932
rect 579344 183540 579396 183592
rect 603080 183540 603132 183592
rect 42156 183404 42208 183456
rect 44180 183404 44232 183456
rect 578240 182180 578292 182232
rect 603080 182180 603132 182232
rect 578332 180888 578384 180940
rect 603172 180888 603224 180940
rect 578424 180820 578476 180872
rect 603080 180820 603132 180872
rect 578792 179392 578844 179444
rect 603080 179392 603132 179444
rect 667940 178780 667992 178832
rect 670056 178780 670108 178832
rect 671528 178304 671580 178356
rect 676036 178304 676088 178356
rect 668768 178168 668820 178220
rect 675944 178168 675996 178220
rect 578700 178032 578752 178084
rect 603080 178032 603132 178084
rect 674656 177284 674708 177336
rect 676036 177284 676088 177336
rect 670240 176808 670292 176860
rect 675944 176808 675996 176860
rect 579436 176740 579488 176792
rect 603172 176740 603224 176792
rect 579344 176672 579396 176724
rect 603080 176672 603132 176724
rect 672908 176672 672960 176724
rect 676036 176672 676088 176724
rect 673184 175992 673236 176044
rect 676036 175992 676088 176044
rect 672632 175652 672684 175704
rect 676036 175652 676088 175704
rect 580264 175244 580316 175296
rect 603080 175244 603132 175296
rect 673276 175176 673328 175228
rect 676036 175176 676088 175228
rect 673368 174836 673420 174888
rect 676036 174836 676088 174888
rect 580356 173884 580408 173936
rect 603080 173884 603132 173936
rect 668308 173748 668360 173800
rect 672724 173748 672776 173800
rect 579160 172524 579212 172576
rect 603080 172524 603132 172576
rect 676220 171232 676272 171284
rect 677048 171232 677100 171284
rect 579252 171096 579304 171148
rect 603080 171096 603132 171148
rect 676220 171096 676272 171148
rect 676864 171096 676916 171148
rect 674656 170280 674708 170332
rect 676036 170280 676088 170332
rect 579068 169804 579120 169856
rect 603172 169804 603224 169856
rect 578884 169736 578936 169788
rect 603080 169736 603132 169788
rect 673000 169464 673052 169516
rect 676036 169464 676088 169516
rect 674564 169056 674616 169108
rect 676036 169056 676088 169108
rect 668308 168648 668360 168700
rect 674196 168648 674248 168700
rect 673092 168580 673144 168632
rect 676036 168580 676088 168632
rect 578976 168376 579028 168428
rect 603080 168376 603132 168428
rect 669964 168240 670016 168292
rect 676036 168240 676088 168292
rect 671528 167832 671580 167884
rect 676036 167832 676088 167884
rect 583116 167016 583168 167068
rect 603080 167016 603132 167068
rect 674196 167016 674248 167068
rect 676036 167016 676088 167068
rect 578608 166948 578660 167000
rect 580264 166948 580316 167000
rect 581644 165588 581696 165640
rect 603080 165588 603132 165640
rect 578240 164432 578292 164484
rect 580356 164432 580408 164484
rect 581736 164228 581788 164280
rect 603080 164228 603132 164280
rect 579528 164160 579580 164212
rect 603724 164160 603776 164212
rect 667940 163820 667992 163872
rect 671344 163820 671396 163872
rect 580264 162868 580316 162920
rect 603080 162868 603132 162920
rect 675760 162800 675812 162852
rect 678244 162800 678296 162852
rect 584496 161440 584548 161492
rect 603080 161440 603132 161492
rect 675760 160964 675812 161016
rect 675760 160760 675812 160812
rect 579160 160080 579212 160132
rect 603080 160080 603132 160132
rect 579344 158720 579396 158772
rect 603080 158720 603132 158772
rect 592684 157428 592736 157480
rect 603172 157428 603224 157480
rect 584404 157360 584456 157412
rect 603080 157360 603132 157412
rect 585784 155932 585836 155984
rect 603080 155932 603132 155984
rect 673000 155456 673052 155508
rect 675484 155456 675536 155508
rect 578332 154844 578384 154896
rect 583116 154844 583168 154896
rect 579252 154572 579304 154624
rect 603080 154572 603132 154624
rect 579068 153280 579120 153332
rect 603172 153280 603224 153332
rect 578884 153212 578936 153264
rect 603080 153212 603132 153264
rect 579528 153144 579580 153196
rect 603816 153144 603868 153196
rect 674564 152532 674616 152584
rect 675392 152532 675444 152584
rect 580356 151784 580408 151836
rect 603080 151784 603132 151836
rect 579436 151580 579488 151632
rect 581644 151580 581696 151632
rect 673092 151376 673144 151428
rect 675392 151376 675444 151428
rect 578976 150424 579028 150476
rect 603080 150424 603132 150476
rect 674656 150356 674708 150408
rect 675392 150356 675444 150408
rect 579436 150220 579488 150272
rect 581736 150220 581788 150272
rect 589924 149064 589976 149116
rect 603080 149064 603132 149116
rect 578516 148588 578568 148640
rect 580264 148588 580316 148640
rect 668308 148384 668360 148436
rect 674288 148384 674340 148436
rect 587256 147636 587308 147688
rect 603080 147636 603132 147688
rect 579528 146956 579580 147008
rect 583024 146956 583076 147008
rect 579620 146888 579672 146940
rect 603724 146888 603776 146940
rect 591304 146276 591356 146328
rect 603080 146276 603132 146328
rect 578700 146140 578752 146192
rect 584496 146140 584548 146192
rect 583024 144916 583076 144968
rect 603172 144916 603224 144968
rect 580264 143556 580316 143608
rect 603080 143556 603132 143608
rect 578700 143488 578752 143540
rect 592684 143488 592736 143540
rect 667940 143420 667992 143472
rect 670148 143420 670200 143472
rect 591488 142128 591540 142180
rect 603080 142128 603132 142180
rect 588636 140768 588688 140820
rect 603080 140768 603132 140820
rect 584680 140020 584732 140072
rect 603908 140020 603960 140072
rect 594156 139408 594208 139460
rect 603080 139408 603132 139460
rect 667940 138184 667992 138236
rect 671436 138184 671488 138236
rect 590108 138048 590160 138100
rect 603080 138048 603132 138100
rect 587164 137980 587216 138032
rect 603172 137980 603224 138032
rect 579528 137912 579580 137964
rect 585784 137912 585836 137964
rect 588544 136620 588596 136672
rect 603080 136620 603132 136672
rect 579528 136484 579580 136536
rect 584404 136484 584456 136536
rect 585784 135260 585836 135312
rect 603080 135260 603132 135312
rect 585968 133968 586020 134020
rect 603172 133968 603224 134020
rect 581828 133900 581880 133952
rect 603080 133900 603132 133952
rect 581644 133152 581696 133204
rect 603724 133152 603776 133204
rect 674104 133016 674156 133068
rect 676036 133016 676088 133068
rect 668584 132948 668636 133000
rect 674380 132948 674432 133000
rect 672816 132744 672868 132796
rect 676220 132744 676272 132796
rect 667204 132608 667256 132660
rect 676128 132608 676180 132660
rect 592776 132472 592828 132524
rect 603080 132472 603132 132524
rect 672908 131384 672960 131436
rect 676220 131384 676272 131436
rect 673184 131248 673236 131300
rect 676036 131248 676088 131300
rect 584588 131112 584640 131164
rect 603080 131112 603132 131164
rect 668676 131112 668728 131164
rect 669044 131112 669096 131164
rect 676128 131112 676180 131164
rect 578332 130500 578384 130552
rect 580356 130500 580408 130552
rect 673276 129956 673328 130008
rect 676220 129956 676272 130008
rect 583116 129820 583168 129872
rect 603172 129820 603224 129872
rect 672724 129820 672776 129872
rect 676128 129820 676180 129872
rect 581736 129752 581788 129804
rect 603080 129752 603132 129804
rect 668584 129752 668636 129804
rect 668952 129752 669004 129804
rect 676220 129752 676272 129804
rect 584496 128324 584548 128376
rect 603080 128324 603132 128376
rect 668768 128324 668820 128376
rect 676220 128324 676272 128376
rect 579528 128256 579580 128308
rect 587256 128256 587308 128308
rect 667940 127916 667992 127968
rect 671620 127916 671672 127968
rect 580356 126964 580408 127016
rect 603080 126964 603132 127016
rect 675116 126964 675168 127016
rect 676036 126964 676088 127016
rect 578700 126012 578752 126064
rect 584680 126012 584732 126064
rect 594064 125672 594116 125724
rect 603080 125672 603132 125724
rect 587256 125604 587308 125656
rect 603172 125604 603224 125656
rect 578424 125536 578476 125588
rect 589924 125536 589976 125588
rect 591396 124176 591448 124228
rect 603080 124176 603132 124228
rect 579252 124108 579304 124160
rect 591304 124108 591356 124160
rect 667940 124040 667992 124092
rect 670332 124040 670384 124092
rect 674656 123904 674708 123956
rect 676036 123904 676088 123956
rect 598204 122884 598256 122936
rect 603172 122884 603224 122936
rect 592684 122816 592736 122868
rect 603080 122816 603132 122868
rect 668860 122816 668912 122868
rect 676220 122816 676272 122868
rect 579436 122068 579488 122120
rect 591488 122068 591540 122120
rect 591304 121456 591356 121508
rect 603080 121456 603132 121508
rect 671344 121456 671396 121508
rect 676128 121456 676180 121508
rect 579528 121388 579580 121440
rect 583024 121388 583076 121440
rect 670056 120708 670108 120760
rect 676220 120708 676272 120760
rect 590016 120096 590068 120148
rect 603080 120096 603132 120148
rect 579252 120028 579304 120080
rect 581644 120028 581696 120080
rect 579160 118668 579212 118720
rect 603080 118668 603132 118720
rect 578516 118532 578568 118584
rect 580264 118532 580316 118584
rect 667940 117716 667992 117768
rect 669964 117716 670016 117768
rect 579068 117308 579120 117360
rect 603080 117308 603132 117360
rect 579528 117240 579580 117292
rect 603816 117240 603868 117292
rect 668400 116968 668452 117020
rect 671528 116968 671580 117020
rect 675484 116696 675536 116748
rect 677600 116696 677652 116748
rect 675208 116560 675260 116612
rect 683304 116560 683356 116612
rect 678244 116152 678296 116204
rect 675484 115744 675536 115796
rect 675116 115540 675168 115592
rect 675392 115540 675444 115592
rect 675116 115404 675168 115456
rect 675208 114792 675260 114844
rect 675392 114792 675444 114844
rect 596824 114588 596876 114640
rect 603172 114588 603224 114640
rect 675116 114588 675168 114640
rect 578976 114520 579028 114572
rect 603080 114520 603132 114572
rect 579252 114452 579304 114504
rect 588636 114452 588688 114504
rect 669228 114316 669280 114368
rect 674196 114316 674248 114368
rect 578884 113160 578936 113212
rect 603080 113160 603132 113212
rect 579528 113092 579580 113144
rect 594156 113092 594208 113144
rect 595444 111800 595496 111852
rect 603080 111800 603132 111852
rect 578700 111732 578752 111784
rect 587164 111732 587216 111784
rect 668308 111732 668360 111784
rect 671344 111732 671396 111784
rect 675208 111120 675260 111172
rect 675392 111120 675444 111172
rect 675116 110644 675168 110696
rect 675392 110644 675444 110696
rect 589924 110440 589976 110492
rect 603080 110440 603132 110492
rect 579528 110372 579580 110424
rect 590108 110372 590160 110424
rect 667940 109284 667992 109336
rect 670056 109284 670108 109336
rect 588636 109012 588688 109064
rect 603080 109012 603132 109064
rect 578792 108944 578844 108996
rect 588544 108944 588596 108996
rect 585876 107652 585928 107704
rect 603080 107652 603132 107704
rect 674656 107516 674708 107568
rect 675392 107516 675444 107568
rect 579436 107040 579488 107092
rect 585784 107040 585836 107092
rect 675116 106700 675168 106752
rect 675392 106700 675444 106752
rect 588544 106360 588596 106412
rect 603172 106360 603224 106412
rect 587164 106292 587216 106344
rect 603080 106292 603132 106344
rect 674748 106224 674800 106276
rect 675392 106224 675444 106276
rect 669228 106088 669280 106140
rect 672724 106088 672776 106140
rect 578240 105136 578292 105188
rect 585968 105136 586020 105188
rect 585784 104864 585836 104916
rect 603080 104864 603132 104916
rect 584404 103504 584456 103556
rect 603080 103504 603132 103556
rect 579344 103436 579396 103488
rect 581828 103436 581880 103488
rect 583024 102212 583076 102264
rect 603172 102212 603224 102264
rect 581644 102144 581696 102196
rect 603080 102144 603132 102196
rect 578332 102076 578384 102128
rect 592776 102076 592828 102128
rect 580264 100716 580316 100768
rect 603080 100716 603132 100768
rect 578700 100308 578752 100360
rect 584588 100308 584640 100360
rect 600964 99356 601016 99408
rect 603448 99356 603500 99408
rect 579528 99084 579580 99136
rect 583116 99084 583168 99136
rect 624608 97928 624660 97980
rect 625804 97928 625856 97980
rect 633808 97928 633860 97980
rect 636384 97928 636436 97980
rect 663064 97928 663116 97980
rect 665364 97928 665416 97980
rect 633072 97860 633124 97912
rect 635280 97860 635332 97912
rect 637488 97860 637540 97912
rect 644664 97860 644716 97912
rect 649448 97860 649500 97912
rect 658832 97860 658884 97912
rect 638316 97792 638368 97844
rect 644756 97792 644808 97844
rect 647516 97792 647568 97844
rect 654784 97792 654836 97844
rect 635096 97724 635148 97776
rect 639052 97724 639104 97776
rect 634452 97656 634504 97708
rect 637580 97656 637632 97708
rect 578700 97588 578752 97640
rect 581736 97588 581788 97640
rect 631140 97588 631192 97640
rect 632152 97588 632204 97640
rect 635740 97588 635792 97640
rect 639880 97588 639932 97640
rect 637028 97520 637080 97572
rect 642180 97520 642232 97572
rect 614856 97452 614908 97504
rect 621664 97452 621716 97504
rect 643560 97452 643612 97504
rect 660396 97452 660448 97504
rect 620744 97384 620796 97436
rect 646044 97384 646096 97436
rect 648160 97384 648212 97436
rect 660120 97384 660172 97436
rect 652024 97316 652076 97368
rect 622032 97248 622084 97300
rect 648620 97248 648672 97300
rect 621388 97180 621440 97232
rect 647424 97180 647476 97232
rect 631784 97112 631836 97164
rect 632980 97112 633032 97164
rect 655980 97316 656032 97368
rect 659568 97316 659620 97368
rect 657728 97248 657780 97300
rect 660672 97248 660724 97300
rect 654692 97180 654744 97232
rect 658372 97180 658424 97232
rect 660580 97180 660632 97232
rect 661408 97180 661460 97232
rect 661960 97112 662012 97164
rect 662328 97112 662380 97164
rect 663984 97112 664036 97164
rect 610072 96908 610124 96960
rect 610900 96908 610952 96960
rect 611360 96908 611412 96960
rect 612188 96908 612240 96960
rect 616144 96908 616196 96960
rect 616788 96908 616840 96960
rect 617432 96908 617484 96960
rect 618168 96908 618220 96960
rect 623688 96908 623740 96960
rect 624424 96908 624476 96960
rect 625896 96908 625948 96960
rect 626448 96908 626500 96960
rect 645492 96908 645544 96960
rect 646504 96908 646556 96960
rect 655428 96908 655480 96960
rect 659292 96908 659344 96960
rect 618720 96840 618772 96892
rect 619548 96840 619600 96892
rect 620008 96840 620060 96892
rect 620928 96840 620980 96892
rect 632428 96840 632480 96892
rect 634084 96840 634136 96892
rect 640984 96840 641036 96892
rect 643284 96840 643336 96892
rect 650736 96840 650788 96892
rect 651288 96840 651340 96892
rect 661868 96840 661920 96892
rect 663064 96840 663116 96892
rect 622676 96772 622728 96824
rect 623688 96772 623740 96824
rect 659200 96772 659252 96824
rect 662512 96772 662564 96824
rect 636108 96704 636160 96756
rect 640984 96704 641036 96756
rect 639604 96568 639656 96620
rect 643100 96568 643152 96620
rect 644848 96568 644900 96620
rect 651932 96568 651984 96620
rect 656808 96568 656860 96620
rect 658280 96568 658332 96620
rect 656624 96160 656676 96212
rect 663892 96160 663944 96212
rect 646780 96024 646832 96076
rect 663800 96024 663852 96076
rect 578516 95956 578568 96008
rect 584496 95956 584548 96008
rect 653312 95956 653364 96008
rect 665272 95956 665324 96008
rect 640064 95888 640116 95940
rect 644572 95888 644624 95940
rect 646136 95888 646188 95940
rect 665180 95888 665232 95940
rect 641628 95616 641680 95668
rect 645952 95616 646004 95668
rect 638868 95548 638920 95600
rect 644480 95548 644532 95600
rect 607220 95480 607272 95532
rect 607680 95480 607732 95532
rect 657268 95208 657320 95260
rect 664076 95208 664128 95260
rect 578608 95140 578660 95192
rect 580356 95140 580408 95192
rect 579528 93780 579580 93832
rect 587256 93780 587308 93832
rect 579528 92420 579580 92472
rect 594064 92420 594116 92472
rect 644388 92420 644440 92472
rect 654324 92420 654376 92472
rect 579528 90992 579580 91044
rect 591396 90992 591448 91044
rect 651932 90924 651984 90976
rect 654324 90924 654376 90976
rect 579528 89632 579580 89684
rect 592684 89632 592736 89684
rect 616696 89632 616748 89684
rect 626448 89632 626500 89684
rect 656808 88816 656860 88868
rect 658096 88816 658148 88868
rect 662328 88816 662380 88868
rect 663984 88816 664036 88868
rect 616788 88272 616840 88324
rect 626448 88272 626500 88324
rect 659476 88272 659528 88324
rect 663156 88272 663208 88324
rect 620928 88204 620980 88256
rect 626356 88204 626408 88256
rect 584496 87592 584548 87644
rect 603724 87592 603776 87644
rect 646504 86980 646556 87032
rect 660120 86980 660172 87032
rect 579528 86912 579580 86964
rect 598204 86912 598256 86964
rect 651196 86912 651248 86964
rect 657176 86912 657228 86964
rect 651288 86844 651340 86896
rect 657728 86844 657780 86896
rect 649908 86776 649960 86828
rect 660672 86776 660724 86828
rect 648528 86708 648580 86760
rect 661408 86708 661460 86760
rect 653956 86640 654008 86692
rect 658832 86640 658884 86692
rect 652668 86572 652720 86624
rect 662512 86572 662564 86624
rect 619456 86232 619508 86284
rect 626448 86232 626500 86284
rect 579528 85484 579580 85536
rect 591304 85484 591356 85536
rect 619548 85484 619600 85536
rect 626448 85484 626500 85536
rect 579528 84124 579580 84176
rect 590016 84124 590068 84176
rect 618168 84124 618220 84176
rect 626080 84124 626132 84176
rect 618076 84056 618128 84108
rect 625620 84056 625672 84108
rect 581736 82084 581788 82136
rect 603816 82084 603868 82136
rect 579528 80860 579580 80912
rect 584496 80860 584548 80912
rect 624424 80656 624476 80708
rect 648712 80656 648764 80708
rect 623596 79296 623648 79348
rect 647332 79296 647384 79348
rect 579528 78616 579580 78668
rect 602344 78616 602396 78668
rect 626448 78140 626500 78192
rect 642456 78140 642508 78192
rect 631048 78072 631100 78124
rect 638960 78072 639012 78124
rect 629208 78004 629260 78056
rect 645308 78004 645360 78056
rect 605748 77936 605800 77988
rect 636752 77936 636804 77988
rect 628380 77596 628432 77648
rect 631508 77596 631560 77648
rect 579068 77324 579120 77376
rect 628380 77324 628432 77376
rect 576124 77256 576176 77308
rect 631048 77256 631100 77308
rect 623688 76508 623740 76560
rect 646136 76508 646188 76560
rect 579528 75828 579580 75880
rect 596824 75828 596876 75880
rect 617524 75216 617576 75268
rect 631140 75216 631192 75268
rect 615408 75148 615460 75200
rect 646872 75148 646924 75200
rect 579528 71680 579580 71732
rect 595444 71680 595496 71732
rect 579252 70252 579304 70304
rect 581736 70252 581788 70304
rect 578700 68960 578752 69012
rect 589924 68960 589976 69012
rect 579528 67532 579580 67584
rect 588636 67532 588688 67584
rect 579528 65900 579580 65952
rect 585876 65900 585928 65952
rect 578700 64812 578752 64864
rect 588544 64812 588596 64864
rect 579528 63452 579580 63504
rect 587164 63452 587216 63504
rect 578700 62024 578752 62076
rect 585784 62024 585836 62076
rect 614764 62024 614816 62076
rect 617524 62092 617576 62144
rect 578884 60664 578936 60716
rect 584404 60664 584456 60716
rect 578884 58760 578936 58812
rect 583024 58760 583076 58812
rect 578884 57876 578936 57928
rect 581644 57876 581696 57928
rect 578332 57196 578384 57248
rect 600964 57196 601016 57248
rect 621664 57196 621716 57248
rect 662420 57196 662472 57248
rect 578240 55632 578292 55684
rect 580264 55632 580316 55684
rect 405096 53116 405148 53168
rect 608784 53116 608836 53168
rect 145380 53048 145432 53100
rect 579068 53048 579120 53100
rect 52276 52436 52328 52488
rect 346814 52436 346866 52488
rect 614764 52436 614816 52488
rect 478144 49716 478196 49768
rect 478788 49716 478840 49768
rect 664260 49512 664312 49564
rect 672080 49512 672132 49564
rect 194048 46180 194100 46232
rect 661472 46180 661524 46232
rect 473176 42476 473228 42528
rect 415124 42340 415176 42392
<< metal2 >>
rect 110170 1029098 110262 1029126
rect 212934 1029098 213026 1029126
rect 264362 1029098 264454 1029126
rect 315974 1029098 316066 1029126
rect 366390 1029098 366482 1029126
rect 433734 1029098 433826 1029126
rect 510738 1029098 510830 1029126
rect 562166 1029098 562258 1029126
rect 110170 1028622 110262 1028650
rect 212934 1028622 213026 1028650
rect 264362 1028622 264454 1028650
rect 315974 1028622 316066 1028650
rect 366390 1028622 366482 1028650
rect 433734 1028622 433826 1028650
rect 510738 1028622 510830 1028650
rect 562166 1028622 562258 1028650
rect 110170 1028177 110262 1028205
rect 212934 1028177 213026 1028205
rect 264362 1028177 264454 1028205
rect 315974 1028177 316066 1028205
rect 366390 1028177 366482 1028205
rect 433734 1028177 433826 1028205
rect 510738 1028177 510830 1028205
rect 562166 1028177 562258 1028205
rect 366284 1027806 366496 1027834
rect 110170 1027738 110262 1027766
rect 212934 1027738 213026 1027766
rect 264362 1027738 264454 1027766
rect 315974 1027738 316066 1027766
rect 366284 1027752 366312 1027806
rect 366468 1027752 366496 1027806
rect 433734 1027738 433826 1027766
rect 510738 1027738 510830 1027766
rect 562166 1027738 562258 1027766
rect 110170 1027262 110262 1027290
rect 212934 1027262 213026 1027290
rect 264362 1027262 264454 1027290
rect 315974 1027262 316066 1027290
rect 366390 1027262 366482 1027290
rect 433734 1027262 433826 1027290
rect 510738 1027262 510830 1027290
rect 562166 1027262 562258 1027290
rect 110170 1026786 110262 1026814
rect 212934 1026786 213026 1026814
rect 264362 1026786 264454 1026814
rect 315974 1026786 316066 1026814
rect 366390 1026786 366482 1026814
rect 433734 1026786 433826 1026814
rect 510738 1026786 510830 1026814
rect 562166 1026786 562258 1026814
rect 110170 1026310 110262 1026338
rect 212934 1026310 213026 1026338
rect 264362 1026310 264454 1026338
rect 315974 1026310 316066 1026338
rect 366284 1026202 366312 1026324
rect 366468 1026202 366496 1026324
rect 433734 1026310 433826 1026338
rect 510738 1026310 510830 1026338
rect 562166 1026310 562258 1026338
rect 366284 1026174 366496 1026202
rect 366284 1026038 366496 1026066
rect 110170 1025902 110262 1025930
rect 212934 1025902 213026 1025930
rect 264362 1025902 264454 1025930
rect 315974 1025902 316066 1025930
rect 366284 1025916 366312 1026038
rect 366468 1025916 366496 1026038
rect 433734 1025902 433826 1025930
rect 510738 1025902 510830 1025930
rect 562166 1025902 562258 1025930
rect 110170 1025426 110262 1025454
rect 212934 1025426 213026 1025454
rect 264362 1025426 264454 1025454
rect 315974 1025426 316066 1025454
rect 366390 1025426 366482 1025454
rect 433734 1025426 433826 1025454
rect 510738 1025426 510830 1025454
rect 562166 1025426 562258 1025454
rect 110170 1024950 110262 1024978
rect 212934 1024950 213026 1024978
rect 264362 1024950 264454 1024978
rect 315974 1024950 316066 1024978
rect 366390 1024950 366482 1024978
rect 433734 1024950 433826 1024978
rect 510738 1024950 510830 1024978
rect 562166 1024950 562258 1024978
rect 110170 1024474 110262 1024502
rect 212934 1024474 213026 1024502
rect 264362 1024474 264454 1024502
rect 315974 1024474 316066 1024502
rect 366284 1024434 366312 1024488
rect 366468 1024434 366496 1024488
rect 433734 1024474 433826 1024502
rect 510738 1024474 510830 1024502
rect 562166 1024474 562258 1024502
rect 366284 1024406 366496 1024434
rect 110170 1024037 110262 1024065
rect 212934 1024037 213026 1024065
rect 264362 1024037 264454 1024065
rect 315974 1024037 316066 1024065
rect 366390 1024037 366482 1024065
rect 433734 1024037 433826 1024065
rect 510738 1024037 510830 1024065
rect 562166 1024037 562258 1024065
rect 110170 1023590 110262 1023618
rect 212934 1023590 213026 1023618
rect 264362 1023590 264454 1023618
rect 315974 1023590 316066 1023618
rect 366390 1023590 366482 1023618
rect 433734 1023590 433826 1023618
rect 510738 1023590 510830 1023618
rect 562166 1023590 562258 1023618
rect 203890 1007176 203946 1007185
rect 195336 1007140 195388 1007146
rect 203890 1007111 203892 1007120
rect 195336 1007082 195388 1007088
rect 203944 1007111 203946 1007120
rect 203892 1007082 203944 1007088
rect 99930 1006632 99986 1006641
rect 92612 1006596 92664 1006602
rect 99930 1006567 99932 1006576
rect 92612 1006538 92664 1006544
rect 99984 1006567 99986 1006576
rect 99932 1006538 99984 1006544
rect 92520 1003332 92572 1003338
rect 92520 1003274 92572 1003280
rect 92336 1002040 92388 1002046
rect 92256 1001988 92336 1001994
rect 92256 1001982 92388 1001988
rect 92256 1001966 92376 1001982
rect 92256 995858 92284 1001966
rect 92428 1001224 92480 1001230
rect 92428 1001166 92480 1001172
rect 92336 999116 92388 999122
rect 92336 999058 92388 999064
rect 85304 995852 85356 995858
rect 85304 995794 85356 995800
rect 92244 995852 92296 995858
rect 92244 995794 92296 995800
rect 85316 995738 85344 995794
rect 92348 995790 92376 999058
rect 91560 995784 91612 995790
rect 86498 995752 86554 995761
rect 85054 995710 85344 995738
rect 86342 995710 86498 995738
rect 89626 995752 89682 995761
rect 87538 995722 87920 995738
rect 87538 995716 87932 995722
rect 87538 995710 87880 995716
rect 86498 995687 86554 995696
rect 89378 995710 89626 995738
rect 91218 995732 91560 995738
rect 91218 995726 91612 995732
rect 92336 995784 92388 995790
rect 92336 995726 92388 995732
rect 91218 995710 91600 995726
rect 92440 995722 92468 1001166
rect 92532 996577 92560 1003274
rect 92624 1002046 92652 1006538
rect 95976 1006528 96028 1006534
rect 104808 1006528 104860 1006534
rect 95976 1006470 96028 1006476
rect 104346 1006496 104402 1006505
rect 93216 1006460 93268 1006466
rect 93216 1006402 93268 1006408
rect 93124 1006324 93176 1006330
rect 93124 1006266 93176 1006272
rect 92612 1002040 92664 1002046
rect 92612 1001982 92664 1001988
rect 92704 1000544 92756 1000550
rect 92704 1000486 92756 1000492
rect 92612 997892 92664 997898
rect 92612 997834 92664 997840
rect 92518 996568 92574 996577
rect 92518 996503 92574 996512
rect 92428 995716 92480 995722
rect 89626 995687 89682 995696
rect 87880 995658 87932 995664
rect 92428 995658 92480 995664
rect 82358 995616 82414 995625
rect 82018 995574 82358 995602
rect 85946 995616 86002 995625
rect 85698 995574 85946 995602
rect 82358 995551 82414 995560
rect 85946 995551 86002 995560
rect 92624 995489 92652 997834
rect 84658 995480 84714 995489
rect 77036 995110 77064 995452
rect 77680 995178 77708 995452
rect 78324 995314 78352 995452
rect 78312 995308 78364 995314
rect 78312 995250 78364 995256
rect 77668 995172 77720 995178
rect 77668 995114 77720 995120
rect 77024 995104 77076 995110
rect 80164 995081 80192 995452
rect 80716 995246 80744 995452
rect 81268 995438 81374 995466
rect 84502 995438 84658 995466
rect 81268 995382 81296 995438
rect 92610 995480 92666 995489
rect 84658 995415 84714 995424
rect 81256 995376 81308 995382
rect 81256 995318 81308 995324
rect 80704 995240 80756 995246
rect 80704 995182 80756 995188
rect 77024 995046 77076 995052
rect 80150 995072 80206 995081
rect 88720 995042 88748 995452
rect 92610 995415 92666 995424
rect 92716 995081 92744 1000486
rect 93136 995625 93164 1006266
rect 93228 996441 93256 1006402
rect 94688 1006188 94740 1006194
rect 94688 1006130 94740 1006136
rect 94504 1006052 94556 1006058
rect 94504 1005994 94556 1006000
rect 94516 997898 94544 1005994
rect 94596 1004692 94648 1004698
rect 94596 1004634 94648 1004640
rect 94608 999122 94636 1004634
rect 94700 1000550 94728 1006130
rect 95884 1002244 95936 1002250
rect 95884 1002186 95936 1002192
rect 94688 1000544 94740 1000550
rect 94688 1000486 94740 1000492
rect 94596 999116 94648 999122
rect 94596 999058 94648 999064
rect 94504 997892 94556 997898
rect 94504 997834 94556 997840
rect 93214 996432 93270 996441
rect 93214 996367 93270 996376
rect 93122 995616 93178 995625
rect 93122 995551 93178 995560
rect 95896 995382 95924 1002186
rect 95884 995376 95936 995382
rect 95884 995318 95936 995324
rect 95988 995314 96016 1006470
rect 104346 1006431 104348 1006440
rect 104400 1006431 104402 1006440
rect 104806 1006496 104808 1006505
rect 104860 1006496 104862 1006505
rect 104806 1006431 104862 1006440
rect 104348 1006402 104400 1006408
rect 99104 1006392 99156 1006398
rect 126244 1006392 126296 1006398
rect 99104 1006334 99156 1006340
rect 100666 1006360 100722 1006369
rect 99116 1006126 99144 1006334
rect 149704 1006392 149756 1006398
rect 126244 1006334 126296 1006340
rect 149702 1006360 149704 1006369
rect 150900 1006392 150952 1006398
rect 149756 1006360 149758 1006369
rect 100666 1006295 100668 1006304
rect 100720 1006295 100722 1006304
rect 100668 1006266 100720 1006272
rect 103610 1006224 103666 1006233
rect 103610 1006159 103612 1006168
rect 103664 1006159 103666 1006168
rect 103612 1006130 103664 1006136
rect 98276 1006120 98328 1006126
rect 98274 1006088 98276 1006097
rect 99104 1006120 99156 1006126
rect 98328 1006088 98330 1006097
rect 98274 1006023 98330 1006032
rect 99102 1006088 99104 1006097
rect 102784 1006120 102836 1006126
rect 99156 1006088 99158 1006097
rect 108856 1006120 108908 1006126
rect 102784 1006062 102836 1006068
rect 103150 1006088 103206 1006097
rect 99102 1006023 99158 1006032
rect 99470 1003368 99526 1003377
rect 99470 1003303 99472 1003312
rect 99524 1003303 99526 1003312
rect 99472 1003274 99524 1003280
rect 101494 1002280 101550 1002289
rect 101494 1002215 101496 1002224
rect 101548 1002215 101550 1002224
rect 101496 1002186 101548 1002192
rect 97356 1002176 97408 1002182
rect 102324 1002176 102376 1002182
rect 97356 1002118 97408 1002124
rect 100298 1002144 100354 1002153
rect 97264 1002108 97316 1002114
rect 97264 1002050 97316 1002056
rect 97276 996305 97304 1002050
rect 97262 996296 97318 996305
rect 97262 996231 97318 996240
rect 95976 995308 96028 995314
rect 95976 995250 96028 995256
rect 97368 995178 97396 1002118
rect 100298 1002079 100300 1002088
rect 100352 1002079 100354 1002088
rect 102322 1002144 102324 1002153
rect 102376 1002144 102378 1002153
rect 102322 1002079 102378 1002088
rect 100300 1002050 100352 1002056
rect 98644 1002040 98696 1002046
rect 101128 1002040 101180 1002046
rect 98644 1001982 98696 1001988
rect 101126 1002008 101128 1002017
rect 101180 1002008 101182 1002017
rect 98656 1001230 98684 1001982
rect 100024 1001972 100076 1001978
rect 101126 1001943 101182 1001952
rect 101954 1002008 102010 1002017
rect 101954 1001943 101956 1001952
rect 100024 1001914 100076 1001920
rect 102008 1001943 102010 1001952
rect 101956 1001914 102008 1001920
rect 98644 1001224 98696 1001230
rect 98644 1001166 98696 1001172
rect 100036 995246 100064 1001914
rect 100024 995240 100076 995246
rect 100024 995182 100076 995188
rect 97356 995172 97408 995178
rect 97356 995114 97408 995120
rect 92702 995072 92758 995081
rect 80150 995007 80206 995016
rect 88708 995036 88760 995042
rect 92702 995007 92758 995016
rect 88708 994978 88760 994984
rect 48964 992928 49016 992934
rect 48964 992870 49016 992876
rect 47584 991568 47636 991574
rect 47584 991510 47636 991516
rect 44824 991500 44876 991506
rect 44824 991442 44876 991448
rect 42708 975724 42760 975730
rect 42708 975666 42760 975672
rect 41800 968833 41828 969272
rect 41786 968824 41842 968833
rect 41786 968759 41842 968768
rect 41800 967337 41828 967405
rect 41786 967328 41842 967337
rect 42720 967298 42748 975666
rect 41786 967263 41842 967272
rect 42156 967292 42208 967298
rect 42156 967234 42208 967240
rect 42708 967292 42760 967298
rect 42708 967234 42760 967240
rect 42168 966756 42196 967234
rect 42076 965161 42104 965565
rect 42062 965152 42118 965161
rect 42062 965087 42118 965096
rect 42168 964034 42196 964376
rect 42156 964028 42208 964034
rect 42156 963970 42208 963976
rect 42800 964028 42852 964034
rect 42800 963970 42852 963976
rect 41800 963393 41828 963725
rect 41786 963384 41842 963393
rect 41786 963319 41842 963328
rect 42168 962878 42196 963084
rect 42156 962872 42208 962878
rect 42156 962814 42208 962820
rect 41800 962169 41828 962540
rect 41786 962160 41842 962169
rect 41786 962095 41842 962104
rect 42076 959750 42104 960024
rect 42064 959744 42116 959750
rect 42064 959686 42116 959692
rect 42168 959138 42196 959412
rect 42156 959132 42208 959138
rect 42156 959074 42208 959080
rect 41800 958361 41828 958732
rect 41786 958352 41842 958361
rect 41786 958287 41842 958296
rect 42076 957817 42104 958188
rect 42062 957808 42118 957817
rect 42062 957743 42118 957752
rect 42182 956338 42380 956366
rect 42168 955482 42196 955740
rect 42352 955602 42380 956338
rect 42340 955596 42392 955602
rect 42340 955538 42392 955544
rect 42708 955596 42760 955602
rect 42708 955538 42760 955544
rect 42168 955454 42380 955482
rect 42168 955182 42288 955210
rect 42168 955060 42196 955182
rect 42260 954394 42288 955182
rect 41892 954366 42288 954394
rect 36544 952264 36596 952270
rect 36544 952206 36596 952212
rect 37922 952232 37978 952241
rect 32402 951688 32458 951697
rect 32402 951623 32458 951632
rect 31024 951516 31076 951522
rect 31024 951458 31076 951464
rect 8588 944180 8616 944316
rect 9048 944180 9076 944316
rect 9508 944180 9536 944316
rect 9968 944180 9996 944316
rect 10428 944180 10456 944316
rect 10888 944180 10916 944316
rect 11348 944180 11376 944316
rect 11808 944180 11836 944316
rect 12268 944180 12296 944316
rect 12728 944180 12756 944316
rect 13188 944180 13216 944316
rect 13648 944180 13676 944316
rect 14108 944180 14136 944316
rect 31036 938233 31064 951458
rect 31022 938224 31078 938233
rect 31022 938159 31078 938168
rect 32416 937417 32444 951623
rect 34520 946008 34572 946014
rect 34520 945950 34572 945956
rect 34532 943809 34560 945950
rect 34518 943800 34574 943809
rect 34518 943735 34574 943744
rect 35808 943288 35860 943294
rect 35808 943230 35860 943236
rect 35716 943220 35768 943226
rect 35716 943162 35768 943168
rect 35728 942721 35756 943162
rect 35820 943129 35848 943230
rect 35806 943120 35862 943129
rect 35806 943055 35862 943064
rect 35714 942712 35770 942721
rect 35714 942647 35770 942656
rect 32402 937408 32458 937417
rect 32402 937343 32458 937352
rect 36556 936601 36584 952206
rect 37922 952167 37978 952176
rect 36542 936592 36598 936601
rect 36542 936527 36598 936536
rect 37936 936193 37964 952167
rect 41786 951688 41842 951697
rect 41786 951623 41842 951632
rect 41800 941866 41828 951623
rect 41892 951522 41920 954366
rect 42248 954304 42300 954310
rect 42248 954246 42300 954252
rect 42260 953578 42288 954246
rect 42168 953550 42288 953578
rect 41970 951824 42026 951833
rect 41970 951759 42026 951768
rect 41880 951516 41932 951522
rect 41880 951458 41932 951464
rect 41984 949454 42012 951759
rect 41892 949426 42012 949454
rect 41892 942018 41920 949426
rect 41892 941990 42012 942018
rect 41878 941896 41934 941905
rect 41788 941860 41840 941866
rect 41878 941831 41934 941840
rect 41788 941802 41840 941808
rect 41786 941080 41842 941089
rect 41786 941015 41842 941024
rect 41694 940128 41750 940137
rect 41524 940086 41694 940114
rect 37922 936184 37978 936193
rect 37922 936119 37978 936128
rect 39946 933328 40002 933337
rect 39946 933263 40002 933272
rect 39960 932142 39988 933263
rect 39948 932136 40000 932142
rect 39948 932078 40000 932084
rect 40684 909492 40736 909498
rect 40684 909434 40736 909440
rect 8588 818380 8616 818516
rect 9048 818380 9076 818516
rect 9508 818380 9536 818516
rect 9968 818380 9996 818516
rect 10428 818380 10456 818516
rect 10888 818380 10916 818516
rect 11348 818380 11376 818516
rect 11808 818380 11836 818516
rect 12268 818380 12296 818516
rect 12728 818380 12756 818516
rect 13188 818380 13216 818516
rect 13648 818380 13676 818516
rect 14108 818380 14136 818516
rect 40696 816921 40724 909434
rect 41234 818000 41290 818009
rect 41234 817935 41290 817944
rect 41248 817426 41276 817935
rect 41328 817556 41380 817562
rect 41328 817498 41380 817504
rect 41236 817420 41288 817426
rect 41236 817362 41288 817368
rect 41340 817329 41368 817498
rect 41326 817320 41382 817329
rect 41326 817255 41382 817264
rect 40682 816912 40738 816921
rect 40682 816847 40738 816856
rect 41524 814910 41552 940086
rect 41694 940063 41750 940072
rect 41694 939312 41750 939321
rect 41616 939270 41694 939298
rect 41616 823874 41644 939270
rect 41694 939247 41750 939256
rect 41800 923234 41828 941015
rect 41892 932894 41920 941831
rect 41984 937825 42012 941990
rect 42064 941860 42116 941866
rect 42064 941802 42116 941808
rect 41970 937816 42026 937825
rect 41970 937751 42026 937760
rect 42076 935377 42104 941802
rect 42168 939049 42196 953550
rect 42352 952270 42380 955454
rect 42720 954310 42748 955538
rect 42708 954304 42760 954310
rect 42708 954246 42760 954252
rect 42340 952264 42392 952270
rect 42340 952206 42392 952212
rect 42154 939040 42210 939049
rect 42154 938975 42210 938984
rect 42062 935368 42118 935377
rect 42062 935303 42118 935312
rect 42812 933745 42840 963970
rect 42892 962872 42944 962878
rect 42892 962814 42944 962820
rect 42904 934153 42932 962814
rect 44180 959744 44232 959750
rect 44180 959686 44232 959692
rect 42984 959132 43036 959138
rect 42984 959074 43036 959080
rect 42996 935785 43024 959074
rect 42982 935776 43038 935785
rect 42982 935711 43038 935720
rect 44192 934561 44220 959686
rect 44836 941497 44864 991442
rect 44822 941488 44878 941497
rect 44822 941423 44878 941432
rect 47596 940681 47624 991510
rect 47676 961920 47728 961926
rect 47676 961862 47728 961868
rect 47688 943226 47716 961862
rect 48412 943288 48464 943294
rect 48412 943230 48464 943236
rect 47676 943220 47728 943226
rect 47676 943162 47728 943168
rect 47582 940672 47638 940681
rect 47582 940607 47638 940616
rect 48424 937038 48452 943230
rect 48976 942313 49004 992870
rect 50344 990140 50396 990146
rect 50344 990082 50396 990088
rect 48962 942304 49018 942313
rect 48962 942239 49018 942248
rect 50356 939865 50384 990082
rect 89628 986060 89680 986066
rect 89628 986002 89680 986008
rect 73436 985992 73488 985998
rect 73436 985934 73488 985940
rect 73448 983620 73476 985934
rect 89640 983620 89668 986002
rect 102796 985998 102824 1006062
rect 103150 1006023 103152 1006032
rect 103204 1006023 103206 1006032
rect 108854 1006088 108856 1006097
rect 108908 1006088 108910 1006097
rect 108854 1006023 108910 1006032
rect 103152 1005994 103204 1006000
rect 103150 1004728 103206 1004737
rect 103150 1004663 103152 1004672
rect 103204 1004663 103206 1004672
rect 103152 1004634 103204 1004640
rect 106830 1002416 106886 1002425
rect 106830 1002351 106832 1002360
rect 106884 1002351 106886 1002360
rect 109868 1002380 109920 1002386
rect 106832 1002322 106884 1002328
rect 109868 1002322 109920 1002328
rect 106188 1002312 106240 1002318
rect 106002 1002280 106058 1002289
rect 108488 1002312 108540 1002318
rect 106188 1002254 106240 1002260
rect 108486 1002280 108488 1002289
rect 108540 1002280 108542 1002289
rect 106002 1002215 106004 1002224
rect 106056 1002215 106058 1002224
rect 106004 1002186 106056 1002192
rect 105636 1002176 105688 1002182
rect 105634 1002144 105636 1002153
rect 105688 1002144 105690 1002153
rect 105634 1002079 105690 1002088
rect 104348 1002040 104400 1002046
rect 104346 1002008 104348 1002017
rect 104400 1002008 104402 1002017
rect 104346 1001943 104402 1001952
rect 102784 985992 102836 985998
rect 102784 985934 102836 985940
rect 106200 983634 106228 1002254
rect 108304 1002244 108356 1002250
rect 108486 1002215 108542 1002224
rect 108304 1002186 108356 1002192
rect 107936 1002176 107988 1002182
rect 107658 1002144 107714 1002153
rect 108028 1002176 108080 1002182
rect 107936 1002118 107988 1002124
rect 108026 1002144 108028 1002153
rect 108080 1002144 108082 1002153
rect 107658 1002079 107660 1002088
rect 107712 1002079 107714 1002088
rect 107660 1002050 107712 1002056
rect 106648 1002040 106700 1002046
rect 106462 1002008 106518 1002017
rect 107200 1002040 107252 1002046
rect 106648 1001982 106700 1001988
rect 107198 1002008 107200 1002017
rect 107252 1002008 107254 1002017
rect 106462 1001943 106464 1001952
rect 106516 1001943 106518 1001952
rect 106464 1001914 106516 1001920
rect 106660 995110 106688 1001982
rect 107198 1001943 107254 1001952
rect 107752 1001972 107804 1001978
rect 107752 1001914 107804 1001920
rect 106648 995104 106700 995110
rect 106648 995046 106700 995052
rect 107764 991574 107792 1001914
rect 107752 991568 107804 991574
rect 107752 991510 107804 991516
rect 107948 990146 107976 1002118
rect 108026 1002079 108082 1002088
rect 108316 996130 108344 1002186
rect 109592 1002108 109644 1002114
rect 109592 1002050 109644 1002056
rect 109040 1002040 109092 1002046
rect 108486 1002008 108542 1002017
rect 109040 1001982 109092 1001988
rect 108486 1001943 108488 1001952
rect 108540 1001943 108542 1001952
rect 108488 1001914 108540 1001920
rect 108304 996124 108356 996130
rect 108304 996066 108356 996072
rect 109052 991506 109080 1001982
rect 109604 996062 109632 1002050
rect 109684 1002040 109736 1002046
rect 109682 1002008 109684 1002017
rect 109736 1002008 109738 1002017
rect 109682 1001943 109738 1001952
rect 109880 997762 109908 1002322
rect 110512 1002176 110564 1002182
rect 110512 1002118 110564 1002124
rect 109868 997756 109920 997762
rect 109868 997698 109920 997704
rect 109592 996056 109644 996062
rect 109592 995998 109644 996004
rect 110524 992934 110552 1002118
rect 111800 1002040 111852 1002046
rect 111800 1001982 111852 1001988
rect 111064 1001972 111116 1001978
rect 111064 1001914 111116 1001920
rect 111076 997694 111104 1001914
rect 111064 997688 111116 997694
rect 111064 997630 111116 997636
rect 110512 992928 110564 992934
rect 110512 992870 110564 992876
rect 109040 991500 109092 991506
rect 109040 991442 109092 991448
rect 107936 990140 107988 990146
rect 107936 990082 107988 990088
rect 111812 986066 111840 1001982
rect 117228 997756 117280 997762
rect 117228 997698 117280 997704
rect 116308 997688 116360 997694
rect 116308 997630 116360 997636
rect 116320 996985 116348 997630
rect 117240 997121 117268 997698
rect 117226 997112 117282 997121
rect 117226 997047 117282 997056
rect 116306 996976 116362 996985
rect 116306 996911 116362 996920
rect 121736 995036 121788 995042
rect 121736 994978 121788 994984
rect 111800 986060 111852 986066
rect 111800 986002 111852 986008
rect 105846 983606 106228 983634
rect 121748 983634 121776 994978
rect 126256 984638 126284 1006334
rect 146944 1006324 146996 1006330
rect 149702 1006295 149758 1006304
rect 150898 1006360 150900 1006369
rect 150952 1006360 150954 1006369
rect 150898 1006295 150954 1006304
rect 154118 1006360 154174 1006369
rect 154118 1006295 154120 1006304
rect 146944 1006266 146996 1006272
rect 154172 1006295 154174 1006304
rect 177304 1006324 177356 1006330
rect 154120 1006266 154172 1006272
rect 177304 1006266 177356 1006272
rect 195152 1006324 195204 1006330
rect 195152 1006266 195204 1006272
rect 145564 1006256 145616 1006262
rect 145564 1006198 145616 1006204
rect 144184 1006052 144236 1006058
rect 144184 1005994 144236 1006000
rect 143724 1005440 143776 1005446
rect 143724 1005382 143776 1005388
rect 143736 995858 143764 1005382
rect 144092 1002584 144144 1002590
rect 144092 1002526 144144 1002532
rect 143816 999796 143868 999802
rect 143816 999738 143868 999744
rect 139216 995852 139268 995858
rect 139216 995794 139268 995800
rect 140504 995852 140556 995858
rect 140504 995794 140556 995800
rect 143724 995852 143776 995858
rect 143724 995794 143776 995800
rect 131762 995752 131818 995761
rect 131606 995710 131762 995738
rect 133050 995752 133106 995761
rect 132802 995710 133050 995738
rect 131762 995687 131818 995696
rect 137926 995752 137982 995761
rect 135930 995722 136312 995738
rect 135930 995716 136324 995722
rect 135930 995710 136272 995716
rect 133050 995687 133106 995696
rect 137770 995710 137926 995738
rect 139228 995738 139256 995794
rect 140516 995738 140544 995794
rect 143828 995790 143856 999738
rect 144000 997348 144052 997354
rect 144000 997290 144052 997296
rect 141056 995784 141108 995790
rect 138966 995710 139256 995738
rect 140162 995710 140544 995738
rect 140806 995732 141056 995738
rect 143816 995784 143868 995790
rect 142894 995752 142950 995761
rect 140806 995726 141108 995732
rect 140806 995710 141096 995726
rect 142646 995710 142894 995738
rect 137926 995687 137982 995696
rect 143816 995726 143868 995732
rect 142894 995687 142950 995696
rect 136272 995658 136324 995664
rect 144012 995489 144040 997290
rect 144104 995722 144132 1002526
rect 144092 995716 144144 995722
rect 144092 995658 144144 995664
rect 144196 995625 144224 1005994
rect 144828 997688 144880 997694
rect 144828 997630 144880 997636
rect 144736 997620 144788 997626
rect 144736 997562 144788 997568
rect 144748 996985 144776 997562
rect 144840 997121 144868 997630
rect 144826 997112 144882 997121
rect 144826 997047 144882 997056
rect 144734 996976 144790 996985
rect 144734 996911 144790 996920
rect 144182 995616 144238 995625
rect 144182 995551 144238 995560
rect 137374 995480 137430 995489
rect 128464 995081 128492 995452
rect 129108 995178 129136 995452
rect 129096 995172 129148 995178
rect 129096 995114 129148 995120
rect 129752 995110 129780 995452
rect 132144 995217 132172 995452
rect 133432 995314 133460 995452
rect 136468 995353 136496 995452
rect 137126 995438 137374 995466
rect 137374 995415 137430 995424
rect 143998 995480 144054 995489
rect 143998 995415 144054 995424
rect 136454 995344 136510 995353
rect 133420 995308 133472 995314
rect 145576 995314 145604 1006198
rect 146956 995761 146984 1006266
rect 151728 1006256 151780 1006262
rect 151726 1006224 151728 1006233
rect 151780 1006224 151782 1006233
rect 147036 1006188 147088 1006194
rect 151726 1006159 151782 1006168
rect 152094 1006224 152150 1006233
rect 152094 1006159 152096 1006168
rect 147036 1006130 147088 1006136
rect 152148 1006159 152150 1006168
rect 152096 1006130 152148 1006136
rect 147048 997354 147076 1006130
rect 154488 1006120 154540 1006126
rect 150898 1006088 150954 1006097
rect 160652 1006120 160704 1006126
rect 154488 1006062 154540 1006068
rect 159086 1006088 159142 1006097
rect 150898 1006023 150900 1006032
rect 150952 1006023 150954 1006032
rect 150900 1005994 150952 1006000
rect 152740 1000544 152792 1000550
rect 152740 1000486 152792 1000492
rect 149060 998096 149112 998102
rect 149060 998038 149112 998044
rect 151266 998064 151322 998073
rect 148324 998028 148376 998034
rect 148324 997970 148376 997976
rect 147036 997348 147088 997354
rect 147036 997290 147088 997296
rect 146942 995752 146998 995761
rect 146942 995687 146998 995696
rect 148336 995353 148364 997970
rect 148874 996296 148930 996305
rect 149072 996282 149100 998038
rect 151266 997999 151268 998008
rect 151320 997999 151322 998008
rect 151268 997970 151320 997976
rect 151084 997960 151136 997966
rect 151084 997902 151136 997908
rect 152554 997928 152610 997937
rect 150348 997892 150400 997898
rect 150348 997834 150400 997840
rect 148930 996254 149100 996282
rect 148874 996231 148930 996240
rect 150360 995926 150388 997834
rect 150348 995920 150400 995926
rect 150348 995862 150400 995868
rect 148322 995344 148378 995353
rect 136454 995279 136510 995288
rect 145564 995308 145616 995314
rect 133420 995250 133472 995256
rect 148322 995279 148378 995288
rect 145564 995250 145616 995256
rect 132130 995208 132186 995217
rect 151096 995178 151124 997902
rect 152554 997863 152556 997872
rect 152608 997863 152610 997872
rect 152556 997834 152608 997840
rect 151268 997824 151320 997830
rect 151268 997766 151320 997772
rect 151280 995217 151308 997766
rect 152752 995897 152780 1000486
rect 152924 998096 152976 998102
rect 152922 998064 152924 998073
rect 152976 998064 152978 998073
rect 152922 997999 152978 998008
rect 153752 997960 153804 997966
rect 153750 997928 153752 997937
rect 153804 997928 153806 997937
rect 153750 997863 153806 997872
rect 153384 997824 153436 997830
rect 153382 997792 153384 997801
rect 153436 997792 153438 997801
rect 153382 997727 153438 997736
rect 152738 995888 152794 995897
rect 152738 995823 152794 995832
rect 151266 995208 151322 995217
rect 132130 995143 132186 995152
rect 151084 995172 151136 995178
rect 151266 995143 151322 995152
rect 151084 995114 151136 995120
rect 129740 995104 129792 995110
rect 128450 995072 128506 995081
rect 129740 995046 129792 995052
rect 128450 995007 128506 995016
rect 138296 991500 138348 991506
rect 138296 991442 138348 991448
rect 126244 984632 126296 984638
rect 126244 984574 126296 984580
rect 121748 983606 122130 983634
rect 138308 983620 138336 991442
rect 154500 983620 154528 1006062
rect 159086 1006023 159088 1006032
rect 159140 1006023 159142 1006032
rect 160650 1006088 160652 1006097
rect 160704 1006088 160706 1006097
rect 160650 1006023 160706 1006032
rect 162124 1006052 162176 1006058
rect 159088 1005994 159140 1006000
rect 162124 1005994 162176 1006000
rect 159824 1004896 159876 1004902
rect 159454 1004864 159510 1004873
rect 159454 1004799 159456 1004808
rect 159508 1004799 159510 1004808
rect 159822 1004864 159824 1004873
rect 159876 1004864 159878 1004873
rect 159822 1004799 159878 1004808
rect 161480 1004828 161532 1004834
rect 159456 1004770 159508 1004776
rect 161480 1004770 161532 1004776
rect 160284 1004760 160336 1004766
rect 160282 1004728 160284 1004737
rect 160336 1004728 160338 1004737
rect 160282 1004663 160338 1004672
rect 160650 1004728 160706 1004737
rect 160650 1004663 160652 1004672
rect 160704 1004663 160706 1004672
rect 160652 1004634 160704 1004640
rect 154580 1002584 154632 1002590
rect 154578 1002552 154580 1002561
rect 154632 1002552 154634 1002561
rect 154578 1002487 154634 1002496
rect 158258 1002280 158314 1002289
rect 158258 1002215 158260 1002224
rect 158312 1002215 158314 1002224
rect 160744 1002244 160796 1002250
rect 158260 1002186 158312 1002192
rect 160744 1002186 160796 1002192
rect 157800 1002176 157852 1002182
rect 157430 1002144 157486 1002153
rect 157430 1002079 157432 1002088
rect 157484 1002079 157486 1002088
rect 157798 1002144 157800 1002153
rect 160192 1002176 160244 1002182
rect 157852 1002144 157854 1002153
rect 160192 1002118 160244 1002124
rect 157798 1002079 157854 1002088
rect 159364 1002108 159416 1002114
rect 157432 1002050 157484 1002056
rect 159364 1002050 159416 1002056
rect 158628 1002040 158680 1002046
rect 156970 1002008 157026 1002017
rect 156970 1001943 156972 1001952
rect 157024 1001943 157026 1001952
rect 158626 1002008 158628 1002017
rect 158680 1002008 158682 1002017
rect 158626 1001943 158682 1001952
rect 158720 1001972 158772 1001978
rect 156972 1001914 157024 1001920
rect 158720 1001914 158772 1001920
rect 154946 1000648 155002 1000657
rect 154946 1000583 155002 1000592
rect 154960 1000550 154988 1000583
rect 154948 1000544 155000 1000550
rect 154948 1000486 155000 1000492
rect 155774 999832 155830 999841
rect 155774 999767 155776 999776
rect 155828 999767 155830 999776
rect 155776 999738 155828 999744
rect 156142 997792 156198 997801
rect 155236 997750 156142 997778
rect 155236 995110 155264 997750
rect 156142 997727 156198 997736
rect 158732 996130 158760 1001914
rect 159376 996198 159404 1002050
rect 160100 1002040 160152 1002046
rect 160100 1001982 160152 1001988
rect 159364 996192 159416 996198
rect 159364 996134 159416 996140
rect 158720 996124 158772 996130
rect 158720 996066 158772 996072
rect 160112 996062 160140 1001982
rect 160204 997694 160232 1002118
rect 160756 997762 160784 1002186
rect 160744 997756 160796 997762
rect 160744 997698 160796 997704
rect 160192 997688 160244 997694
rect 160192 997630 160244 997636
rect 161492 997626 161520 1004770
rect 161480 997620 161532 997626
rect 161480 997562 161532 997568
rect 162136 996130 162164 1005994
rect 169024 1005440 169076 1005446
rect 169024 1005382 169076 1005388
rect 162308 1004896 162360 1004902
rect 162308 1004838 162360 1004844
rect 162320 997694 162348 1004838
rect 163504 1004760 163556 1004766
rect 163504 1004702 163556 1004708
rect 162952 1004692 163004 1004698
rect 162952 1004634 163004 1004640
rect 162308 997688 162360 997694
rect 162308 997630 162360 997636
rect 162124 996124 162176 996130
rect 162124 996066 162176 996072
rect 160100 996056 160152 996062
rect 160100 995998 160152 996004
rect 155224 995104 155276 995110
rect 155224 995046 155276 995052
rect 162964 991506 162992 1004634
rect 162952 991500 163004 991506
rect 162952 991442 163004 991448
rect 163516 985930 163544 1004702
rect 167552 997756 167604 997762
rect 167552 997698 167604 997704
rect 167564 996985 167592 997698
rect 167644 997688 167696 997694
rect 167644 997630 167696 997636
rect 167656 997257 167684 997630
rect 167642 997248 167698 997257
rect 167642 997183 167698 997192
rect 167550 996976 167606 996985
rect 167550 996911 167606 996920
rect 169036 995654 169064 1005382
rect 169024 995648 169076 995654
rect 169024 995590 169076 995596
rect 163504 985924 163556 985930
rect 163504 985866 163556 985872
rect 170772 985924 170824 985930
rect 170772 985866 170824 985872
rect 170784 983620 170812 985866
rect 177316 984706 177344 1006266
rect 195164 1002130 195192 1006266
rect 195072 1002102 195192 1002130
rect 192484 995852 192536 995858
rect 192484 995794 192536 995800
rect 190460 995784 190512 995790
rect 184938 995752 184994 995761
rect 184828 995710 184938 995738
rect 188802 995752 188858 995761
rect 188508 995710 188802 995738
rect 184938 995687 184994 995696
rect 189446 995752 189502 995761
rect 189152 995710 189446 995738
rect 188802 995687 188858 995696
rect 190348 995732 190460 995738
rect 192496 995738 192524 995794
rect 195072 995761 195100 1002102
rect 195152 1001972 195204 1001978
rect 195152 1001914 195204 1001920
rect 195164 995858 195192 1001914
rect 195244 997756 195296 997762
rect 195244 997698 195296 997704
rect 195256 996985 195284 997698
rect 195242 996976 195298 996985
rect 195242 996911 195298 996920
rect 195244 996872 195296 996878
rect 195244 996814 195296 996820
rect 195256 995897 195284 996814
rect 195242 995888 195298 995897
rect 195152 995852 195204 995858
rect 195242 995823 195298 995832
rect 195152 995794 195204 995800
rect 195348 995790 195376 1007082
rect 249064 1006528 249116 1006534
rect 258172 1006528 258224 1006534
rect 249064 1006470 249116 1006476
rect 258170 1006496 258172 1006505
rect 302884 1006528 302936 1006534
rect 258224 1006496 258226 1006505
rect 201868 1006392 201920 1006398
rect 228364 1006392 228416 1006398
rect 201868 1006334 201920 1006340
rect 202694 1006360 202750 1006369
rect 196624 1006256 196676 1006262
rect 196624 1006198 196676 1006204
rect 195428 1001224 195480 1001230
rect 195428 1001166 195480 1001172
rect 195440 996033 195468 1001166
rect 195980 996804 196032 996810
rect 195980 996746 196032 996752
rect 195426 996024 195482 996033
rect 195426 995959 195482 995968
rect 195336 995784 195388 995790
rect 190348 995726 190512 995732
rect 190348 995710 190500 995726
rect 192188 995710 192524 995738
rect 195058 995752 195114 995761
rect 189446 995687 189502 995696
rect 195336 995726 195388 995732
rect 195058 995687 195114 995696
rect 184296 995648 184348 995654
rect 188158 995616 188214 995625
rect 184296 995590 184348 995596
rect 183834 995480 183890 995489
rect 179846 995353 179874 995452
rect 180504 995438 180748 995466
rect 181148 995438 181484 995466
rect 179832 995344 179888 995353
rect 179832 995279 179888 995288
rect 180720 995042 180748 995438
rect 181456 995110 181484 995438
rect 182974 995217 183002 995452
rect 183540 995438 183834 995466
rect 183834 995415 183890 995424
rect 184170 995246 184198 995452
rect 184158 995240 184210 995246
rect 182960 995208 183016 995217
rect 184158 995182 184210 995188
rect 182960 995143 183016 995152
rect 181444 995104 181496 995110
rect 181444 995046 181496 995052
rect 180708 995036 180760 995042
rect 180708 994978 180760 994984
rect 184308 990894 184336 995590
rect 187864 995574 188158 995602
rect 194322 995616 194378 995625
rect 194028 995574 194322 995602
rect 188158 995551 188214 995560
rect 194322 995551 194378 995560
rect 195992 995489 196020 996746
rect 195978 995480 196034 995489
rect 187312 995438 187648 995466
rect 191544 995438 191788 995466
rect 187620 995178 187648 995438
rect 187608 995172 187660 995178
rect 187608 995114 187660 995120
rect 191760 995081 191788 995438
rect 195978 995415 196034 995424
rect 196636 995246 196664 1006198
rect 197360 1006188 197412 1006194
rect 197360 1006130 197412 1006136
rect 197372 1001978 197400 1006130
rect 201880 1006126 201908 1006334
rect 210054 1006360 210110 1006369
rect 202694 1006295 202696 1006304
rect 202748 1006295 202750 1006304
rect 207664 1006324 207716 1006330
rect 202696 1006266 202748 1006272
rect 228364 1006334 228416 1006340
rect 248328 1006392 248380 1006398
rect 248328 1006334 248380 1006340
rect 210054 1006295 210056 1006304
rect 207664 1006266 207716 1006272
rect 210108 1006295 210110 1006304
rect 210056 1006266 210108 1006272
rect 204352 1006256 204404 1006262
rect 204350 1006224 204352 1006233
rect 204404 1006224 204406 1006233
rect 204350 1006159 204406 1006168
rect 204996 1006188 205048 1006194
rect 204996 1006130 205048 1006136
rect 198004 1006120 198056 1006126
rect 201040 1006120 201092 1006126
rect 198004 1006062 198056 1006068
rect 201038 1006088 201040 1006097
rect 201868 1006120 201920 1006126
rect 201092 1006088 201094 1006097
rect 197360 1001972 197412 1001978
rect 197360 1001914 197412 1001920
rect 196624 995240 196676 995246
rect 196624 995182 196676 995188
rect 198016 995110 198044 1006062
rect 201038 1006023 201094 1006032
rect 201866 1006088 201868 1006097
rect 201920 1006088 201922 1006097
rect 201866 1006023 201922 1006032
rect 202234 1004728 202290 1004737
rect 199384 1004692 199436 1004698
rect 202234 1004663 202236 1004672
rect 199384 1004634 199436 1004640
rect 202288 1004663 202290 1004672
rect 202236 1004634 202288 1004640
rect 199396 996878 199424 1004634
rect 202144 1002244 202196 1002250
rect 202144 1002186 202196 1002192
rect 200948 1002176 201000 1002182
rect 200948 1002118 201000 1002124
rect 200304 1002040 200356 1002046
rect 200304 1001982 200356 1001988
rect 200212 997280 200264 997286
rect 200210 997248 200212 997257
rect 200264 997248 200266 997257
rect 200210 997183 200266 997192
rect 199384 996872 199436 996878
rect 199384 996814 199436 996820
rect 200210 996296 200266 996305
rect 200316 996282 200344 1001982
rect 200960 1001230 200988 1002118
rect 200948 1001224 201000 1001230
rect 200948 1001166 201000 1001172
rect 201408 997688 201460 997694
rect 201408 997630 201460 997636
rect 200266 996254 200344 996282
rect 200210 996231 200266 996240
rect 201420 995178 201448 997630
rect 202052 997348 202104 997354
rect 202052 997290 202104 997296
rect 202064 995353 202092 997290
rect 202050 995344 202106 995353
rect 202050 995279 202106 995288
rect 201408 995172 201460 995178
rect 201408 995114 201460 995120
rect 198004 995104 198056 995110
rect 191746 995072 191802 995081
rect 198004 995046 198056 995052
rect 202156 995042 202184 1002186
rect 203524 1002176 203576 1002182
rect 203522 1002144 203524 1002153
rect 203576 1002144 203578 1002153
rect 203522 1002079 203578 1002088
rect 203708 1002108 203760 1002114
rect 203708 1002050 203760 1002056
rect 203064 1002040 203116 1002046
rect 203062 1002008 203064 1002017
rect 203524 1002040 203576 1002046
rect 203116 1002008 203118 1002017
rect 202328 1001972 202380 1001978
rect 203524 1001982 203576 1001988
rect 203062 1001943 203118 1001952
rect 202328 1001914 202380 1001920
rect 202340 996810 202368 1001914
rect 202328 996804 202380 996810
rect 202328 996746 202380 996752
rect 203536 995625 203564 1001982
rect 203720 997694 203748 1002050
rect 204718 1002008 204774 1002017
rect 204718 1001943 204720 1001952
rect 204772 1001943 204774 1001952
rect 204904 1001972 204956 1001978
rect 204720 1001914 204772 1001920
rect 204904 1001914 204956 1001920
rect 203708 997688 203760 997694
rect 203708 997630 203760 997636
rect 204916 997354 204944 1001914
rect 204904 997348 204956 997354
rect 204904 997290 204956 997296
rect 205008 997286 205036 1006130
rect 207204 1006120 207256 1006126
rect 207202 1006088 207204 1006097
rect 207256 1006088 207258 1006097
rect 207202 1006023 207258 1006032
rect 207570 1006088 207626 1006097
rect 207570 1006023 207572 1006032
rect 207624 1006023 207626 1006032
rect 207572 1005994 207624 1006000
rect 205178 1002280 205234 1002289
rect 205178 1002215 205180 1002224
rect 205232 1002215 205234 1002224
rect 205180 1002186 205232 1002192
rect 205914 1002144 205970 1002153
rect 205914 1002079 205916 1002088
rect 205968 1002079 205970 1002088
rect 205916 1002050 205968 1002056
rect 205548 1002040 205600 1002046
rect 205546 1002008 205548 1002017
rect 205600 1002008 205602 1002017
rect 205546 1001943 205602 1001952
rect 206742 1002008 206798 1002017
rect 206742 1001943 206744 1001952
rect 206796 1001943 206798 1001952
rect 206744 1001914 206796 1001920
rect 204996 997280 205048 997286
rect 204996 997222 205048 997228
rect 207676 996130 207704 1006266
rect 210422 1006224 210478 1006233
rect 210422 1006159 210424 1006168
rect 210476 1006159 210478 1006168
rect 210424 1006130 210476 1006136
rect 209596 1006120 209648 1006126
rect 209594 1006088 209596 1006097
rect 209648 1006088 209650 1006097
rect 209594 1006023 209650 1006032
rect 208766 1004864 208822 1004873
rect 208766 1004799 208768 1004808
rect 208820 1004799 208822 1004808
rect 211804 1004828 211856 1004834
rect 208768 1004770 208820 1004776
rect 211804 1004770 211856 1004776
rect 209228 1004760 209280 1004766
rect 208398 1004728 208454 1004737
rect 208398 1004663 208400 1004672
rect 208452 1004663 208454 1004672
rect 209226 1004728 209228 1004737
rect 211160 1004760 211212 1004766
rect 209280 1004728 209282 1004737
rect 211160 1004702 211212 1004708
rect 209226 1004663 209282 1004672
rect 209780 1004692 209832 1004698
rect 208400 1004634 208452 1004640
rect 209780 1004634 209832 1004640
rect 209792 996198 209820 1004634
rect 210424 1002176 210476 1002182
rect 210422 1002144 210424 1002153
rect 210476 1002144 210478 1002153
rect 210422 1002079 210478 1002088
rect 211172 997762 211200 1004702
rect 211618 1002280 211674 1002289
rect 211618 1002215 211620 1002224
rect 211672 1002215 211674 1002224
rect 211620 1002186 211672 1002192
rect 211250 1002144 211306 1002153
rect 211250 1002079 211252 1002088
rect 211304 1002079 211306 1002088
rect 211252 1002050 211304 1002056
rect 211160 997756 211212 997762
rect 211160 997698 211212 997704
rect 209780 996192 209832 996198
rect 209780 996134 209832 996140
rect 211816 996130 211844 1004770
rect 215944 1002244 215996 1002250
rect 215944 1002186 215996 1002192
rect 213184 1002176 213236 1002182
rect 213184 1002118 213236 1002124
rect 212540 1002040 212592 1002046
rect 212078 1002008 212134 1002017
rect 212078 1001943 212080 1001952
rect 212132 1001943 212134 1001952
rect 212538 1002008 212540 1002017
rect 212592 1002008 212594 1002017
rect 212538 1001943 212594 1001952
rect 212080 1001914 212132 1001920
rect 207664 996124 207716 996130
rect 207664 996066 207716 996072
rect 211804 996124 211856 996130
rect 211804 996066 211856 996072
rect 213196 995926 213224 1002118
rect 213368 1002108 213420 1002114
rect 213368 1002050 213420 1002056
rect 213380 997762 213408 1002050
rect 214564 1002040 214616 1002046
rect 214564 1001982 214616 1001988
rect 213920 1001972 213972 1001978
rect 213920 1001914 213972 1001920
rect 213368 997756 213420 997762
rect 213368 997698 213420 997704
rect 213184 995920 213236 995926
rect 213184 995862 213236 995868
rect 203522 995616 203578 995625
rect 203522 995551 203578 995560
rect 191746 995007 191802 995016
rect 202144 995036 202196 995042
rect 202144 994978 202196 994984
rect 213932 991506 213960 1001914
rect 203156 991500 203208 991506
rect 203156 991442 203208 991448
rect 213920 991500 213972 991506
rect 213920 991442 213972 991448
rect 184296 990888 184348 990894
rect 184296 990830 184348 990836
rect 186964 990888 187016 990894
rect 186964 990830 187016 990836
rect 177304 984700 177356 984706
rect 177304 984642 177356 984648
rect 186976 983620 187004 990830
rect 203168 983620 203196 991442
rect 214576 991234 214604 1001982
rect 215298 995072 215354 995081
rect 215298 995007 215354 995016
rect 215312 992934 215340 995007
rect 215300 992928 215352 992934
rect 215300 992870 215352 992876
rect 214564 991228 214616 991234
rect 214564 991170 214616 991176
rect 215956 985998 215984 1002186
rect 218888 997756 218940 997762
rect 218888 997698 218940 997704
rect 218900 996985 218928 997698
rect 218886 996976 218942 996985
rect 218886 996911 218942 996920
rect 219440 991228 219492 991234
rect 219440 991170 219492 991176
rect 215944 985992 215996 985998
rect 215944 985934 215996 985940
rect 219452 983620 219480 991170
rect 228376 984774 228404 1006334
rect 247684 1006188 247736 1006194
rect 247684 1006130 247736 1006136
rect 228456 1006120 228508 1006126
rect 228456 1006062 228508 1006068
rect 228468 996062 228496 1006062
rect 247040 1000000 247092 1000006
rect 247040 999942 247092 999948
rect 246672 997960 246724 997966
rect 246672 997902 246724 997908
rect 246580 997756 246632 997762
rect 246580 997698 246632 997704
rect 246592 996985 246620 997698
rect 246578 996976 246634 996985
rect 246578 996911 246634 996920
rect 228456 996056 228508 996062
rect 228456 995998 228508 996004
rect 242072 995852 242124 995858
rect 242072 995794 242124 995800
rect 238574 995752 238630 995761
rect 234968 995722 235304 995738
rect 234968 995716 235316 995722
rect 234968 995710 235264 995716
rect 240230 995752 240286 995761
rect 238630 995710 238740 995738
rect 239936 995710 240230 995738
rect 238574 995687 238630 995696
rect 242084 995738 242112 995794
rect 246684 995790 246712 997902
rect 246764 997824 246816 997830
rect 246764 997766 246816 997772
rect 245568 995784 245620 995790
rect 243818 995752 243874 995761
rect 241776 995710 242112 995738
rect 243616 995710 243818 995738
rect 240230 995687 240286 995696
rect 245456 995732 245568 995738
rect 245456 995726 245620 995732
rect 246672 995784 246724 995790
rect 246672 995726 246724 995732
rect 245456 995710 245608 995726
rect 243818 995687 243874 995696
rect 235264 995658 235316 995664
rect 246776 995654 246804 997766
rect 247052 996305 247080 999942
rect 247132 999524 247184 999530
rect 247132 999466 247184 999472
rect 247038 996296 247094 996305
rect 247038 996231 247094 996240
rect 247144 995722 247172 999466
rect 247696 995858 247724 1006130
rect 248340 997393 248368 1006334
rect 248420 1006120 248472 1006126
rect 248420 1006062 248472 1006068
rect 248432 997966 248460 1006062
rect 248420 997960 248472 997966
rect 248420 997902 248472 997908
rect 248326 997384 248382 997393
rect 248326 997319 248382 997328
rect 247684 995852 247736 995858
rect 247684 995794 247736 995800
rect 247132 995716 247184 995722
rect 247132 995658 247184 995664
rect 240876 995648 240928 995654
rect 236550 995616 236606 995625
rect 236256 995574 236550 995602
rect 240580 995596 240876 995602
rect 240580 995590 240928 995596
rect 246764 995648 246816 995654
rect 246764 995590 246816 995596
rect 240580 995574 240916 995590
rect 236550 995551 236606 995560
rect 231288 995438 231624 995466
rect 231932 995438 232268 995466
rect 232576 995438 232912 995466
rect 231596 995178 231624 995438
rect 231584 995172 231636 995178
rect 231584 995114 231636 995120
rect 232240 995110 232268 995438
rect 232228 995104 232280 995110
rect 232884 995081 232912 995438
rect 234402 995217 234430 995452
rect 235598 995246 235626 995452
rect 239278 995314 239306 995452
rect 242972 995438 243308 995466
rect 239266 995308 239318 995314
rect 239266 995250 239318 995256
rect 235586 995240 235638 995246
rect 234388 995208 234444 995217
rect 235586 995182 235638 995188
rect 234388 995143 234444 995152
rect 232228 995046 232280 995052
rect 232870 995072 232926 995081
rect 243280 995042 243308 995438
rect 249076 995178 249104 1006470
rect 253296 1006460 253348 1006466
rect 308128 1006528 308180 1006534
rect 302884 1006470 302936 1006476
rect 307298 1006496 307354 1006505
rect 258170 1006431 258226 1006440
rect 301504 1006460 301556 1006466
rect 253296 1006402 253348 1006408
rect 301504 1006402 301556 1006408
rect 249156 1006256 249208 1006262
rect 249156 1006198 249208 1006204
rect 249168 997257 249196 1006198
rect 253308 1006097 253336 1006402
rect 254860 1006392 254912 1006398
rect 254858 1006360 254860 1006369
rect 254912 1006360 254914 1006369
rect 254858 1006295 254914 1006304
rect 280804 1006324 280856 1006330
rect 280804 1006266 280856 1006272
rect 298744 1006324 298796 1006330
rect 298744 1006266 298796 1006272
rect 257344 1006256 257396 1006262
rect 255318 1006224 255374 1006233
rect 255318 1006159 255320 1006168
rect 255372 1006159 255374 1006168
rect 257342 1006224 257344 1006233
rect 257396 1006224 257398 1006233
rect 257342 1006159 257398 1006168
rect 255320 1006130 255372 1006136
rect 254676 1006120 254728 1006126
rect 252466 1006088 252522 1006097
rect 252466 1006023 252468 1006032
rect 252520 1006023 252522 1006032
rect 253294 1006088 253350 1006097
rect 258540 1006120 258592 1006126
rect 254676 1006062 254728 1006068
rect 256974 1006088 257030 1006097
rect 253294 1006023 253296 1006032
rect 252468 1005994 252520 1006000
rect 253348 1006023 253350 1006032
rect 253296 1005994 253348 1006000
rect 254490 1002280 254546 1002289
rect 252468 1002244 252520 1002250
rect 254490 1002215 254492 1002224
rect 252468 1002186 252520 1002192
rect 254544 1002215 254546 1002224
rect 254492 1002186 254544 1002192
rect 251824 1001972 251876 1001978
rect 251824 1001914 251876 1001920
rect 249708 999184 249760 999190
rect 249708 999126 249760 999132
rect 249154 997248 249210 997257
rect 249154 997183 249210 997192
rect 249720 996441 249748 999126
rect 250720 999116 250772 999122
rect 250720 999058 250772 999064
rect 249706 996432 249762 996441
rect 249706 996367 249762 996376
rect 250732 995246 250760 999058
rect 251836 995314 251864 1001914
rect 252480 1000006 252508 1002186
rect 253756 1002176 253808 1002182
rect 253756 1002118 253808 1002124
rect 252468 1000000 252520 1000006
rect 252468 999942 252520 999948
rect 253768 999530 253796 1002118
rect 253848 1002108 253900 1002114
rect 253848 1002050 253900 1002056
rect 253756 999524 253808 999530
rect 253756 999466 253808 999472
rect 253860 999122 253888 1002050
rect 254122 1002008 254178 1002017
rect 254122 1001943 254124 1001952
rect 254176 1001943 254178 1001952
rect 254584 1001972 254636 1001978
rect 254124 1001914 254176 1001920
rect 254584 1001914 254636 1001920
rect 253848 999116 253900 999122
rect 253848 999058 253900 999064
rect 253664 997824 253716 997830
rect 253662 997792 253664 997801
rect 253716 997792 253718 997801
rect 253662 997727 253718 997736
rect 251824 995308 251876 995314
rect 251824 995250 251876 995256
rect 250720 995240 250772 995246
rect 250720 995182 250772 995188
rect 249064 995172 249116 995178
rect 249064 995114 249116 995120
rect 254596 995110 254624 1001914
rect 254688 999190 254716 1006062
rect 258538 1006088 258540 1006097
rect 258592 1006088 258594 1006097
rect 256974 1006023 256976 1006032
rect 257028 1006023 257030 1006032
rect 257344 1006052 257396 1006058
rect 256976 1005994 257028 1006000
rect 258538 1006023 258594 1006032
rect 258998 1006088 259054 1006097
rect 258998 1006023 259000 1006032
rect 257344 1005994 257396 1006000
rect 259052 1006023 259054 1006032
rect 261022 1006088 261078 1006097
rect 261022 1006023 261024 1006032
rect 259000 1005994 259052 1006000
rect 261076 1006023 261078 1006032
rect 269764 1006052 269816 1006058
rect 261024 1005994 261076 1006000
rect 269764 1005994 269816 1006000
rect 256148 1002176 256200 1002182
rect 255686 1002144 255742 1002153
rect 255686 1002079 255688 1002088
rect 255740 1002079 255742 1002088
rect 256146 1002144 256148 1002153
rect 256200 1002144 256202 1002153
rect 256146 1002079 256202 1002088
rect 255688 1002050 255740 1002056
rect 256514 1002008 256570 1002017
rect 256514 1001943 256516 1001952
rect 256568 1001943 256570 1001952
rect 256516 1001914 256568 1001920
rect 254676 999184 254728 999190
rect 254676 999126 254728 999132
rect 254584 995104 254636 995110
rect 257356 995081 257384 1005994
rect 261852 1002312 261904 1002318
rect 261482 1002280 261538 1002289
rect 261482 1002215 261484 1002224
rect 261536 1002215 261538 1002224
rect 261850 1002280 261852 1002289
rect 264244 1002312 264296 1002318
rect 261904 1002280 261906 1002289
rect 264244 1002254 264296 1002260
rect 261850 1002215 261906 1002224
rect 263600 1002244 263652 1002250
rect 261484 1002186 261536 1002192
rect 263600 1002186 263652 1002192
rect 260840 1002176 260892 1002182
rect 259826 1002144 259882 1002153
rect 261852 1002176 261904 1002182
rect 260840 1002118 260892 1002124
rect 261850 1002144 261852 1002153
rect 262680 1002176 262732 1002182
rect 261904 1002144 261906 1002153
rect 259826 1002079 259828 1002088
rect 259880 1002079 259882 1002088
rect 259828 1002050 259880 1002056
rect 260196 1002040 260248 1002046
rect 260194 1002008 260196 1002017
rect 260248 1002008 260250 1002017
rect 260194 1001943 260250 1001952
rect 260654 1002008 260710 1002017
rect 260654 1001943 260656 1001952
rect 260708 1001943 260710 1001952
rect 260656 1001914 260708 1001920
rect 260852 997762 260880 1002118
rect 261484 1002108 261536 1002114
rect 261850 1002079 261906 1002088
rect 262678 1002144 262680 1002153
rect 262732 1002144 262734 1002153
rect 262678 1002079 262734 1002088
rect 263506 1002144 263562 1002153
rect 263506 1002079 263508 1002088
rect 261484 1002050 261536 1002056
rect 263560 1002079 263562 1002088
rect 263508 1002050 263560 1002056
rect 260840 997756 260892 997762
rect 260840 997698 260892 997704
rect 261496 996130 261524 1002050
rect 262864 1002040 262916 1002046
rect 263048 1002040 263100 1002046
rect 262864 1001982 262916 1001988
rect 263046 1002008 263048 1002017
rect 263100 1002008 263102 1002017
rect 262220 1001972 262272 1001978
rect 262220 1001914 262272 1001920
rect 261484 996124 261536 996130
rect 261484 996066 261536 996072
rect 262232 996062 262260 1001914
rect 262876 996198 262904 1001982
rect 263046 1001943 263102 1001952
rect 262864 996192 262916 996198
rect 262864 996134 262916 996140
rect 262220 996056 262272 996062
rect 262220 995998 262272 996004
rect 263612 995926 263640 1002186
rect 263874 1002008 263930 1002017
rect 263874 1001943 263876 1001952
rect 263928 1001943 263930 1001952
rect 263876 1001914 263928 1001920
rect 264256 996130 264284 1002254
rect 265808 1002176 265860 1002182
rect 265808 1002118 265860 1002124
rect 265624 1002040 265676 1002046
rect 265624 1001982 265676 1001988
rect 264244 996124 264296 996130
rect 264244 996066 264296 996072
rect 263600 995920 263652 995926
rect 263600 995862 263652 995868
rect 254584 995046 254636 995052
rect 257342 995072 257398 995081
rect 232870 995007 232926 995016
rect 243268 995036 243320 995042
rect 257342 995007 257398 995016
rect 243268 994978 243320 994984
rect 265636 992934 265664 1001982
rect 265820 997762 265848 1002118
rect 267004 1002108 267056 1002114
rect 267004 1002050 267056 1002056
rect 265808 997756 265860 997762
rect 265808 997698 265860 997704
rect 251456 992928 251508 992934
rect 251456 992870 251508 992876
rect 265624 992928 265676 992934
rect 265624 992870 265676 992876
rect 235632 985992 235684 985998
rect 235632 985934 235684 985940
rect 228364 984768 228416 984774
rect 228364 984710 228416 984716
rect 235644 983620 235672 985934
rect 251468 983634 251496 992870
rect 267016 986678 267044 1002050
rect 267096 1001972 267148 1001978
rect 267096 1001914 267148 1001920
rect 267108 990894 267136 1001914
rect 269776 996062 269804 1005994
rect 270408 997756 270460 997762
rect 270408 997698 270460 997704
rect 270420 996985 270448 997698
rect 270406 996976 270462 996985
rect 270406 996911 270462 996920
rect 269764 996056 269816 996062
rect 269764 995998 269816 996004
rect 267096 990888 267148 990894
rect 267096 990830 267148 990836
rect 268752 990888 268804 990894
rect 268752 990830 268804 990836
rect 267004 986672 267056 986678
rect 267004 986614 267056 986620
rect 268108 986672 268160 986678
rect 268108 986614 268160 986620
rect 251468 983606 251850 983634
rect 268120 983620 268148 986614
rect 268764 985998 268792 990830
rect 268752 985992 268804 985998
rect 268752 985934 268804 985940
rect 280816 984842 280844 1006266
rect 298376 1001904 298428 1001910
rect 298756 1001894 298784 1006266
rect 300308 1006256 300360 1006262
rect 300308 1006198 300360 1006204
rect 298836 1006052 298888 1006058
rect 298836 1005994 298888 1006000
rect 298376 1001846 298428 1001852
rect 298664 1001866 298784 1001894
rect 298284 997892 298336 997898
rect 298284 997834 298336 997840
rect 298190 997792 298246 997801
rect 298060 997750 298190 997778
rect 290648 995852 290700 995858
rect 290648 995794 290700 995800
rect 291108 995852 291160 995858
rect 291108 995794 291160 995800
rect 292488 995852 292540 995858
rect 292488 995794 292540 995800
rect 290660 995738 290688 995794
rect 291120 995738 291148 995794
rect 292500 995738 292528 995794
rect 298060 995790 298088 997750
rect 298190 997727 298246 997736
rect 297272 995784 297324 995790
rect 293498 995752 293554 995761
rect 290306 995710 290688 995738
rect 290858 995710 291148 995738
rect 292146 995710 292528 995738
rect 293342 995710 293498 995738
rect 294538 995722 294920 995738
rect 297022 995732 297272 995738
rect 297022 995726 297324 995732
rect 298048 995784 298100 995790
rect 298048 995726 298100 995732
rect 294538 995716 294932 995722
rect 294538 995710 294880 995716
rect 293498 995687 293554 995696
rect 297022 995710 297312 995726
rect 298296 995722 298324 997834
rect 298284 995716 298336 995722
rect 294880 995658 294932 995664
rect 298284 995658 298336 995664
rect 298388 995654 298416 1001846
rect 298560 1000544 298612 1000550
rect 298560 1000486 298612 1000492
rect 298466 998200 298522 998209
rect 298466 998135 298522 998144
rect 298480 995926 298508 998135
rect 298468 995920 298520 995926
rect 298468 995862 298520 995868
rect 295432 995648 295484 995654
rect 291750 995616 291806 995625
rect 291502 995574 291750 995602
rect 295182 995596 295432 995602
rect 295182 995590 295484 995596
rect 298376 995648 298428 995654
rect 298572 995625 298600 1000486
rect 298376 995590 298428 995596
rect 298558 995616 298614 995625
rect 295182 995574 295472 995590
rect 291750 995551 291806 995560
rect 298558 995551 298614 995560
rect 288072 995512 288124 995518
rect 282840 995110 282868 995452
rect 283484 995178 283512 995452
rect 284128 995246 284156 995452
rect 284116 995240 284168 995246
rect 284116 995182 284168 995188
rect 283472 995172 283524 995178
rect 283472 995114 283524 995120
rect 282828 995104 282880 995110
rect 285968 995081 285996 995452
rect 286534 995450 286824 995466
rect 286534 995444 286836 995450
rect 286534 995438 286784 995444
rect 287178 995438 287560 995466
rect 287822 995460 288072 995466
rect 287822 995454 288124 995460
rect 287822 995438 288112 995454
rect 286784 995386 286836 995392
rect 287532 995382 287560 995438
rect 287520 995376 287572 995382
rect 287520 995318 287572 995324
rect 298664 995246 298692 1001866
rect 298744 997756 298796 997762
rect 298744 997698 298796 997704
rect 298756 996985 298784 997698
rect 298742 996976 298798 996985
rect 298742 996911 298798 996920
rect 298848 995858 298876 1005994
rect 298928 1004624 298980 1004630
rect 298928 1004566 298980 1004572
rect 298940 995994 298968 1004566
rect 300124 1002040 300176 1002046
rect 300124 1001982 300176 1001988
rect 299388 1000612 299440 1000618
rect 299388 1000554 299440 1000560
rect 299296 996396 299348 996402
rect 299296 996338 299348 996344
rect 298928 995988 298980 995994
rect 298928 995930 298980 995936
rect 298836 995852 298888 995858
rect 298836 995794 298888 995800
rect 299308 995450 299336 996338
rect 299296 995444 299348 995450
rect 299296 995386 299348 995392
rect 298652 995240 298704 995246
rect 298652 995182 298704 995188
rect 299400 995178 299428 1000554
rect 300136 995518 300164 1001982
rect 300216 1001972 300268 1001978
rect 300216 1001914 300268 1001920
rect 300228 998209 300256 1001914
rect 300320 1000550 300348 1006198
rect 300308 1000544 300360 1000550
rect 300308 1000486 300360 1000492
rect 300214 998200 300270 998209
rect 300214 998135 300270 998144
rect 300124 995512 300176 995518
rect 300124 995454 300176 995460
rect 301516 995382 301544 1006402
rect 302896 1000618 302924 1006470
rect 307298 1006431 307300 1006440
rect 307352 1006431 307354 1006440
rect 308126 1006496 308128 1006505
rect 428372 1006528 428424 1006534
rect 308180 1006496 308182 1006505
rect 308126 1006431 308182 1006440
rect 358174 1006496 358230 1006505
rect 427542 1006496 427598 1006505
rect 358174 1006431 358176 1006440
rect 307300 1006402 307352 1006408
rect 358228 1006431 358230 1006440
rect 369124 1006460 369176 1006466
rect 358176 1006402 358228 1006408
rect 427542 1006431 427544 1006440
rect 369124 1006402 369176 1006408
rect 427596 1006431 427598 1006440
rect 428370 1006496 428372 1006505
rect 428424 1006496 428426 1006505
rect 428370 1006431 428426 1006440
rect 427544 1006402 427596 1006408
rect 356060 1006392 356112 1006398
rect 310610 1006360 310666 1006369
rect 310610 1006295 310612 1006304
rect 310664 1006295 310666 1006304
rect 356058 1006360 356060 1006369
rect 356112 1006360 356114 1006369
rect 356058 1006295 356114 1006304
rect 357714 1006360 357770 1006369
rect 357714 1006295 357716 1006304
rect 310612 1006266 310664 1006272
rect 357768 1006295 357770 1006304
rect 357716 1006266 357768 1006272
rect 306472 1006256 306524 1006262
rect 306470 1006224 306472 1006233
rect 358912 1006256 358964 1006262
rect 306524 1006224 306526 1006233
rect 306470 1006159 306526 1006168
rect 358910 1006224 358912 1006233
rect 358964 1006224 358966 1006233
rect 358910 1006159 358966 1006168
rect 369136 1006126 369164 1006402
rect 380164 1006392 380216 1006398
rect 504548 1006392 504600 1006398
rect 380164 1006334 380216 1006340
rect 504546 1006360 504548 1006369
rect 514208 1006392 514260 1006398
rect 504600 1006360 504602 1006369
rect 374644 1006324 374696 1006330
rect 374644 1006266 374696 1006272
rect 303528 1006120 303580 1006126
rect 304080 1006120 304132 1006126
rect 303528 1006062 303580 1006068
rect 304078 1006088 304080 1006097
rect 304908 1006120 304960 1006126
rect 304132 1006088 304134 1006097
rect 302884 1000612 302936 1000618
rect 302884 1000554 302936 1000560
rect 303252 997824 303304 997830
rect 303250 997792 303252 997801
rect 303304 997792 303306 997801
rect 303250 997727 303306 997736
rect 303252 996464 303304 996470
rect 303250 996432 303252 996441
rect 303304 996432 303306 996441
rect 303250 996367 303306 996376
rect 301504 995376 301556 995382
rect 301504 995318 301556 995324
rect 299388 995172 299440 995178
rect 299388 995114 299440 995120
rect 282828 995046 282880 995052
rect 285954 995072 286010 995081
rect 285954 995007 286010 995016
rect 300032 992928 300084 992934
rect 300032 992870 300084 992876
rect 284300 985992 284352 985998
rect 284300 985934 284352 985940
rect 280804 984836 280856 984842
rect 280804 984778 280856 984784
rect 284312 983620 284340 985934
rect 300044 983634 300072 992870
rect 303540 984910 303568 1006062
rect 304078 1006023 304134 1006032
rect 304906 1006088 304908 1006097
rect 356888 1006120 356940 1006126
rect 304960 1006088 304962 1006097
rect 304906 1006023 304962 1006032
rect 305274 1006088 305330 1006097
rect 305274 1006023 305276 1006032
rect 305328 1006023 305330 1006032
rect 315118 1006088 315174 1006097
rect 354494 1006088 354550 1006097
rect 315118 1006023 315120 1006032
rect 305276 1005994 305328 1006000
rect 315172 1006023 315174 1006032
rect 319444 1006052 319496 1006058
rect 315120 1005994 315172 1006000
rect 319444 1005994 319496 1006000
rect 353116 1006052 353168 1006058
rect 355230 1006088 355286 1006097
rect 354550 1006046 355230 1006074
rect 354494 1006023 354496 1006032
rect 353116 1005994 353168 1006000
rect 354548 1006023 354550 1006032
rect 355230 1006023 355286 1006032
rect 356886 1006088 356888 1006097
rect 360844 1006120 360896 1006126
rect 356940 1006088 356942 1006097
rect 356886 1006023 356942 1006032
rect 358542 1006088 358598 1006097
rect 361396 1006120 361448 1006126
rect 360844 1006062 360896 1006068
rect 361394 1006088 361396 1006097
rect 368480 1006120 368532 1006126
rect 361448 1006088 361450 1006097
rect 358542 1006023 358544 1006032
rect 354496 1005994 354548 1006000
rect 358596 1006023 358598 1006032
rect 358544 1005994 358596 1006000
rect 306930 1004864 306986 1004873
rect 304264 1004828 304316 1004834
rect 306930 1004799 306932 1004808
rect 304264 1004770 304316 1004776
rect 306984 1004799 306986 1004808
rect 313830 1004864 313886 1004873
rect 313830 1004799 313832 1004808
rect 306932 1004770 306984 1004776
rect 313884 1004799 313886 1004808
rect 316040 1004828 316092 1004834
rect 313832 1004770 313884 1004776
rect 316040 1004770 316092 1004776
rect 304276 996470 304304 1004770
rect 305828 1004760 305880 1004766
rect 308588 1004760 308640 1004766
rect 305828 1004702 305880 1004708
rect 307758 1004728 307814 1004737
rect 305644 1004692 305696 1004698
rect 305644 1004634 305696 1004640
rect 304264 996464 304316 996470
rect 304264 996406 304316 996412
rect 305656 996402 305684 1004634
rect 305734 1002008 305790 1002017
rect 305734 1001943 305736 1001952
rect 305788 1001943 305790 1001952
rect 305736 1001914 305788 1001920
rect 305840 997830 305868 1004702
rect 307758 1004663 307760 1004672
rect 307812 1004663 307814 1004672
rect 308586 1004728 308588 1004737
rect 314660 1004760 314712 1004766
rect 308640 1004728 308642 1004737
rect 308586 1004663 308642 1004672
rect 314658 1004728 314660 1004737
rect 314712 1004728 314714 1004737
rect 314658 1004663 314714 1004672
rect 315486 1004728 315542 1004737
rect 315486 1004663 315488 1004672
rect 307760 1004634 307812 1004640
rect 315540 1004663 315542 1004672
rect 315488 1004634 315540 1004640
rect 308956 1004624 309008 1004630
rect 308954 1004592 308956 1004601
rect 309008 1004592 309010 1004601
rect 308954 1004527 309010 1004536
rect 310150 1002144 310206 1002153
rect 310150 1002079 310152 1002088
rect 310204 1002079 310206 1002088
rect 311900 1002108 311952 1002114
rect 310152 1002050 310204 1002056
rect 311900 1002050 311952 1002056
rect 306104 1002040 306156 1002046
rect 306102 1002008 306104 1002017
rect 307024 1002040 307076 1002046
rect 306156 1002008 306158 1002017
rect 309324 1002040 309376 1002046
rect 307024 1001982 307076 1001988
rect 309322 1002008 309324 1002017
rect 309376 1002008 309378 1002017
rect 306102 1001943 306158 1001952
rect 305828 997824 305880 997830
rect 305828 997766 305880 997772
rect 305644 996396 305696 996402
rect 305644 996338 305696 996344
rect 307036 995081 307064 1001982
rect 309322 1001943 309378 1001952
rect 310150 1002008 310206 1002017
rect 310150 1001943 310206 1001952
rect 311438 1002008 311494 1002017
rect 311438 1001943 311440 1001952
rect 310164 1001910 310192 1001943
rect 311492 1001943 311494 1001952
rect 311440 1001914 311492 1001920
rect 310152 1001904 310204 1001910
rect 310152 1001846 310204 1001852
rect 311912 995110 311940 1002050
rect 312268 1002040 312320 1002046
rect 312266 1002008 312268 1002017
rect 314660 1002040 314712 1002046
rect 312320 1002008 312322 1002017
rect 312266 1001943 312322 1001952
rect 313002 1002008 313058 1002017
rect 313058 1001966 313412 1001994
rect 314660 1001982 314712 1001988
rect 313002 1001943 313058 1001952
rect 313384 996130 313412 1001966
rect 313556 1001972 313608 1001978
rect 313556 1001914 313608 1001920
rect 313568 996198 313596 1001914
rect 313556 996192 313608 996198
rect 313556 996134 313608 996140
rect 313372 996124 313424 996130
rect 313372 996066 313424 996072
rect 314672 996062 314700 1001982
rect 316052 997762 316080 1004770
rect 316684 1004760 316736 1004766
rect 316684 1004702 316736 1004708
rect 316040 997756 316092 997762
rect 316040 997698 316092 997704
rect 314660 996056 314712 996062
rect 314660 995998 314712 996004
rect 311900 995104 311952 995110
rect 307022 995072 307078 995081
rect 311900 995046 311952 995052
rect 307022 995007 307078 995016
rect 316408 995036 316460 995042
rect 316408 994978 316460 994984
rect 303528 984904 303580 984910
rect 303528 984846 303580 984852
rect 316420 983634 316448 994978
rect 316696 992934 316724 1004702
rect 318064 1004692 318116 1004698
rect 318064 1004634 318116 1004640
rect 316684 992928 316736 992934
rect 316684 992870 316736 992876
rect 318076 985998 318104 1004634
rect 319456 993002 319484 1005994
rect 328368 997824 328420 997830
rect 328368 997766 328420 997772
rect 328380 997082 328408 997766
rect 328368 997076 328420 997082
rect 328368 997018 328420 997024
rect 319444 992996 319496 993002
rect 319444 992938 319496 992944
rect 332600 992996 332652 993002
rect 332600 992938 332652 992944
rect 318064 985992 318116 985998
rect 318064 985934 318116 985940
rect 332612 983634 332640 992938
rect 353128 990146 353156 1005994
rect 354508 1005963 354536 1005994
rect 360566 1005408 360622 1005417
rect 360566 1005343 360568 1005352
rect 360620 1005343 360622 1005352
rect 360568 1005314 360620 1005320
rect 360200 1005304 360252 1005310
rect 360198 1005272 360200 1005281
rect 360252 1005272 360254 1005281
rect 360198 1005207 360254 1005216
rect 354312 1004760 354364 1004766
rect 356888 1004760 356940 1004766
rect 354312 1004702 354364 1004708
rect 356058 1004728 356114 1004737
rect 354324 995178 354352 1004702
rect 354588 1004692 354640 1004698
rect 356058 1004663 356060 1004672
rect 354588 1004634 354640 1004640
rect 356112 1004663 356114 1004672
rect 356886 1004728 356888 1004737
rect 356940 1004728 356942 1004737
rect 356886 1004663 356942 1004672
rect 356060 1004634 356112 1004640
rect 354600 1002590 354628 1004634
rect 354588 1002584 354640 1002590
rect 354588 1002526 354640 1002532
rect 359188 1002584 359240 1002590
rect 359188 1002526 359240 1002532
rect 357164 1002040 357216 1002046
rect 357164 1001982 357216 1001988
rect 358910 1002008 358966 1002017
rect 357176 999054 357204 1001982
rect 357348 1001972 357400 1001978
rect 358910 1001943 358912 1001952
rect 357348 1001914 357400 1001920
rect 358964 1001943 358966 1001952
rect 358912 1001914 358964 1001920
rect 357164 999048 357216 999054
rect 357164 998990 357216 998996
rect 354312 995172 354364 995178
rect 354312 995114 354364 995120
rect 357360 995042 357388 1001914
rect 359200 995314 359228 1002526
rect 359372 1002040 359424 1002046
rect 359370 1002008 359372 1002017
rect 359424 1002008 359426 1002017
rect 359370 1001943 359426 1001952
rect 360856 998442 360884 1006062
rect 368480 1006062 368532 1006068
rect 369124 1006120 369176 1006126
rect 369124 1006062 369176 1006068
rect 361394 1006023 361450 1006032
rect 362224 1006052 362276 1006058
rect 362224 1005994 362276 1006000
rect 361028 1005440 361080 1005446
rect 361026 1005408 361028 1005417
rect 361080 1005408 361082 1005417
rect 361026 1005343 361082 1005352
rect 361856 1004760 361908 1004766
rect 361854 1004728 361856 1004737
rect 361908 1004728 361910 1004737
rect 361854 1004663 361910 1004672
rect 361580 999048 361632 999054
rect 361580 998990 361632 998996
rect 360844 998436 360896 998442
rect 360844 998378 360896 998384
rect 361592 996062 361620 998990
rect 362236 997762 362264 1005994
rect 363420 1004896 363472 1004902
rect 363418 1004864 363420 1004873
rect 366364 1004896 366416 1004902
rect 363472 1004864 363474 1004873
rect 363418 1004799 363474 1004808
rect 364246 1004864 364302 1004873
rect 366364 1004838 366416 1004844
rect 364246 1004799 364248 1004808
rect 364300 1004799 364302 1004808
rect 364248 1004770 364300 1004776
rect 364984 1004760 365036 1004766
rect 362590 1004728 362646 1004737
rect 364984 1004702 365036 1004708
rect 362590 1004663 362592 1004672
rect 362644 1004663 362646 1004672
rect 362592 1004634 362644 1004640
rect 362224 997756 362276 997762
rect 362224 997698 362276 997704
rect 364996 996198 365024 1004702
rect 365168 1004692 365220 1004698
rect 365168 1004634 365220 1004640
rect 365074 1002144 365130 1002153
rect 365074 1002079 365076 1002088
rect 365128 1002079 365130 1002088
rect 365076 1002050 365128 1002056
rect 365180 997626 365208 1004634
rect 365904 1002040 365956 1002046
rect 365442 1002008 365498 1002017
rect 365442 1001943 365444 1001952
rect 365496 1001943 365498 1001952
rect 365902 1002008 365904 1002017
rect 365956 1002008 365958 1002017
rect 365902 1001943 365958 1001952
rect 365444 1001914 365496 1001920
rect 365168 997620 365220 997626
rect 365168 997562 365220 997568
rect 364984 996192 365036 996198
rect 364984 996134 365036 996140
rect 366376 996130 366404 1004838
rect 366548 1004828 366600 1004834
rect 366548 1004770 366600 1004776
rect 366560 997694 366588 1004770
rect 367928 1002108 367980 1002114
rect 367928 1002050 367980 1002056
rect 367744 1001972 367796 1001978
rect 367744 1001914 367796 1001920
rect 366548 997688 366600 997694
rect 366548 997630 366600 997636
rect 366364 996124 366416 996130
rect 366364 996066 366416 996072
rect 361580 996056 361632 996062
rect 361580 995998 361632 996004
rect 359188 995308 359240 995314
rect 359188 995250 359240 995256
rect 357348 995036 357400 995042
rect 357348 994978 357400 994984
rect 364984 992928 365036 992934
rect 364984 992870 365036 992876
rect 353116 990140 353168 990146
rect 353116 990082 353168 990088
rect 349160 985992 349212 985998
rect 349160 985934 349212 985940
rect 300044 983606 300518 983634
rect 316420 983606 316802 983634
rect 332612 983606 332994 983634
rect 349172 983620 349200 985934
rect 364996 983634 365024 992870
rect 367756 991506 367784 1001914
rect 367940 993002 367968 1002050
rect 368492 998510 368520 1006062
rect 371884 1005440 371936 1005446
rect 371884 1005382 371936 1005388
rect 369124 1002040 369176 1002046
rect 369124 1001982 369176 1001988
rect 368480 998504 368532 998510
rect 368480 998446 368532 998452
rect 367928 992996 367980 993002
rect 367928 992938 367980 992944
rect 367744 991500 367796 991506
rect 367744 991442 367796 991448
rect 369136 985998 369164 1001982
rect 371896 995110 371924 1005382
rect 372344 997756 372396 997762
rect 372344 997698 372396 997704
rect 372356 996441 372384 997698
rect 372436 997688 372488 997694
rect 372436 997630 372488 997636
rect 372448 997121 372476 997630
rect 372528 997620 372580 997626
rect 372528 997562 372580 997568
rect 372434 997112 372490 997121
rect 372434 997047 372490 997056
rect 372540 996985 372568 997562
rect 372526 996976 372582 996985
rect 372526 996911 372582 996920
rect 372342 996432 372398 996441
rect 372342 996367 372398 996376
rect 374656 995625 374684 1006266
rect 376024 1006256 376076 1006262
rect 376024 1006198 376076 1006204
rect 374642 995616 374698 995625
rect 374642 995551 374698 995560
rect 376036 995353 376064 1006198
rect 378784 1005372 378836 1005378
rect 378784 1005314 378836 1005320
rect 378796 997830 378824 1005314
rect 378784 997824 378836 997830
rect 378784 997766 378836 997772
rect 376022 995344 376078 995353
rect 376022 995279 376078 995288
rect 380176 995217 380204 1006334
rect 445760 1006324 445812 1006330
rect 514208 1006334 514260 1006340
rect 555974 1006360 556030 1006369
rect 504546 1006295 504602 1006304
rect 445760 1006266 445812 1006272
rect 425150 1006224 425206 1006233
rect 425150 1006159 425152 1006168
rect 425204 1006159 425206 1006168
rect 425152 1006130 425204 1006136
rect 380900 1006120 380952 1006126
rect 380900 1006062 380952 1006068
rect 420828 1006120 420880 1006126
rect 422668 1006120 422720 1006126
rect 420828 1006062 420880 1006068
rect 422666 1006088 422668 1006097
rect 428004 1006120 428056 1006126
rect 422720 1006088 422722 1006097
rect 380912 1003338 380940 1006062
rect 381544 1005304 381596 1005310
rect 381544 1005246 381596 1005252
rect 380900 1003332 380952 1003338
rect 380900 1003274 380952 1003280
rect 380900 998436 380952 998442
rect 380900 998378 380952 998384
rect 380912 995489 380940 998378
rect 381176 997076 381228 997082
rect 381176 997018 381228 997024
rect 380898 995480 380954 995489
rect 380898 995415 380954 995424
rect 380162 995208 380218 995217
rect 380162 995143 380218 995152
rect 371884 995104 371936 995110
rect 371884 995046 371936 995052
rect 369124 985992 369176 985998
rect 369124 985934 369176 985940
rect 381188 983634 381216 997018
rect 381556 995761 381584 1005246
rect 383568 1003332 383620 1003338
rect 383568 1003274 383620 1003280
rect 383384 998504 383436 998510
rect 383384 998446 383436 998452
rect 383396 995858 383424 998446
rect 383476 997824 383528 997830
rect 383476 997766 383528 997772
rect 383488 997098 383516 997766
rect 383580 997529 383608 1003274
rect 420840 1001978 420868 1006062
rect 422666 1006023 422722 1006032
rect 423494 1006088 423550 1006097
rect 428002 1006088 428004 1006097
rect 428056 1006088 428058 1006097
rect 423494 1006023 423496 1006032
rect 423548 1006023 423550 1006032
rect 426348 1006052 426400 1006058
rect 423496 1005994 423548 1006000
rect 428002 1006023 428058 1006032
rect 430026 1006088 430082 1006097
rect 430026 1006023 430028 1006032
rect 426348 1005994 426400 1006000
rect 430080 1006023 430082 1006032
rect 430028 1005994 430080 1006000
rect 426360 1005310 426388 1005994
rect 426348 1005304 426400 1005310
rect 426348 1005246 426400 1005252
rect 422024 1004624 422076 1004630
rect 423864 1004624 423916 1004630
rect 422024 1004566 422076 1004572
rect 423862 1004592 423864 1004601
rect 423916 1004592 423918 1004601
rect 421470 1002008 421526 1002017
rect 420828 1001972 420880 1001978
rect 421470 1001943 421472 1001952
rect 420828 1001914 420880 1001920
rect 421524 1001943 421526 1001952
rect 421472 1001914 421524 1001920
rect 399944 997756 399996 997762
rect 399944 997698 399996 997704
rect 383566 997520 383622 997529
rect 383566 997455 383622 997464
rect 383658 997384 383714 997393
rect 383714 997342 383772 997370
rect 383658 997319 383714 997328
rect 383488 997070 383680 997098
rect 383384 995852 383436 995858
rect 383384 995794 383436 995800
rect 383652 995790 383680 997070
rect 383640 995784 383692 995790
rect 381542 995752 381598 995761
rect 383640 995726 383692 995732
rect 383744 995722 383772 997342
rect 399956 997121 399984 997698
rect 400036 997688 400088 997694
rect 400036 997630 400088 997636
rect 399942 997112 399998 997121
rect 399942 997047 399998 997056
rect 400048 996985 400076 997630
rect 400034 996976 400090 996985
rect 400034 996911 400090 996920
rect 385684 995852 385736 995858
rect 385684 995794 385736 995800
rect 391756 995852 391808 995858
rect 391756 995794 391808 995800
rect 384396 995784 384448 995790
rect 385696 995738 385724 995794
rect 387890 995752 387946 995761
rect 384448 995732 384698 995738
rect 384396 995726 384698 995732
rect 381542 995687 381598 995696
rect 383732 995716 383784 995722
rect 384408 995710 384698 995726
rect 385696 995710 385986 995738
rect 387826 995710 387890 995738
rect 387890 995687 387946 995696
rect 388166 995752 388222 995761
rect 391768 995738 391796 995794
rect 396630 995752 396686 995761
rect 388222 995710 388378 995738
rect 388640 995722 389022 995738
rect 388628 995716 389022 995722
rect 388166 995687 388222 995696
rect 383732 995658 383784 995664
rect 388680 995710 389022 995716
rect 391768 995710 392150 995738
rect 396382 995710 396630 995738
rect 396630 995687 396686 995696
rect 388628 995658 388680 995664
rect 394882 995616 394938 995625
rect 394938 995574 395186 995602
rect 394882 995551 394938 995560
rect 389362 995480 389418 995489
rect 385328 995353 385356 995452
rect 389418 995438 389666 995466
rect 389362 995415 389418 995424
rect 385314 995344 385370 995353
rect 392688 995314 392716 995452
rect 393240 995438 393346 995466
rect 385314 995279 385370 995288
rect 392676 995308 392728 995314
rect 392676 995250 392728 995256
rect 393240 995178 393268 995438
rect 393976 995217 394004 995452
rect 393962 995208 394018 995217
rect 393228 995172 393280 995178
rect 393962 995143 394018 995152
rect 393228 995114 393280 995120
rect 397012 995110 397040 995452
rect 397000 995104 397052 995110
rect 397000 995046 397052 995052
rect 398852 995042 398880 995452
rect 398840 995036 398892 995042
rect 398840 994978 398892 994984
rect 420840 992934 420868 1001914
rect 422036 998442 422064 1004566
rect 423862 1004527 423918 1004536
rect 424692 1004080 424744 1004086
rect 424690 1004048 424692 1004057
rect 424744 1004048 424746 1004057
rect 424690 1003983 424746 1003992
rect 423496 1003944 423548 1003950
rect 423494 1003912 423496 1003921
rect 423548 1003912 423550 1003921
rect 423494 1003847 423550 1003856
rect 445772 1003270 445800 1006266
rect 456064 1006256 456116 1006262
rect 505376 1006256 505428 1006262
rect 456064 1006198 456116 1006204
rect 505006 1006224 505062 1006233
rect 449256 1006188 449308 1006194
rect 449256 1006130 449308 1006136
rect 445760 1003264 445812 1003270
rect 445760 1003206 445812 1003212
rect 425980 1002584 426032 1002590
rect 425978 1002552 425980 1002561
rect 426032 1002552 426034 1002561
rect 425978 1002487 426034 1002496
rect 425978 1002144 426034 1002153
rect 423312 1002108 423364 1002114
rect 425978 1002079 425980 1002088
rect 423312 1002050 423364 1002056
rect 426032 1002079 426034 1002088
rect 425980 1002050 426032 1002056
rect 423324 1001230 423352 1002050
rect 424968 1002040 425020 1002046
rect 426348 1002040 426400 1002046
rect 424968 1001982 425020 1001988
rect 425150 1002008 425206 1002017
rect 423404 1001972 423456 1001978
rect 423404 1001914 423456 1001920
rect 423312 1001224 423364 1001230
rect 423312 1001166 423364 1001172
rect 423416 998578 423444 1001914
rect 424980 1001298 425008 1001982
rect 426346 1002008 426348 1002017
rect 426400 1002008 426402 1002017
rect 425150 1001943 425152 1001952
rect 425204 1001943 425206 1001952
rect 425704 1001972 425756 1001978
rect 425152 1001914 425204 1001920
rect 426346 1001943 426402 1001952
rect 426806 1002008 426862 1002017
rect 426806 1001943 426808 1001952
rect 425704 1001914 425756 1001920
rect 426860 1001943 426862 1001952
rect 426808 1001914 426860 1001920
rect 424968 1001292 425020 1001298
rect 424968 1001234 425020 1001240
rect 423404 998572 423456 998578
rect 423404 998514 423456 998520
rect 425716 998510 425744 1001914
rect 449268 1001842 449296 1006130
rect 451280 1004080 451332 1004086
rect 451280 1004022 451332 1004028
rect 449808 1003264 449860 1003270
rect 449808 1003206 449860 1003212
rect 449256 1001836 449308 1001842
rect 449256 1001778 449308 1001784
rect 447140 1001292 447192 1001298
rect 447140 1001234 447192 1001240
rect 428830 999832 428886 999841
rect 428830 999767 428832 999776
rect 428884 999767 428886 999776
rect 428832 999738 428884 999744
rect 425704 998504 425756 998510
rect 425704 998446 425756 998452
rect 422024 998436 422076 998442
rect 422024 998378 422076 998384
rect 430854 998200 430910 998209
rect 430854 998135 430856 998144
rect 430908 998135 430910 998144
rect 433984 998164 434036 998170
rect 430856 998106 430908 998112
rect 433984 998106 434036 998112
rect 431684 998096 431736 998102
rect 429658 998064 429714 998073
rect 429658 997999 429660 998008
rect 429712 997999 429714 998008
rect 431682 998064 431684 998073
rect 431736 998064 431738 998073
rect 431682 997999 431738 998008
rect 431960 998028 432012 998034
rect 429660 997970 429712 997976
rect 431960 997970 432012 997976
rect 428464 997960 428516 997966
rect 430856 997960 430908 997966
rect 428464 997902 428516 997908
rect 430394 997928 430450 997937
rect 428476 996130 428504 997902
rect 430394 997863 430396 997872
rect 430448 997863 430450 997872
rect 430854 997928 430856 997937
rect 430908 997928 430910 997937
rect 430854 997863 430910 997872
rect 430396 997834 430448 997840
rect 429200 997824 429252 997830
rect 429198 997792 429200 997801
rect 431224 997824 431276 997830
rect 429252 997792 429254 997801
rect 431224 997766 431276 997772
rect 429198 997727 429254 997736
rect 431236 996130 431264 997766
rect 431972 996198 432000 997970
rect 432880 997960 432932 997966
rect 432418 997928 432474 997937
rect 432144 997892 432196 997898
rect 432418 997863 432420 997872
rect 432144 997834 432196 997840
rect 432472 997863 432474 997872
rect 432878 997928 432880 997937
rect 432932 997928 432934 997937
rect 432878 997863 432934 997872
rect 432420 997834 432472 997840
rect 432052 997824 432104 997830
rect 432050 997792 432052 997801
rect 432104 997792 432106 997801
rect 432050 997727 432106 997736
rect 432156 997694 432184 997834
rect 433340 997824 433392 997830
rect 433392 997772 433472 997778
rect 433340 997766 433472 997772
rect 433352 997762 433472 997766
rect 433352 997756 433484 997762
rect 433352 997750 433432 997756
rect 433432 997698 433484 997704
rect 432144 997688 432196 997694
rect 432144 997630 432196 997636
rect 433996 996198 434024 998106
rect 434168 998096 434220 998102
rect 434168 998038 434220 998044
rect 434180 997762 434208 998038
rect 436744 997960 436796 997966
rect 436744 997902 436796 997908
rect 435548 997892 435600 997898
rect 435548 997834 435600 997840
rect 435362 997792 435418 997801
rect 434168 997756 434220 997762
rect 435362 997727 435418 997736
rect 434168 997698 434220 997704
rect 431960 996192 432012 996198
rect 431960 996134 432012 996140
rect 433984 996192 434036 996198
rect 433984 996134 434036 996140
rect 428464 996124 428516 996130
rect 428464 996066 428516 996072
rect 431224 996124 431276 996130
rect 431224 996066 431276 996072
rect 432050 995888 432106 995897
rect 432050 995823 432106 995832
rect 432064 995790 432092 995823
rect 432052 995784 432104 995790
rect 432052 995726 432104 995732
rect 429936 992996 429988 993002
rect 429936 992938 429988 992944
rect 420828 992928 420880 992934
rect 420828 992870 420880 992876
rect 397828 991500 397880 991506
rect 397828 991442 397880 991448
rect 364996 983606 365470 983634
rect 381188 983606 381662 983634
rect 397840 983620 397868 991442
rect 414112 985992 414164 985998
rect 414112 985934 414164 985940
rect 414124 983620 414152 985934
rect 429948 983634 429976 992938
rect 435376 987426 435404 997727
rect 435560 991506 435588 997834
rect 435548 991500 435600 991506
rect 435548 991442 435600 991448
rect 435364 987420 435416 987426
rect 435364 987362 435416 987368
rect 436756 985998 436784 997902
rect 439688 997756 439740 997762
rect 439688 997698 439740 997704
rect 439700 996985 439728 997698
rect 439686 996976 439742 996985
rect 439686 996911 439742 996920
rect 439780 995784 439832 995790
rect 439778 995752 439780 995761
rect 439832 995752 439834 995761
rect 439778 995687 439834 995696
rect 447152 995042 447180 1001234
rect 449820 995081 449848 1003206
rect 451292 1000278 451320 1004022
rect 454316 1003944 454368 1003950
rect 454316 1003886 454368 1003892
rect 452568 1001836 452620 1001842
rect 452568 1001778 452620 1001784
rect 451280 1000272 451332 1000278
rect 451280 1000214 451332 1000220
rect 452580 998646 452608 1001778
rect 452568 998640 452620 998646
rect 452568 998582 452620 998588
rect 454328 995217 454356 1003886
rect 456076 995489 456104 1006198
rect 505006 1006159 505008 1006168
rect 505060 1006159 505062 1006168
rect 505374 1006224 505376 1006233
rect 514116 1006256 514168 1006262
rect 505428 1006224 505430 1006233
rect 514116 1006198 514168 1006204
rect 505374 1006159 505430 1006168
rect 505008 1006130 505060 1006136
rect 465724 1006120 465776 1006126
rect 502524 1006120 502576 1006126
rect 465724 1006062 465776 1006068
rect 499670 1006088 499726 1006097
rect 462964 1005304 463016 1005310
rect 462964 1005246 463016 1005252
rect 459560 1000272 459612 1000278
rect 459560 1000214 459612 1000220
rect 459572 998345 459600 1000214
rect 459652 998640 459704 998646
rect 459652 998582 459704 998588
rect 459558 998336 459614 998345
rect 459558 998271 459614 998280
rect 456062 995480 456118 995489
rect 456062 995415 456118 995424
rect 459664 995353 459692 998582
rect 462976 996305 463004 1005246
rect 465736 998442 465764 1006062
rect 468484 1006052 468536 1006058
rect 468484 1005994 468536 1006000
rect 498108 1006052 498160 1006058
rect 499670 1006023 499672 1006032
rect 498108 1005994 498160 1006000
rect 499724 1006023 499726 1006032
rect 500498 1006088 500554 1006097
rect 500498 1006023 500500 1006032
rect 499672 1005994 499724 1006000
rect 500552 1006023 500554 1006032
rect 502522 1006088 502524 1006097
rect 502576 1006088 502578 1006097
rect 502522 1006023 502578 1006032
rect 504364 1006052 504416 1006058
rect 500500 1005994 500552 1006000
rect 504364 1005994 504416 1006000
rect 465724 998436 465776 998442
rect 465724 998378 465776 998384
rect 462962 996296 463018 996305
rect 462962 996231 463018 996240
rect 468496 996062 468524 1005994
rect 469312 1002584 469364 1002590
rect 469312 1002526 469364 1002532
rect 469220 1001224 469272 1001230
rect 469220 1001166 469272 1001172
rect 469232 998918 469260 1001166
rect 469324 999190 469352 1002526
rect 498120 1001994 498148 1005994
rect 503352 1005304 503404 1005310
rect 503350 1005272 503352 1005281
rect 503404 1005272 503406 1005281
rect 503350 1005207 503406 1005216
rect 501326 1004864 501382 1004873
rect 499488 1004828 499540 1004834
rect 501326 1004799 501328 1004808
rect 499488 1004770 499540 1004776
rect 501380 1004799 501382 1004808
rect 501328 1004770 501380 1004776
rect 499028 1004760 499080 1004766
rect 499028 1004702 499080 1004708
rect 498474 1002008 498530 1002017
rect 498120 1001966 498474 1001994
rect 469404 999796 469456 999802
rect 469404 999738 469456 999744
rect 469312 999184 469364 999190
rect 469312 999126 469364 999132
rect 469220 998912 469272 998918
rect 469220 998854 469272 998860
rect 469416 998481 469444 999738
rect 472072 999184 472124 999190
rect 472072 999126 472124 999132
rect 469402 998472 469458 998481
rect 469402 998407 469458 998416
rect 468484 996056 468536 996062
rect 468484 995998 468536 996004
rect 472084 995586 472112 999126
rect 472256 998912 472308 998918
rect 472256 998854 472308 998860
rect 472164 998572 472216 998578
rect 472164 998514 472216 998520
rect 472176 995654 472204 998514
rect 472268 995722 472296 998854
rect 472624 998504 472676 998510
rect 472438 998472 472494 998481
rect 472624 998446 472676 998452
rect 472438 998407 472494 998416
rect 472532 998436 472584 998442
rect 472348 998232 472400 998238
rect 472348 998174 472400 998180
rect 472360 995926 472388 998174
rect 472348 995920 472400 995926
rect 472348 995862 472400 995868
rect 472452 995790 472480 998407
rect 472532 998378 472584 998384
rect 472544 995858 472572 998378
rect 472636 997257 472664 998446
rect 472714 998336 472770 998345
rect 472714 998271 472770 998280
rect 472622 997248 472678 997257
rect 472622 997183 472678 997192
rect 472728 996441 472756 998271
rect 488908 997756 488960 997762
rect 488908 997698 488960 997704
rect 488920 996985 488948 997698
rect 488906 996976 488962 996985
rect 488906 996911 488962 996920
rect 472714 996432 472770 996441
rect 472714 996367 472770 996376
rect 472532 995852 472584 995858
rect 472532 995794 472584 995800
rect 473360 995852 473412 995858
rect 473360 995794 473412 995800
rect 478236 995852 478288 995858
rect 478236 995794 478288 995800
rect 472440 995784 472492 995790
rect 472440 995726 472492 995732
rect 473372 995738 473400 995794
rect 474740 995784 474792 995790
rect 472256 995716 472308 995722
rect 473372 995710 473662 995738
rect 474016 995722 474306 995738
rect 478248 995738 478276 995794
rect 480810 995752 480866 995761
rect 474792 995732 474950 995738
rect 474740 995726 474950 995732
rect 474004 995716 474306 995722
rect 472256 995658 472308 995664
rect 474056 995710 474306 995716
rect 474752 995710 474950 995726
rect 478248 995710 478630 995738
rect 482006 995752 482062 995761
rect 480866 995710 481114 995738
rect 480810 995687 480866 995696
rect 485594 995752 485650 995761
rect 482062 995710 482310 995738
rect 485346 995710 485594 995738
rect 482006 995687 482062 995696
rect 485594 995687 485650 995696
rect 474004 995658 474056 995664
rect 472164 995648 472216 995654
rect 477684 995648 477736 995654
rect 472164 995590 472216 995596
rect 476960 995586 477342 995602
rect 482650 995616 482706 995625
rect 477736 995596 477986 995602
rect 477684 995590 477986 995596
rect 472072 995580 472124 995586
rect 472072 995522 472124 995528
rect 476948 995580 477342 995586
rect 477000 995574 477342 995580
rect 477696 995574 477986 995590
rect 482706 995574 482954 995602
rect 482650 995551 482706 995560
rect 476948 995522 477000 995528
rect 476394 995480 476450 995489
rect 476450 995438 476790 995466
rect 476394 995415 476450 995424
rect 459650 995344 459706 995353
rect 459650 995279 459706 995288
rect 481652 995217 481680 995452
rect 484136 995353 484164 995452
rect 484122 995344 484178 995353
rect 484122 995279 484178 995288
rect 454314 995208 454370 995217
rect 454314 995143 454370 995152
rect 481638 995208 481694 995217
rect 481638 995143 481694 995152
rect 485976 995081 486004 995452
rect 449806 995072 449862 995081
rect 447140 995036 447192 995042
rect 449806 995007 449862 995016
rect 485962 995072 486018 995081
rect 487816 995042 487844 995452
rect 485962 995007 486018 995016
rect 487804 995036 487856 995042
rect 447140 994978 447192 994984
rect 487804 994978 487856 994984
rect 446494 991536 446550 991545
rect 498120 991506 498148 1001966
rect 498474 1001943 498530 1001952
rect 499040 998646 499068 1004702
rect 499212 1004692 499264 1004698
rect 499212 1004634 499264 1004640
rect 499028 998640 499080 998646
rect 499028 998582 499080 998588
rect 499224 998578 499252 1004634
rect 499500 999802 499528 1004770
rect 500868 1004760 500920 1004766
rect 500498 1004728 500554 1004737
rect 500498 1004663 500500 1004672
rect 500552 1004663 500554 1004672
rect 500866 1004728 500868 1004737
rect 500920 1004728 500922 1004737
rect 500866 1004663 500922 1004672
rect 500500 1004634 500552 1004640
rect 503720 1003944 503772 1003950
rect 503718 1003912 503720 1003921
rect 503772 1003912 503774 1003921
rect 503718 1003847 503774 1003856
rect 502522 1002280 502578 1002289
rect 501984 1002238 502522 1002266
rect 501694 1002008 501750 1002017
rect 501694 1001943 501750 1001952
rect 499488 999796 499540 999802
rect 499488 999738 499540 999744
rect 499212 998572 499264 998578
rect 499212 998514 499264 998520
rect 501708 995042 501736 1001943
rect 501984 995110 502012 1002238
rect 502522 1002215 502578 1002224
rect 503718 1002144 503774 1002153
rect 502156 1002108 502208 1002114
rect 503718 1002079 503720 1002088
rect 502156 1002050 502208 1002056
rect 503772 1002079 503774 1002088
rect 503720 1002050 503772 1002056
rect 502168 998442 502196 1002050
rect 504272 999796 504324 999802
rect 504272 999738 504324 999744
rect 502156 998436 502208 998442
rect 502156 998378 502208 998384
rect 504284 995994 504312 999738
rect 504376 998510 504404 1005994
rect 508686 1005136 508742 1005145
rect 508686 1005071 508688 1005080
rect 508740 1005071 508742 1005080
rect 511264 1005100 511316 1005106
rect 508688 1005042 508740 1005048
rect 511264 1005042 511316 1005048
rect 507032 1005032 507084 1005038
rect 507030 1005000 507032 1005009
rect 509792 1005032 509844 1005038
rect 507084 1005000 507086 1005009
rect 507030 1004935 507086 1004944
rect 508226 1005000 508282 1005009
rect 509792 1004974 509844 1004980
rect 508226 1004935 508228 1004944
rect 508280 1004935 508282 1004944
rect 508228 1004906 508280 1004912
rect 507858 1004864 507914 1004873
rect 507858 1004799 507860 1004808
rect 507912 1004799 507914 1004808
rect 507860 1004770 507912 1004776
rect 509056 1004760 509108 1004766
rect 507398 1004728 507454 1004737
rect 507398 1004663 507400 1004672
rect 507452 1004663 507454 1004672
rect 509054 1004728 509056 1004737
rect 509108 1004728 509110 1004737
rect 509054 1004663 509110 1004672
rect 509240 1004692 509292 1004698
rect 507400 1004634 507452 1004640
rect 509240 1004634 509292 1004640
rect 505836 1002040 505888 1002046
rect 505834 1002008 505836 1002017
rect 508688 1002040 508740 1002046
rect 505888 1002008 505890 1002017
rect 505834 1001943 505890 1001952
rect 506202 1002008 506258 1002017
rect 506202 1001943 506204 1001952
rect 506256 1001943 506258 1001952
rect 506570 1002008 506626 1002017
rect 508688 1001982 508740 1001988
rect 506570 1001943 506626 1001952
rect 508504 1001972 508556 1001978
rect 506204 1001914 506256 1001920
rect 504364 998504 504416 998510
rect 504364 998446 504416 998452
rect 506584 996130 506612 1001943
rect 508504 1001914 508556 1001920
rect 508516 996130 508544 1001914
rect 508700 999802 508728 1001982
rect 508688 999796 508740 999802
rect 508688 999738 508740 999744
rect 506572 996124 506624 996130
rect 506572 996066 506624 996072
rect 508504 996124 508556 996130
rect 508504 996066 508556 996072
rect 509252 996062 509280 1004634
rect 509514 1002144 509570 1002153
rect 509514 1002079 509516 1002088
rect 509568 1002079 509570 1002088
rect 509516 1002050 509568 1002056
rect 509240 996056 509292 996062
rect 509240 995998 509292 996004
rect 504272 995988 504324 995994
rect 504272 995930 504324 995936
rect 509804 995926 509832 1004974
rect 510620 1004964 510672 1004970
rect 510620 1004906 510672 1004912
rect 510068 1004828 510120 1004834
rect 510068 1004770 510120 1004776
rect 509884 1002040 509936 1002046
rect 509882 1002008 509884 1002017
rect 509936 1002008 509938 1002017
rect 509882 1001943 509938 1001952
rect 510080 996062 510108 1004770
rect 510342 1002008 510398 1002017
rect 510342 1001943 510344 1001952
rect 510396 1001943 510398 1001952
rect 510344 1001914 510396 1001920
rect 510632 996198 510660 1004906
rect 510712 1004760 510764 1004766
rect 510712 1004702 510764 1004708
rect 510724 997762 510752 1004702
rect 510712 997756 510764 997762
rect 510712 997698 510764 997704
rect 511276 997694 511304 1005042
rect 514024 1002108 514076 1002114
rect 514024 1002050 514076 1002056
rect 512828 1002040 512880 1002046
rect 512828 1001982 512880 1001988
rect 512644 1001972 512696 1001978
rect 512644 1001914 512696 1001920
rect 511264 997688 511316 997694
rect 511264 997630 511316 997636
rect 510620 996192 510672 996198
rect 510620 996134 510672 996140
rect 510068 996056 510120 996062
rect 510068 995998 510120 996004
rect 509792 995920 509844 995926
rect 509792 995862 509844 995868
rect 501972 995104 502024 995110
rect 501972 995046 502024 995052
rect 501696 995036 501748 995042
rect 501696 994978 501748 994984
rect 511078 992352 511134 992361
rect 511078 992287 511134 992296
rect 446494 991471 446550 991480
rect 495164 991500 495216 991506
rect 436744 985992 436796 985998
rect 436744 985934 436796 985940
rect 429948 983606 430330 983634
rect 446508 983620 446536 991471
rect 495164 991442 495216 991448
rect 498108 991500 498160 991506
rect 498108 991442 498160 991448
rect 478972 987420 479024 987426
rect 478972 987362 479024 987368
rect 462780 985992 462832 985998
rect 462780 985934 462832 985940
rect 462792 983620 462820 985934
rect 478984 983620 479012 987362
rect 495176 983620 495204 991442
rect 511092 983634 511120 992287
rect 512656 988786 512684 1001914
rect 512840 991574 512868 1001982
rect 513932 999796 513984 999802
rect 513932 999738 513984 999744
rect 513944 997762 513972 999738
rect 513932 997756 513984 997762
rect 513932 997698 513984 997704
rect 512828 991568 512880 991574
rect 512828 991510 512880 991516
rect 512644 988780 512696 988786
rect 512644 988722 512696 988728
rect 514036 985998 514064 1002050
rect 514128 999122 514156 1006198
rect 514220 1000482 514248 1006334
rect 555974 1006295 555976 1006304
rect 556028 1006295 556030 1006304
rect 555976 1006266 556028 1006272
rect 557170 1006224 557226 1006233
rect 516784 1006188 516836 1006194
rect 557170 1006159 557172 1006168
rect 516784 1006130 516836 1006136
rect 557224 1006159 557226 1006168
rect 565176 1006188 565228 1006194
rect 557172 1006130 557224 1006136
rect 565176 1006130 565228 1006136
rect 514208 1000476 514260 1000482
rect 514208 1000418 514260 1000424
rect 514116 999116 514168 999122
rect 514116 999058 514168 999064
rect 516796 998714 516824 1006130
rect 550270 1006088 550326 1006097
rect 518900 1006052 518952 1006058
rect 518900 1005994 518952 1006000
rect 549168 1006052 549220 1006058
rect 550270 1006023 550272 1006032
rect 549168 1005994 549220 1006000
rect 550324 1006023 550326 1006032
rect 551098 1006088 551154 1006097
rect 551098 1006023 551100 1006032
rect 550272 1005994 550324 1006000
rect 551152 1006023 551154 1006032
rect 552294 1006088 552350 1006097
rect 556802 1006088 556858 1006097
rect 552294 1006023 552296 1006032
rect 551100 1005994 551152 1006000
rect 552348 1006023 552350 1006032
rect 556712 1006052 556764 1006058
rect 552296 1005994 552348 1006000
rect 556802 1006023 556804 1006032
rect 556712 1005994 556764 1006000
rect 556856 1006023 556858 1006032
rect 556804 1005994 556856 1006000
rect 518912 1001910 518940 1005994
rect 518992 1005304 519044 1005310
rect 518992 1005246 519044 1005252
rect 518900 1001904 518952 1001910
rect 518900 1001846 518952 1001852
rect 516784 998708 516836 998714
rect 516784 998650 516836 998656
rect 516876 998640 516928 998646
rect 516876 998582 516928 998588
rect 516692 997756 516744 997762
rect 516692 997698 516744 997704
rect 516704 996441 516732 997698
rect 516784 997688 516836 997694
rect 516784 997630 516836 997636
rect 516796 996985 516824 997630
rect 516782 996976 516838 996985
rect 516782 996911 516838 996920
rect 516690 996432 516746 996441
rect 516690 996367 516746 996376
rect 516888 995625 516916 998582
rect 516968 998572 517020 998578
rect 516968 998514 517020 998520
rect 516874 995616 516930 995625
rect 516874 995551 516930 995560
rect 516980 995217 517008 998514
rect 519004 997966 519032 1005246
rect 519268 1003944 519320 1003950
rect 519268 1003886 519320 1003892
rect 518992 997960 519044 997966
rect 518992 997902 519044 997908
rect 519280 995489 519308 1003886
rect 549076 1001972 549128 1001978
rect 549076 1001914 549128 1001920
rect 523868 1001904 523920 1001910
rect 523868 1001846 523920 1001852
rect 520188 1000476 520240 1000482
rect 520188 1000418 520240 1000424
rect 520096 999116 520148 999122
rect 520096 999058 520148 999064
rect 519266 995480 519322 995489
rect 519266 995415 519322 995424
rect 516966 995208 517022 995217
rect 520108 995178 520136 999058
rect 520200 996577 520228 1000418
rect 522396 998504 522448 998510
rect 522396 998446 522448 998452
rect 520186 996568 520242 996577
rect 520186 996503 520242 996512
rect 522408 995353 522436 998446
rect 523880 995722 523908 1001846
rect 524052 998708 524104 998714
rect 524052 998650 524104 998656
rect 524064 998594 524092 998650
rect 524064 998566 524184 998594
rect 524052 998436 524104 998442
rect 524052 998378 524104 998384
rect 523960 997960 524012 997966
rect 523960 997902 524012 997908
rect 523972 995858 524000 997902
rect 524064 997257 524092 998378
rect 524050 997248 524106 997257
rect 524050 997183 524106 997192
rect 523960 995852 524012 995858
rect 523960 995794 524012 995800
rect 524156 995790 524184 998566
rect 549088 998442 549116 1001914
rect 549076 998436 549128 998442
rect 549076 998378 549128 998384
rect 540888 997756 540940 997762
rect 540888 997698 540940 997704
rect 540900 996985 540928 997698
rect 540886 996976 540942 996985
rect 540886 996911 540942 996920
rect 525340 995852 525392 995858
rect 525340 995794 525392 995800
rect 533436 995852 533488 995858
rect 533436 995794 533488 995800
rect 524144 995784 524196 995790
rect 524144 995726 524196 995732
rect 524788 995784 524840 995790
rect 525352 995738 525380 995794
rect 526166 995752 526222 995761
rect 524840 995732 525090 995738
rect 524788 995726 525090 995732
rect 523868 995716 523920 995722
rect 524800 995710 525090 995726
rect 525352 995710 525734 995738
rect 528006 995752 528062 995761
rect 526222 995710 526378 995738
rect 526166 995687 526222 995696
rect 532146 995752 532202 995761
rect 528062 995710 528218 995738
rect 529032 995722 529414 995738
rect 529020 995716 529414 995722
rect 528006 995687 528062 995696
rect 523868 995658 523920 995664
rect 529072 995710 529414 995716
rect 533448 995738 533476 995794
rect 536562 995752 536618 995761
rect 532202 995710 532542 995738
rect 533448 995710 533738 995738
rect 532146 995687 532202 995696
rect 536618 995710 536774 995738
rect 536562 995687 536618 995696
rect 529020 995658 529072 995664
rect 529846 995616 529902 995625
rect 529902 995574 530058 995602
rect 529846 995551 529902 995560
rect 538954 995480 539010 995489
rect 522394 995344 522450 995353
rect 522394 995279 522450 995288
rect 516966 995143 517022 995152
rect 520096 995172 520148 995178
rect 520096 995114 520148 995120
rect 528756 995110 528784 995452
rect 533080 995217 533108 995452
rect 534368 995353 534396 995452
rect 534354 995344 534410 995353
rect 534354 995279 534410 995288
rect 533066 995208 533122 995217
rect 533066 995143 533122 995152
rect 528744 995104 528796 995110
rect 528744 995046 528796 995052
rect 535564 995042 535592 995452
rect 537404 995178 537432 995452
rect 539010 995438 539258 995466
rect 538954 995415 539010 995424
rect 537392 995172 537444 995178
rect 537392 995114 537444 995120
rect 535552 995036 535604 995042
rect 535552 994978 535604 994984
rect 527640 991568 527692 991574
rect 527640 991510 527692 991516
rect 514024 985992 514076 985998
rect 514024 985934 514076 985940
rect 511092 983606 511474 983634
rect 527652 983620 527680 991510
rect 543832 988780 543884 988786
rect 543832 988722 543884 988728
rect 543844 983620 543872 988722
rect 549180 984978 549208 1005994
rect 556344 1004760 556396 1004766
rect 556342 1004728 556344 1004737
rect 556396 1004728 556398 1004737
rect 556342 1004663 556398 1004672
rect 554778 1003368 554834 1003377
rect 554700 1003338 554778 1003354
rect 553400 1003332 553452 1003338
rect 553400 1003274 553452 1003280
rect 554688 1003332 554778 1003338
rect 554740 1003326 554778 1003332
rect 554778 1003303 554834 1003312
rect 554688 1003274 554740 1003280
rect 550272 1002176 550324 1002182
rect 553124 1002176 553176 1002182
rect 550272 1002118 550324 1002124
rect 552294 1002144 552350 1002153
rect 550284 999802 550312 1002118
rect 550364 1002108 550416 1002114
rect 552294 1002079 552296 1002088
rect 550364 1002050 550416 1002056
rect 552348 1002079 552350 1002088
rect 553122 1002144 553124 1002153
rect 553176 1002144 553178 1002153
rect 553122 1002079 553178 1002088
rect 552296 1002050 552348 1002056
rect 550272 999796 550324 999802
rect 550272 999738 550324 999744
rect 550376 997626 550404 1002050
rect 550456 1002040 550508 1002046
rect 552664 1002040 552716 1002046
rect 550456 1001982 550508 1001988
rect 551466 1002008 551522 1002017
rect 550364 997620 550416 997626
rect 550364 997562 550416 997568
rect 550468 997082 550496 1001982
rect 552662 1002008 552664 1002017
rect 553124 1002040 553176 1002046
rect 552716 1002008 552718 1002017
rect 551466 1001943 551468 1001952
rect 551520 1001943 551522 1001952
rect 551928 1001972 551980 1001978
rect 551468 1001914 551520 1001920
rect 553124 1001982 553176 1001988
rect 552662 1001943 552718 1001952
rect 551928 1001914 551980 1001920
rect 551940 999870 551968 1001914
rect 551928 999864 551980 999870
rect 551928 999806 551980 999812
rect 550456 997076 550508 997082
rect 550456 997018 550508 997024
rect 553136 995110 553164 1001982
rect 553124 995104 553176 995110
rect 553124 995046 553176 995052
rect 553412 995042 553440 1003274
rect 553950 1002688 554006 1002697
rect 553950 1002623 553952 1002632
rect 554004 1002623 554006 1002632
rect 553952 1002594 554004 1002600
rect 554320 1002584 554372 1002590
rect 554318 1002552 554320 1002561
rect 554372 1002552 554374 1002561
rect 554318 1002487 554374 1002496
rect 555148 1002040 555200 1002046
rect 553490 1002008 553546 1002017
rect 553490 1001943 553492 1001952
rect 553544 1001943 553546 1001952
rect 555146 1002008 555148 1002017
rect 555200 1002008 555202 1002017
rect 555146 1001943 555202 1001952
rect 553492 1001914 553544 1001920
rect 556724 996198 556752 1005994
rect 559748 1004760 559800 1004766
rect 557630 1004728 557686 1004737
rect 559748 1004702 559800 1004708
rect 557630 1004663 557632 1004672
rect 557684 1004663 557686 1004672
rect 559564 1004692 559616 1004698
rect 557632 1004634 557684 1004640
rect 559564 1004634 559616 1004640
rect 559196 1002448 559248 1002454
rect 559194 1002416 559196 1002425
rect 559248 1002416 559250 1002425
rect 559194 1002351 559250 1002360
rect 558460 1002312 558512 1002318
rect 558458 1002280 558460 1002289
rect 558512 1002280 558514 1002289
rect 558458 1002215 558514 1002224
rect 558000 1002040 558052 1002046
rect 557998 1002008 558000 1002017
rect 558052 1002008 558054 1002017
rect 557998 1001943 558054 1001952
rect 558826 1002008 558882 1002017
rect 558826 1001943 558828 1001952
rect 558880 1001943 558882 1001952
rect 558828 1001914 558880 1001920
rect 556712 996192 556764 996198
rect 556712 996134 556764 996140
rect 557538 995888 557594 995897
rect 557538 995823 557540 995832
rect 557592 995823 557594 995832
rect 557540 995794 557592 995800
rect 553400 995036 553452 995042
rect 553400 994978 553452 994984
rect 559576 991574 559604 1004634
rect 559654 1002280 559710 1002289
rect 559654 1002215 559656 1002224
rect 559708 1002215 559710 1002224
rect 559656 1002186 559708 1002192
rect 559760 997150 559788 1004702
rect 564992 1002652 565044 1002658
rect 564992 1002594 565044 1002600
rect 562508 1002448 562560 1002454
rect 560850 1002416 560906 1002425
rect 562508 1002390 562560 1002396
rect 560850 1002351 560852 1002360
rect 560904 1002351 560906 1002360
rect 560852 1002322 560904 1002328
rect 560944 1002312 560996 1002318
rect 560944 1002254 560996 1002260
rect 560484 1002176 560536 1002182
rect 560022 1002144 560078 1002153
rect 560022 1002079 560024 1002088
rect 560076 1002079 560078 1002088
rect 560482 1002144 560484 1002153
rect 560536 1002144 560538 1002153
rect 560482 1002079 560538 1002088
rect 560024 1002050 560076 1002056
rect 560576 1002040 560628 1002046
rect 560576 1001982 560628 1001988
rect 560300 1001972 560352 1001978
rect 560300 1001914 560352 1001920
rect 559748 997144 559800 997150
rect 559748 997086 559800 997092
rect 560312 995926 560340 1001914
rect 560588 996130 560616 1001982
rect 560576 996124 560628 996130
rect 560576 996066 560628 996072
rect 560300 995920 560352 995926
rect 560300 995862 560352 995868
rect 559564 991568 559616 991574
rect 559564 991510 559616 991516
rect 560956 990282 560984 1002254
rect 561772 1002244 561824 1002250
rect 561772 1002186 561824 1002192
rect 561680 1002040 561732 1002046
rect 561310 1002008 561366 1002017
rect 561310 1001943 561312 1001952
rect 561364 1001943 561366 1001952
rect 561678 1002008 561680 1002017
rect 561732 1002008 561734 1002017
rect 561678 1001943 561734 1001952
rect 561312 1001914 561364 1001920
rect 561784 996062 561812 1002186
rect 562324 1002108 562376 1002114
rect 562324 1002050 562376 1002056
rect 561772 996056 561824 996062
rect 561772 995998 561824 996004
rect 560944 990276 560996 990282
rect 560944 990218 560996 990224
rect 562336 990214 562364 1002050
rect 562520 993002 562548 1002390
rect 563060 1002176 563112 1002182
rect 563060 1002118 563112 1002124
rect 563072 997762 563100 1002118
rect 563704 1002040 563756 1002046
rect 563704 1001982 563756 1001988
rect 563060 997756 563112 997762
rect 563060 997698 563112 997704
rect 562508 992996 562560 993002
rect 562508 992938 562560 992944
rect 562324 990208 562376 990214
rect 562324 990150 562376 990156
rect 563716 987426 563744 1001982
rect 563888 1001972 563940 1001978
rect 563888 1001914 563940 1001920
rect 563900 988786 563928 1001914
rect 565004 997558 565032 1002594
rect 565084 1002380 565136 1002386
rect 565084 1002322 565136 1002328
rect 564992 997552 565044 997558
rect 564992 997494 565044 997500
rect 563888 988780 563940 988786
rect 563888 988722 563940 988728
rect 563704 987420 563756 987426
rect 563704 987362 563756 987368
rect 565096 985998 565124 1002322
rect 565188 997490 565216 1006130
rect 570604 1006052 570656 1006058
rect 570604 1005994 570656 1006000
rect 573364 1006052 573416 1006058
rect 573364 1005994 573416 1006000
rect 567292 1002584 567344 1002590
rect 567292 1002526 567344 1002532
rect 567304 997762 567332 1002526
rect 568212 999864 568264 999870
rect 568212 999806 568264 999812
rect 567936 999796 567988 999802
rect 567936 999738 567988 999744
rect 567292 997756 567344 997762
rect 567292 997698 567344 997704
rect 565176 997484 565228 997490
rect 565176 997426 565228 997432
rect 567948 995246 567976 999738
rect 568224 997694 568252 999806
rect 568212 997688 568264 997694
rect 568212 997630 568264 997636
rect 568212 995852 568264 995858
rect 568212 995794 568264 995800
rect 568224 995761 568252 995794
rect 568210 995752 568266 995761
rect 568210 995687 568266 995696
rect 567936 995240 567988 995246
rect 567936 995182 567988 995188
rect 570616 995178 570644 1005994
rect 572720 998436 572772 998442
rect 572720 998378 572772 998384
rect 572732 995314 572760 998378
rect 573376 997218 573404 1005994
rect 611360 1000544 611412 1000550
rect 611360 1000486 611412 1000492
rect 625712 1000544 625764 1000550
rect 625712 1000486 625764 1000492
rect 611372 997694 611400 1000486
rect 611360 997688 611412 997694
rect 611360 997630 611412 997636
rect 590476 997532 590528 997538
rect 590476 997474 590528 997480
rect 590384 997336 590436 997342
rect 590384 997278 590436 997284
rect 573364 997212 573416 997218
rect 573364 997154 573416 997160
rect 590396 996418 590424 997278
rect 590488 996554 590516 997474
rect 590568 997444 590620 997450
rect 590568 997386 590620 997392
rect 590580 996713 590608 997386
rect 620284 997212 620336 997218
rect 620284 997154 620336 997160
rect 618168 997144 618220 997150
rect 618168 997086 618220 997092
rect 590566 996704 590622 996713
rect 590566 996639 590622 996648
rect 590566 996568 590622 996577
rect 590488 996526 590566 996554
rect 590566 996503 590622 996512
rect 590566 996432 590622 996441
rect 590396 996390 590566 996418
rect 590566 996367 590622 996376
rect 572720 995308 572772 995314
rect 572720 995250 572772 995256
rect 618180 995217 618208 997086
rect 618166 995208 618222 995217
rect 570604 995172 570656 995178
rect 618166 995143 618222 995152
rect 570604 995114 570656 995120
rect 620296 995081 620324 997154
rect 622400 997076 622452 997082
rect 622400 997018 622452 997024
rect 622412 996169 622440 997018
rect 622398 996160 622454 996169
rect 622398 996095 622454 996104
rect 625724 995722 625752 1000486
rect 625804 997824 625856 997830
rect 625804 997766 625856 997772
rect 625816 995790 625844 997766
rect 634728 995852 634780 995858
rect 634728 995794 634780 995800
rect 625804 995784 625856 995790
rect 625804 995726 625856 995732
rect 627184 995784 627236 995790
rect 627918 995752 627974 995761
rect 627236 995732 627532 995738
rect 627184 995726 627532 995732
rect 625712 995716 625764 995722
rect 627196 995710 627532 995726
rect 630310 995752 630366 995761
rect 627974 995710 628176 995738
rect 627918 995687 627974 995696
rect 631598 995752 631654 995761
rect 630366 995710 630568 995738
rect 630876 995722 631212 995738
rect 630864 995716 631212 995722
rect 630310 995687 630366 995696
rect 625712 995658 625764 995664
rect 630916 995710 631212 995716
rect 634740 995738 634768 995794
rect 631654 995710 631856 995738
rect 634740 995710 634892 995738
rect 631598 995687 631654 995696
rect 630864 995658 630916 995664
rect 635186 995616 635242 995625
rect 635242 995574 635536 995602
rect 635186 995551 635242 995560
rect 626874 995217 626902 995452
rect 629680 995438 630016 995466
rect 634004 995438 634340 995466
rect 626860 995208 626916 995217
rect 626860 995143 626916 995152
rect 629680 995081 629708 995438
rect 634004 995110 634032 995438
rect 636166 995314 636194 995452
rect 636154 995308 636206 995314
rect 636154 995250 636206 995256
rect 637362 995246 637390 995452
rect 638572 995438 638908 995466
rect 637350 995240 637402 995246
rect 637350 995182 637402 995188
rect 633992 995104 634044 995110
rect 620282 995072 620338 995081
rect 620282 995007 620338 995016
rect 629666 995072 629722 995081
rect 633992 995046 634044 995052
rect 638880 995042 638908 995438
rect 638972 995438 639216 995466
rect 640720 995438 641056 995466
rect 638972 995178 639000 995438
rect 638960 995172 639012 995178
rect 638960 995114 639012 995120
rect 640720 995110 640748 995438
rect 640708 995104 640760 995110
rect 640708 995046 640760 995052
rect 629666 995007 629722 995016
rect 638868 995036 638920 995042
rect 638868 994978 638920 994984
rect 640800 995036 640852 995042
rect 640800 994978 640852 994984
rect 576306 990992 576362 991001
rect 576306 990927 576362 990936
rect 560116 985992 560168 985998
rect 560116 985934 560168 985940
rect 565084 985992 565136 985998
rect 565084 985934 565136 985940
rect 549168 984972 549220 984978
rect 549168 984914 549220 984920
rect 560128 983620 560156 985934
rect 576320 983620 576348 990927
rect 592500 988780 592552 988786
rect 592500 988722 592552 988728
rect 592512 983620 592540 988722
rect 608784 987420 608836 987426
rect 608784 987362 608836 987368
rect 608796 983620 608824 987362
rect 624976 985992 625028 985998
rect 624976 985934 625028 985940
rect 624988 983620 625016 985934
rect 640812 983634 640840 994978
rect 661684 992996 661736 993002
rect 661684 992938 661736 992944
rect 660304 991568 660356 991574
rect 660304 991510 660356 991516
rect 658924 990276 658976 990282
rect 658924 990218 658976 990224
rect 650092 984836 650144 984842
rect 650092 984778 650144 984784
rect 650000 984700 650052 984706
rect 650000 984642 650052 984648
rect 640812 983606 641194 983634
rect 62118 976032 62174 976041
rect 62118 975967 62174 975976
rect 62132 975730 62160 975967
rect 62120 975724 62172 975730
rect 62120 975666 62172 975672
rect 62118 962976 62174 962985
rect 62118 962911 62174 962920
rect 62132 961926 62160 962911
rect 62120 961920 62172 961926
rect 62120 961862 62172 961868
rect 62118 949920 62174 949929
rect 62118 949855 62174 949864
rect 62132 946014 62160 949855
rect 62120 946008 62172 946014
rect 62120 945950 62172 945956
rect 50342 939856 50398 939865
rect 50342 939791 50398 939800
rect 48412 937032 48464 937038
rect 62120 937032 62172 937038
rect 48412 936974 48464 936980
rect 62118 937000 62120 937009
rect 62172 937000 62174 937009
rect 62118 936935 62174 936944
rect 44178 934552 44234 934561
rect 44178 934487 44234 934496
rect 42890 934144 42946 934153
rect 42890 934079 42946 934088
rect 42798 933736 42854 933745
rect 42798 933671 42854 933680
rect 41892 932866 42012 932894
rect 41880 932136 41932 932142
rect 41878 932104 41880 932113
rect 41932 932104 41934 932113
rect 41878 932039 41934 932048
rect 41708 923206 41828 923234
rect 41708 828014 41736 923206
rect 41708 827986 41828 828014
rect 41616 823846 41736 823874
rect 41708 814994 41736 823846
rect 41800 815697 41828 827986
rect 41984 816513 42012 932866
rect 43442 932104 43498 932113
rect 43442 932039 43498 932048
rect 41970 816504 42026 816513
rect 41970 816439 42026 816448
rect 41786 815688 41842 815697
rect 41786 815623 41842 815632
rect 41708 814966 41920 814994
rect 41512 814904 41564 814910
rect 41788 814904 41840 814910
rect 41512 814846 41564 814852
rect 41786 814872 41788 814881
rect 41840 814872 41842 814881
rect 41786 814807 41842 814816
rect 41892 814065 41920 814966
rect 41878 814056 41934 814065
rect 41878 813991 41934 814000
rect 42154 812832 42210 812841
rect 42154 812767 42210 812776
rect 33782 812424 33838 812433
rect 33782 812359 33838 812368
rect 33046 810384 33102 810393
rect 33046 810319 33102 810328
rect 32402 809160 32458 809169
rect 32402 809095 32458 809104
rect 32416 801106 32444 809095
rect 33060 802505 33088 810319
rect 33046 802496 33102 802505
rect 33046 802431 33102 802440
rect 32404 801100 32456 801106
rect 32404 801042 32456 801048
rect 33796 801009 33824 812359
rect 35162 812016 35218 812025
rect 35162 811951 35218 811960
rect 34426 810792 34482 810801
rect 34426 810727 34482 810736
rect 34440 802641 34468 810727
rect 35176 802777 35204 811951
rect 40682 811608 40738 811617
rect 40682 811543 40738 811552
rect 35254 808752 35310 808761
rect 35254 808687 35310 808696
rect 35162 802768 35218 802777
rect 35162 802703 35218 802712
rect 34426 802632 34482 802641
rect 34426 802567 34482 802576
rect 35268 801174 35296 808687
rect 35806 807328 35862 807337
rect 35806 807263 35862 807272
rect 35820 806478 35848 807263
rect 35808 806472 35860 806478
rect 35808 806414 35860 806420
rect 35256 801168 35308 801174
rect 35256 801110 35308 801116
rect 33782 801000 33838 801009
rect 33782 800935 33838 800944
rect 40696 800562 40724 811543
rect 42062 809568 42118 809577
rect 42062 809503 42118 809512
rect 41786 807936 41842 807945
rect 41786 807871 41842 807880
rect 41800 804817 41828 807871
rect 41880 806472 41932 806478
rect 41880 806414 41932 806420
rect 41892 806313 41920 806414
rect 41878 806304 41934 806313
rect 41878 806239 41934 806248
rect 41786 804808 41842 804817
rect 41786 804743 41842 804752
rect 42076 803826 42104 809503
rect 42168 803894 42196 812767
rect 42338 811200 42394 811209
rect 42338 811135 42394 811144
rect 42156 803888 42208 803894
rect 42156 803830 42208 803836
rect 42064 803820 42116 803826
rect 42064 803762 42116 803768
rect 40684 800556 40736 800562
rect 40684 800498 40736 800504
rect 42352 800018 42380 811135
rect 42616 803888 42668 803894
rect 42616 803830 42668 803836
rect 42156 800012 42208 800018
rect 42156 799954 42208 799960
rect 42340 800012 42392 800018
rect 42340 799954 42392 799960
rect 42168 799445 42196 799954
rect 42628 798182 42656 803830
rect 42708 803820 42760 803826
rect 42708 803762 42760 803768
rect 42720 799218 42748 803762
rect 43076 801168 43128 801174
rect 43076 801110 43128 801116
rect 42892 801100 42944 801106
rect 42892 801042 42944 801048
rect 42720 799190 42840 799218
rect 42708 799128 42760 799134
rect 42708 799070 42760 799076
rect 42156 798176 42208 798182
rect 42156 798118 42208 798124
rect 42616 798176 42668 798182
rect 42616 798118 42668 798124
rect 42168 797605 42196 798118
rect 42720 797298 42748 799070
rect 42156 797292 42208 797298
rect 42156 797234 42208 797240
rect 42708 797292 42760 797298
rect 42708 797234 42760 797240
rect 42168 796960 42196 797234
rect 42812 797178 42840 799190
rect 42720 797150 42840 797178
rect 42430 796784 42486 796793
rect 42430 796719 42486 796728
rect 42156 796340 42208 796346
rect 42156 796282 42208 796288
rect 42168 795765 42196 796282
rect 42444 795054 42472 796719
rect 42720 796346 42748 797150
rect 42708 796340 42760 796346
rect 42708 796282 42760 796288
rect 42904 796226 42932 801042
rect 42984 800556 43036 800562
rect 42984 800498 43036 800504
rect 42720 796198 42932 796226
rect 42156 795048 42208 795054
rect 42156 794990 42208 794996
rect 42432 795048 42484 795054
rect 42432 794990 42484 794996
rect 42168 794580 42196 794990
rect 42432 794912 42484 794918
rect 42432 794854 42484 794860
rect 42156 794300 42208 794306
rect 42156 794242 42208 794248
rect 42168 793900 42196 794242
rect 42156 793824 42208 793830
rect 42156 793766 42208 793772
rect 42168 793288 42196 793766
rect 42444 793218 42472 794854
rect 42720 794306 42748 796198
rect 42996 794918 43024 800498
rect 42984 794912 43036 794918
rect 42984 794854 43036 794860
rect 43088 794594 43116 801110
rect 43168 794912 43220 794918
rect 43168 794854 43220 794860
rect 42812 794566 43116 794594
rect 42708 794300 42760 794306
rect 42708 794242 42760 794248
rect 42812 794186 42840 794566
rect 42720 794158 42840 794186
rect 42156 793212 42208 793218
rect 42156 793154 42208 793160
rect 42432 793212 42484 793218
rect 42432 793154 42484 793160
rect 42168 792744 42196 793154
rect 42432 793076 42484 793082
rect 42432 793018 42484 793024
rect 42338 792024 42394 792033
rect 42338 791959 42394 791968
rect 42156 790696 42208 790702
rect 42156 790638 42208 790644
rect 42168 790228 42196 790638
rect 42156 790152 42208 790158
rect 42156 790094 42208 790100
rect 42168 789616 42196 790094
rect 42352 789478 42380 791959
rect 42444 790158 42472 793018
rect 42720 790702 42748 794158
rect 43180 793830 43208 794854
rect 43168 793824 43220 793830
rect 43168 793766 43220 793772
rect 42708 790696 42760 790702
rect 42708 790638 42760 790644
rect 42432 790152 42484 790158
rect 42432 790094 42484 790100
rect 42156 789472 42208 789478
rect 42156 789414 42208 789420
rect 42340 789472 42392 789478
rect 42340 789414 42392 789420
rect 42168 788936 42196 789414
rect 42154 788760 42210 788769
rect 42154 788695 42210 788704
rect 42168 788392 42196 788695
rect 42706 788216 42762 788225
rect 42706 788151 42762 788160
rect 42430 788080 42486 788089
rect 42430 788015 42486 788024
rect 41878 786992 41934 787001
rect 41878 786927 41934 786936
rect 41892 786556 41920 786927
rect 42444 786486 42472 788015
rect 42064 786480 42116 786486
rect 42064 786422 42116 786428
rect 42432 786480 42484 786486
rect 42432 786422 42484 786428
rect 42076 785944 42104 786422
rect 42720 785670 42748 788151
rect 42156 785664 42208 785670
rect 42156 785606 42208 785612
rect 42708 785664 42760 785670
rect 42708 785606 42760 785612
rect 42168 785264 42196 785606
rect 8588 775132 8616 775268
rect 9048 775132 9076 775268
rect 9508 775132 9536 775268
rect 9968 775132 9996 775268
rect 10428 775132 10456 775268
rect 10888 775132 10916 775268
rect 11348 775132 11376 775268
rect 11808 775132 11836 775268
rect 12268 775132 12296 775268
rect 12728 775132 12756 775268
rect 13188 775132 13216 775268
rect 13648 775132 13676 775268
rect 14108 775132 14136 775268
rect 35806 774344 35862 774353
rect 35806 774279 35862 774288
rect 35820 774246 35848 774279
rect 35808 774240 35860 774246
rect 35808 774182 35860 774188
rect 42798 772032 42854 772041
rect 42798 771967 42854 771976
rect 33782 769448 33838 769457
rect 33782 769383 33838 769392
rect 32402 768632 32458 768641
rect 32402 768567 32458 768576
rect 31022 767816 31078 767825
rect 31022 767751 31078 767760
rect 30378 764144 30434 764153
rect 30378 764079 30434 764088
rect 30392 763337 30420 764079
rect 30378 763328 30434 763337
rect 30378 763263 30434 763272
rect 31036 759694 31064 767751
rect 31024 759688 31076 759694
rect 31024 759630 31076 759636
rect 32416 758334 32444 768567
rect 32494 766592 32550 766601
rect 32494 766527 32550 766536
rect 32508 758402 32536 766527
rect 33796 758538 33824 769383
rect 40682 769040 40738 769049
rect 40682 768975 40738 768984
rect 33874 767408 33930 767417
rect 33874 767343 33930 767352
rect 33784 758532 33836 758538
rect 33784 758474 33836 758480
rect 32496 758396 32548 758402
rect 32496 758338 32548 758344
rect 32404 758328 32456 758334
rect 33888 758305 33916 767343
rect 32404 758270 32456 758276
rect 33874 758296 33930 758305
rect 33874 758231 33930 758240
rect 40696 757761 40724 768975
rect 41510 762920 41566 762929
rect 41510 762855 41566 762864
rect 41524 761802 41552 762855
rect 41512 761796 41564 761802
rect 41512 761738 41564 761744
rect 41880 759688 41932 759694
rect 41880 759630 41932 759636
rect 41788 758532 41840 758538
rect 41788 758474 41840 758480
rect 40682 757752 40738 757761
rect 40682 757687 40738 757696
rect 41800 757081 41828 758474
rect 41786 757072 41842 757081
rect 41892 757042 41920 759630
rect 42708 758396 42760 758402
rect 42708 758338 42760 758344
rect 42432 758328 42484 758334
rect 42432 758270 42484 758276
rect 42444 757081 42472 758270
rect 42430 757072 42486 757081
rect 41786 757007 41842 757016
rect 41880 757036 41932 757042
rect 42430 757007 42486 757016
rect 41880 756978 41932 756984
rect 42432 756900 42484 756906
rect 42432 756842 42484 756848
rect 41880 756764 41932 756770
rect 41880 756706 41932 756712
rect 41892 756228 41920 756706
rect 42444 755546 42472 756842
rect 42720 756566 42748 758338
rect 42708 756560 42760 756566
rect 42708 756502 42760 756508
rect 42432 755540 42484 755546
rect 42432 755482 42484 755488
rect 42616 755268 42668 755274
rect 42616 755210 42668 755216
rect 41878 754896 41934 754905
rect 41878 754831 41934 754840
rect 41892 754392 41920 754831
rect 42628 754322 42656 755210
rect 42064 754316 42116 754322
rect 42064 754258 42116 754264
rect 42616 754316 42668 754322
rect 42616 754258 42668 754264
rect 42076 753780 42104 754258
rect 42614 754216 42670 754225
rect 42614 754151 42670 754160
rect 41786 753128 41842 753137
rect 41786 753063 41842 753072
rect 41800 752556 41828 753063
rect 42628 751806 42656 754151
rect 42156 751800 42208 751806
rect 42156 751742 42208 751748
rect 42616 751800 42668 751806
rect 42616 751742 42668 751748
rect 42168 751369 42196 751742
rect 42616 751664 42668 751670
rect 42616 751606 42668 751612
rect 42156 751120 42208 751126
rect 42156 751062 42208 751068
rect 42168 750720 42196 751062
rect 41786 750408 41842 750417
rect 41786 750343 41842 750352
rect 41800 750108 41828 750343
rect 42156 749828 42208 749834
rect 42156 749770 42208 749776
rect 42168 749529 42196 749770
rect 42076 746978 42104 747048
rect 42628 746978 42656 751606
rect 42706 749320 42762 749329
rect 42706 749255 42762 749264
rect 42064 746972 42116 746978
rect 42064 746914 42116 746920
rect 42156 746972 42208 746978
rect 42156 746914 42208 746920
rect 42616 746972 42668 746978
rect 42616 746914 42668 746920
rect 42168 746401 42196 746914
rect 42614 746600 42670 746609
rect 42614 746535 42670 746544
rect 42156 746088 42208 746094
rect 42156 746030 42208 746036
rect 42168 745756 42196 746030
rect 42156 745680 42208 745686
rect 42156 745622 42208 745628
rect 42168 745212 42196 745622
rect 42156 743776 42208 743782
rect 42156 743718 42208 743724
rect 42168 743376 42196 743718
rect 42628 743306 42656 746535
rect 42720 745686 42748 749255
rect 42708 745680 42760 745686
rect 42708 745622 42760 745628
rect 42708 745544 42760 745550
rect 42708 745486 42760 745492
rect 42720 743782 42748 745486
rect 42708 743776 42760 743782
rect 42708 743718 42760 743724
rect 42156 743300 42208 743306
rect 42156 743242 42208 743248
rect 42616 743300 42668 743306
rect 42616 743242 42668 743248
rect 42168 742696 42196 743242
rect 41786 742384 41842 742393
rect 41786 742319 41842 742328
rect 41800 742084 41828 742319
rect 8588 731884 8616 732020
rect 9048 731884 9076 732020
rect 9508 731884 9536 732020
rect 9968 731884 9996 732020
rect 10428 731884 10456 732020
rect 10888 731884 10916 732020
rect 11348 731884 11376 732020
rect 11808 731884 11836 732020
rect 12268 731884 12296 732020
rect 12728 731884 12756 732020
rect 13188 731884 13216 732020
rect 13648 731884 13676 732020
rect 14108 731884 14136 732020
rect 31392 731400 31444 731406
rect 31392 731342 31444 731348
rect 31404 730289 31432 731342
rect 31484 731264 31536 731270
rect 31484 731206 31536 731212
rect 31496 731105 31524 731206
rect 31576 731128 31628 731134
rect 31482 731096 31538 731105
rect 31576 731070 31628 731076
rect 31666 731096 31722 731105
rect 31482 731031 31538 731040
rect 31588 730697 31616 731070
rect 31666 731031 31722 731040
rect 31680 730998 31708 731031
rect 31668 730992 31720 730998
rect 31668 730934 31720 730940
rect 31574 730688 31630 730697
rect 31574 730623 31630 730632
rect 31390 730280 31446 730289
rect 31390 730215 31446 730224
rect 42812 729337 42840 771967
rect 42890 769992 42946 770001
rect 42890 769927 42946 769936
rect 42904 745550 42932 769927
rect 42982 768360 43038 768369
rect 42982 768295 43038 768304
rect 42996 757058 43024 768295
rect 43258 765912 43314 765921
rect 43258 765847 43314 765856
rect 42996 757030 43208 757058
rect 42984 756560 43036 756566
rect 42984 756502 43036 756508
rect 42996 751670 43024 756502
rect 42984 751664 43036 751670
rect 42984 751606 43036 751612
rect 43180 749834 43208 757030
rect 43272 751126 43300 765847
rect 43260 751120 43312 751126
rect 43260 751062 43312 751068
rect 43168 749828 43220 749834
rect 43168 749770 43220 749776
rect 42984 749420 43036 749426
rect 42984 749362 43036 749368
rect 42996 747046 43024 749362
rect 43076 747992 43128 747998
rect 43076 747934 43128 747940
rect 42984 747040 43036 747046
rect 42984 746982 43036 746988
rect 43088 746094 43116 747934
rect 43076 746088 43128 746094
rect 43076 746030 43128 746036
rect 42892 745544 42944 745550
rect 42892 745486 42944 745492
rect 42798 729328 42854 729337
rect 42798 729263 42854 729272
rect 31022 726608 31078 726617
rect 31022 726543 31078 726552
rect 31036 715465 31064 726543
rect 40682 726200 40738 726209
rect 40682 726135 40738 726144
rect 39302 725792 39358 725801
rect 39302 725727 39358 725736
rect 35806 723752 35862 723761
rect 35806 723687 35862 723696
rect 35714 723344 35770 723353
rect 35714 723279 35770 723288
rect 35728 715562 35756 723279
rect 35820 716922 35848 723687
rect 35808 716916 35860 716922
rect 35808 716858 35860 716864
rect 39316 716145 39344 725727
rect 39302 716136 39358 716145
rect 39302 716071 39358 716080
rect 35716 715556 35768 715562
rect 35716 715498 35768 715504
rect 31022 715456 31078 715465
rect 31022 715391 31078 715400
rect 40696 714270 40724 726135
rect 42062 725248 42118 725257
rect 42062 725183 42118 725192
rect 40774 724568 40830 724577
rect 40774 724503 40830 724512
rect 40788 716242 40816 724503
rect 40866 723344 40922 723353
rect 40866 723279 40922 723288
rect 40776 716236 40828 716242
rect 40776 716178 40828 716184
rect 40684 714264 40736 714270
rect 40684 714206 40736 714212
rect 40880 714202 40908 723279
rect 41510 720896 41566 720905
rect 41510 720831 41566 720840
rect 41524 719710 41552 720831
rect 41512 719704 41564 719710
rect 41510 719672 41512 719681
rect 41564 719672 41566 719681
rect 41510 719607 41566 719616
rect 41880 716236 41932 716242
rect 41880 716178 41932 716184
rect 40868 714196 40920 714202
rect 40868 714138 40920 714144
rect 41892 713862 41920 716178
rect 41880 713856 41932 713862
rect 42076 713833 42104 725183
rect 42982 722800 43038 722809
rect 42982 722735 43038 722744
rect 42432 716916 42484 716922
rect 42432 716858 42484 716864
rect 41880 713798 41932 713804
rect 42062 713824 42118 713833
rect 42062 713759 42118 713768
rect 41880 713584 41932 713590
rect 41880 713526 41932 713532
rect 41892 713048 41920 713526
rect 42444 713289 42472 716858
rect 42524 715556 42576 715562
rect 42524 715498 42576 715504
rect 42430 713280 42486 713289
rect 42430 713215 42486 713224
rect 42156 711680 42208 711686
rect 42156 711622 42208 711628
rect 42168 711212 42196 711622
rect 42536 711006 42564 715498
rect 42800 714264 42852 714270
rect 42800 714206 42852 714212
rect 42812 711686 42840 714206
rect 42892 714196 42944 714202
rect 42892 714138 42944 714144
rect 42800 711680 42852 711686
rect 42800 711622 42852 711628
rect 42524 711000 42576 711006
rect 42524 710942 42576 710948
rect 42800 711000 42852 711006
rect 42800 710942 42852 710948
rect 42156 710932 42208 710938
rect 42156 710874 42208 710880
rect 42168 710561 42196 710874
rect 42522 710832 42578 710841
rect 42522 710767 42578 710776
rect 42156 709912 42208 709918
rect 42156 709854 42208 709860
rect 42168 709376 42196 709854
rect 42536 708626 42564 710767
rect 42156 708620 42208 708626
rect 42156 708562 42208 708568
rect 42524 708620 42576 708626
rect 42524 708562 42576 708568
rect 42168 708152 42196 708562
rect 42522 708520 42578 708529
rect 42522 708455 42578 708464
rect 42156 708076 42208 708082
rect 42156 708018 42208 708024
rect 42168 707540 42196 708018
rect 42156 707260 42208 707266
rect 42156 707202 42208 707208
rect 42168 706860 42196 707202
rect 42062 706752 42118 706761
rect 42062 706687 42118 706696
rect 42076 706316 42104 706687
rect 42432 706104 42484 706110
rect 42432 706046 42484 706052
rect 42246 705120 42302 705129
rect 42246 705055 42302 705064
rect 42064 704268 42116 704274
rect 42064 704210 42116 704216
rect 42076 703868 42104 704210
rect 42156 703724 42208 703730
rect 42156 703666 42208 703672
rect 42168 703188 42196 703666
rect 42168 702522 42196 702576
rect 42260 702522 42288 705055
rect 42444 704274 42472 706046
rect 42536 705129 42564 708455
rect 42522 705120 42578 705129
rect 42522 705055 42578 705064
rect 42432 704268 42484 704274
rect 42432 704210 42484 704216
rect 42430 703760 42486 703769
rect 42812 703730 42840 710942
rect 42904 709918 42932 714138
rect 42892 709912 42944 709918
rect 42892 709854 42944 709860
rect 42892 709368 42944 709374
rect 42892 709310 42944 709316
rect 42904 707266 42932 709310
rect 42996 708082 43024 722735
rect 43076 712156 43128 712162
rect 43076 712098 43128 712104
rect 43088 710938 43116 712098
rect 43076 710932 43128 710938
rect 43076 710874 43128 710880
rect 42984 708076 43036 708082
rect 42984 708018 43036 708024
rect 42892 707260 42944 707266
rect 42892 707202 42944 707208
rect 42430 703695 42486 703704
rect 42800 703724 42852 703730
rect 42168 702494 42288 702522
rect 41786 702400 41842 702409
rect 41786 702335 41842 702344
rect 41800 702032 41828 702335
rect 42444 700466 42472 703695
rect 42800 703666 42852 703672
rect 42800 701072 42852 701078
rect 42800 701014 42852 701020
rect 42812 700754 42840 701014
rect 42720 700726 42840 700754
rect 42156 700460 42208 700466
rect 42156 700402 42208 700408
rect 42432 700460 42484 700466
rect 42432 700402 42484 700408
rect 42168 700165 42196 700402
rect 42720 699922 42748 700726
rect 42156 699916 42208 699922
rect 42156 699858 42208 699864
rect 42708 699916 42760 699922
rect 42708 699858 42760 699864
rect 42168 699516 42196 699858
rect 41786 699408 41842 699417
rect 41786 699343 41842 699352
rect 41800 698904 41828 699343
rect 30288 696244 30340 696250
rect 30288 696186 30340 696192
rect 8588 688772 8616 688908
rect 9048 688772 9076 688908
rect 9508 688772 9536 688908
rect 9968 688772 9996 688908
rect 10428 688772 10456 688908
rect 10888 688772 10916 688908
rect 11348 688772 11376 688908
rect 11808 688772 11836 688908
rect 12268 688772 12296 688908
rect 12728 688772 12756 688908
rect 13188 688772 13216 688908
rect 13648 688772 13676 688908
rect 14108 688772 14136 688908
rect 30300 687313 30328 696186
rect 35622 688392 35678 688401
rect 35622 688327 35678 688336
rect 35636 687818 35664 688327
rect 35808 687948 35860 687954
rect 35808 687890 35860 687896
rect 35624 687812 35676 687818
rect 35624 687754 35676 687760
rect 35820 687721 35848 687890
rect 35806 687712 35862 687721
rect 35806 687647 35862 687656
rect 30286 687304 30342 687313
rect 30286 687239 30342 687248
rect 39302 683632 39358 683641
rect 39302 683567 39358 683576
rect 32402 682816 32458 682825
rect 32402 682751 32458 682760
rect 31022 681592 31078 681601
rect 31022 681527 31078 681536
rect 30470 676866 30526 676875
rect 30470 676801 30526 676810
rect 31036 672790 31064 681527
rect 31024 672784 31076 672790
rect 31024 672726 31076 672732
rect 32416 671401 32444 682751
rect 35162 680368 35218 680377
rect 35162 680303 35218 680312
rect 35176 672858 35204 680303
rect 35164 672852 35216 672858
rect 35164 672794 35216 672800
rect 32402 671392 32458 671401
rect 32402 671327 32458 671336
rect 39316 670993 39344 683567
rect 41694 683088 41750 683097
rect 40684 683052 40736 683058
rect 41694 683023 41696 683032
rect 40684 682994 40736 683000
rect 41748 683023 41750 683032
rect 41696 682994 41748 683000
rect 39302 670984 39358 670993
rect 40696 670954 40724 682994
rect 41694 681864 41750 681873
rect 40776 681828 40828 681834
rect 41694 681799 41696 681808
rect 40776 681770 40828 681776
rect 41748 681799 41750 681808
rect 41696 681770 41748 681776
rect 40788 671022 40816 681770
rect 42798 681184 42854 681193
rect 42798 681119 42854 681128
rect 41970 680776 42026 680785
rect 41970 680711 42026 680720
rect 41880 672784 41932 672790
rect 41880 672726 41932 672732
rect 40776 671016 40828 671022
rect 40776 670958 40828 670964
rect 39302 670919 39358 670928
rect 40684 670948 40736 670954
rect 40684 670890 40736 670896
rect 41788 670948 41840 670954
rect 41788 670890 41840 670896
rect 41800 670721 41828 670890
rect 41786 670712 41842 670721
rect 41786 670647 41842 670656
rect 41892 670614 41920 672726
rect 41984 670614 42012 680711
rect 42432 672852 42484 672858
rect 42432 672794 42484 672800
rect 42064 671016 42116 671022
rect 42064 670958 42116 670964
rect 42076 670721 42104 670958
rect 42062 670712 42118 670721
rect 42062 670647 42118 670656
rect 41880 670608 41932 670614
rect 41880 670550 41932 670556
rect 41972 670608 42024 670614
rect 41972 670550 42024 670556
rect 41880 670404 41932 670410
rect 41880 670346 41932 670352
rect 41892 669868 41920 670346
rect 42444 670177 42472 672794
rect 42430 670168 42486 670177
rect 42430 670103 42486 670112
rect 42708 670064 42760 670070
rect 42708 670006 42760 670012
rect 41878 668536 41934 668545
rect 41878 668471 41934 668480
rect 41892 668032 41920 668471
rect 42720 667894 42748 670006
rect 42156 667888 42208 667894
rect 42156 667830 42208 667836
rect 42708 667888 42760 667894
rect 42708 667830 42760 667836
rect 42168 667352 42196 667830
rect 42812 667826 42840 681119
rect 42890 679144 42946 679153
rect 42890 679079 42946 679088
rect 42904 673454 42932 679079
rect 42904 673426 43024 673454
rect 42892 670608 42944 670614
rect 42892 670550 42944 670556
rect 42800 667820 42852 667826
rect 42800 667762 42852 667768
rect 42904 667706 42932 670550
rect 42720 667678 42932 667706
rect 42156 666732 42208 666738
rect 42156 666674 42208 666680
rect 42168 666165 42196 666674
rect 41786 665408 41842 665417
rect 41786 665343 41842 665352
rect 41800 664972 41828 665343
rect 41786 664592 41842 664601
rect 41786 664527 41842 664536
rect 41800 664325 41828 664527
rect 42156 664012 42208 664018
rect 42156 663954 42208 663960
rect 42168 663680 42196 663954
rect 42720 663814 42748 667678
rect 42800 667616 42852 667622
rect 42800 667558 42852 667564
rect 42708 663808 42760 663814
rect 42708 663750 42760 663756
rect 42062 663368 42118 663377
rect 42062 663303 42118 663312
rect 42076 663136 42104 663303
rect 42812 662658 42840 667558
rect 42892 665236 42944 665242
rect 42892 665178 42944 665184
rect 42904 664018 42932 665178
rect 42892 664012 42944 664018
rect 42892 663954 42944 663960
rect 42892 663808 42944 663814
rect 42892 663750 42944 663756
rect 42800 662652 42852 662658
rect 42800 662594 42852 662600
rect 42708 662448 42760 662454
rect 42708 662390 42760 662396
rect 42720 661450 42748 662390
rect 42720 661422 42840 661450
rect 42706 661328 42762 661337
rect 42706 661263 42762 661272
rect 42156 661088 42208 661094
rect 42156 661030 42208 661036
rect 42168 660620 42196 661030
rect 42154 660512 42210 660521
rect 42154 660447 42210 660456
rect 42168 660008 42196 660447
rect 42522 660376 42578 660385
rect 42522 660311 42578 660320
rect 42156 659728 42208 659734
rect 42156 659670 42208 659676
rect 42168 659357 42196 659670
rect 42156 659048 42208 659054
rect 42156 658990 42208 658996
rect 42168 658784 42196 658990
rect 42338 658336 42394 658345
rect 42338 658271 42394 658280
rect 42156 657280 42208 657286
rect 42156 657222 42208 657228
rect 42168 656948 42196 657222
rect 42156 656872 42208 656878
rect 42156 656814 42208 656820
rect 42168 656336 42196 656814
rect 42352 656198 42380 658271
rect 42536 657286 42564 660311
rect 42720 659054 42748 661263
rect 42812 661094 42840 661422
rect 42800 661088 42852 661094
rect 42800 661030 42852 661036
rect 42904 659734 42932 663750
rect 42996 662454 43024 673426
rect 43076 662652 43128 662658
rect 43076 662594 43128 662600
rect 42984 662448 43036 662454
rect 42984 662390 43036 662396
rect 42892 659728 42944 659734
rect 42892 659670 42944 659676
rect 42708 659048 42760 659054
rect 42708 658990 42760 658996
rect 42524 657280 42576 657286
rect 42524 657222 42576 657228
rect 43088 656878 43116 662594
rect 43076 656872 43128 656878
rect 43076 656814 43128 656820
rect 42156 656192 42208 656198
rect 42156 656134 42208 656140
rect 42340 656192 42392 656198
rect 42340 656134 42392 656140
rect 42168 655656 42196 656134
rect 8588 645524 8616 645660
rect 9048 645524 9076 645660
rect 9508 645524 9536 645660
rect 9968 645524 9996 645660
rect 10428 645524 10456 645660
rect 10888 645524 10916 645660
rect 11348 645524 11376 645660
rect 11808 645524 11836 645660
rect 12268 645524 12296 645660
rect 12728 645524 12756 645660
rect 13188 645524 13216 645660
rect 13648 645524 13676 645660
rect 14108 645524 14136 645660
rect 35622 644736 35678 644745
rect 35622 644671 35678 644680
rect 35806 644736 35862 644745
rect 35806 644671 35862 644680
rect 35636 644638 35664 644671
rect 35624 644632 35676 644638
rect 35624 644574 35676 644580
rect 35820 644570 35848 644671
rect 35808 644564 35860 644570
rect 35808 644506 35860 644512
rect 35162 640248 35218 640257
rect 35162 640183 35218 640192
rect 32402 638208 32458 638217
rect 32402 638143 32458 638152
rect 32416 629950 32444 638143
rect 33782 637800 33838 637809
rect 33782 637735 33838 637744
rect 32404 629944 32456 629950
rect 33796 629921 33824 637735
rect 32404 629886 32456 629892
rect 33782 629912 33838 629921
rect 33782 629847 33838 629856
rect 35176 628561 35204 640183
rect 39302 639840 39358 639849
rect 39302 639775 39358 639784
rect 39316 629270 39344 639775
rect 40682 639024 40738 639033
rect 40682 638959 40738 638968
rect 39304 629264 39356 629270
rect 39304 629206 39356 629212
rect 40696 629105 40724 638959
rect 42890 638616 42946 638625
rect 42890 638551 42946 638560
rect 40866 637392 40922 637401
rect 40866 637327 40922 637336
rect 40880 629241 40908 637327
rect 42798 635760 42854 635769
rect 42798 635695 42854 635704
rect 41788 629944 41840 629950
rect 41788 629886 41840 629892
rect 40866 629232 40922 629241
rect 40866 629167 40922 629176
rect 40682 629096 40738 629105
rect 40682 629031 40738 629040
rect 35162 628552 35218 628561
rect 35162 628487 35218 628496
rect 41800 627434 41828 629886
rect 42524 629264 42576 629270
rect 42524 629206 42576 629212
rect 41788 627428 41840 627434
rect 41788 627370 41840 627376
rect 41788 627088 41840 627094
rect 41788 627030 41840 627036
rect 41800 626620 41828 627030
rect 42536 625326 42564 629206
rect 42156 625320 42208 625326
rect 42156 625262 42208 625268
rect 42524 625320 42576 625326
rect 42524 625262 42576 625268
rect 42168 624784 42196 625262
rect 42522 625152 42578 625161
rect 42522 625087 42578 625096
rect 42156 624708 42208 624714
rect 42156 624650 42208 624656
rect 42168 624172 42196 624650
rect 42536 623898 42564 625087
rect 42524 623892 42576 623898
rect 42524 623834 42576 623840
rect 42522 623792 42578 623801
rect 42522 623727 42578 623736
rect 42156 623484 42208 623490
rect 42156 623426 42208 623432
rect 42168 622948 42196 623426
rect 42536 622198 42564 623727
rect 42064 622192 42116 622198
rect 42064 622134 42116 622140
rect 42524 622192 42576 622198
rect 42524 622134 42576 622140
rect 42076 621792 42104 622134
rect 42524 622056 42576 622062
rect 42524 621998 42576 622004
rect 41786 621480 41842 621489
rect 41786 621415 41842 621424
rect 41800 621112 41828 621415
rect 42536 621110 42564 621998
rect 42524 621104 42576 621110
rect 42524 621046 42576 621052
rect 42812 620974 42840 635695
rect 42904 634814 42932 638551
rect 42904 634786 43024 634814
rect 42892 627224 42944 627230
rect 42892 627166 42944 627172
rect 42904 624714 42932 627166
rect 42892 624708 42944 624714
rect 42892 624650 42944 624656
rect 42524 620968 42576 620974
rect 42524 620910 42576 620916
rect 42800 620968 42852 620974
rect 42800 620910 42852 620916
rect 42064 620832 42116 620838
rect 42064 620774 42116 620780
rect 42076 620500 42104 620774
rect 42064 620356 42116 620362
rect 42064 620298 42116 620304
rect 42076 619956 42104 620298
rect 42246 619032 42302 619041
rect 42246 618967 42302 618976
rect 42156 617908 42208 617914
rect 42156 617850 42208 617856
rect 42168 617440 42196 617850
rect 42064 617160 42116 617166
rect 42064 617102 42116 617108
rect 42076 616828 42104 617102
rect 42154 616720 42210 616729
rect 42154 616655 42210 616664
rect 42168 616148 42196 616655
rect 42260 615618 42288 618967
rect 42536 617914 42564 620910
rect 42996 620362 43024 634786
rect 42984 620356 43036 620362
rect 42984 620298 43036 620304
rect 42524 617908 42576 617914
rect 42524 617850 42576 617856
rect 42524 617772 42576 617778
rect 42524 617714 42576 617720
rect 42536 617166 42564 617714
rect 42524 617160 42576 617166
rect 42524 617102 42576 617108
rect 42522 616856 42578 616865
rect 42522 616791 42578 616800
rect 42182 615590 42288 615618
rect 42536 614242 42564 616791
rect 42156 614236 42208 614242
rect 42156 614178 42208 614184
rect 42524 614236 42576 614242
rect 42524 614178 42576 614184
rect 42168 613768 42196 614178
rect 42522 614136 42578 614145
rect 42522 614071 42578 614080
rect 41786 613456 41842 613465
rect 41786 613391 41842 613400
rect 41800 613121 41828 613391
rect 42536 612814 42564 614071
rect 42156 612808 42208 612814
rect 42156 612750 42208 612756
rect 42524 612808 42576 612814
rect 42524 612750 42576 612756
rect 42168 612476 42196 612750
rect 8588 602276 8616 602412
rect 9048 602276 9076 602412
rect 9508 602276 9536 602412
rect 9968 602276 9996 602412
rect 10428 602276 10456 602412
rect 10888 602276 10916 602412
rect 11348 602276 11376 602412
rect 11808 602276 11836 602412
rect 12268 602276 12296 602412
rect 12728 602276 12756 602412
rect 13188 602276 13216 602412
rect 13648 602276 13676 602412
rect 14108 602276 14136 602412
rect 35806 601896 35862 601905
rect 35806 601831 35862 601840
rect 35820 601730 35848 601831
rect 35808 601724 35860 601730
rect 35808 601666 35860 601672
rect 35716 601656 35768 601662
rect 35716 601598 35768 601604
rect 35624 601520 35676 601526
rect 35624 601462 35676 601468
rect 35636 600681 35664 601462
rect 35728 601089 35756 601598
rect 35806 601488 35862 601497
rect 35806 601423 35862 601432
rect 35820 601390 35848 601423
rect 35808 601384 35860 601390
rect 35808 601326 35860 601332
rect 35714 601080 35770 601089
rect 35714 601015 35770 601024
rect 35622 600672 35678 600681
rect 35622 600607 35678 600616
rect 42798 599312 42854 599321
rect 42798 599247 42854 599256
rect 39302 597000 39358 597009
rect 39302 596935 39358 596944
rect 31666 594960 31722 594969
rect 31666 594895 31722 594904
rect 33782 594960 33838 594969
rect 33782 594895 33838 594904
rect 31680 587217 31708 594895
rect 32402 593328 32458 593337
rect 32402 593263 32458 593272
rect 31666 587208 31722 587217
rect 31666 587143 31722 587152
rect 32416 585818 32444 593263
rect 33796 585954 33824 594895
rect 33784 585948 33836 585954
rect 33784 585890 33836 585896
rect 32404 585812 32456 585818
rect 32404 585754 32456 585760
rect 39316 585177 39344 596935
rect 40866 596592 40922 596601
rect 40866 596527 40922 596536
rect 40682 596184 40738 596193
rect 40682 596119 40738 596128
rect 39302 585168 39358 585177
rect 39302 585103 39358 585112
rect 40696 584653 40724 596119
rect 40880 585449 40908 596527
rect 42062 596048 42118 596057
rect 42062 595983 42118 595992
rect 41510 591288 41566 591297
rect 41510 591223 41566 591232
rect 41524 590073 41552 591223
rect 41510 590064 41566 590073
rect 41510 589999 41566 590008
rect 41524 589966 41552 589999
rect 41512 589960 41564 589966
rect 41512 589902 41564 589908
rect 41880 585948 41932 585954
rect 41880 585890 41932 585896
rect 41604 585812 41656 585818
rect 41604 585754 41656 585760
rect 40866 585440 40922 585449
rect 40866 585375 40922 585384
rect 40682 584644 40738 584653
rect 40682 584579 40738 584588
rect 41616 584517 41644 585754
rect 41602 584508 41658 584517
rect 41602 584443 41658 584452
rect 41892 584254 41920 585890
rect 42076 584254 42104 595983
rect 42154 594008 42210 594017
rect 42154 593943 42210 593952
rect 41880 584248 41932 584254
rect 41880 584190 41932 584196
rect 42064 584248 42116 584254
rect 42168 584225 42196 593943
rect 42708 584248 42760 584254
rect 42064 584190 42116 584196
rect 42154 584216 42210 584225
rect 42708 584190 42760 584196
rect 42154 584151 42210 584160
rect 41880 583976 41932 583982
rect 41880 583918 41932 583924
rect 41892 583440 41920 583918
rect 41786 581768 41842 581777
rect 41786 581703 41842 581712
rect 41800 581604 41828 581703
rect 42156 581324 42208 581330
rect 42156 581266 42208 581272
rect 42168 580961 42196 581266
rect 41786 580272 41842 580281
rect 41786 580207 41842 580216
rect 41800 579768 41828 580207
rect 41786 579048 41842 579057
rect 41786 578983 41842 578992
rect 41800 578544 41828 578983
rect 42156 578468 42208 578474
rect 42156 578410 42208 578416
rect 42168 577932 42196 578410
rect 41786 577552 41842 577561
rect 41786 577487 41842 577496
rect 41800 577281 41828 577487
rect 42156 576972 42208 576978
rect 42156 576914 42208 576920
rect 42168 576708 42196 576914
rect 42156 576632 42208 576638
rect 42156 576574 42208 576580
rect 42168 576230 42196 576574
rect 42720 576434 42748 584190
rect 42708 576428 42760 576434
rect 42708 576370 42760 576376
rect 42432 576360 42484 576366
rect 42432 576302 42484 576308
rect 42156 576224 42208 576230
rect 42156 576166 42208 576172
rect 42340 576020 42392 576026
rect 42340 575962 42392 575968
rect 42352 574734 42380 575962
rect 42156 574728 42208 574734
rect 42156 574670 42208 574676
rect 42340 574728 42392 574734
rect 42340 574670 42392 574676
rect 42168 574260 42196 574670
rect 42444 574546 42472 576302
rect 42352 574518 42472 574546
rect 42352 574190 42380 574518
rect 42340 574184 42392 574190
rect 42340 574126 42392 574132
rect 42708 574184 42760 574190
rect 42708 574126 42760 574132
rect 42338 574016 42394 574025
rect 42338 573951 42394 573960
rect 42154 573880 42210 573889
rect 42154 573815 42210 573824
rect 42168 573580 42196 573815
rect 42156 573504 42208 573510
rect 42156 573446 42208 573452
rect 42168 572968 42196 573446
rect 41972 572756 42024 572762
rect 41972 572698 42024 572704
rect 41984 572424 42012 572698
rect 42352 571538 42380 573951
rect 42720 572762 42748 574126
rect 42708 572756 42760 572762
rect 42708 572698 42760 572704
rect 42706 571568 42762 571577
rect 42340 571532 42392 571538
rect 42706 571503 42762 571512
rect 42340 571474 42392 571480
rect 42064 570920 42116 570926
rect 42064 570862 42116 570868
rect 42076 570588 42104 570862
rect 42154 570480 42210 570489
rect 42154 570415 42210 570424
rect 42168 569908 42196 570415
rect 42720 569634 42748 571503
rect 42064 569628 42116 569634
rect 42064 569570 42116 569576
rect 42708 569628 42760 569634
rect 42708 569570 42760 569576
rect 42076 569296 42104 569570
rect 35624 566500 35676 566506
rect 35624 566442 35676 566448
rect 8588 559164 8616 559300
rect 9048 559164 9076 559300
rect 9508 559164 9536 559300
rect 9968 559164 9996 559300
rect 10428 559164 10456 559300
rect 10888 559164 10916 559300
rect 11348 559164 11376 559300
rect 11808 559164 11836 559300
rect 12268 559164 12296 559300
rect 12728 559164 12756 559300
rect 13188 559164 13216 559300
rect 13648 559164 13676 559300
rect 14108 559164 14136 559300
rect 35636 558385 35664 566442
rect 35622 558376 35678 558385
rect 35806 558376 35862 558385
rect 35622 558311 35678 558320
rect 35716 558340 35768 558346
rect 35806 558311 35862 558320
rect 35716 558282 35768 558288
rect 35728 557977 35756 558282
rect 35820 558210 35848 558311
rect 35808 558204 35860 558210
rect 35808 558146 35860 558152
rect 35714 557968 35770 557977
rect 35714 557903 35770 557912
rect 42812 556481 42840 599247
rect 42890 594416 42946 594425
rect 42890 594351 42946 594360
rect 42904 573510 42932 594351
rect 42984 579692 43036 579698
rect 42984 579634 43036 579640
rect 42996 578474 43024 579634
rect 42984 578468 43036 578474
rect 42984 578410 43036 578416
rect 42984 578264 43036 578270
rect 42984 578206 43036 578212
rect 42996 576978 43024 578206
rect 42984 576972 43036 576978
rect 42984 576914 43036 576920
rect 42892 573504 42944 573510
rect 42892 573446 42944 573452
rect 42798 556472 42854 556481
rect 42798 556407 42854 556416
rect 42798 556064 42854 556073
rect 42798 555999 42854 556008
rect 40866 553888 40922 553897
rect 40866 553823 40922 553832
rect 40682 553480 40738 553489
rect 40682 553415 40738 553424
rect 32402 552664 32458 552673
rect 32402 552599 32458 552608
rect 31022 551848 31078 551857
rect 31022 551783 31078 551792
rect 31036 543046 31064 551783
rect 31666 548176 31722 548185
rect 31666 548111 31722 548120
rect 31680 547194 31708 548111
rect 31668 547188 31720 547194
rect 31668 547130 31720 547136
rect 31024 543040 31076 543046
rect 31024 542982 31076 542988
rect 32416 542881 32444 552599
rect 35808 547188 35860 547194
rect 35808 547130 35860 547136
rect 35820 546961 35848 547130
rect 35806 546952 35862 546961
rect 35806 546887 35862 546896
rect 32402 542872 32458 542881
rect 32402 542807 32458 542816
rect 40696 542366 40724 553415
rect 40774 552256 40830 552265
rect 40774 552191 40830 552200
rect 40684 542360 40736 542366
rect 40788 542337 40816 552191
rect 40880 545193 40908 553823
rect 40958 553072 41014 553081
rect 40958 553007 41014 553016
rect 40866 545184 40922 545193
rect 40866 545119 40922 545128
rect 40972 543017 41000 553007
rect 41788 543040 41840 543046
rect 40958 543008 41014 543017
rect 41788 542982 41840 542988
rect 40958 542943 41014 542952
rect 40684 542302 40736 542308
rect 40774 542328 40830 542337
rect 40774 542263 40830 542272
rect 41800 541074 41828 542982
rect 42708 542360 42760 542366
rect 42708 542302 42760 542308
rect 41788 541068 41840 541074
rect 41788 541010 41840 541016
rect 41788 540796 41840 540802
rect 41788 540738 41840 540744
rect 41800 540260 41828 540738
rect 42720 538966 42748 542302
rect 42064 538960 42116 538966
rect 42064 538902 42116 538908
rect 42708 538960 42760 538966
rect 42708 538902 42760 538908
rect 42076 538424 42104 538902
rect 42156 538280 42208 538286
rect 42156 538222 42208 538228
rect 42168 537744 42196 538222
rect 42064 537124 42116 537130
rect 42064 537066 42116 537072
rect 42076 536588 42104 537066
rect 42616 536852 42668 536858
rect 42616 536794 42668 536800
rect 42628 536042 42656 536794
rect 42616 536036 42668 536042
rect 42616 535978 42668 535984
rect 42614 535936 42670 535945
rect 42614 535871 42670 535880
rect 42156 535832 42208 535838
rect 42156 535774 42208 535780
rect 42168 535364 42196 535774
rect 42064 535288 42116 535294
rect 42064 535230 42116 535236
rect 42076 534752 42104 535230
rect 41786 534576 41842 534585
rect 41786 534511 41842 534520
rect 41800 534072 41828 534511
rect 42628 534002 42656 535871
rect 42156 533996 42208 534002
rect 42156 533938 42208 533944
rect 42616 533996 42668 534002
rect 42616 533938 42668 533944
rect 42168 533528 42196 533938
rect 42614 533896 42670 533905
rect 42614 533831 42670 533840
rect 42338 532672 42394 532681
rect 42338 532607 42394 532616
rect 41786 531448 41842 531457
rect 41786 531383 41842 531392
rect 41800 531045 41828 531383
rect 42156 530936 42208 530942
rect 42156 530878 42208 530884
rect 42168 530400 42196 530878
rect 42156 530120 42208 530126
rect 42156 530062 42208 530068
rect 42168 529757 42196 530062
rect 42352 529650 42380 532607
rect 42628 530942 42656 533831
rect 42616 530936 42668 530942
rect 42616 530878 42668 530884
rect 42616 530800 42668 530806
rect 42616 530742 42668 530748
rect 42628 530126 42656 530742
rect 42616 530120 42668 530126
rect 42616 530062 42668 530068
rect 42340 529644 42392 529650
rect 42340 529586 42392 529592
rect 42338 529544 42394 529553
rect 42156 529508 42208 529514
rect 42338 529479 42394 529488
rect 42156 529450 42208 529456
rect 42168 529205 42196 529450
rect 42076 527270 42104 527340
rect 42352 527270 42380 529479
rect 42614 529408 42670 529417
rect 42614 529343 42670 529352
rect 42064 527264 42116 527270
rect 42064 527206 42116 527212
rect 42340 527264 42392 527270
rect 42340 527206 42392 527212
rect 42156 527196 42208 527202
rect 42156 527138 42208 527144
rect 42168 526728 42196 527138
rect 42628 526658 42656 529343
rect 42156 526652 42208 526658
rect 42156 526594 42208 526600
rect 42616 526652 42668 526658
rect 42616 526594 42668 526600
rect 42168 526077 42196 526594
rect 40684 518968 40736 518974
rect 40684 518910 40736 518916
rect 40696 432614 40724 518910
rect 40684 432608 40736 432614
rect 40684 432550 40736 432556
rect 41788 432608 41840 432614
rect 41788 432550 41840 432556
rect 8588 431596 8616 431664
rect 9048 431596 9076 431664
rect 9508 431596 9536 431664
rect 9968 431596 9996 431664
rect 10428 431596 10456 431664
rect 10888 431596 10916 431664
rect 11348 431596 11376 431664
rect 11808 431596 11836 431664
rect 12268 431596 12296 431664
rect 12728 431596 12756 431664
rect 13188 431596 13216 431664
rect 13648 431596 13676 431664
rect 14108 431596 14136 431664
rect 41800 430545 41828 432550
rect 41786 430536 41842 430545
rect 41786 430471 41842 430480
rect 42812 428913 42840 555999
rect 42890 551576 42946 551585
rect 42890 551511 42946 551520
rect 42904 527202 42932 551511
rect 43074 549944 43130 549953
rect 43074 549879 43130 549888
rect 42984 540252 43036 540258
rect 42984 540194 43036 540200
rect 42996 538422 43024 540194
rect 42984 538416 43036 538422
rect 42984 538358 43036 538364
rect 42984 538280 43036 538286
rect 42984 538222 43036 538228
rect 42996 537130 43024 538222
rect 42984 537124 43036 537130
rect 42984 537066 43036 537072
rect 43088 535294 43116 549879
rect 43076 535288 43128 535294
rect 43076 535230 43128 535236
rect 42892 527196 42944 527202
rect 42892 527138 42944 527144
rect 43166 430944 43222 430953
rect 43166 430879 43222 430888
rect 43180 430642 43208 430879
rect 43168 430636 43220 430642
rect 43168 430578 43220 430584
rect 42798 428904 42854 428913
rect 42798 428839 42854 428848
rect 42798 428496 42854 428505
rect 42798 428431 42854 428440
rect 32402 426048 32458 426057
rect 32402 425983 32458 425992
rect 31022 422376 31078 422385
rect 31022 422311 31078 422320
rect 31036 414730 31064 422311
rect 31024 414724 31076 414730
rect 31024 414666 31076 414672
rect 32416 414633 32444 425983
rect 35162 425232 35218 425241
rect 35162 425167 35218 425176
rect 32494 424416 32550 424425
rect 32494 424351 32550 424360
rect 32508 414866 32536 424351
rect 32496 414860 32548 414866
rect 32496 414802 32548 414808
rect 35176 414769 35204 425167
rect 41786 419520 41842 419529
rect 41786 419455 41788 419464
rect 41840 419455 41842 419464
rect 41788 419426 41840 419432
rect 41880 414860 41932 414866
rect 41880 414802 41932 414808
rect 35162 414760 35218 414769
rect 35162 414695 35218 414704
rect 32402 414624 32458 414633
rect 32402 414559 32458 414568
rect 41892 413438 41920 414802
rect 42524 414724 42576 414730
rect 42524 414666 42576 414672
rect 41880 413432 41932 413438
rect 41880 413374 41932 413380
rect 41880 413160 41932 413166
rect 41880 413102 41932 413108
rect 41892 412624 41920 413102
rect 41878 411224 41934 411233
rect 41878 411159 41934 411168
rect 41892 410788 41920 411159
rect 42156 410712 42208 410718
rect 42156 410654 42208 410660
rect 42168 410176 42196 410654
rect 41786 409456 41842 409465
rect 41786 409391 41842 409400
rect 41800 408952 41828 409391
rect 42064 408196 42116 408202
rect 42064 408138 42116 408144
rect 42076 407796 42104 408138
rect 42536 407658 42564 414666
rect 42156 407652 42208 407658
rect 42156 407594 42208 407600
rect 42524 407652 42576 407658
rect 42524 407594 42576 407600
rect 42168 407116 42196 407594
rect 42064 406836 42116 406842
rect 42064 406778 42116 406784
rect 42076 406504 42104 406778
rect 41786 406328 41842 406337
rect 41786 406263 41842 406272
rect 41800 405929 41828 406263
rect 42156 403912 42208 403918
rect 42156 403854 42208 403860
rect 42168 403444 42196 403854
rect 42156 402960 42208 402966
rect 42156 402902 42208 402908
rect 42168 402801 42196 402902
rect 42062 402520 42118 402529
rect 42062 402455 42118 402464
rect 42076 402152 42104 402455
rect 41786 401840 41842 401849
rect 41786 401775 41842 401784
rect 41800 401608 41828 401775
rect 41786 400072 41842 400081
rect 41786 400007 41842 400016
rect 41800 399772 41828 400007
rect 41786 399664 41842 399673
rect 41786 399599 41842 399608
rect 41800 399121 41828 399599
rect 41786 398848 41842 398857
rect 41786 398783 41842 398792
rect 41800 398480 41828 398783
rect 8588 388348 8616 388484
rect 9048 388348 9076 388484
rect 9508 388348 9536 388484
rect 9968 388348 9996 388484
rect 10428 388348 10456 388484
rect 10888 388348 10916 388484
rect 11348 388348 11376 388484
rect 11808 388348 11836 388484
rect 12268 388348 12296 388484
rect 12728 388348 12756 388484
rect 13188 388348 13216 388484
rect 13648 388348 13676 388484
rect 14108 388348 14136 388484
rect 35716 387796 35768 387802
rect 35716 387738 35768 387744
rect 35624 387524 35676 387530
rect 35624 387466 35676 387472
rect 35636 387161 35664 387466
rect 35622 387152 35678 387161
rect 35622 387087 35678 387096
rect 35728 386753 35756 387738
rect 35808 387660 35860 387666
rect 35808 387602 35860 387608
rect 35820 387569 35848 387602
rect 35806 387560 35862 387569
rect 35806 387495 35862 387504
rect 35808 387388 35860 387394
rect 35808 387330 35860 387336
rect 35820 387161 35848 387330
rect 35806 387152 35862 387161
rect 35806 387087 35862 387096
rect 35714 386744 35770 386753
rect 35714 386679 35770 386688
rect 42812 385665 42840 428431
rect 42890 423192 42946 423201
rect 42890 423127 42946 423136
rect 42904 402966 42932 423127
rect 42982 421560 43038 421569
rect 42982 421495 43038 421504
rect 42996 406842 43024 421495
rect 42984 406836 43036 406842
rect 42984 406778 43036 406784
rect 42892 402960 42944 402966
rect 42892 402902 42944 402908
rect 42798 385656 42854 385665
rect 42798 385591 42854 385600
rect 42798 383616 42854 383625
rect 42798 383551 42854 383560
rect 40866 382664 40922 382673
rect 40866 382599 40922 382608
rect 37922 381440 37978 381449
rect 37922 381375 37978 381384
rect 31022 381032 31078 381041
rect 31022 380967 31078 380976
rect 31036 371890 31064 380967
rect 33782 378176 33838 378185
rect 33782 378111 33838 378120
rect 33796 371929 33824 378111
rect 35806 377360 35862 377369
rect 35806 377295 35862 377304
rect 35820 376106 35848 377295
rect 35808 376100 35860 376106
rect 35808 376042 35860 376048
rect 33782 371920 33838 371929
rect 31024 371884 31076 371890
rect 33782 371855 33838 371864
rect 31024 371826 31076 371832
rect 37936 371385 37964 381375
rect 40682 379400 40738 379409
rect 40682 379335 40738 379344
rect 37922 371376 37978 371385
rect 37922 371311 37978 371320
rect 40696 370598 40724 379335
rect 40880 371278 40908 382599
rect 41510 376136 41566 376145
rect 41510 376071 41512 376080
rect 41564 376071 41566 376080
rect 41512 376042 41564 376048
rect 42340 371884 42392 371890
rect 42340 371826 42392 371832
rect 40868 371272 40920 371278
rect 40868 371214 40920 371220
rect 40684 370592 40736 370598
rect 40684 370534 40736 370540
rect 41788 370592 41840 370598
rect 41788 370534 41840 370540
rect 41800 370297 41828 370534
rect 41786 370288 41842 370297
rect 41786 370223 41842 370232
rect 42352 369714 42380 371826
rect 42708 371272 42760 371278
rect 42708 371214 42760 371220
rect 42156 369708 42208 369714
rect 42156 369650 42208 369656
rect 42340 369708 42392 369714
rect 42340 369650 42392 369656
rect 42168 369444 42196 369650
rect 42720 368150 42748 371214
rect 42156 368144 42208 368150
rect 42156 368086 42208 368092
rect 42708 368144 42760 368150
rect 42708 368086 42760 368092
rect 42168 367608 42196 368086
rect 42168 366858 42196 366961
rect 42156 366852 42208 366858
rect 42156 366794 42208 366800
rect 42708 366852 42760 366858
rect 42708 366794 42760 366800
rect 41878 366344 41934 366353
rect 41878 366279 41934 366288
rect 41892 365772 41920 366279
rect 42156 365016 42208 365022
rect 42156 364958 42208 364964
rect 42168 364548 42196 364958
rect 42156 364336 42208 364342
rect 42156 364278 42208 364284
rect 42168 363936 42196 364278
rect 42720 364274 42748 366794
rect 42708 364268 42760 364274
rect 42708 364210 42760 364216
rect 41970 363760 42026 363769
rect 41970 363695 42026 363704
rect 41984 363256 42012 363695
rect 41786 362944 41842 362953
rect 41786 362879 41842 362888
rect 41800 362712 41828 362879
rect 42064 360732 42116 360738
rect 42064 360674 42116 360680
rect 42076 360264 42104 360674
rect 41786 360088 41842 360097
rect 41786 360023 41842 360032
rect 41800 359584 41828 360023
rect 42156 359508 42208 359514
rect 42156 359450 42208 359456
rect 42168 358972 42196 359450
rect 41786 358728 41842 358737
rect 41786 358663 41842 358672
rect 41800 358428 41828 358663
rect 41786 356960 41842 356969
rect 41786 356895 41842 356904
rect 41800 356592 41828 356895
rect 42156 356040 42208 356046
rect 42156 355982 42208 355988
rect 42168 355912 42196 355982
rect 41786 355736 41842 355745
rect 41786 355671 41842 355680
rect 41800 355300 41828 355671
rect 27620 351212 27672 351218
rect 27620 351154 27672 351160
rect 8588 345100 8616 345236
rect 9048 345100 9076 345236
rect 9508 345100 9536 345236
rect 9968 345100 9996 345236
rect 10428 345100 10456 345236
rect 10888 345100 10916 345236
rect 11348 345100 11376 345236
rect 11808 345100 11836 345236
rect 12268 345100 12296 345236
rect 12728 345100 12756 345236
rect 13188 345100 13216 345236
rect 13648 345100 13676 345236
rect 14108 345100 14136 345236
rect 27632 344729 27660 351154
rect 27618 344720 27674 344729
rect 27618 344655 27674 344664
rect 35716 344344 35768 344350
rect 35716 344286 35768 344292
rect 35806 344312 35862 344321
rect 35728 343913 35756 344286
rect 35806 344247 35862 344256
rect 35820 344214 35848 344247
rect 35808 344208 35860 344214
rect 35808 344150 35860 344156
rect 35714 343904 35770 343913
rect 35714 343839 35770 343848
rect 42812 340921 42840 383551
rect 43166 380760 43222 380769
rect 43166 380695 43222 380704
rect 42982 380352 43038 380361
rect 42982 380287 43038 380296
rect 42996 359514 43024 380287
rect 43074 378720 43130 378729
rect 43074 378655 43130 378664
rect 43088 360738 43116 378655
rect 43076 360732 43128 360738
rect 43076 360674 43128 360680
rect 42984 359508 43036 359514
rect 42984 359450 43036 359456
rect 43180 356046 43208 380695
rect 43168 356040 43220 356046
rect 43168 355982 43220 355988
rect 42890 341320 42946 341329
rect 42890 341255 42946 341264
rect 42798 340912 42854 340921
rect 42798 340847 42854 340856
rect 42798 340504 42854 340513
rect 42798 340439 42854 340448
rect 31022 339416 31078 339425
rect 31022 339351 31078 339360
rect 30378 334112 30434 334121
rect 30378 334047 30434 334056
rect 30392 333305 30420 334047
rect 30378 333296 30434 333305
rect 30378 333231 30380 333240
rect 30432 333231 30434 333240
rect 30380 333202 30432 333208
rect 30392 333171 30420 333202
rect 31036 327729 31064 339351
rect 32402 338192 32458 338201
rect 32402 338127 32458 338136
rect 32416 327865 32444 338127
rect 32402 327856 32458 327865
rect 32402 327791 32458 327800
rect 31022 327720 31078 327729
rect 31022 327655 31078 327664
rect 42064 326800 42116 326806
rect 42064 326742 42116 326748
rect 42076 326264 42104 326742
rect 41786 324864 41842 324873
rect 41786 324799 41842 324808
rect 41800 324428 41828 324799
rect 42168 323338 42196 323748
rect 42156 323332 42208 323338
rect 42156 323274 42208 323280
rect 42616 323332 42668 323338
rect 42616 323274 42668 323280
rect 42064 322924 42116 322930
rect 42064 322866 42116 322872
rect 42076 322592 42104 322866
rect 42628 321570 42656 323274
rect 42616 321564 42668 321570
rect 42616 321506 42668 321512
rect 42156 321496 42208 321502
rect 42156 321438 42208 321444
rect 42168 321368 42196 321438
rect 41786 321192 41842 321201
rect 41786 321127 41842 321136
rect 41800 320725 41828 321127
rect 42168 320006 42196 320076
rect 42156 320000 42208 320006
rect 41786 319968 41842 319977
rect 42156 319942 42208 319948
rect 41786 319903 41842 319912
rect 41800 319532 41828 319903
rect 41786 317384 41842 317393
rect 41786 317319 41842 317328
rect 41800 317045 41828 317319
rect 42156 316736 42208 316742
rect 42156 316678 42208 316684
rect 42168 316404 42196 316678
rect 41786 315888 41842 315897
rect 41786 315823 41842 315832
rect 41800 315757 41828 315823
rect 41970 315480 42026 315489
rect 41970 315415 42026 315424
rect 41984 315180 42012 315415
rect 41878 313848 41934 313857
rect 41878 313783 41934 313792
rect 41892 313344 41920 313783
rect 41786 313168 41842 313177
rect 41786 313103 41842 313112
rect 41800 312732 41828 313103
rect 41786 312352 41842 312361
rect 41786 312287 41842 312296
rect 41800 312052 41828 312287
rect 8588 301988 8616 302124
rect 9048 301988 9076 302124
rect 9508 301988 9536 302124
rect 9968 301988 9996 302124
rect 10428 301988 10456 302124
rect 10888 301988 10916 302124
rect 11348 301988 11376 302124
rect 11808 301988 11836 302124
rect 12268 301988 12296 302124
rect 12728 301988 12756 302124
rect 13188 301988 13216 302124
rect 13648 301988 13676 302124
rect 14108 301988 14136 302124
rect 35806 301608 35862 301617
rect 35806 301543 35862 301552
rect 35820 301102 35848 301543
rect 35808 301096 35860 301102
rect 35808 301038 35860 301044
rect 35808 300960 35860 300966
rect 35806 300928 35808 300937
rect 35860 300928 35862 300937
rect 35806 300863 35862 300872
rect 42812 297673 42840 340439
rect 42904 298489 42932 341255
rect 42982 336832 43038 336841
rect 42982 336767 43038 336776
rect 42996 316742 43024 336767
rect 43074 335200 43130 335209
rect 43074 335135 43130 335144
rect 43088 320006 43116 335135
rect 43076 320000 43128 320006
rect 43076 319942 43128 319948
rect 42984 316736 43036 316742
rect 42984 316678 43036 316684
rect 42890 298480 42946 298489
rect 42890 298415 42946 298424
rect 42798 297664 42854 297673
rect 42798 297599 42854 297608
rect 42798 297256 42854 297265
rect 42798 297191 42854 297200
rect 35162 296440 35218 296449
rect 35162 296375 35218 296384
rect 32402 294808 32458 294817
rect 32402 294743 32458 294752
rect 32416 284986 32444 294743
rect 32404 284980 32456 284986
rect 32404 284922 32456 284928
rect 35176 284889 35204 296375
rect 41880 284980 41932 284986
rect 41880 284922 41932 284928
rect 35162 284880 35218 284889
rect 35162 284815 35218 284824
rect 41892 283830 41920 284922
rect 41880 283824 41932 283830
rect 41880 283766 41932 283772
rect 41880 283620 41932 283626
rect 41880 283562 41932 283568
rect 41892 283045 41920 283562
rect 41786 281480 41842 281489
rect 41786 281415 41842 281424
rect 41800 281180 41828 281415
rect 42168 280226 42196 280568
rect 42156 280220 42208 280226
rect 42156 280162 42208 280168
rect 41786 279848 41842 279857
rect 41786 279783 41842 279792
rect 41800 279344 41828 279783
rect 42064 278656 42116 278662
rect 42064 278598 42116 278604
rect 42076 278188 42104 278598
rect 41786 278080 41842 278089
rect 41786 278015 41842 278024
rect 41800 277508 41828 278015
rect 42156 277160 42208 277166
rect 42156 277102 42208 277108
rect 42168 276896 42196 277102
rect 42064 276752 42116 276758
rect 42064 276694 42116 276700
rect 42076 276352 42104 276694
rect 42156 274304 42208 274310
rect 42156 274246 42208 274252
rect 42168 273836 42196 274246
rect 42168 273086 42196 273224
rect 42156 273080 42208 273086
rect 41786 273048 41842 273057
rect 42156 273022 42208 273028
rect 41786 272983 41842 272992
rect 41800 272544 41828 272983
rect 41786 272232 41842 272241
rect 41786 272167 41842 272176
rect 41800 272000 41828 272167
rect 41970 270464 42026 270473
rect 41970 270399 42026 270408
rect 41984 270164 42012 270399
rect 41786 269784 41842 269793
rect 41786 269719 41842 269728
rect 41800 269521 41828 269719
rect 41786 269104 41842 269113
rect 41786 269039 41842 269048
rect 41800 268872 41828 269039
rect 28356 265668 28408 265674
rect 28356 265610 28408 265616
rect 8588 258740 8616 258876
rect 9048 258740 9076 258876
rect 9508 258740 9536 258876
rect 9968 258740 9996 258876
rect 10428 258740 10456 258876
rect 10888 258740 10916 258876
rect 11348 258740 11376 258876
rect 11808 258740 11836 258876
rect 12268 258740 12296 258876
rect 12728 258740 12756 258876
rect 13188 258740 13216 258876
rect 13648 258740 13676 258876
rect 14108 258740 14136 258876
rect 28368 258369 28396 265610
rect 28354 258360 28410 258369
rect 28354 258295 28410 258304
rect 31576 258052 31628 258058
rect 31576 257994 31628 258000
rect 31484 257916 31536 257922
rect 31484 257858 31536 257864
rect 31496 257553 31524 257858
rect 31482 257544 31538 257553
rect 31482 257479 31538 257488
rect 31588 257145 31616 257994
rect 31668 257780 31720 257786
rect 31668 257722 31720 257728
rect 31680 257553 31708 257722
rect 31666 257544 31722 257553
rect 31666 257479 31722 257488
rect 31574 257136 31630 257145
rect 31574 257071 31630 257080
rect 42812 254425 42840 297191
rect 42890 295216 42946 295225
rect 42890 295151 42946 295160
rect 42904 276758 42932 295151
rect 42982 292360 43038 292369
rect 42982 292295 43038 292304
rect 42892 276752 42944 276758
rect 42892 276694 42944 276700
rect 42996 274310 43024 292295
rect 43166 291952 43222 291961
rect 43166 291887 43222 291896
rect 43180 277166 43208 291887
rect 43456 278254 43484 932039
rect 62118 923808 62174 923817
rect 62118 923743 62174 923752
rect 62132 923302 62160 923743
rect 51724 923296 51776 923302
rect 51724 923238 51776 923244
rect 62120 923296 62172 923302
rect 62120 923238 62172 923244
rect 44824 884672 44876 884678
rect 44824 884614 44876 884620
rect 43628 858424 43680 858430
rect 43628 858366 43680 858372
rect 43534 806304 43590 806313
rect 43534 806239 43590 806248
rect 43444 278248 43496 278254
rect 43444 278190 43496 278196
rect 43168 277160 43220 277166
rect 43168 277102 43220 277108
rect 42984 274304 43036 274310
rect 42984 274246 43036 274252
rect 42890 256456 42946 256465
rect 42890 256391 42946 256400
rect 42798 254416 42854 254425
rect 42798 254351 42854 254360
rect 31022 253464 31078 253473
rect 31022 253399 31078 253408
rect 31036 242214 31064 253399
rect 32402 253056 32458 253065
rect 32402 252991 32458 253000
rect 31114 252240 31170 252249
rect 31114 252175 31170 252184
rect 31128 242282 31156 252175
rect 32416 242350 32444 252991
rect 35806 246528 35862 246537
rect 35806 246463 35862 246472
rect 35820 245682 35848 246463
rect 35808 245676 35860 245682
rect 35808 245618 35860 245624
rect 32404 242344 32456 242350
rect 32404 242286 32456 242292
rect 41972 242344 42024 242350
rect 41972 242286 42024 242292
rect 31116 242276 31168 242282
rect 31116 242218 31168 242224
rect 31024 242208 31076 242214
rect 31024 242150 31076 242156
rect 41984 240689 42012 242286
rect 42432 242276 42484 242282
rect 42432 242218 42484 242224
rect 41970 240680 42026 240689
rect 41970 240615 42026 240624
rect 42444 240106 42472 242218
rect 42708 242208 42760 242214
rect 42708 242150 42760 242156
rect 42432 240100 42484 240106
rect 42432 240042 42484 240048
rect 42156 240032 42208 240038
rect 42156 239974 42208 239980
rect 42168 239836 42196 239974
rect 42720 238785 42748 242150
rect 42800 240100 42852 240106
rect 42800 240042 42852 240048
rect 42706 238776 42762 238785
rect 42706 238711 42762 238720
rect 42812 238626 42840 240042
rect 42720 238598 42840 238626
rect 41970 238504 42026 238513
rect 41970 238439 42026 238448
rect 41984 238000 42012 238439
rect 42720 237425 42748 238598
rect 42706 237416 42762 237425
rect 42706 237351 42762 237360
rect 41786 236736 41842 236745
rect 41786 236671 41842 236680
rect 41800 236164 41828 236671
rect 42156 235408 42208 235414
rect 42156 235350 42208 235356
rect 42168 234969 42196 235350
rect 42156 234592 42208 234598
rect 42156 234534 42208 234540
rect 42168 234328 42196 234534
rect 42156 234048 42208 234054
rect 42156 233990 42208 233996
rect 42168 233681 42196 233990
rect 42156 233300 42208 233306
rect 42156 233242 42208 233248
rect 42168 233104 42196 233242
rect 42430 232928 42486 232937
rect 42430 232863 42486 232872
rect 42156 231124 42208 231130
rect 42156 231066 42208 231072
rect 42168 230656 42196 231066
rect 42444 230586 42472 232863
rect 42156 230580 42208 230586
rect 42156 230522 42208 230528
rect 42432 230580 42484 230586
rect 42432 230522 42484 230528
rect 42168 229976 42196 230522
rect 42156 229900 42208 229906
rect 42156 229842 42208 229848
rect 42168 229364 42196 229842
rect 42154 228984 42210 228993
rect 42154 228919 42210 228928
rect 42168 228820 42196 228919
rect 41970 227352 42026 227361
rect 41970 227287 42026 227296
rect 41984 226984 42012 227287
rect 42156 226704 42208 226710
rect 42156 226646 42208 226652
rect 42168 226304 42196 226646
rect 42156 226228 42208 226234
rect 42156 226170 42208 226176
rect 42168 225692 42196 226170
rect 28724 221468 28776 221474
rect 28724 221410 28776 221416
rect 8588 215492 8616 215628
rect 9048 215492 9076 215628
rect 9508 215492 9536 215628
rect 9968 215492 9996 215628
rect 10428 215492 10456 215628
rect 10888 215492 10916 215628
rect 11348 215492 11376 215628
rect 11808 215492 11836 215628
rect 12268 215492 12296 215628
rect 12728 215492 12756 215628
rect 13188 215492 13216 215628
rect 13648 215492 13676 215628
rect 14108 215492 14136 215628
rect 28736 215121 28764 221410
rect 35808 217320 35860 217326
rect 35808 217262 35860 217268
rect 28722 215112 28778 215121
rect 28722 215047 28778 215056
rect 35820 214713 35848 217262
rect 35806 214704 35862 214713
rect 35806 214639 35862 214648
rect 35808 214600 35860 214606
rect 35808 214542 35860 214548
rect 35820 214305 35848 214542
rect 35806 214296 35862 214305
rect 35806 214231 35862 214240
rect 41328 214192 41380 214198
rect 41328 214134 41380 214140
rect 31116 214124 31168 214130
rect 31116 214066 31168 214072
rect 31022 210216 31078 210225
rect 31022 210151 31078 210160
rect 31036 199345 31064 210151
rect 31128 204513 31156 214066
rect 31300 214056 31352 214062
rect 31300 213998 31352 214004
rect 31312 204921 31340 213998
rect 41340 211857 41368 214134
rect 41512 213988 41564 213994
rect 41512 213930 41564 213936
rect 41524 213489 41552 213930
rect 42904 213761 42932 256391
rect 43350 255640 43406 255649
rect 43350 255575 43406 255584
rect 42982 252784 43038 252793
rect 42982 252719 43038 252728
rect 42996 226234 43024 252719
rect 43166 251968 43222 251977
rect 43166 251903 43222 251912
rect 43074 250744 43130 250753
rect 43074 250679 43130 250688
rect 43088 229906 43116 250679
rect 43180 233306 43208 251903
rect 43258 249112 43314 249121
rect 43258 249047 43314 249056
rect 43168 233300 43220 233306
rect 43168 233242 43220 233248
rect 43272 231130 43300 249047
rect 43260 231124 43312 231130
rect 43260 231066 43312 231072
rect 43076 229900 43128 229906
rect 43076 229842 43128 229848
rect 42984 226228 43036 226234
rect 42984 226170 43036 226176
rect 42890 213752 42946 213761
rect 42890 213687 42946 213696
rect 41510 213480 41566 213489
rect 41510 213415 41566 213424
rect 43364 212945 43392 255575
rect 43548 231169 43576 806239
rect 43640 773673 43668 858366
rect 44836 817562 44864 884614
rect 50436 832176 50488 832182
rect 50436 832118 50488 832124
rect 47584 818372 47636 818378
rect 47584 818314 47636 818320
rect 44824 817556 44876 817562
rect 44824 817498 44876 817504
rect 44178 815280 44234 815289
rect 44178 815215 44234 815224
rect 43626 773664 43682 773673
rect 43626 773599 43682 773608
rect 44192 772449 44220 815215
rect 44270 813648 44326 813657
rect 44270 813583 44326 813592
rect 44178 772440 44234 772449
rect 44178 772375 44234 772384
rect 44284 770817 44312 813583
rect 44362 809976 44418 809985
rect 44362 809911 44418 809920
rect 44376 793082 44404 809911
rect 44454 808344 44510 808353
rect 44454 808279 44510 808288
rect 44468 794918 44496 808279
rect 44456 794912 44508 794918
rect 44456 794854 44508 794860
rect 44824 793552 44876 793558
rect 44824 793494 44876 793500
rect 44364 793076 44416 793082
rect 44364 793018 44416 793024
rect 44546 772848 44602 772857
rect 44546 772783 44602 772792
rect 44270 770808 44326 770817
rect 44270 770743 44326 770752
rect 44362 767136 44418 767145
rect 44362 767071 44418 767080
rect 43628 753568 43680 753574
rect 43628 753510 43680 753516
rect 43640 696250 43668 753510
rect 44376 747998 44404 767071
rect 44454 765504 44510 765513
rect 44454 765439 44510 765448
rect 44468 749426 44496 765439
rect 44456 749420 44508 749426
rect 44456 749362 44508 749368
rect 44364 747992 44416 747998
rect 44364 747934 44416 747940
rect 44560 731406 44588 772783
rect 44730 770400 44786 770409
rect 44730 770335 44786 770344
rect 44548 731400 44600 731406
rect 44548 731342 44600 731348
rect 44270 728920 44326 728929
rect 44270 728855 44326 728864
rect 44178 721984 44234 721993
rect 44178 721919 44234 721928
rect 44192 709374 44220 721919
rect 44180 709368 44232 709374
rect 44180 709310 44232 709316
rect 43628 696244 43680 696250
rect 43628 696186 43680 696192
rect 43720 688696 43772 688702
rect 43720 688638 43772 688644
rect 43628 647896 43680 647902
rect 43628 647838 43680 647844
rect 43640 601662 43668 647838
rect 43732 644638 43760 688638
rect 44284 686089 44312 728855
rect 44744 727705 44772 770335
rect 44836 731270 44864 793494
rect 44824 731264 44876 731270
rect 44824 731206 44876 731212
rect 44730 727696 44786 727705
rect 44730 727631 44786 727640
rect 44546 727288 44602 727297
rect 44546 727223 44602 727232
rect 44362 724432 44418 724441
rect 44362 724367 44418 724376
rect 44376 701078 44404 724367
rect 44454 722392 44510 722401
rect 44454 722327 44510 722336
rect 44468 706654 44496 722327
rect 44456 706648 44508 706654
rect 44456 706590 44508 706596
rect 44364 701072 44416 701078
rect 44364 701014 44416 701020
rect 44270 686080 44326 686089
rect 44270 686015 44326 686024
rect 44270 685672 44326 685681
rect 44270 685607 44326 685616
rect 44178 679960 44234 679969
rect 44178 679895 44234 679904
rect 44192 666738 44220 679895
rect 44180 666732 44232 666738
rect 44180 666674 44232 666680
rect 43720 644632 43772 644638
rect 43720 644574 43772 644580
rect 44178 643240 44234 643249
rect 44178 643175 44234 643184
rect 43628 601656 43680 601662
rect 43628 601598 43680 601604
rect 44192 601526 44220 643175
rect 44284 643113 44312 685607
rect 44560 684457 44588 727223
rect 47596 712162 47624 818314
rect 50344 805996 50396 806002
rect 50344 805938 50396 805944
rect 48964 767372 49016 767378
rect 48964 767314 49016 767320
rect 47584 712156 47636 712162
rect 47584 712098 47636 712104
rect 44638 686488 44694 686497
rect 44638 686423 44694 686432
rect 44546 684448 44602 684457
rect 44546 684383 44602 684392
rect 44362 684040 44418 684049
rect 44362 683975 44418 683984
rect 44270 643104 44326 643113
rect 44270 643039 44326 643048
rect 44376 641481 44404 683975
rect 44454 678736 44510 678745
rect 44454 678671 44510 678680
rect 44468 665242 44496 678671
rect 44456 665236 44508 665242
rect 44456 665178 44508 665184
rect 44652 643793 44680 686423
rect 48976 670070 49004 767314
rect 50356 731134 50384 805938
rect 50448 773945 50476 832118
rect 51736 799746 51764 923238
rect 62118 910752 62174 910761
rect 62118 910687 62174 910696
rect 62132 909498 62160 910687
rect 62120 909492 62172 909498
rect 62120 909434 62172 909440
rect 62118 897832 62174 897841
rect 62118 897767 62174 897776
rect 62132 897054 62160 897767
rect 53104 897048 53156 897054
rect 53104 896990 53156 896996
rect 62120 897048 62172 897054
rect 62120 896990 62172 896996
rect 53116 817426 53144 896990
rect 62118 884776 62174 884785
rect 62118 884711 62174 884720
rect 62132 884678 62160 884711
rect 62120 884672 62172 884678
rect 62120 884614 62172 884620
rect 62118 871720 62174 871729
rect 62118 871655 62174 871664
rect 62132 870874 62160 871655
rect 55956 870868 56008 870874
rect 55956 870810 56008 870816
rect 62120 870868 62172 870874
rect 62120 870810 62172 870816
rect 54484 844620 54536 844626
rect 54484 844562 54536 844568
rect 53104 817420 53156 817426
rect 53104 817362 53156 817368
rect 51724 799740 51776 799746
rect 51724 799682 51776 799688
rect 51724 779748 51776 779754
rect 51724 779690 51776 779696
rect 50434 773936 50490 773945
rect 50434 773871 50490 773880
rect 50344 731128 50396 731134
rect 50344 731070 50396 731076
rect 51736 730998 51764 779690
rect 54496 774246 54524 844562
rect 54484 774240 54536 774246
rect 54484 774182 54536 774188
rect 55864 761796 55916 761802
rect 55864 761738 55916 761744
rect 54484 741124 54536 741130
rect 54484 741066 54536 741072
rect 51724 730992 51776 730998
rect 51724 730934 51776 730940
rect 51724 727320 51776 727326
rect 51724 727262 51776 727268
rect 50344 719704 50396 719710
rect 50344 719646 50396 719652
rect 48964 670064 49016 670070
rect 48964 670006 49016 670012
rect 47584 662448 47636 662454
rect 47584 662390 47636 662396
rect 44638 643784 44694 643793
rect 44638 643719 44694 643728
rect 44638 642288 44694 642297
rect 44638 642223 44694 642232
rect 44362 641472 44418 641481
rect 44362 641407 44418 641416
rect 44454 636984 44510 636993
rect 44454 636919 44510 636928
rect 44468 618322 44496 636919
rect 44546 635352 44602 635361
rect 44546 635287 44602 635296
rect 44560 622470 44588 635287
rect 44548 622464 44600 622470
rect 44548 622406 44600 622412
rect 44456 618316 44508 618322
rect 44456 618258 44508 618264
rect 44180 601520 44232 601526
rect 44180 601462 44232 601468
rect 44178 600128 44234 600137
rect 44178 600063 44234 600072
rect 43720 571396 43772 571402
rect 43720 571338 43772 571344
rect 43732 566506 43760 571338
rect 43720 566500 43772 566506
rect 43720 566442 43772 566448
rect 44192 557297 44220 600063
rect 44652 599729 44680 642223
rect 44730 640656 44786 640665
rect 44730 640591 44786 640600
rect 44638 599720 44694 599729
rect 44638 599655 44694 599664
rect 44744 598097 44772 640591
rect 44730 598088 44786 598097
rect 44730 598023 44786 598032
rect 44270 597680 44326 597689
rect 44270 597615 44326 597624
rect 44178 557288 44234 557297
rect 44178 557223 44234 557232
rect 44284 554849 44312 597615
rect 44362 595640 44418 595649
rect 44362 595575 44418 595584
rect 44376 578270 44404 595575
rect 44638 593192 44694 593201
rect 44638 593127 44694 593136
rect 44454 592784 44510 592793
rect 44454 592719 44510 592728
rect 44364 578264 44416 578270
rect 44364 578206 44416 578212
rect 44468 576910 44496 592719
rect 44652 579698 44680 593127
rect 47596 581330 47624 662390
rect 48964 610020 49016 610026
rect 48964 609962 49016 609968
rect 47584 581324 47636 581330
rect 47584 581266 47636 581272
rect 44640 579692 44692 579698
rect 44640 579634 44692 579640
rect 44456 576904 44508 576910
rect 44456 576846 44508 576852
rect 47584 557592 47636 557598
rect 47584 557534 47636 557540
rect 44638 556880 44694 556889
rect 44638 556815 44694 556824
rect 44362 555248 44418 555257
rect 44362 555183 44418 555192
rect 44270 554840 44326 554849
rect 44270 554775 44326 554784
rect 44270 554432 44326 554441
rect 44270 554367 44326 554376
rect 44178 550352 44234 550361
rect 44178 550287 44234 550296
rect 43628 545148 43680 545154
rect 43628 545090 43680 545096
rect 43640 430137 43668 545090
rect 44192 538286 44220 550287
rect 44180 538280 44232 538286
rect 44180 538222 44232 538228
rect 43720 440292 43772 440298
rect 43720 440234 43772 440240
rect 43626 430128 43682 430137
rect 43626 430063 43682 430072
rect 43628 419484 43680 419490
rect 43628 419426 43680 419432
rect 43640 278050 43668 419426
rect 43732 344350 43760 440234
rect 44178 429312 44234 429321
rect 44178 429247 44234 429256
rect 44192 387802 44220 429247
rect 44284 427281 44312 554367
rect 44376 428097 44404 555183
rect 44454 551168 44510 551177
rect 44454 551103 44510 551112
rect 44468 531350 44496 551103
rect 44546 548720 44602 548729
rect 44546 548655 44602 548664
rect 44560 536858 44588 548655
rect 44548 536852 44600 536858
rect 44548 536794 44600 536800
rect 44456 531344 44508 531350
rect 44456 531286 44508 531292
rect 44652 429729 44680 556815
rect 46204 491972 46256 491978
rect 46204 491914 46256 491920
rect 44824 480276 44876 480282
rect 44824 480218 44876 480224
rect 44638 429720 44694 429729
rect 44638 429655 44694 429664
rect 44362 428088 44418 428097
rect 44362 428023 44418 428032
rect 44362 427680 44418 427689
rect 44362 427615 44418 427624
rect 44270 427272 44326 427281
rect 44270 427207 44326 427216
rect 44180 387796 44232 387802
rect 44180 387738 44232 387744
rect 44178 385248 44234 385257
rect 44178 385183 44234 385192
rect 43720 344344 43772 344350
rect 43720 344286 43772 344292
rect 44192 342553 44220 385183
rect 44376 384849 44404 427615
rect 44546 426864 44602 426873
rect 44546 426799 44602 426808
rect 44454 421968 44510 421977
rect 44454 421903 44510 421912
rect 44468 403918 44496 421903
rect 44456 403912 44508 403918
rect 44456 403854 44508 403860
rect 44362 384840 44418 384849
rect 44362 384775 44418 384784
rect 44560 384033 44588 426799
rect 44638 421152 44694 421161
rect 44638 421087 44694 421096
rect 44652 408202 44680 421087
rect 44640 408196 44692 408202
rect 44640 408138 44692 408144
rect 44836 387666 44864 480218
rect 45008 389224 45060 389230
rect 45008 389166 45060 389172
rect 44824 387660 44876 387666
rect 44824 387602 44876 387608
rect 44638 386064 44694 386073
rect 44638 385999 44694 386008
rect 44546 384024 44602 384033
rect 44546 383959 44602 383968
rect 44454 379128 44510 379137
rect 44454 379063 44510 379072
rect 44468 364342 44496 379063
rect 44546 377904 44602 377913
rect 44546 377839 44602 377848
rect 44560 365022 44588 377839
rect 44548 365016 44600 365022
rect 44548 364958 44600 364964
rect 44456 364336 44508 364342
rect 44456 364278 44508 364284
rect 44652 343369 44680 385999
rect 44730 384432 44786 384441
rect 44730 384367 44786 384376
rect 44638 343360 44694 343369
rect 44638 343295 44694 343304
rect 44270 342952 44326 342961
rect 44270 342887 44326 342896
rect 44178 342544 44234 342553
rect 44178 342479 44234 342488
rect 44178 338056 44234 338065
rect 44178 337991 44234 338000
rect 44192 326806 44220 337991
rect 44180 326800 44232 326806
rect 44180 326742 44232 326748
rect 44284 300121 44312 342887
rect 44546 342136 44602 342145
rect 44546 342071 44602 342080
rect 44362 336424 44418 336433
rect 44362 336359 44418 336368
rect 44376 322930 44404 336359
rect 44454 334792 44510 334801
rect 44454 334727 44510 334736
rect 44364 322924 44416 322930
rect 44364 322866 44416 322872
rect 44468 321502 44496 334727
rect 44456 321496 44508 321502
rect 44456 321438 44508 321444
rect 44270 300112 44326 300121
rect 44270 300047 44326 300056
rect 44362 299704 44418 299713
rect 44362 299639 44418 299648
rect 44270 298888 44326 298897
rect 44270 298823 44326 298832
rect 43720 298172 43772 298178
rect 43720 298114 43772 298120
rect 43628 278044 43680 278050
rect 43628 277986 43680 277992
rect 43534 231160 43590 231169
rect 43534 231095 43590 231104
rect 43732 221474 43760 298114
rect 44178 298072 44234 298081
rect 44178 298007 44234 298016
rect 43902 290728 43958 290737
rect 43902 290663 43958 290672
rect 43812 284368 43864 284374
rect 43812 284310 43864 284316
rect 43720 221468 43772 221474
rect 43720 221410 43772 221416
rect 43824 217326 43852 284310
rect 43916 231130 43944 290663
rect 44192 255241 44220 298007
rect 44284 256057 44312 298823
rect 44376 258058 44404 299639
rect 44560 299305 44588 342071
rect 44744 341737 44772 384367
rect 44824 376100 44876 376106
rect 44824 376042 44876 376048
rect 44730 341728 44786 341737
rect 44730 341663 44786 341672
rect 44546 299296 44602 299305
rect 44546 299231 44602 299240
rect 44454 293584 44510 293593
rect 44454 293519 44510 293528
rect 44468 273086 44496 293519
rect 44546 291544 44602 291553
rect 44546 291479 44602 291488
rect 44560 278662 44588 291479
rect 44548 278656 44600 278662
rect 44548 278598 44600 278604
rect 44456 273080 44508 273086
rect 44456 273022 44508 273028
rect 44364 258052 44416 258058
rect 44364 257994 44416 258000
rect 44270 256048 44326 256057
rect 44270 255983 44326 255992
rect 44178 255232 44234 255241
rect 44178 255167 44234 255176
rect 44270 254824 44326 254833
rect 44270 254759 44326 254768
rect 44178 251560 44234 251569
rect 44178 251495 44234 251504
rect 44192 240038 44220 251495
rect 44180 240032 44232 240038
rect 44180 239974 44232 239980
rect 43904 231124 43956 231130
rect 43904 231066 43956 231072
rect 43812 217320 43864 217326
rect 43812 217262 43864 217268
rect 43350 212936 43406 212945
rect 43350 212871 43406 212880
rect 44284 212129 44312 254759
rect 44730 254008 44786 254017
rect 44730 253943 44786 253952
rect 44362 251152 44418 251161
rect 44362 251087 44418 251096
rect 44376 226710 44404 251087
rect 44546 249520 44602 249529
rect 44546 249455 44602 249464
rect 44560 234598 44588 249455
rect 44638 248296 44694 248305
rect 44638 248231 44694 248240
rect 44652 235414 44680 248231
rect 44640 235408 44692 235414
rect 44640 235350 44692 235356
rect 44548 234592 44600 234598
rect 44548 234534 44600 234540
rect 44364 226704 44416 226710
rect 44364 226646 44416 226652
rect 44270 212120 44326 212129
rect 44270 212055 44326 212064
rect 41326 211848 41382 211857
rect 41326 211783 41382 211792
rect 44744 211313 44772 253943
rect 44836 218754 44864 376042
rect 44916 347064 44968 347070
rect 44916 347006 44968 347012
rect 44928 257922 44956 347006
rect 45020 300529 45048 389166
rect 46216 387530 46244 491914
rect 46296 427848 46348 427854
rect 46296 427790 46348 427796
rect 46204 387524 46256 387530
rect 46204 387466 46256 387472
rect 46308 351218 46336 427790
rect 47596 410718 47624 557534
rect 48976 540258 49004 609962
rect 48964 540252 49016 540258
rect 48964 540194 49016 540200
rect 48964 506524 49016 506530
rect 48964 506466 49016 506472
rect 47584 410712 47636 410718
rect 47584 410654 47636 410660
rect 47584 401668 47636 401674
rect 47584 401610 47636 401616
rect 46296 351212 46348 351218
rect 46296 351154 46348 351160
rect 46296 336796 46348 336802
rect 46296 336738 46348 336744
rect 46204 310548 46256 310554
rect 46204 310490 46256 310496
rect 45006 300520 45062 300529
rect 45006 300455 45062 300464
rect 45006 291136 45062 291145
rect 45006 291071 45062 291080
rect 45020 264246 45048 291071
rect 45008 264240 45060 264246
rect 45008 264182 45060 264188
rect 44916 257916 44968 257922
rect 44916 257858 44968 257864
rect 44914 248704 44970 248713
rect 44914 248639 44970 248648
rect 44928 234054 44956 248639
rect 44916 234048 44968 234054
rect 44916 233990 44968 233996
rect 44824 218748 44876 218754
rect 44824 218690 44876 218696
rect 46216 214606 46244 310490
rect 46308 265674 46336 336738
rect 47596 280226 47624 401610
rect 48976 364274 49004 506466
rect 49056 375420 49108 375426
rect 49056 375362 49108 375368
rect 48964 364268 49016 364274
rect 48964 364210 49016 364216
rect 47676 322992 47728 322998
rect 47676 322934 47728 322940
rect 47584 280220 47636 280226
rect 47584 280162 47636 280168
rect 46296 265668 46348 265674
rect 46296 265610 46348 265616
rect 47688 257786 47716 322934
rect 49068 301034 49096 375362
rect 49056 301028 49108 301034
rect 49056 300970 49108 300976
rect 47676 257780 47728 257786
rect 47676 257722 47728 257728
rect 50356 231334 50384 719646
rect 50436 714876 50488 714882
rect 50436 714818 50488 714824
rect 50448 627230 50476 714818
rect 51736 687954 51764 727262
rect 51724 687948 51776 687954
rect 51724 687890 51776 687896
rect 54496 687818 54524 741066
rect 54484 687812 54536 687818
rect 54484 687754 54536 687760
rect 51724 676864 51776 676870
rect 51724 676806 51776 676812
rect 50436 627224 50488 627230
rect 50436 627166 50488 627172
rect 50436 597576 50488 597582
rect 50436 597518 50488 597524
rect 50448 558346 50476 597518
rect 50436 558340 50488 558346
rect 50436 558282 50488 558288
rect 50436 454096 50488 454102
rect 50436 454038 50488 454044
rect 50448 321570 50476 454038
rect 50436 321564 50488 321570
rect 50436 321506 50488 321512
rect 50344 231328 50396 231334
rect 50344 231270 50396 231276
rect 51736 231266 51764 676806
rect 54482 633448 54538 633457
rect 54482 633383 54538 633392
rect 51816 623824 51868 623830
rect 51816 623766 51868 623772
rect 51828 601390 51856 623766
rect 51816 601384 51868 601390
rect 51816 601326 51868 601332
rect 53104 589960 53156 589966
rect 53104 589902 53156 589908
rect 51816 583772 51868 583778
rect 51816 583714 51868 583720
rect 51828 558210 51856 583714
rect 51816 558204 51868 558210
rect 51816 558146 51868 558152
rect 51816 466472 51868 466478
rect 51816 466414 51868 466420
rect 51828 387394 51856 466414
rect 51816 387388 51868 387394
rect 51816 387330 51868 387336
rect 51814 289912 51870 289921
rect 51814 289847 51870 289856
rect 51828 278118 51856 289847
rect 51816 278112 51868 278118
rect 51816 278054 51868 278060
rect 51724 231260 51776 231266
rect 51724 231202 51776 231208
rect 53116 231198 53144 589902
rect 53196 547188 53248 547194
rect 53196 547130 53248 547136
rect 53208 278186 53236 547130
rect 53196 278180 53248 278186
rect 53196 278122 53248 278128
rect 54496 231402 54524 633383
rect 55876 231538 55904 761738
rect 55968 756906 55996 870810
rect 62118 858664 62174 858673
rect 62118 858599 62174 858608
rect 62132 858430 62160 858599
rect 62120 858424 62172 858430
rect 62120 858366 62172 858372
rect 62118 845608 62174 845617
rect 62118 845543 62174 845552
rect 62132 844626 62160 845543
rect 62120 844620 62172 844626
rect 62120 844562 62172 844568
rect 62118 832552 62174 832561
rect 62118 832487 62174 832496
rect 62132 832182 62160 832487
rect 62120 832176 62172 832182
rect 62120 832118 62172 832124
rect 62118 819496 62174 819505
rect 62118 819431 62174 819440
rect 62132 818378 62160 819431
rect 62120 818372 62172 818378
rect 62120 818314 62172 818320
rect 62118 806576 62174 806585
rect 62118 806511 62174 806520
rect 62132 806002 62160 806511
rect 62120 805996 62172 806002
rect 62120 805938 62172 805944
rect 62118 793656 62174 793665
rect 62118 793591 62174 793600
rect 62132 793558 62160 793591
rect 62120 793552 62172 793558
rect 62120 793494 62172 793500
rect 62118 780464 62174 780473
rect 62118 780399 62174 780408
rect 62132 779754 62160 780399
rect 62120 779748 62172 779754
rect 62120 779690 62172 779696
rect 62118 767408 62174 767417
rect 62118 767343 62120 767352
rect 62172 767343 62174 767352
rect 62120 767314 62172 767320
rect 55956 756900 56008 756906
rect 55956 756842 56008 756848
rect 62118 754352 62174 754361
rect 62118 754287 62174 754296
rect 62132 753574 62160 754287
rect 62120 753568 62172 753574
rect 62120 753510 62172 753516
rect 62118 741296 62174 741305
rect 62118 741231 62174 741240
rect 62132 741130 62160 741231
rect 62120 741124 62172 741130
rect 62120 741066 62172 741072
rect 62118 728240 62174 728249
rect 62118 728175 62174 728184
rect 62132 727326 62160 728175
rect 62120 727320 62172 727326
rect 62120 727262 62172 727268
rect 62118 715320 62174 715329
rect 62118 715255 62174 715264
rect 62132 714882 62160 715255
rect 62120 714876 62172 714882
rect 62120 714818 62172 714824
rect 62762 702264 62818 702273
rect 62762 702199 62818 702208
rect 62118 689208 62174 689217
rect 62118 689143 62174 689152
rect 62132 688702 62160 689143
rect 62120 688696 62172 688702
rect 62120 688638 62172 688644
rect 62118 676152 62174 676161
rect 62118 676087 62174 676096
rect 62132 674898 62160 676087
rect 55956 674892 56008 674898
rect 55956 674834 56008 674840
rect 62120 674892 62172 674898
rect 62120 674834 62172 674840
rect 55968 644570 55996 674834
rect 62118 663096 62174 663105
rect 62118 663031 62174 663040
rect 62132 662454 62160 663031
rect 62120 662448 62172 662454
rect 62120 662390 62172 662396
rect 62118 650040 62174 650049
rect 62118 649975 62174 649984
rect 62132 647902 62160 649975
rect 62120 647896 62172 647902
rect 62120 647838 62172 647844
rect 55956 644564 56008 644570
rect 55956 644506 56008 644512
rect 62776 643521 62804 702199
rect 62762 643512 62818 643521
rect 62762 643447 62818 643456
rect 62118 637120 62174 637129
rect 62118 637055 62174 637064
rect 62132 636274 62160 637055
rect 55956 636268 56008 636274
rect 55956 636210 56008 636216
rect 62120 636268 62172 636274
rect 62120 636210 62172 636216
rect 55968 601730 55996 636210
rect 62118 624064 62174 624073
rect 62118 623999 62174 624008
rect 62132 623830 62160 623999
rect 62120 623824 62172 623830
rect 62120 623766 62172 623772
rect 62118 611008 62174 611017
rect 62118 610943 62174 610952
rect 62132 610026 62160 610943
rect 62120 610020 62172 610026
rect 62120 609962 62172 609968
rect 55956 601724 56008 601730
rect 55956 601666 56008 601672
rect 62118 597952 62174 597961
rect 62118 597887 62174 597896
rect 62132 597582 62160 597887
rect 62120 597576 62172 597582
rect 62120 597518 62172 597524
rect 62118 584896 62174 584905
rect 62118 584831 62174 584840
rect 62132 583778 62160 584831
rect 62120 583772 62172 583778
rect 62120 583714 62172 583720
rect 62118 571840 62174 571849
rect 62118 571775 62174 571784
rect 62132 571402 62160 571775
rect 62120 571396 62172 571402
rect 62120 571338 62172 571344
rect 62118 558784 62174 558793
rect 62118 558719 62174 558728
rect 62132 557598 62160 558719
rect 62120 557592 62172 557598
rect 62120 557534 62172 557540
rect 62118 545864 62174 545873
rect 62118 545799 62174 545808
rect 62132 545154 62160 545799
rect 62120 545148 62172 545154
rect 62120 545090 62172 545096
rect 62118 532808 62174 532817
rect 55956 532772 56008 532778
rect 62118 532743 62120 532752
rect 55956 532714 56008 532720
rect 62172 532743 62174 532752
rect 62120 532714 62172 532720
rect 55968 430642 55996 532714
rect 62118 519752 62174 519761
rect 62118 519687 62174 519696
rect 62132 518974 62160 519687
rect 62120 518968 62172 518974
rect 62120 518910 62172 518916
rect 62118 506696 62174 506705
rect 62118 506631 62174 506640
rect 62132 506530 62160 506631
rect 62120 506524 62172 506530
rect 62120 506466 62172 506472
rect 62118 493640 62174 493649
rect 62118 493575 62174 493584
rect 62132 491978 62160 493575
rect 62120 491972 62172 491978
rect 62120 491914 62172 491920
rect 62118 480584 62174 480593
rect 62118 480519 62174 480528
rect 62132 480282 62160 480519
rect 62120 480276 62172 480282
rect 62120 480218 62172 480224
rect 62118 467528 62174 467537
rect 62118 467463 62174 467472
rect 62132 466478 62160 467463
rect 62120 466472 62172 466478
rect 62120 466414 62172 466420
rect 62118 454608 62174 454617
rect 62118 454543 62174 454552
rect 62132 454102 62160 454543
rect 62120 454096 62172 454102
rect 62120 454038 62172 454044
rect 62118 441552 62174 441561
rect 62118 441487 62174 441496
rect 62132 440298 62160 441487
rect 62120 440292 62172 440298
rect 62120 440234 62172 440240
rect 55956 430636 56008 430642
rect 55956 430578 56008 430584
rect 62118 428496 62174 428505
rect 62118 428431 62174 428440
rect 62132 427854 62160 428431
rect 62120 427848 62172 427854
rect 62120 427790 62172 427796
rect 55956 415472 56008 415478
rect 62120 415472 62172 415478
rect 55956 415414 56008 415420
rect 62118 415440 62120 415449
rect 62172 415440 62174 415449
rect 55968 344214 55996 415414
rect 62118 415375 62174 415384
rect 62118 402384 62174 402393
rect 62118 402319 62174 402328
rect 62132 401674 62160 402319
rect 62120 401668 62172 401674
rect 62120 401610 62172 401616
rect 62118 389328 62174 389337
rect 62118 389263 62174 389272
rect 62132 389230 62160 389263
rect 62120 389224 62172 389230
rect 62120 389166 62172 389172
rect 62118 376272 62174 376281
rect 62118 376207 62174 376216
rect 62132 375426 62160 376207
rect 62120 375420 62172 375426
rect 62120 375362 62172 375368
rect 62118 363352 62174 363361
rect 62118 363287 62174 363296
rect 62132 362982 62160 363287
rect 56048 362976 56100 362982
rect 56048 362918 56100 362924
rect 62120 362976 62172 362982
rect 62120 362918 62172 362924
rect 55956 344208 56008 344214
rect 55956 344150 56008 344156
rect 56060 300966 56088 362918
rect 62118 350296 62174 350305
rect 62118 350231 62174 350240
rect 62132 347070 62160 350231
rect 62120 347064 62172 347070
rect 62120 347006 62172 347012
rect 62118 337240 62174 337249
rect 62118 337175 62174 337184
rect 62132 336802 62160 337175
rect 62120 336796 62172 336802
rect 62120 336738 62172 336744
rect 64144 333260 64196 333266
rect 64144 333202 64196 333208
rect 62118 324184 62174 324193
rect 62118 324119 62174 324128
rect 62132 322998 62160 324119
rect 62120 322992 62172 322998
rect 62120 322934 62172 322940
rect 62118 311128 62174 311137
rect 62118 311063 62174 311072
rect 62132 310554 62160 311063
rect 62120 310548 62172 310554
rect 62120 310490 62172 310496
rect 56048 300960 56100 300966
rect 56048 300902 56100 300908
rect 62118 298208 62174 298217
rect 62118 298143 62120 298152
rect 62172 298143 62174 298152
rect 62120 298114 62172 298120
rect 62118 285152 62174 285161
rect 62118 285087 62174 285096
rect 62132 284374 62160 285087
rect 62120 284368 62172 284374
rect 62120 284310 62172 284316
rect 55864 231532 55916 231538
rect 55864 231474 55916 231480
rect 64156 231470 64184 333202
rect 645872 278310 646346 278338
rect 332508 277976 332560 277982
rect 332508 277918 332560 277924
rect 436652 277976 436704 277982
rect 436704 277924 437046 277930
rect 436652 277918 437046 277924
rect 65918 277766 66208 277794
rect 66180 268394 66208 277766
rect 67008 275398 67036 277780
rect 66996 275392 67048 275398
rect 66996 275334 67048 275340
rect 68204 272542 68232 277780
rect 68192 272536 68244 272542
rect 68192 272478 68244 272484
rect 69400 268462 69428 277780
rect 70596 270502 70624 277780
rect 71792 275330 71820 277780
rect 71780 275324 71832 275330
rect 71780 275266 71832 275272
rect 72988 273970 73016 277780
rect 74092 274718 74120 277780
rect 75302 277766 75868 277794
rect 76498 277766 77248 277794
rect 74080 274712 74132 274718
rect 74080 274654 74132 274660
rect 72976 273964 73028 273970
rect 72976 273906 73028 273912
rect 70584 270496 70636 270502
rect 70584 270438 70636 270444
rect 71780 270496 71832 270502
rect 71780 270438 71832 270444
rect 69388 268456 69440 268462
rect 69388 268398 69440 268404
rect 66168 268388 66220 268394
rect 66168 268330 66220 268336
rect 71792 267034 71820 270438
rect 75840 268530 75868 277766
rect 76012 274712 76064 274718
rect 76012 274654 76064 274660
rect 76024 272610 76052 274654
rect 76012 272604 76064 272610
rect 76012 272546 76064 272552
rect 77220 269890 77248 277766
rect 77208 269884 77260 269890
rect 77208 269826 77260 269832
rect 77680 268598 77708 277780
rect 78876 271522 78904 277780
rect 78864 271516 78916 271522
rect 78864 271458 78916 271464
rect 80072 268666 80100 277780
rect 81268 275466 81296 277780
rect 82386 277766 82768 277794
rect 81256 275460 81308 275466
rect 81256 275402 81308 275408
rect 82740 268734 82768 277766
rect 83568 275534 83596 277780
rect 83556 275528 83608 275534
rect 83556 275470 83608 275476
rect 84764 274038 84792 277780
rect 84752 274032 84804 274038
rect 84752 273974 84804 273980
rect 85960 269958 85988 277780
rect 85948 269952 86000 269958
rect 85948 269894 86000 269900
rect 87156 268802 87184 277780
rect 88352 274718 88380 277780
rect 88340 274712 88392 274718
rect 88340 274654 88392 274660
rect 89548 272678 89576 277780
rect 90652 275602 90680 277780
rect 91862 277766 92428 277794
rect 90640 275596 90692 275602
rect 90640 275538 90692 275544
rect 89536 272672 89588 272678
rect 89536 272614 89588 272620
rect 92400 268870 92428 277766
rect 93044 271726 93072 277780
rect 93124 274712 93176 274718
rect 93124 274654 93176 274660
rect 93032 271720 93084 271726
rect 93032 271662 93084 271668
rect 92388 268864 92440 268870
rect 92388 268806 92440 268812
rect 87144 268796 87196 268802
rect 87144 268738 87196 268744
rect 82728 268728 82780 268734
rect 82728 268670 82780 268676
rect 80060 268660 80112 268666
rect 80060 268602 80112 268608
rect 77668 268592 77720 268598
rect 77668 268534 77720 268540
rect 75828 268524 75880 268530
rect 75828 268466 75880 268472
rect 93136 267102 93164 274654
rect 94240 274106 94268 277780
rect 94228 274100 94280 274106
rect 94228 274042 94280 274048
rect 95436 268938 95464 277780
rect 96632 271386 96660 277780
rect 97736 274174 97764 277780
rect 98946 277766 99328 277794
rect 97724 274168 97776 274174
rect 97724 274110 97776 274116
rect 96620 271380 96672 271386
rect 96620 271322 96672 271328
rect 99300 269006 99328 277766
rect 100128 275670 100156 277780
rect 100116 275664 100168 275670
rect 100116 275606 100168 275612
rect 101324 272746 101352 277780
rect 101312 272740 101364 272746
rect 101312 272682 101364 272688
rect 102520 269074 102548 277780
rect 103716 270162 103744 277780
rect 104912 271182 104940 277780
rect 106030 277766 106228 277794
rect 104900 271176 104952 271182
rect 104900 271118 104952 271124
rect 103704 270156 103756 270162
rect 103704 270098 103756 270104
rect 102508 269068 102560 269074
rect 102508 269010 102560 269016
rect 99288 269000 99340 269006
rect 99288 268942 99340 268948
rect 95424 268932 95476 268938
rect 95424 268874 95476 268880
rect 106200 268326 106228 277766
rect 107212 275738 107240 277780
rect 107200 275732 107252 275738
rect 107200 275674 107252 275680
rect 108408 272814 108436 277780
rect 109618 277766 110368 277794
rect 108396 272808 108448 272814
rect 108396 272750 108448 272756
rect 110340 269822 110368 277766
rect 110800 270026 110828 277780
rect 111996 274242 112024 277780
rect 111984 274236 112036 274242
rect 111984 274178 112036 274184
rect 113192 272882 113220 277780
rect 113180 272876 113232 272882
rect 113180 272818 113232 272824
rect 114296 271250 114324 277780
rect 115506 277766 115888 277794
rect 114284 271244 114336 271250
rect 114284 271186 114336 271192
rect 110788 270020 110840 270026
rect 110788 269962 110840 269968
rect 110512 269952 110564 269958
rect 110512 269894 110564 269900
rect 110328 269816 110380 269822
rect 110328 269758 110380 269764
rect 106188 268320 106240 268326
rect 106188 268262 106240 268268
rect 110524 267238 110552 269894
rect 115860 269890 115888 277766
rect 116688 274310 116716 277780
rect 117898 277766 118648 277794
rect 116676 274304 116728 274310
rect 116676 274246 116728 274252
rect 118620 269958 118648 277766
rect 119080 270094 119108 277780
rect 120276 272950 120304 277780
rect 121380 274378 121408 277780
rect 122590 277766 122788 277794
rect 121368 274372 121420 274378
rect 121368 274314 121420 274320
rect 120264 272944 120316 272950
rect 120264 272886 120316 272892
rect 122760 270094 122788 277766
rect 123772 274446 123800 277780
rect 123760 274440 123812 274446
rect 123760 274382 123812 274388
rect 124968 271318 124996 277780
rect 126178 277766 126928 277794
rect 124956 271312 125008 271318
rect 124956 271254 125008 271260
rect 126900 270162 126928 277766
rect 127360 273018 127388 277780
rect 128556 275262 128584 277780
rect 128544 275256 128596 275262
rect 128544 275198 128596 275204
rect 127348 273012 127400 273018
rect 127348 272954 127400 272960
rect 129660 270230 129688 277780
rect 130870 277766 131068 277794
rect 129648 270224 129700 270230
rect 129648 270166 129700 270172
rect 125968 270156 126020 270162
rect 125968 270098 126020 270104
rect 126888 270156 126940 270162
rect 126888 270098 126940 270104
rect 119068 270088 119120 270094
rect 119068 270030 119120 270036
rect 122748 270088 122800 270094
rect 122748 270030 122800 270036
rect 119620 270020 119672 270026
rect 119620 269962 119672 269968
rect 118608 269952 118660 269958
rect 118608 269894 118660 269900
rect 113180 269884 113232 269890
rect 113180 269826 113232 269832
rect 115848 269884 115900 269890
rect 115848 269826 115900 269832
rect 113192 267306 113220 269826
rect 113180 267300 113232 267306
rect 113180 267242 113232 267248
rect 110512 267232 110564 267238
rect 110512 267174 110564 267180
rect 119632 267170 119660 269962
rect 125980 267374 126008 270098
rect 131040 268258 131068 277766
rect 131120 275256 131172 275262
rect 131120 275198 131172 275204
rect 131132 273086 131160 275198
rect 132052 273834 132080 277780
rect 133262 277766 133828 277794
rect 134458 277766 135208 277794
rect 132040 273828 132092 273834
rect 132040 273770 132092 273776
rect 131120 273080 131172 273086
rect 131120 273022 131172 273028
rect 133800 270298 133828 277766
rect 133788 270292 133840 270298
rect 133788 270234 133840 270240
rect 131028 268252 131080 268258
rect 131028 268194 131080 268200
rect 135180 268190 135208 277766
rect 135640 269550 135668 277780
rect 136836 274650 136864 277780
rect 136824 274644 136876 274650
rect 136824 274586 136876 274592
rect 137940 274514 137968 277780
rect 139136 275194 139164 277780
rect 140346 277766 140728 277794
rect 139124 275188 139176 275194
rect 139124 275130 139176 275136
rect 137928 274508 137980 274514
rect 137928 274450 137980 274456
rect 140700 270366 140728 277766
rect 141528 273154 141556 277780
rect 141516 273148 141568 273154
rect 141516 273090 141568 273096
rect 142724 271794 142752 277780
rect 142712 271788 142764 271794
rect 142712 271730 142764 271736
rect 143920 271454 143948 277780
rect 145024 274582 145052 277780
rect 146220 276010 146248 277780
rect 146208 276004 146260 276010
rect 146208 275946 146260 275952
rect 145012 274576 145064 274582
rect 145012 274518 145064 274524
rect 147416 271454 147444 277780
rect 148612 273222 148640 277780
rect 149808 275806 149836 277780
rect 149796 275800 149848 275806
rect 149796 275742 149848 275748
rect 148600 273216 148652 273222
rect 148600 273158 148652 273164
rect 151004 271590 151032 277780
rect 152200 271658 152228 277780
rect 153304 272270 153332 277780
rect 153292 272264 153344 272270
rect 153292 272206 153344 272212
rect 153844 271720 153896 271726
rect 153844 271662 153896 271668
rect 152188 271652 152240 271658
rect 152188 271594 152240 271600
rect 150992 271584 151044 271590
rect 150992 271526 151044 271532
rect 152464 271516 152516 271522
rect 152464 271458 152516 271464
rect 143908 271448 143960 271454
rect 143908 271390 143960 271396
rect 147404 271448 147456 271454
rect 147404 271390 147456 271396
rect 144184 271380 144236 271386
rect 144184 271322 144236 271328
rect 140688 270360 140740 270366
rect 140688 270302 140740 270308
rect 135628 269544 135680 269550
rect 135628 269486 135680 269492
rect 135168 268184 135220 268190
rect 135168 268126 135220 268132
rect 144196 267578 144224 271322
rect 144184 267572 144236 267578
rect 144184 267514 144236 267520
rect 125968 267368 126020 267374
rect 125968 267310 126020 267316
rect 119620 267164 119672 267170
rect 119620 267106 119672 267112
rect 93124 267096 93176 267102
rect 93124 267038 93176 267044
rect 71780 267028 71832 267034
rect 71780 266970 71832 266976
rect 152476 266830 152504 271458
rect 153856 266898 153884 271662
rect 154500 271522 154528 277780
rect 155696 273902 155724 277780
rect 156892 275262 156920 277780
rect 156880 275256 156932 275262
rect 156880 275198 156932 275204
rect 155684 273896 155736 273902
rect 155684 273838 155736 273844
rect 158088 271726 158116 277780
rect 159284 272474 159312 277780
rect 160480 274718 160508 277780
rect 160468 274712 160520 274718
rect 160468 274654 160520 274660
rect 161388 274712 161440 274718
rect 161388 274654 161440 274660
rect 159272 272468 159324 272474
rect 159272 272410 159324 272416
rect 158076 271720 158128 271726
rect 158076 271662 158128 271668
rect 154488 271516 154540 271522
rect 154488 271458 154540 271464
rect 161400 267442 161428 274654
rect 161584 271862 161612 277780
rect 161572 271856 161624 271862
rect 161572 271798 161624 271804
rect 162780 271794 162808 277780
rect 163976 275942 164004 277780
rect 163964 275936 164016 275942
rect 163964 275878 164016 275884
rect 162124 271788 162176 271794
rect 162124 271730 162176 271736
rect 162768 271788 162820 271794
rect 162768 271730 162820 271736
rect 162136 267646 162164 271730
rect 165172 271114 165200 277780
rect 166382 277766 166948 277794
rect 167578 277766 168328 277794
rect 165160 271108 165212 271114
rect 165160 271050 165212 271056
rect 166920 270434 166948 277766
rect 166908 270428 166960 270434
rect 166908 270370 166960 270376
rect 162124 267640 162176 267646
rect 162124 267582 162176 267588
rect 168300 267510 168328 277766
rect 168668 271046 168696 277780
rect 168656 271040 168708 271046
rect 168656 270982 168708 270988
rect 169864 270502 169892 277780
rect 171060 275874 171088 277780
rect 171048 275868 171100 275874
rect 171048 275810 171100 275816
rect 172256 270978 172284 277780
rect 173466 277766 173848 277794
rect 174662 277766 175228 277794
rect 172244 270972 172296 270978
rect 172244 270914 172296 270920
rect 169852 270496 169904 270502
rect 169852 270438 169904 270444
rect 173820 269754 173848 277766
rect 173808 269748 173860 269754
rect 173808 269690 173860 269696
rect 175200 267714 175228 277766
rect 175844 270910 175872 277780
rect 175832 270904 175884 270910
rect 175832 270846 175884 270852
rect 176948 269686 176976 277780
rect 178144 275126 178172 277780
rect 178132 275120 178184 275126
rect 178132 275062 178184 275068
rect 179340 272406 179368 277780
rect 180550 277766 180748 277794
rect 181746 277766 182128 277794
rect 179328 272400 179380 272406
rect 179328 272342 179380 272348
rect 176936 269680 176988 269686
rect 176936 269622 176988 269628
rect 180720 269618 180748 277766
rect 180708 269612 180760 269618
rect 180708 269554 180760 269560
rect 175188 267708 175240 267714
rect 175188 267650 175240 267656
rect 168288 267504 168340 267510
rect 168288 267446 168340 267452
rect 161388 267436 161440 267442
rect 161388 267378 161440 267384
rect 182100 266966 182128 277766
rect 182928 273766 182956 277780
rect 184138 277766 184888 277794
rect 182916 273760 182968 273766
rect 182916 273702 182968 273708
rect 184860 269550 184888 277766
rect 185032 275188 185084 275194
rect 185032 275130 185084 275136
rect 184756 269544 184808 269550
rect 184756 269486 184808 269492
rect 184848 269544 184900 269550
rect 184848 269486 184900 269492
rect 182088 266960 182140 266966
rect 182088 266902 182140 266908
rect 153844 266892 153896 266898
rect 153844 266834 153896 266840
rect 152464 266824 152516 266830
rect 152464 266766 152516 266772
rect 184768 266762 184796 269486
rect 185044 268054 185072 275130
rect 185228 275058 185256 277780
rect 185216 275052 185268 275058
rect 185216 274994 185268 275000
rect 186424 268122 186452 277780
rect 187620 277394 187648 277780
rect 187528 277366 187648 277394
rect 187528 269482 187556 277366
rect 187700 275392 187752 275398
rect 187700 275334 187752 275340
rect 187712 273562 187740 275334
rect 188816 275194 188844 277780
rect 188804 275188 188856 275194
rect 188804 275130 188856 275136
rect 187700 273556 187752 273562
rect 187700 273498 187752 273504
rect 190012 270842 190040 277780
rect 191208 272338 191236 277780
rect 192326 277766 192616 277794
rect 192392 273556 192444 273562
rect 192392 273498 192444 273504
rect 191196 272332 191248 272338
rect 191196 272274 191248 272280
rect 190000 270836 190052 270842
rect 190000 270778 190052 270784
rect 187516 269476 187568 269482
rect 187516 269418 187568 269424
rect 192116 268388 192168 268394
rect 192116 268330 192168 268336
rect 186412 268116 186464 268122
rect 186412 268058 186464 268064
rect 185032 268048 185084 268054
rect 185032 267990 185084 267996
rect 184756 266756 184808 266762
rect 184756 266698 184808 266704
rect 192128 264330 192156 268330
rect 192404 264738 192432 273498
rect 192588 272270 192616 277766
rect 193508 272542 193536 277780
rect 194600 273964 194652 273970
rect 194600 273906 194652 273912
rect 193220 272536 193272 272542
rect 193220 272478 193272 272484
rect 193496 272536 193548 272542
rect 193496 272478 193548 272484
rect 192484 272264 192536 272270
rect 192484 272206 192536 272212
rect 192576 272264 192628 272270
rect 192576 272206 192628 272212
rect 192496 266694 192524 272206
rect 192484 266688 192536 266694
rect 192484 266630 192536 266636
rect 192404 264710 192524 264738
rect 192496 264330 192524 264710
rect 192128 264302 192418 264330
rect 192496 264302 192786 264330
rect 193232 264316 193260 272478
rect 193680 268456 193732 268462
rect 193680 268398 193732 268404
rect 193692 264316 193720 268398
rect 194140 267028 194192 267034
rect 194140 266970 194192 266976
rect 194152 264316 194180 266970
rect 194612 265538 194640 273906
rect 194704 273698 194732 277780
rect 194876 275324 194928 275330
rect 194876 275266 194928 275272
rect 194692 273692 194744 273698
rect 194692 273634 194744 273640
rect 194784 272604 194836 272610
rect 194784 272546 194836 272552
rect 194796 265606 194824 272546
rect 194784 265600 194836 265606
rect 194784 265542 194836 265548
rect 194600 265532 194652 265538
rect 194600 265474 194652 265480
rect 194888 264194 194916 275266
rect 195900 273970 195928 277780
rect 195980 276004 196032 276010
rect 195980 275946 196032 275952
rect 195888 273964 195940 273970
rect 195888 273906 195940 273912
rect 195428 268524 195480 268530
rect 195428 268466 195480 268472
rect 194968 265532 195020 265538
rect 194968 265474 195020 265480
rect 194980 264330 195008 265474
rect 194980 264302 195086 264330
rect 195440 264316 195468 268466
rect 195992 267986 196020 275946
rect 197096 273834 197124 277780
rect 197820 275460 197872 275466
rect 197820 275402 197872 275408
rect 196624 273828 196676 273834
rect 196624 273770 196676 273776
rect 197084 273828 197136 273834
rect 197084 273770 197136 273776
rect 195980 267980 196032 267986
rect 195980 267922 196032 267928
rect 196636 267306 196664 273770
rect 197268 268660 197320 268666
rect 197268 268602 197320 268608
rect 196808 268592 196860 268598
rect 196808 268534 196860 268540
rect 196348 267300 196400 267306
rect 196348 267242 196400 267248
rect 196624 267300 196676 267306
rect 196624 267242 196676 267248
rect 195612 265600 195664 265606
rect 195612 265542 195664 265548
rect 195624 264330 195652 265542
rect 195624 264302 195914 264330
rect 196360 264316 196388 267242
rect 196820 264316 196848 268534
rect 197280 264316 197308 268602
rect 197728 266824 197780 266830
rect 197728 266766 197780 266772
rect 197740 264316 197768 266766
rect 197832 264330 197860 275402
rect 198292 272610 198320 277780
rect 199108 275528 199160 275534
rect 199108 275470 199160 275476
rect 198832 274032 198884 274038
rect 198832 273974 198884 273980
rect 198280 272604 198332 272610
rect 198280 272546 198332 272552
rect 198556 268728 198608 268734
rect 198556 268670 198608 268676
rect 197832 264302 198122 264330
rect 198568 264316 198596 268670
rect 198844 264330 198872 273974
rect 199120 264330 199148 275470
rect 199488 272202 199516 277780
rect 200592 272678 200620 277780
rect 201684 275596 201736 275602
rect 201684 275538 201736 275544
rect 201592 274100 201644 274106
rect 201592 274042 201644 274048
rect 200488 272672 200540 272678
rect 200488 272614 200540 272620
rect 200580 272672 200632 272678
rect 200580 272614 200632 272620
rect 199476 272196 199528 272202
rect 199476 272138 199528 272144
rect 200396 268796 200448 268802
rect 200396 268738 200448 268744
rect 199936 267232 199988 267238
rect 199936 267174 199988 267180
rect 198844 264302 199042 264330
rect 199120 264302 199502 264330
rect 199948 264316 199976 267174
rect 200408 264316 200436 268738
rect 200500 264330 200528 272614
rect 201224 267096 201276 267102
rect 201224 267038 201276 267044
rect 200500 264302 200790 264330
rect 201236 264316 201264 267038
rect 201604 265606 201632 274042
rect 201592 265600 201644 265606
rect 201592 265542 201644 265548
rect 201696 264316 201724 275538
rect 201788 274038 201816 277780
rect 202984 274106 203012 277780
rect 203616 274168 203668 274174
rect 203616 274110 203668 274116
rect 202972 274100 203024 274106
rect 202972 274042 203024 274048
rect 201776 274032 201828 274038
rect 201776 273974 201828 273980
rect 203524 268932 203576 268938
rect 203524 268874 203576 268880
rect 202144 268864 202196 268870
rect 202144 268806 202196 268812
rect 202156 264316 202184 268806
rect 203064 266892 203116 266898
rect 203064 266834 203116 266840
rect 202236 265600 202288 265606
rect 202236 265542 202288 265548
rect 202248 264330 202276 265542
rect 202248 264302 202630 264330
rect 203076 264316 203104 266834
rect 203536 264316 203564 268874
rect 203628 264330 203656 274110
rect 204180 273630 204208 277780
rect 204904 275256 204956 275262
rect 204904 275198 204956 275204
rect 204168 273624 204220 273630
rect 204168 273566 204220 273572
rect 204812 272740 204864 272746
rect 204812 272682 204864 272688
rect 204444 269000 204496 269006
rect 204444 268942 204496 268948
rect 204352 267572 204404 267578
rect 204352 267514 204404 267520
rect 203628 264302 203918 264330
rect 204364 264316 204392 267514
rect 204456 264330 204484 268942
rect 204824 267734 204852 272682
rect 204916 268802 204944 275198
rect 205376 274174 205404 277780
rect 205824 275664 205876 275670
rect 205824 275606 205876 275612
rect 205364 274168 205416 274174
rect 205364 274110 205416 274116
rect 204904 268796 204956 268802
rect 204904 268738 204956 268744
rect 204824 267706 204944 267734
rect 204916 264330 204944 267706
rect 205836 264330 205864 275606
rect 206572 275330 206600 277780
rect 207768 275670 207796 277780
rect 208308 275732 208360 275738
rect 208308 275674 208360 275680
rect 207756 275664 207808 275670
rect 207756 275606 207808 275612
rect 206560 275324 206612 275330
rect 206560 275266 206612 275272
rect 207572 272808 207624 272814
rect 207572 272750 207624 272756
rect 206284 271176 206336 271182
rect 206284 271118 206336 271124
rect 206192 269068 206244 269074
rect 206192 269010 206244 269016
rect 204456 264302 204838 264330
rect 204916 264302 205298 264330
rect 205758 264302 205864 264330
rect 206204 264316 206232 269010
rect 206296 264330 206324 271118
rect 207480 268320 207532 268326
rect 207480 268262 207532 268268
rect 207020 267368 207072 267374
rect 207020 267310 207072 267316
rect 206296 264302 206586 264330
rect 207032 264316 207060 267310
rect 207492 264316 207520 268262
rect 207584 264330 207612 272750
rect 208320 267734 208348 275674
rect 208872 275398 208900 277780
rect 210068 275534 210096 277780
rect 210056 275528 210108 275534
rect 210056 275470 210108 275476
rect 208860 275392 208912 275398
rect 208860 275334 208912 275340
rect 210424 275188 210476 275194
rect 210424 275130 210476 275136
rect 208952 274236 209004 274242
rect 208952 274178 209004 274184
rect 208860 269816 208912 269822
rect 208860 269758 208912 269764
rect 208320 267706 208440 267734
rect 207584 264302 207966 264330
rect 208412 264316 208440 267706
rect 208872 264316 208900 269758
rect 208964 264330 208992 274178
rect 209964 272876 210016 272882
rect 209964 272818 210016 272824
rect 209872 271244 209924 271250
rect 209872 271186 209924 271192
rect 209688 267164 209740 267170
rect 209688 267106 209740 267112
rect 208964 264302 209254 264330
rect 209700 264316 209728 267106
rect 209884 265606 209912 271186
rect 209872 265600 209924 265606
rect 209872 265542 209924 265548
rect 209976 264330 210004 272818
rect 210436 267034 210464 275130
rect 210608 269884 210660 269890
rect 210608 269826 210660 269832
rect 210424 267028 210476 267034
rect 210424 266970 210476 266976
rect 209976 264302 210174 264330
rect 210620 264316 210648 269826
rect 211264 268394 211292 277780
rect 212460 275602 212488 277780
rect 213460 275664 213512 275670
rect 213460 275606 213512 275612
rect 212448 275596 212500 275602
rect 212448 275538 212500 275544
rect 213092 274372 213144 274378
rect 213092 274314 213144 274320
rect 211344 274304 211396 274310
rect 211344 274246 211396 274252
rect 211252 268388 211304 268394
rect 211252 268330 211304 268336
rect 210700 265600 210752 265606
rect 210700 265542 210752 265548
rect 210712 264330 210740 265542
rect 211356 264330 211384 274246
rect 212632 272944 212684 272950
rect 212632 272886 212684 272892
rect 211896 270020 211948 270026
rect 211896 269962 211948 269968
rect 210712 264302 211094 264330
rect 211356 264302 211554 264330
rect 211908 264316 211936 269962
rect 212356 269952 212408 269958
rect 212356 269894 212408 269900
rect 212368 264316 212396 269894
rect 212644 264330 212672 272886
rect 212908 270088 212960 270094
rect 212908 270030 212960 270036
rect 212920 264330 212948 270030
rect 213104 267734 213132 274314
rect 213472 268462 213500 275606
rect 213656 275466 213684 277780
rect 214852 275738 214880 277780
rect 215970 277766 216628 277794
rect 214840 275732 214892 275738
rect 214840 275674 214892 275680
rect 213644 275460 213696 275466
rect 213644 275402 213696 275408
rect 214564 275052 214616 275058
rect 214564 274994 214616 275000
rect 214104 274440 214156 274446
rect 214104 274382 214156 274388
rect 214012 271312 214064 271318
rect 214012 271254 214064 271260
rect 213460 268456 213512 268462
rect 213460 268398 213512 268404
rect 213104 267706 213408 267734
rect 213380 264330 213408 267706
rect 214024 265606 214052 271254
rect 214012 265600 214064 265606
rect 214012 265542 214064 265548
rect 214116 264330 214144 274382
rect 214576 267102 214604 274994
rect 216036 273080 216088 273086
rect 216036 273022 216088 273028
rect 215392 273012 215444 273018
rect 215392 272954 215444 272960
rect 214656 270156 214708 270162
rect 214656 270098 214708 270104
rect 214564 267096 214616 267102
rect 214564 267038 214616 267044
rect 212644 264302 212842 264330
rect 212920 264302 213302 264330
rect 213380 264302 213762 264330
rect 214116 264302 214222 264330
rect 214668 264316 214696 270098
rect 214748 265600 214800 265606
rect 214748 265542 214800 265548
rect 214760 264330 214788 265542
rect 215404 264330 215432 272954
rect 215944 270224 215996 270230
rect 215944 270166 215996 270172
rect 214760 264302 215050 264330
rect 215404 264302 215510 264330
rect 215956 264316 215984 270166
rect 216048 264330 216076 273022
rect 216600 268530 216628 277766
rect 216680 275936 216732 275942
rect 216680 275878 216732 275884
rect 216692 269822 216720 275878
rect 216956 270292 217008 270298
rect 216956 270234 217008 270240
rect 216680 269816 216732 269822
rect 216680 269758 216732 269764
rect 216588 268524 216640 268530
rect 216588 268466 216640 268472
rect 216864 268252 216916 268258
rect 216864 268194 216916 268200
rect 216048 264302 216430 264330
rect 216876 264316 216904 268194
rect 216968 264330 216996 270234
rect 217152 268598 217180 277780
rect 218244 274644 218296 274650
rect 218244 274586 218296 274592
rect 217140 268592 217192 268598
rect 217140 268534 217192 268540
rect 218152 268184 218204 268190
rect 218152 268126 218204 268132
rect 217692 267300 217744 267306
rect 217692 267242 217744 267248
rect 216968 264302 217350 264330
rect 217704 264316 217732 267242
rect 218164 264316 218192 268126
rect 218256 264330 218284 274586
rect 218348 268734 218376 277780
rect 218336 268728 218388 268734
rect 218336 268670 218388 268676
rect 219544 268666 219572 277780
rect 220636 275800 220688 275806
rect 220636 275742 220688 275748
rect 219624 274508 219676 274514
rect 219624 274450 219676 274456
rect 219532 268660 219584 268666
rect 219532 268602 219584 268608
rect 219072 266756 219124 266762
rect 219072 266698 219124 266704
rect 218256 264302 218638 264330
rect 219084 264316 219112 266698
rect 219636 264330 219664 274450
rect 220648 270366 220676 275742
rect 220740 274718 220768 277780
rect 221464 275120 221516 275126
rect 221464 275062 221516 275068
rect 220728 274712 220780 274718
rect 220728 274654 220780 274660
rect 220820 273148 220872 273154
rect 220820 273090 220872 273096
rect 219992 270360 220044 270366
rect 219992 270302 220044 270308
rect 220636 270360 220688 270366
rect 220636 270302 220688 270308
rect 219558 264302 219664 264330
rect 220004 264316 220032 270302
rect 220360 268048 220412 268054
rect 220360 267990 220412 267996
rect 220372 264316 220400 267990
rect 220832 264316 220860 273090
rect 220912 271380 220964 271386
rect 220912 271322 220964 271328
rect 220924 264330 220952 271322
rect 221476 267238 221504 275062
rect 221936 270774 221964 277780
rect 223132 275670 223160 277780
rect 223120 275664 223172 275670
rect 223120 275606 223172 275612
rect 224236 275602 224264 277780
rect 222476 275596 222528 275602
rect 222476 275538 222528 275544
rect 224224 275596 224276 275602
rect 224224 275538 224276 275544
rect 222200 274576 222252 274582
rect 222200 274518 222252 274524
rect 221924 270768 221976 270774
rect 221924 270710 221976 270716
rect 221740 267640 221792 267646
rect 221740 267582 221792 267588
rect 221464 267232 221516 267238
rect 221464 267174 221516 267180
rect 220924 264302 221306 264330
rect 221752 264316 221780 267582
rect 222212 264316 222240 274518
rect 222292 273216 222344 273222
rect 222292 273158 222344 273164
rect 222304 265606 222332 273158
rect 222488 272746 222516 275538
rect 224960 275528 225012 275534
rect 224960 275470 225012 275476
rect 223580 274712 223632 274718
rect 223580 274654 223632 274660
rect 222476 272740 222528 272746
rect 222476 272682 222528 272688
rect 222476 271448 222528 271454
rect 222476 271390 222528 271396
rect 222292 265600 222344 265606
rect 222292 265542 222344 265548
rect 222488 264330 222516 271390
rect 223592 271182 223620 274654
rect 224500 271652 224552 271658
rect 224500 271594 224552 271600
rect 223672 271584 223724 271590
rect 223672 271526 223724 271532
rect 223580 271176 223632 271182
rect 223580 271118 223632 271124
rect 223028 267980 223080 267986
rect 223028 267922 223080 267928
rect 222488 264302 222686 264330
rect 223040 264316 223068 267922
rect 223212 265600 223264 265606
rect 223212 265542 223264 265548
rect 223224 264330 223252 265542
rect 223684 264330 223712 271526
rect 224408 270360 224460 270366
rect 224408 270302 224460 270308
rect 223224 264302 223514 264330
rect 223684 264302 223974 264330
rect 224420 264316 224448 270302
rect 224512 264330 224540 271594
rect 224972 271454 225000 275470
rect 225432 274718 225460 277780
rect 225420 274712 225472 274718
rect 225420 274654 225472 274660
rect 225880 273896 225932 273902
rect 225880 273838 225932 273844
rect 225052 271516 225104 271522
rect 225052 271458 225104 271464
rect 224960 271448 225012 271454
rect 224960 271390 225012 271396
rect 225064 264330 225092 271458
rect 225788 266688 225840 266694
rect 225788 266630 225840 266636
rect 224512 264302 224894 264330
rect 225064 264302 225354 264330
rect 225800 264316 225828 266630
rect 225892 264330 225920 273838
rect 226432 271720 226484 271726
rect 226432 271662 226484 271668
rect 226444 264330 226472 271662
rect 226628 271250 226656 277780
rect 226984 275868 227036 275874
rect 226984 275810 227036 275816
rect 226892 272468 226944 272474
rect 226892 272410 226944 272416
rect 226616 271244 226668 271250
rect 226616 271186 226668 271192
rect 226708 268796 226760 268802
rect 226708 268738 226760 268744
rect 226720 264330 226748 268738
rect 226904 264602 226932 272410
rect 226996 267170 227024 275810
rect 227720 275732 227772 275738
rect 227720 275674 227772 275680
rect 227732 269890 227760 275674
rect 227824 275534 227852 277780
rect 227812 275528 227864 275534
rect 227812 275470 227864 275476
rect 229020 274242 229048 277780
rect 229836 274712 229888 274718
rect 229836 274654 229888 274660
rect 229008 274236 229060 274242
rect 229008 274178 229060 274184
rect 227812 271856 227864 271862
rect 227812 271798 227864 271804
rect 227720 269884 227772 269890
rect 227720 269826 227772 269832
rect 226984 267164 227036 267170
rect 226984 267106 227036 267112
rect 226904 264574 227208 264602
rect 227180 264330 227208 264574
rect 227824 264330 227852 271798
rect 228272 271788 228324 271794
rect 228272 271730 228324 271736
rect 228284 267734 228312 271730
rect 229284 271108 229336 271114
rect 229284 271050 229336 271056
rect 228284 267706 228588 267734
rect 228456 267436 228508 267442
rect 228456 267378 228508 267384
rect 225892 264302 226182 264330
rect 226444 264302 226642 264330
rect 226720 264302 227102 264330
rect 227180 264302 227562 264330
rect 227824 264302 228022 264330
rect 228468 264316 228496 267378
rect 228560 264330 228588 267706
rect 228560 264302 228850 264330
rect 229296 264316 229324 271050
rect 229848 269822 229876 274654
rect 230216 271318 230244 277780
rect 231124 273760 231176 273766
rect 231124 273702 231176 273708
rect 230204 271312 230256 271318
rect 230204 271254 230256 271260
rect 230664 271040 230716 271046
rect 230664 270982 230716 270988
rect 230204 270428 230256 270434
rect 230204 270370 230256 270376
rect 229468 269816 229520 269822
rect 229468 269758 229520 269764
rect 229836 269816 229888 269822
rect 229836 269758 229888 269764
rect 229480 264330 229508 269758
rect 229480 264302 229770 264330
rect 230216 264316 230244 270370
rect 230676 264316 230704 270982
rect 231136 267646 231164 273702
rect 231412 271386 231440 277780
rect 232530 277766 233188 277794
rect 231400 271380 231452 271386
rect 231400 271322 231452 271328
rect 232044 270972 232096 270978
rect 232044 270914 232096 270920
rect 231492 270496 231544 270502
rect 231492 270438 231544 270444
rect 231124 267640 231176 267646
rect 231124 267582 231176 267588
rect 231124 267504 231176 267510
rect 231124 267446 231176 267452
rect 231136 264316 231164 267446
rect 231504 264316 231532 270438
rect 232056 264330 232084 270914
rect 232872 269748 232924 269754
rect 232872 269690 232924 269696
rect 232412 267164 232464 267170
rect 232412 267106 232464 267112
rect 231978 264302 232084 264330
rect 232424 264316 232452 267106
rect 232884 264316 232912 269690
rect 233160 267170 233188 277766
rect 233712 272814 233740 277780
rect 234620 275460 234672 275466
rect 234620 275402 234672 275408
rect 233884 275392 233936 275398
rect 233884 275334 233936 275340
rect 233700 272808 233752 272814
rect 233700 272750 233752 272756
rect 233792 272400 233844 272406
rect 233792 272342 233844 272348
rect 233804 271402 233832 272342
rect 233896 271522 233924 275334
rect 233884 271516 233936 271522
rect 233884 271458 233936 271464
rect 233804 271374 233924 271402
rect 233424 270904 233476 270910
rect 233424 270846 233476 270852
rect 233148 267164 233200 267170
rect 233148 267106 233200 267112
rect 233436 264330 233464 270846
rect 233792 267708 233844 267714
rect 233792 267650 233844 267656
rect 233358 264302 233464 264330
rect 233804 264316 233832 267650
rect 233896 266422 233924 271374
rect 234632 270094 234660 275402
rect 234908 275262 234936 277780
rect 234896 275256 234948 275262
rect 234896 275198 234948 275204
rect 235908 275256 235960 275262
rect 235908 275198 235960 275204
rect 235356 270836 235408 270842
rect 235356 270778 235408 270784
rect 234620 270088 234672 270094
rect 234620 270030 234672 270036
rect 234160 269680 234212 269686
rect 234160 269622 234212 269628
rect 233884 266416 233936 266422
rect 233884 266358 233936 266364
rect 234172 264316 234200 269622
rect 235080 267232 235132 267238
rect 235080 267174 235132 267180
rect 234620 266416 234672 266422
rect 234620 266358 234672 266364
rect 234632 264316 234660 266358
rect 235092 264316 235120 267174
rect 235368 266422 235396 270778
rect 235540 269612 235592 269618
rect 235540 269554 235592 269560
rect 235356 266416 235408 266422
rect 235356 266358 235408 266364
rect 235552 264316 235580 269554
rect 235920 267238 235948 275198
rect 236104 269958 236132 277780
rect 237300 274310 237328 277780
rect 238510 277766 238708 277794
rect 237380 275324 237432 275330
rect 237380 275266 237432 275272
rect 237288 274304 237340 274310
rect 237288 274246 237340 274252
rect 236644 273828 236696 273834
rect 236644 273770 236696 273776
rect 236092 269952 236144 269958
rect 236092 269894 236144 269900
rect 236000 267640 236052 267646
rect 236000 267582 236052 267588
rect 235908 267232 235960 267238
rect 235908 267174 235960 267180
rect 236012 264316 236040 267582
rect 236656 267442 236684 273770
rect 237392 270026 237420 275266
rect 238116 270768 238168 270774
rect 238116 270710 238168 270716
rect 237380 270020 237432 270026
rect 237380 269962 237432 269968
rect 236920 269544 236972 269550
rect 236920 269486 236972 269492
rect 236644 267436 236696 267442
rect 236644 267378 236696 267384
rect 236460 266960 236512 266966
rect 236460 266902 236512 266908
rect 236472 264316 236500 266902
rect 236932 264316 236960 269486
rect 237288 268116 237340 268122
rect 237288 268058 237340 268064
rect 237300 264316 237328 268058
rect 238128 267306 238156 270710
rect 238208 269476 238260 269482
rect 238208 269418 238260 269424
rect 238116 267300 238168 267306
rect 238116 267242 238168 267248
rect 237748 267096 237800 267102
rect 237748 267038 237800 267044
rect 237760 264316 237788 267038
rect 238220 264316 238248 269418
rect 238680 267102 238708 277766
rect 239600 275466 239628 277780
rect 239588 275460 239640 275466
rect 239588 275402 239640 275408
rect 240796 275330 240824 277780
rect 241428 275664 241480 275670
rect 241428 275606 241480 275612
rect 240784 275324 240836 275330
rect 240784 275266 240836 275272
rect 240232 273964 240284 273970
rect 240232 273906 240284 273912
rect 240140 273692 240192 273698
rect 240140 273634 240192 273640
rect 239404 273624 239456 273630
rect 239404 273566 239456 273572
rect 239220 272332 239272 272338
rect 239220 272274 239272 272280
rect 238852 272264 238904 272270
rect 238852 272206 238904 272212
rect 238668 267096 238720 267102
rect 238668 267038 238720 267044
rect 238668 266416 238720 266422
rect 238668 266358 238720 266364
rect 238680 264316 238708 266358
rect 238864 265606 238892 272206
rect 239128 267028 239180 267034
rect 239128 266970 239180 266976
rect 238852 265600 238904 265606
rect 238852 265542 238904 265548
rect 239140 264316 239168 266970
rect 239232 264330 239260 272274
rect 239416 266490 239444 273566
rect 239404 266484 239456 266490
rect 239404 266426 239456 266432
rect 240152 265606 240180 273634
rect 239680 265600 239732 265606
rect 239680 265542 239732 265548
rect 240140 265600 240192 265606
rect 240140 265542 240192 265548
rect 239692 264330 239720 265542
rect 240244 265538 240272 273906
rect 240324 272536 240376 272542
rect 240324 272478 240376 272484
rect 240232 265532 240284 265538
rect 240232 265474 240284 265480
rect 240336 264330 240364 272478
rect 241440 271590 241468 275606
rect 241888 272604 241940 272610
rect 241888 272546 241940 272552
rect 241612 272196 241664 272202
rect 241612 272138 241664 272144
rect 241428 271584 241480 271590
rect 241428 271526 241480 271532
rect 241624 265606 241652 272138
rect 241796 267436 241848 267442
rect 241796 267378 241848 267384
rect 240508 265600 240560 265606
rect 240508 265542 240560 265548
rect 241612 265600 241664 265606
rect 241612 265542 241664 265548
rect 240520 264330 240548 265542
rect 241060 265532 241112 265538
rect 241060 265474 241112 265480
rect 241072 264330 241100 265474
rect 239232 264302 239614 264330
rect 239692 264302 239982 264330
rect 240336 264302 240442 264330
rect 240520 264302 240902 264330
rect 241072 264302 241362 264330
rect 241808 264316 241836 267378
rect 241900 264330 241928 272546
rect 241992 272542 242020 277780
rect 243188 274854 243216 277780
rect 243544 275596 243596 275602
rect 243544 275538 243596 275544
rect 243176 274848 243228 274854
rect 243176 274790 243228 274796
rect 242900 274100 242952 274106
rect 242900 274042 242952 274048
rect 241980 272536 242032 272542
rect 241980 272478 242032 272484
rect 242808 268728 242860 268734
rect 242808 268670 242860 268676
rect 242820 266422 242848 268670
rect 242808 266416 242860 266422
rect 242808 266358 242860 266364
rect 242348 265600 242400 265606
rect 242348 265542 242400 265548
rect 242360 264330 242388 265542
rect 242912 265538 242940 274042
rect 243556 274038 243584 275538
rect 242992 274032 243044 274038
rect 242992 273974 243044 273980
rect 243544 274032 243596 274038
rect 243544 273974 243596 273980
rect 243004 265606 243032 273974
rect 243084 272672 243136 272678
rect 243084 272614 243136 272620
rect 242992 265600 243044 265606
rect 242992 265542 243044 265548
rect 242900 265532 242952 265538
rect 242900 265474 242952 265480
rect 241900 264302 242282 264330
rect 242360 264302 242650 264330
rect 243096 264316 243124 272614
rect 244384 270026 244412 277780
rect 244556 274168 244608 274174
rect 244556 274110 244608 274116
rect 244372 270020 244424 270026
rect 244372 269962 244424 269968
rect 244464 266484 244516 266490
rect 244464 266426 244516 266432
rect 243268 265600 243320 265606
rect 243268 265542 243320 265548
rect 243280 264330 243308 265542
rect 243636 265532 243688 265538
rect 243636 265474 243688 265480
rect 243648 264330 243676 265474
rect 243280 264302 243570 264330
rect 243648 264302 244030 264330
rect 244476 264316 244504 266426
rect 244568 264330 244596 274110
rect 245580 273902 245608 277780
rect 245844 274848 245896 274854
rect 245844 274790 245896 274796
rect 245568 273896 245620 273902
rect 245568 273838 245620 273844
rect 245292 270088 245344 270094
rect 245292 270030 245344 270036
rect 244568 264302 244950 264330
rect 245304 264316 245332 270030
rect 245856 268462 245884 274790
rect 246776 272610 246804 277780
rect 247894 277766 248368 277794
rect 247224 272740 247276 272746
rect 247224 272682 247276 272688
rect 246764 272604 246816 272610
rect 246764 272546 246816 272552
rect 246028 271516 246080 271522
rect 246028 271458 246080 271464
rect 245936 271448 245988 271454
rect 245936 271390 245988 271396
rect 245752 268456 245804 268462
rect 245752 268398 245804 268404
rect 245844 268456 245896 268462
rect 245844 268398 245896 268404
rect 245764 264316 245792 268398
rect 245948 268274 245976 271390
rect 245856 268246 245976 268274
rect 245856 264994 245884 268246
rect 245844 264988 245896 264994
rect 245844 264930 245896 264936
rect 246040 264330 246068 271458
rect 247132 268388 247184 268394
rect 247132 268330 247184 268336
rect 246396 264988 246448 264994
rect 246396 264930 246448 264936
rect 246408 264330 246436 264930
rect 246040 264302 246238 264330
rect 246408 264302 246698 264330
rect 247144 264316 247172 268330
rect 247236 264330 247264 272682
rect 248052 270156 248104 270162
rect 248052 270098 248104 270104
rect 247236 264302 247618 264330
rect 248064 264316 248092 270098
rect 248340 270094 248368 277766
rect 249076 275398 249104 277780
rect 249616 275528 249668 275534
rect 249616 275470 249668 275476
rect 249064 275392 249116 275398
rect 249064 275334 249116 275340
rect 248328 270088 248380 270094
rect 248328 270030 248380 270036
rect 248420 269884 248472 269890
rect 248420 269826 248472 269832
rect 248432 264316 248460 269826
rect 249628 269074 249656 275470
rect 249708 275460 249760 275466
rect 249708 275402 249760 275408
rect 249616 269068 249668 269074
rect 249616 269010 249668 269016
rect 249720 269006 249748 275402
rect 250272 274854 250300 277780
rect 251468 275738 251496 277780
rect 252678 277766 252968 277794
rect 251456 275732 251508 275738
rect 251456 275674 251508 275680
rect 252376 275732 252428 275738
rect 252376 275674 252428 275680
rect 250260 274848 250312 274854
rect 250260 274790 250312 274796
rect 251640 274032 251692 274038
rect 251640 273974 251692 273980
rect 251272 271584 251324 271590
rect 251272 271526 251324 271532
rect 250352 271176 250404 271182
rect 250352 271118 250404 271124
rect 249708 269000 249760 269006
rect 249708 268942 249760 268948
rect 250260 268660 250312 268666
rect 250260 268602 250312 268608
rect 249340 268592 249392 268598
rect 249340 268534 249392 268540
rect 248880 268524 248932 268530
rect 248880 268466 248932 268472
rect 248892 264316 248920 268466
rect 249352 264316 249380 268534
rect 249800 266416 249852 266422
rect 249800 266358 249852 266364
rect 249812 264316 249840 266358
rect 250272 264316 250300 268602
rect 250364 264330 250392 271118
rect 251088 267300 251140 267306
rect 251088 267242 251140 267248
rect 250364 264302 250746 264330
rect 251100 264316 251128 267242
rect 251284 264330 251312 271526
rect 251652 264330 251680 273974
rect 252388 267034 252416 275674
rect 252652 271244 252704 271250
rect 252652 271186 252704 271192
rect 252468 269816 252520 269822
rect 252468 269758 252520 269764
rect 252376 267028 252428 267034
rect 252376 266970 252428 266976
rect 251284 264302 251574 264330
rect 251652 264302 252034 264330
rect 252480 264316 252508 269758
rect 252664 264330 252692 271186
rect 252940 271182 252968 277766
rect 253480 274236 253532 274242
rect 253480 274178 253532 274184
rect 252928 271176 252980 271182
rect 252928 271118 252980 271124
rect 253388 269068 253440 269074
rect 253388 269010 253440 269016
rect 252664 264302 252954 264330
rect 253400 264316 253428 269010
rect 253492 264330 253520 274178
rect 253860 274038 253888 277780
rect 255070 277766 255268 277794
rect 254216 274848 254268 274854
rect 254216 274790 254268 274796
rect 253848 274032 253900 274038
rect 253848 273974 253900 273980
rect 254228 271318 254256 274790
rect 254308 271380 254360 271386
rect 254308 271322 254360 271328
rect 254032 271312 254084 271318
rect 254032 271254 254084 271260
rect 254216 271312 254268 271318
rect 254216 271254 254268 271260
rect 254044 264330 254072 271254
rect 254320 264330 254348 271322
rect 255240 267170 255268 277766
rect 255504 272808 255556 272814
rect 255504 272750 255556 272756
rect 255136 267164 255188 267170
rect 255136 267106 255188 267112
rect 255228 267164 255280 267170
rect 255228 267106 255280 267112
rect 253492 264302 253782 264330
rect 254044 264302 254242 264330
rect 254320 264302 254702 264330
rect 255148 264316 255176 267106
rect 255516 264330 255544 272750
rect 256160 271250 256188 277780
rect 257370 277766 258028 277794
rect 256884 274304 256936 274310
rect 256884 274246 256936 274252
rect 256148 271244 256200 271250
rect 256148 271186 256200 271192
rect 256424 269952 256476 269958
rect 256424 269894 256476 269900
rect 256056 267232 256108 267238
rect 256056 267174 256108 267180
rect 255516 264302 255622 264330
rect 256068 264316 256096 267174
rect 256436 264316 256464 269894
rect 256896 264316 256924 274246
rect 257804 269000 257856 269006
rect 257804 268942 257856 268948
rect 257344 267096 257396 267102
rect 257344 267038 257396 267044
rect 257356 264316 257384 267038
rect 257816 264316 257844 268942
rect 258000 268394 258028 277766
rect 258552 275806 258580 277780
rect 258540 275800 258592 275806
rect 258540 275742 258592 275748
rect 258264 275324 258316 275330
rect 258264 275266 258316 275272
rect 257988 268388 258040 268394
rect 257988 268330 258040 268336
rect 258276 264316 258304 275266
rect 259748 275262 259776 277780
rect 260748 275392 260800 275398
rect 260748 275334 260800 275340
rect 259736 275256 259788 275262
rect 259736 275198 259788 275204
rect 260760 274530 260788 275334
rect 260944 274990 260972 277780
rect 260932 274984 260984 274990
rect 260932 274926 260984 274932
rect 262140 274786 262168 277780
rect 263244 275330 263272 277780
rect 263232 275324 263284 275330
rect 263232 275266 263284 275272
rect 262128 274780 262180 274786
rect 262128 274722 262180 274728
rect 264440 274718 264468 277780
rect 265650 277766 266308 277794
rect 264612 275800 264664 275806
rect 264612 275742 264664 275748
rect 264428 274712 264480 274718
rect 264428 274654 264480 274660
rect 260760 274502 261064 274530
rect 259644 273896 259696 273902
rect 259644 273838 259696 273844
rect 258356 272536 258408 272542
rect 258356 272478 258408 272484
rect 258368 264330 258396 272478
rect 259552 270020 259604 270026
rect 259552 269962 259604 269968
rect 259184 268456 259236 268462
rect 259184 268398 259236 268404
rect 258368 264302 258750 264330
rect 259196 264316 259224 268398
rect 259564 264316 259592 269962
rect 259656 264330 259684 273838
rect 260104 272604 260156 272610
rect 260104 272546 260156 272552
rect 260116 264330 260144 272546
rect 260932 270088 260984 270094
rect 260932 270030 260984 270036
rect 259656 264302 260038 264330
rect 260116 264302 260498 264330
rect 260944 264316 260972 270030
rect 261036 264330 261064 274502
rect 262772 274032 262824 274038
rect 262772 273974 262824 273980
rect 261484 271312 261536 271318
rect 261484 271254 261536 271260
rect 261496 264330 261524 271254
rect 262312 271176 262364 271182
rect 262312 271118 262364 271124
rect 262220 267028 262272 267034
rect 262220 266970 262272 266976
rect 261036 264302 261418 264330
rect 261496 264302 261878 264330
rect 262232 264316 262260 266970
rect 262324 264330 262352 271118
rect 262784 264330 262812 273974
rect 263692 271244 263744 271250
rect 263692 271186 263744 271192
rect 263600 267164 263652 267170
rect 263600 267106 263652 267112
rect 262324 264302 262706 264330
rect 262784 264302 263166 264330
rect 263612 264316 263640 267106
rect 263704 264330 263732 271186
rect 264520 268388 264572 268394
rect 264520 268330 264572 268336
rect 263704 264302 264086 264330
rect 264532 264316 264560 268330
rect 264624 264330 264652 275742
rect 264980 275256 265032 275262
rect 264980 275198 265032 275204
rect 264992 264330 265020 275198
rect 265072 274984 265124 274990
rect 265072 274926 265124 274932
rect 265084 267734 265112 274926
rect 265900 274780 265952 274786
rect 265900 274722 265952 274728
rect 265084 267706 265480 267734
rect 265452 264330 265480 267706
rect 265912 264330 265940 274722
rect 266280 274666 266308 277766
rect 266544 275324 266596 275330
rect 266544 275266 266596 275272
rect 266280 274638 266400 274666
rect 266372 265606 266400 274638
rect 266360 265600 266412 265606
rect 266360 265542 266412 265548
rect 266556 264330 266584 275266
rect 266832 274718 266860 277780
rect 268042 277766 268148 277794
rect 266728 274712 266780 274718
rect 266728 274654 266780 274660
rect 266820 274712 266872 274718
rect 266820 274654 266872 274660
rect 267740 274712 267792 274718
rect 267740 274654 267792 274660
rect 266740 267734 266768 274654
rect 266740 267706 266860 267734
rect 266832 264330 266860 267706
rect 267280 265600 267332 265606
rect 267280 265542 267332 265548
rect 267292 264330 267320 265542
rect 267752 264330 267780 274654
rect 268120 264330 268148 277766
rect 269224 267734 269252 277780
rect 269040 267706 269252 267734
rect 269408 277766 270434 277794
rect 270512 277766 271538 277794
rect 272076 277766 272734 277794
rect 273272 277766 273930 277794
rect 274652 277766 275126 277794
rect 269040 264330 269068 267706
rect 264624 264302 264914 264330
rect 264992 264302 265374 264330
rect 265452 264302 265834 264330
rect 265912 264302 266294 264330
rect 266556 264302 266754 264330
rect 266832 264302 267214 264330
rect 267292 264302 267582 264330
rect 267752 264302 268042 264330
rect 268120 264302 268502 264330
rect 268962 264302 269068 264330
rect 269408 264316 269436 277766
rect 270512 267734 270540 277766
rect 270236 267706 270540 267734
rect 270236 264330 270264 267706
rect 271604 266620 271656 266626
rect 271604 266562 271656 266568
rect 271144 266552 271196 266558
rect 271144 266494 271196 266500
rect 270684 266484 270736 266490
rect 270684 266426 270736 266432
rect 270316 266416 270368 266422
rect 270316 266358 270368 266364
rect 269882 264302 270264 264330
rect 270328 264316 270356 266358
rect 270696 264316 270724 266426
rect 271156 264316 271184 266494
rect 271616 264316 271644 266562
rect 272076 266422 272104 277766
rect 273168 273624 273220 273630
rect 273168 273566 273220 273572
rect 272524 267232 272576 267238
rect 272524 267174 272576 267180
rect 272432 267028 272484 267034
rect 272432 266970 272484 266976
rect 272064 266416 272116 266422
rect 272064 266358 272116 266364
rect 272444 264330 272472 266970
rect 272090 264302 272472 264330
rect 272536 264316 272564 267174
rect 273180 264330 273208 273566
rect 273272 266490 273300 277766
rect 273812 271924 273864 271930
rect 273812 271866 273864 271872
rect 273352 271312 273404 271318
rect 273352 271254 273404 271260
rect 273260 266484 273312 266490
rect 273260 266426 273312 266432
rect 273010 264302 273208 264330
rect 273364 264316 273392 271254
rect 273824 264316 273852 271866
rect 274272 269952 274324 269958
rect 274272 269894 274324 269900
rect 274284 264316 274312 269894
rect 274652 266558 274680 277766
rect 275928 274032 275980 274038
rect 275928 273974 275980 273980
rect 275940 273254 275968 273974
rect 275572 273226 275968 273254
rect 274732 272536 274784 272542
rect 274732 272478 274784 272484
rect 274640 266552 274692 266558
rect 274640 266494 274692 266500
rect 274744 264316 274772 272478
rect 275572 264330 275600 273226
rect 275652 271380 275704 271386
rect 275652 271322 275704 271328
rect 275218 264302 275600 264330
rect 275664 264316 275692 271322
rect 276020 267368 276072 267374
rect 276020 267310 276072 267316
rect 276032 264316 276060 267310
rect 276308 266626 276336 277780
rect 277518 277766 277808 277794
rect 277308 273964 277360 273970
rect 277308 273906 277360 273912
rect 276940 269884 276992 269890
rect 276940 269826 276992 269832
rect 276480 267708 276532 267714
rect 276480 267650 276532 267656
rect 276296 266620 276348 266626
rect 276296 266562 276348 266568
rect 276492 264316 276520 267650
rect 276952 264316 276980 269826
rect 277320 267714 277348 273906
rect 277400 268728 277452 268734
rect 277400 268670 277452 268676
rect 277308 267708 277360 267714
rect 277308 267650 277360 267656
rect 277412 264316 277440 268670
rect 277780 267034 277808 277766
rect 277872 277766 278714 277794
rect 277872 267238 277900 277766
rect 279424 274100 279476 274106
rect 279424 274042 279476 274048
rect 279148 271244 279200 271250
rect 279148 271186 279200 271192
rect 278688 269816 278740 269822
rect 278688 269758 278740 269764
rect 278320 267436 278372 267442
rect 278320 267378 278372 267384
rect 277860 267232 277912 267238
rect 277860 267174 277912 267180
rect 277768 267028 277820 267034
rect 277768 266970 277820 266976
rect 277860 266620 277912 266626
rect 277860 266562 277912 266568
rect 277872 264316 277900 266562
rect 278332 264316 278360 267378
rect 278700 264316 278728 269758
rect 279160 264316 279188 271186
rect 279436 267374 279464 274042
rect 279804 273630 279832 277780
rect 279792 273624 279844 273630
rect 279792 273566 279844 273572
rect 281000 271318 281028 277780
rect 282196 271930 282224 277780
rect 282932 277766 283406 277794
rect 282736 272808 282788 272814
rect 282736 272750 282788 272756
rect 282184 271924 282236 271930
rect 282184 271866 282236 271872
rect 281540 271448 281592 271454
rect 281540 271390 281592 271396
rect 280988 271312 281040 271318
rect 280988 271254 281040 271260
rect 280528 271176 280580 271182
rect 280528 271118 280580 271124
rect 280068 268660 280120 268666
rect 280068 268602 280120 268608
rect 279424 267368 279476 267374
rect 279424 267310 279476 267316
rect 279608 267028 279660 267034
rect 279608 266970 279660 266976
rect 279620 264316 279648 266970
rect 280080 264316 280108 268602
rect 280540 264316 280568 271118
rect 280988 271040 281040 271046
rect 280988 270982 281040 270988
rect 281000 264316 281028 270982
rect 281448 268456 281500 268462
rect 281448 268398 281500 268404
rect 281460 264316 281488 268398
rect 281552 267442 281580 271390
rect 281540 267436 281592 267442
rect 281540 267378 281592 267384
rect 281816 267300 281868 267306
rect 281816 267242 281868 267248
rect 281828 264316 281856 267242
rect 282276 266756 282328 266762
rect 282276 266698 282328 266704
rect 282288 264316 282316 266698
rect 282748 264316 282776 272750
rect 282932 269958 282960 277766
rect 284588 272542 284616 277780
rect 285784 274038 285812 277780
rect 286520 277766 286902 277794
rect 285772 274032 285824 274038
rect 285772 273974 285824 273980
rect 285588 272740 285640 272746
rect 285588 272682 285640 272688
rect 285404 272672 285456 272678
rect 285404 272614 285456 272620
rect 284576 272536 284628 272542
rect 284576 272478 284628 272484
rect 282920 269952 282972 269958
rect 282920 269894 282972 269900
rect 283564 269952 283616 269958
rect 283564 269894 283616 269900
rect 283196 268524 283248 268530
rect 283196 268466 283248 268472
rect 283208 264316 283236 268466
rect 283576 266626 283604 269894
rect 284116 268388 284168 268394
rect 284116 268330 284168 268336
rect 283656 267436 283708 267442
rect 283656 267378 283708 267384
rect 283564 266620 283616 266626
rect 283564 266562 283616 266568
rect 283668 264316 283696 267378
rect 284128 264316 284156 268330
rect 284944 267572 284996 267578
rect 284944 267514 284996 267520
rect 284484 266416 284536 266422
rect 284484 266358 284536 266364
rect 284496 264316 284524 266358
rect 284956 264316 284984 267514
rect 285416 264316 285444 272614
rect 285600 267442 285628 272682
rect 285864 272604 285916 272610
rect 285864 272546 285916 272552
rect 285588 267436 285640 267442
rect 285588 267378 285640 267384
rect 285876 264316 285904 272546
rect 286520 271386 286548 277766
rect 288084 274106 288112 277780
rect 288348 274304 288400 274310
rect 288348 274246 288400 274252
rect 288072 274100 288124 274106
rect 288072 274042 288124 274048
rect 287704 274032 287756 274038
rect 287704 273974 287756 273980
rect 286784 272536 286836 272542
rect 286784 272478 286836 272484
rect 286508 271380 286560 271386
rect 286508 271322 286560 271328
rect 286324 267164 286376 267170
rect 286324 267106 286376 267112
rect 286336 264316 286364 267106
rect 286796 264316 286824 272478
rect 286968 270972 287020 270978
rect 286968 270914 287020 270920
rect 286980 267306 287008 270914
rect 287612 267708 287664 267714
rect 287612 267650 287664 267656
rect 287152 267504 287204 267510
rect 287152 267446 287204 267452
rect 286968 267300 287020 267306
rect 286968 267242 287020 267248
rect 287164 264316 287192 267446
rect 287624 264316 287652 267650
rect 287716 267034 287744 273974
rect 287796 271312 287848 271318
rect 287796 271254 287848 271260
rect 287808 270978 287836 271254
rect 287796 270972 287848 270978
rect 287796 270914 287848 270920
rect 288360 267714 288388 274246
rect 289280 273970 289308 277780
rect 289832 277766 290490 277794
rect 291212 277766 291686 277794
rect 292592 277766 292882 277794
rect 289636 274508 289688 274514
rect 289636 274450 289688 274456
rect 289268 273964 289320 273970
rect 289268 273906 289320 273912
rect 288440 272876 288492 272882
rect 288440 272818 288492 272824
rect 288348 267708 288400 267714
rect 288348 267650 288400 267656
rect 288072 267368 288124 267374
rect 288072 267310 288124 267316
rect 287704 267028 287756 267034
rect 287704 266970 287756 266976
rect 288084 264316 288112 267310
rect 288452 266762 288480 272818
rect 289648 267306 289676 274450
rect 289728 274100 289780 274106
rect 289728 274042 289780 274048
rect 288532 267300 288584 267306
rect 288532 267242 288584 267248
rect 289636 267300 289688 267306
rect 289636 267242 289688 267248
rect 288440 266756 288492 266762
rect 288440 266698 288492 266704
rect 288544 264316 288572 267242
rect 289740 267186 289768 274042
rect 289832 269890 289860 277766
rect 291108 273964 291160 273970
rect 291108 273906 291160 273912
rect 289820 269884 289872 269890
rect 289820 269826 289872 269832
rect 290740 269544 290792 269550
rect 290740 269486 290792 269492
rect 289912 268592 289964 268598
rect 289912 268534 289964 268540
rect 289820 267708 289872 267714
rect 289820 267650 289872 267656
rect 289372 267158 289768 267186
rect 289372 264330 289400 267158
rect 289452 267096 289504 267102
rect 289452 267038 289504 267044
rect 289018 264302 289400 264330
rect 289464 264316 289492 267038
rect 289832 264316 289860 267650
rect 289924 266422 289952 268534
rect 290280 267232 290332 267238
rect 290280 267174 290332 267180
rect 289912 266416 289964 266422
rect 289912 266358 289964 266364
rect 290292 264316 290320 267174
rect 290752 264316 290780 269486
rect 291120 267714 291148 273906
rect 291212 268734 291240 277766
rect 291844 274440 291896 274446
rect 291844 274382 291896 274388
rect 291200 268728 291252 268734
rect 291200 268670 291252 268676
rect 291108 267708 291160 267714
rect 291108 267650 291160 267656
rect 291856 267578 291884 274382
rect 292592 269958 292620 277766
rect 293684 274236 293736 274242
rect 293684 274178 293736 274184
rect 293408 270088 293460 270094
rect 293408 270030 293460 270036
rect 292580 269952 292632 269958
rect 292580 269894 292632 269900
rect 292580 269680 292632 269686
rect 292580 269622 292632 269628
rect 292120 269612 292172 269618
rect 292120 269554 292172 269560
rect 291844 267572 291896 267578
rect 291844 267514 291896 267520
rect 291200 267028 291252 267034
rect 291200 266970 291252 266976
rect 291212 264316 291240 266970
rect 291660 266484 291712 266490
rect 291660 266426 291712 266432
rect 291672 264316 291700 266426
rect 292132 264316 292160 269554
rect 292592 264316 292620 269622
rect 292948 267300 293000 267306
rect 292948 267242 293000 267248
rect 292960 264316 292988 267242
rect 293420 264316 293448 270030
rect 293696 264330 293724 274178
rect 294064 271454 294092 277780
rect 294156 277766 295182 277794
rect 294052 271448 294104 271454
rect 294052 271390 294104 271396
rect 294156 269822 294184 277766
rect 295984 274372 296036 274378
rect 295984 274314 296036 274320
rect 295248 271856 295300 271862
rect 295248 271798 295300 271804
rect 294788 269884 294840 269890
rect 294788 269826 294840 269832
rect 294144 269816 294196 269822
rect 294144 269758 294196 269764
rect 294328 266416 294380 266422
rect 294328 266358 294380 266364
rect 293696 264302 293894 264330
rect 294340 264316 294368 266358
rect 294800 264316 294828 269826
rect 295156 267572 295208 267578
rect 295156 267514 295208 267520
rect 295168 264330 295196 267514
rect 295260 266422 295288 271798
rect 295996 266490 296024 274314
rect 296364 271386 296392 277780
rect 297364 274644 297416 274650
rect 297364 274586 297416 274592
rect 296444 271788 296496 271794
rect 296444 271730 296496 271736
rect 296352 271380 296404 271386
rect 296352 271322 296404 271328
rect 296076 269748 296128 269754
rect 296076 269690 296128 269696
rect 295984 266484 296036 266490
rect 295984 266426 296036 266432
rect 295248 266416 295300 266422
rect 295248 266358 295300 266364
rect 295616 266416 295668 266422
rect 295616 266358 295668 266364
rect 295168 264302 295274 264330
rect 295628 264316 295656 266358
rect 296088 264316 296116 269690
rect 296456 266422 296484 271730
rect 296536 270496 296588 270502
rect 296536 270438 296588 270444
rect 296444 266416 296496 266422
rect 296444 266358 296496 266364
rect 296548 264316 296576 270438
rect 297376 267374 297404 274586
rect 297560 274038 297588 277780
rect 298112 277766 298770 277794
rect 298008 274168 298060 274174
rect 298008 274110 298060 274116
rect 297548 274032 297600 274038
rect 297548 273974 297600 273980
rect 297456 270428 297508 270434
rect 297456 270370 297508 270376
rect 297364 267368 297416 267374
rect 297364 267310 297416 267316
rect 296996 266824 297048 266830
rect 296996 266766 297048 266772
rect 297008 264316 297036 266766
rect 297468 264316 297496 270370
rect 298020 264330 298048 274110
rect 298112 268666 298140 277766
rect 299952 271250 299980 277780
rect 300768 271720 300820 271726
rect 300768 271662 300820 271668
rect 299940 271244 299992 271250
rect 299940 271186 299992 271192
rect 298744 270360 298796 270366
rect 298744 270302 298796 270308
rect 298100 268660 298152 268666
rect 298100 268602 298152 268608
rect 298284 267436 298336 267442
rect 298284 267378 298336 267384
rect 297942 264302 298048 264330
rect 298296 264316 298324 267378
rect 298756 264316 298784 270302
rect 300124 270292 300176 270298
rect 300124 270234 300176 270240
rect 299204 267708 299256 267714
rect 299204 267650 299256 267656
rect 299216 264316 299244 267650
rect 299664 266416 299716 266422
rect 299664 266358 299716 266364
rect 299676 264316 299704 266358
rect 300136 264316 300164 270234
rect 300584 267640 300636 267646
rect 300584 267582 300636 267588
rect 300596 264316 300624 267582
rect 300780 266422 300808 271662
rect 301148 271182 301176 277780
rect 302344 277394 302372 277780
rect 302252 277366 302372 277394
rect 301504 272468 301556 272474
rect 301504 272410 301556 272416
rect 301136 271176 301188 271182
rect 301136 271118 301188 271124
rect 301412 270224 301464 270230
rect 301412 270166 301464 270172
rect 300952 267368 301004 267374
rect 300952 267310 301004 267316
rect 300768 266416 300820 266422
rect 300768 266358 300820 266364
rect 300964 264316 300992 267310
rect 301424 264316 301452 270166
rect 301516 267510 301544 272410
rect 301872 270156 301924 270162
rect 301872 270098 301924 270104
rect 301504 267504 301556 267510
rect 301504 267446 301556 267452
rect 301884 264316 301912 270098
rect 302252 268462 302280 277366
rect 303344 274032 303396 274038
rect 303344 273974 303396 273980
rect 303160 271652 303212 271658
rect 303160 271594 303212 271600
rect 302240 268456 302292 268462
rect 302240 268398 302292 268404
rect 302332 266416 302384 266422
rect 302332 266358 302384 266364
rect 302344 264316 302372 266358
rect 303172 264330 303200 271594
rect 303356 270026 303384 273974
rect 303448 271318 303476 277780
rect 303528 273216 303580 273222
rect 303528 273158 303580 273164
rect 303436 271312 303488 271318
rect 303436 271254 303488 271260
rect 303540 270484 303568 273158
rect 304644 272882 304672 277780
rect 305644 273828 305696 273834
rect 305644 273770 305696 273776
rect 304632 272876 304684 272882
rect 304632 272818 304684 272824
rect 304448 271584 304500 271590
rect 304448 271526 304500 271532
rect 303448 270456 303568 270484
rect 303344 270020 303396 270026
rect 303344 269962 303396 269968
rect 303448 266422 303476 270456
rect 303528 270020 303580 270026
rect 303528 269962 303580 269968
rect 303436 266416 303488 266422
rect 303436 266358 303488 266364
rect 303540 264330 303568 269962
rect 303712 269068 303764 269074
rect 303712 269010 303764 269016
rect 302818 264302 303200 264330
rect 303278 264302 303568 264330
rect 303724 264316 303752 269010
rect 304460 264330 304488 271526
rect 304540 270020 304592 270026
rect 304540 269962 304592 269968
rect 304106 264302 304488 264330
rect 304552 264316 304580 269962
rect 305656 267170 305684 273770
rect 305840 272814 305868 277780
rect 306392 277766 307050 277794
rect 306288 273148 306340 273154
rect 306288 273090 306340 273096
rect 305828 272808 305880 272814
rect 305828 272750 305880 272756
rect 306196 271516 306248 271522
rect 306196 271458 306248 271464
rect 305644 267164 305696 267170
rect 305644 267106 305696 267112
rect 305920 266688 305972 266694
rect 305920 266630 305972 266636
rect 305000 266484 305052 266490
rect 305000 266426 305052 266432
rect 305012 264316 305040 266426
rect 305460 266416 305512 266422
rect 305460 266358 305512 266364
rect 305472 264316 305500 266358
rect 305932 264316 305960 266630
rect 306208 266422 306236 271458
rect 306300 266490 306328 273090
rect 306392 268530 306420 277766
rect 307024 273896 307076 273902
rect 307024 273838 307076 273844
rect 306656 268932 306708 268938
rect 306656 268874 306708 268880
rect 306380 268524 306432 268530
rect 306380 268466 306432 268472
rect 306380 267504 306432 267510
rect 306380 267446 306432 267452
rect 306392 267102 306420 267446
rect 306380 267096 306432 267102
rect 306380 267038 306432 267044
rect 306288 266484 306340 266490
rect 306288 266426 306340 266432
rect 306196 266416 306248 266422
rect 306196 266358 306248 266364
rect 306668 264330 306696 268874
rect 307036 267238 307064 273838
rect 308232 272746 308260 277780
rect 309152 277766 309442 277794
rect 308220 272740 308272 272746
rect 308220 272682 308272 272688
rect 307484 271448 307536 271454
rect 307484 271390 307536 271396
rect 307024 267232 307076 267238
rect 307024 267174 307076 267180
rect 307496 266422 307524 271390
rect 307576 271380 307628 271386
rect 307576 271322 307628 271328
rect 306748 266416 306800 266422
rect 306748 266358 306800 266364
rect 307484 266416 307536 266422
rect 307484 266358 307536 266364
rect 306406 264302 306696 264330
rect 306760 264316 306788 266358
rect 307588 264330 307616 271322
rect 308956 271312 309008 271318
rect 308956 271254 309008 271260
rect 308864 269000 308916 269006
rect 308864 268942 308916 268948
rect 307668 268320 307720 268326
rect 307668 268262 307720 268268
rect 307234 264302 307616 264330
rect 307680 264316 307708 268262
rect 308588 266620 308640 266626
rect 308588 266562 308640 266568
rect 308128 266416 308180 266422
rect 308128 266358 308180 266364
rect 308140 264316 308168 266358
rect 308600 264316 308628 266562
rect 308876 264330 308904 268942
rect 308968 266422 308996 271254
rect 309152 268394 309180 277766
rect 309784 274576 309836 274582
rect 309784 274518 309836 274524
rect 309140 268388 309192 268394
rect 309140 268330 309192 268336
rect 309324 267708 309376 267714
rect 309324 267650 309376 267656
rect 309336 267306 309364 267650
rect 309324 267300 309376 267306
rect 309324 267242 309376 267248
rect 309796 267238 309824 274518
rect 310336 271244 310388 271250
rect 310336 271186 310388 271192
rect 309784 267232 309836 267238
rect 309784 267174 309836 267180
rect 309876 266484 309928 266490
rect 309876 266426 309928 266432
rect 308956 266416 309008 266422
rect 308956 266358 309008 266364
rect 309416 266416 309468 266422
rect 309416 266358 309468 266364
rect 308876 264302 309074 264330
rect 309428 264316 309456 266358
rect 309888 264316 309916 266426
rect 310348 266422 310376 271186
rect 310428 268796 310480 268802
rect 310428 268738 310480 268744
rect 310336 266416 310388 266422
rect 310336 266358 310388 266364
rect 310440 264330 310468 268738
rect 310532 268598 310560 277780
rect 311728 274446 311756 277780
rect 311716 274440 311768 274446
rect 311716 274382 311768 274388
rect 311164 273760 311216 273766
rect 311164 273702 311216 273708
rect 310520 268592 310572 268598
rect 310520 268534 310572 268540
rect 311176 267510 311204 273702
rect 312924 272678 312952 277780
rect 313096 273080 313148 273086
rect 313096 273022 313148 273028
rect 312912 272672 312964 272678
rect 312912 272614 312964 272620
rect 311808 271176 311860 271182
rect 311808 271118 311860 271124
rect 311716 267708 311768 267714
rect 311716 267650 311768 267656
rect 311164 267504 311216 267510
rect 311164 267446 311216 267452
rect 311256 267504 311308 267510
rect 311256 267446 311308 267452
rect 310796 266416 310848 266422
rect 310796 266358 310848 266364
rect 310362 264302 310468 264330
rect 310808 264316 310836 266358
rect 311268 264316 311296 267446
rect 311728 264316 311756 267650
rect 311820 266422 311848 271118
rect 312452 271108 312504 271114
rect 312452 271050 312504 271056
rect 312464 267034 312492 271050
rect 313004 268728 313056 268734
rect 313004 268670 313056 268676
rect 312452 267028 312504 267034
rect 312452 266970 312504 266976
rect 312544 266756 312596 266762
rect 312544 266698 312596 266704
rect 311808 266416 311860 266422
rect 311808 266358 311860 266364
rect 312084 266416 312136 266422
rect 312084 266358 312136 266364
rect 312096 264316 312124 266358
rect 312556 264316 312584 266698
rect 313016 264316 313044 268670
rect 313108 266422 313136 273022
rect 314120 272610 314148 277780
rect 315316 273834 315344 277780
rect 315304 273828 315356 273834
rect 315304 273770 315356 273776
rect 315396 273828 315448 273834
rect 315396 273770 315448 273776
rect 314476 273012 314528 273018
rect 314476 272954 314528 272960
rect 314108 272604 314160 272610
rect 314108 272546 314160 272552
rect 314292 269952 314344 269958
rect 314292 269894 314344 269900
rect 313924 267232 313976 267238
rect 313924 267174 313976 267180
rect 313096 266416 313148 266422
rect 313096 266358 313148 266364
rect 313464 266416 313516 266422
rect 313464 266358 313516 266364
rect 313476 264316 313504 266358
rect 313936 264316 313964 267174
rect 314304 266490 314332 269894
rect 314384 268660 314436 268666
rect 314384 268602 314436 268608
rect 314292 266484 314344 266490
rect 314292 266426 314344 266432
rect 314396 264316 314424 268602
rect 314488 266422 314516 272954
rect 315212 267164 315264 267170
rect 315212 267106 315264 267112
rect 314476 266416 314528 266422
rect 314476 266358 314528 266364
rect 314844 266416 314896 266422
rect 314844 266358 314896 266364
rect 314856 264316 314884 266358
rect 315224 264316 315252 267106
rect 315408 267102 315436 273770
rect 315856 272944 315908 272950
rect 315856 272886 315908 272892
rect 315672 268592 315724 268598
rect 315672 268534 315724 268540
rect 315396 267096 315448 267102
rect 315396 267038 315448 267044
rect 315684 264316 315712 268534
rect 315868 266422 315896 272886
rect 316512 272542 316540 277780
rect 317236 272876 317288 272882
rect 317236 272818 317288 272824
rect 316500 272536 316552 272542
rect 316500 272478 316552 272484
rect 317052 268524 317104 268530
rect 317052 268466 317104 268472
rect 316040 267504 316092 267510
rect 316092 267452 316172 267458
rect 316040 267446 316172 267452
rect 316052 267430 316172 267446
rect 316144 267238 316172 267430
rect 316040 267232 316092 267238
rect 316040 267174 316092 267180
rect 316132 267232 316184 267238
rect 316132 267174 316184 267180
rect 316052 267102 316080 267174
rect 316040 267096 316092 267102
rect 316040 267038 316092 267044
rect 316592 267028 316644 267034
rect 316592 266970 316644 266976
rect 315856 266416 315908 266422
rect 315856 266358 315908 266364
rect 316132 266416 316184 266422
rect 316132 266358 316184 266364
rect 316144 264316 316172 266358
rect 316604 264316 316632 266970
rect 317064 264316 317092 268466
rect 317248 266422 317276 272818
rect 317708 272474 317736 277780
rect 317788 274440 317840 274446
rect 317788 274382 317840 274388
rect 317696 272468 317748 272474
rect 317696 272410 317748 272416
rect 317800 267306 317828 274382
rect 318812 274310 318840 277780
rect 320008 274650 320036 277780
rect 319996 274644 320048 274650
rect 319996 274586 320048 274592
rect 320088 274644 320140 274650
rect 320088 274586 320140 274592
rect 318800 274304 318852 274310
rect 318800 274246 318852 274252
rect 319444 274304 319496 274310
rect 319444 274246 319496 274252
rect 318616 272808 318668 272814
rect 318616 272750 318668 272756
rect 318340 268388 318392 268394
rect 318340 268330 318392 268336
rect 317788 267300 317840 267306
rect 317788 267242 317840 267248
rect 317880 267300 317932 267306
rect 317880 267242 317932 267248
rect 317236 266416 317288 266422
rect 317236 266358 317288 266364
rect 317512 266416 317564 266422
rect 317512 266358 317564 266364
rect 317524 264316 317552 266358
rect 317892 264316 317920 267242
rect 318352 264316 318380 268330
rect 318628 266422 318656 272750
rect 319260 269816 319312 269822
rect 319260 269758 319312 269764
rect 318616 266416 318668 266422
rect 318616 266358 318668 266364
rect 318800 266416 318852 266422
rect 318800 266358 318852 266364
rect 318812 264316 318840 266358
rect 319272 264316 319300 269758
rect 319456 267646 319484 274246
rect 320100 273290 320128 274586
rect 321204 274514 321232 277780
rect 321192 274508 321244 274514
rect 321192 274450 321244 274456
rect 322400 274106 322428 277780
rect 322388 274100 322440 274106
rect 322388 274042 322440 274048
rect 323596 273766 323624 277780
rect 324044 276276 324096 276282
rect 324044 276218 324096 276224
rect 323676 274100 323728 274106
rect 323676 274042 323728 274048
rect 323584 273760 323636 273766
rect 323584 273702 323636 273708
rect 322204 273420 322256 273426
rect 322204 273362 322256 273368
rect 319536 273284 319588 273290
rect 319536 273226 319588 273232
rect 320088 273284 320140 273290
rect 320088 273226 320140 273232
rect 319444 267640 319496 267646
rect 319444 267582 319496 267588
rect 319548 267578 319576 273226
rect 321284 272740 321336 272746
rect 321284 272682 321336 272688
rect 319904 272672 319956 272678
rect 319904 272614 319956 272620
rect 319720 268456 319772 268462
rect 319720 268398 319772 268404
rect 319536 267572 319588 267578
rect 319536 267514 319588 267520
rect 319732 264316 319760 268398
rect 319916 266422 319944 272614
rect 321192 272536 321244 272542
rect 321192 272478 321244 272484
rect 321008 268864 321060 268870
rect 321008 268806 321060 268812
rect 320180 266484 320232 266490
rect 320180 266426 320232 266432
rect 319904 266416 319956 266422
rect 319904 266358 319956 266364
rect 320192 264316 320220 266426
rect 320548 266416 320600 266422
rect 320548 266358 320600 266364
rect 320560 264316 320588 266358
rect 321020 264316 321048 268806
rect 321204 264330 321232 272478
rect 321296 266422 321324 272682
rect 321376 272604 321428 272610
rect 321376 272546 321428 272552
rect 321388 266490 321416 272546
rect 322216 266966 322244 273362
rect 322664 272264 322716 272270
rect 322664 272206 322716 272212
rect 322388 267980 322440 267986
rect 322388 267922 322440 267928
rect 322204 266960 322256 266966
rect 322204 266902 322256 266908
rect 321376 266484 321428 266490
rect 321376 266426 321428 266432
rect 321284 266416 321336 266422
rect 321284 266358 321336 266364
rect 321928 266416 321980 266422
rect 321928 266358 321980 266364
rect 321204 264302 321494 264330
rect 321940 264316 321968 266358
rect 322400 264316 322428 267922
rect 322676 264330 322704 272206
rect 322756 272128 322808 272134
rect 322756 272070 322808 272076
rect 322768 266422 322796 272070
rect 323688 266898 323716 274042
rect 323676 266892 323728 266898
rect 323676 266834 323728 266840
rect 323216 266552 323268 266558
rect 323216 266494 323268 266500
rect 322756 266416 322808 266422
rect 322756 266358 322808 266364
rect 322676 264302 322874 264330
rect 323228 264316 323256 266494
rect 324056 264330 324084 276218
rect 324792 273970 324820 277780
rect 324780 273964 324832 273970
rect 324780 273906 324832 273912
rect 325988 273902 326016 277780
rect 326712 276344 326764 276350
rect 326712 276286 326764 276292
rect 326344 273964 326396 273970
rect 326344 273906 326396 273912
rect 325976 273896 326028 273902
rect 325976 273838 326028 273844
rect 325608 272196 325660 272202
rect 325608 272138 325660 272144
rect 324136 267640 324188 267646
rect 324136 267582 324188 267588
rect 323702 264302 324084 264330
rect 324148 264316 324176 267582
rect 324596 266960 324648 266966
rect 324596 266902 324648 266908
rect 324608 264316 324636 266902
rect 325056 265192 325108 265198
rect 325056 265134 325108 265140
rect 325068 264316 325096 265134
rect 325620 264330 325648 272138
rect 326356 266694 326384 273906
rect 326344 266688 326396 266694
rect 326344 266630 326396 266636
rect 325976 266620 326028 266626
rect 325976 266562 326028 266568
rect 325542 264302 325648 264330
rect 325988 264316 326016 266562
rect 326724 264330 326752 276286
rect 327092 269550 327120 277780
rect 328288 273834 328316 277780
rect 329484 274378 329512 277780
rect 329852 277766 330694 277794
rect 331232 277766 331890 277794
rect 329748 276412 329800 276418
rect 329748 276354 329800 276360
rect 329656 275052 329708 275058
rect 329656 274994 329708 275000
rect 329472 274372 329524 274378
rect 329472 274314 329524 274320
rect 328276 273828 328328 273834
rect 328276 273770 328328 273776
rect 327724 273556 327776 273562
rect 327724 273498 327776 273504
rect 327080 269544 327132 269550
rect 327080 269486 327132 269492
rect 326804 267572 326856 267578
rect 326804 267514 326856 267520
rect 326370 264302 326752 264330
rect 326816 264316 326844 267514
rect 327736 266966 327764 273498
rect 327816 270972 327868 270978
rect 327816 270914 327868 270920
rect 327828 267442 327856 270914
rect 329564 270700 329616 270706
rect 329564 270642 329616 270648
rect 327816 267436 327868 267442
rect 327816 267378 327868 267384
rect 327724 266960 327776 266966
rect 327724 266902 327776 266908
rect 328184 266960 328236 266966
rect 328184 266902 328236 266908
rect 327264 266416 327316 266422
rect 327264 266358 327316 266364
rect 327276 264316 327304 266358
rect 327724 265260 327776 265266
rect 327724 265202 327776 265208
rect 327736 264316 327764 265202
rect 328196 264316 328224 266902
rect 328644 266484 328696 266490
rect 328644 266426 328696 266432
rect 328656 264316 328684 266426
rect 329012 266416 329064 266422
rect 329012 266358 329064 266364
rect 329024 264316 329052 266358
rect 329576 264330 329604 270642
rect 329668 266490 329696 274994
rect 329656 266484 329708 266490
rect 329656 266426 329708 266432
rect 329760 266422 329788 276354
rect 329852 269618 329880 277766
rect 331232 269686 331260 277766
rect 332416 276480 332468 276486
rect 332416 276422 332468 276428
rect 332324 270632 332376 270638
rect 332324 270574 332376 270580
rect 331220 269680 331272 269686
rect 331220 269622 331272 269628
rect 329840 269612 329892 269618
rect 329840 269554 329892 269560
rect 331128 268116 331180 268122
rect 331128 268058 331180 268064
rect 329932 266688 329984 266694
rect 329932 266630 329984 266636
rect 329748 266416 329800 266422
rect 329748 266358 329800 266364
rect 329498 264302 329604 264330
rect 329944 264316 329972 266630
rect 331140 266626 331168 268058
rect 331128 266620 331180 266626
rect 331128 266562 331180 266568
rect 332336 266422 332364 270574
rect 331312 266416 331364 266422
rect 331312 266358 331364 266364
rect 332324 266416 332376 266422
rect 332324 266358 332376 266364
rect 330852 265396 330904 265402
rect 330852 265338 330904 265344
rect 330392 265328 330444 265334
rect 330392 265270 330444 265276
rect 330404 264316 330432 265270
rect 330864 264316 330892 265338
rect 331324 264316 331352 266358
rect 332428 264602 332456 276422
rect 332060 264574 332456 264602
rect 332060 264330 332088 264574
rect 332520 264330 332548 277918
rect 333888 277908 333940 277914
rect 436664 277902 437046 277918
rect 440344 277914 440634 277930
rect 440332 277908 440634 277914
rect 333888 277850 333940 277856
rect 440384 277902 440634 277908
rect 440332 277850 440384 277856
rect 333072 274582 333100 277780
rect 333060 274576 333112 274582
rect 333060 274518 333112 274524
rect 333244 271040 333296 271046
rect 333244 270982 333296 270988
rect 333256 267374 333284 270982
rect 333244 267368 333296 267374
rect 333244 267310 333296 267316
rect 332600 266688 332652 266694
rect 332600 266630 332652 266636
rect 331706 264302 332088 264330
rect 332166 264302 332548 264330
rect 332612 264316 332640 266630
rect 333060 265464 333112 265470
rect 333060 265406 333112 265412
rect 333072 264316 333100 265406
rect 333900 264330 333928 277850
rect 335084 277840 335136 277846
rect 333992 277766 334190 277794
rect 443828 277840 443880 277846
rect 335084 277782 335136 277788
rect 333992 270094 334020 277766
rect 333980 270088 334032 270094
rect 333980 270030 334032 270036
rect 334348 269340 334400 269346
rect 334348 269282 334400 269288
rect 333980 266416 334032 266422
rect 333980 266358 334032 266364
rect 333546 264302 333928 264330
rect 333992 264316 334020 266358
rect 334360 264316 334388 269282
rect 335096 264330 335124 277782
rect 335176 275120 335228 275126
rect 335176 275062 335228 275068
rect 335188 266422 335216 275062
rect 335372 274242 335400 277780
rect 336372 277772 336424 277778
rect 336372 277714 336424 277720
rect 335360 274236 335412 274242
rect 335360 274178 335412 274184
rect 335728 269408 335780 269414
rect 335728 269350 335780 269356
rect 335268 266756 335320 266762
rect 335268 266698 335320 266704
rect 335176 266416 335228 266422
rect 335176 266358 335228 266364
rect 334834 264302 335124 264330
rect 335280 264316 335308 266698
rect 335740 264316 335768 269350
rect 336384 264330 336412 277714
rect 336568 271862 336596 277780
rect 336752 277766 337778 277794
rect 336648 275392 336700 275398
rect 336648 275334 336700 275340
rect 336556 271856 336608 271862
rect 336556 271798 336608 271804
rect 336214 264302 336412 264330
rect 336660 264316 336688 275334
rect 336752 269890 336780 277766
rect 338028 277704 338080 277710
rect 338028 277646 338080 277652
rect 336740 269884 336792 269890
rect 336740 269826 336792 269832
rect 337108 269884 337160 269890
rect 337108 269826 337160 269832
rect 337120 264316 337148 269826
rect 337476 264580 337528 264586
rect 337476 264522 337528 264528
rect 337488 264316 337516 264522
rect 338040 264330 338068 277646
rect 338960 274650 338988 277780
rect 339224 277636 339276 277642
rect 339224 277578 339276 277584
rect 338948 274644 339000 274650
rect 338948 274586 339000 274592
rect 338396 269476 338448 269482
rect 338396 269418 338448 269424
rect 337962 264302 338068 264330
rect 338408 264316 338436 269418
rect 339236 264330 339264 277578
rect 340156 271794 340184 277780
rect 340892 277766 341366 277794
rect 342272 277766 342470 277794
rect 340604 275460 340656 275466
rect 340604 275402 340656 275408
rect 340144 271788 340196 271794
rect 340144 271730 340196 271736
rect 339776 270088 339828 270094
rect 339776 270030 339828 270036
rect 339408 268252 339460 268258
rect 339408 268194 339460 268200
rect 339420 267510 339448 268194
rect 339408 267504 339460 267510
rect 339408 267446 339460 267452
rect 339316 266824 339368 266830
rect 339316 266766 339368 266772
rect 338882 264302 339264 264330
rect 339328 264316 339356 266766
rect 339788 264316 339816 270030
rect 340144 266416 340196 266422
rect 340144 266358 340196 266364
rect 340156 264316 340184 266358
rect 340616 264316 340644 275402
rect 340696 273488 340748 273494
rect 340696 273430 340748 273436
rect 340708 266422 340736 273430
rect 340892 269754 340920 277766
rect 341892 273624 341944 273630
rect 341892 273566 341944 273572
rect 340880 269748 340932 269754
rect 340880 269690 340932 269696
rect 341064 269544 341116 269550
rect 341064 269486 341116 269492
rect 340696 266416 340748 266422
rect 340696 266358 340748 266364
rect 341076 264316 341104 269486
rect 341904 264330 341932 273566
rect 342272 270502 342300 277766
rect 343364 275188 343416 275194
rect 343364 275130 343416 275136
rect 342260 270496 342312 270502
rect 342260 270438 342312 270444
rect 342444 269612 342496 269618
rect 342444 269554 342496 269560
rect 341984 266892 342036 266898
rect 341984 266834 342036 266840
rect 341550 264302 341932 264330
rect 341996 264316 342024 266834
rect 342456 264316 342484 269554
rect 342812 266416 342864 266422
rect 342812 266358 342864 266364
rect 342824 264316 342852 266358
rect 343376 264330 343404 275130
rect 343456 273692 343508 273698
rect 343456 273634 343508 273640
rect 343468 266422 343496 273634
rect 343652 271114 343680 277780
rect 343836 277766 344862 277794
rect 343640 271108 343692 271114
rect 343640 271050 343692 271056
rect 343836 270434 343864 277766
rect 346044 274174 346072 277780
rect 346124 275256 346176 275262
rect 346124 275198 346176 275204
rect 346032 274168 346084 274174
rect 346032 274110 346084 274116
rect 344560 273760 344612 273766
rect 344560 273702 344612 273708
rect 343824 270428 343876 270434
rect 343824 270370 343876 270376
rect 343732 269680 343784 269686
rect 343732 269622 343784 269628
rect 343640 267912 343692 267918
rect 343640 267854 343692 267860
rect 343652 266966 343680 267854
rect 343640 266960 343692 266966
rect 343640 266902 343692 266908
rect 343456 266416 343508 266422
rect 343456 266358 343508 266364
rect 343298 264302 343404 264330
rect 343744 264316 343772 269622
rect 344572 264330 344600 273702
rect 345112 269748 345164 269754
rect 345112 269690 345164 269696
rect 344652 267708 344704 267714
rect 344652 267650 344704 267656
rect 344218 264302 344600 264330
rect 344664 264316 344692 267650
rect 345124 264316 345152 269690
rect 345480 266416 345532 266422
rect 345480 266358 345532 266364
rect 345492 264316 345520 266358
rect 346136 264330 346164 275198
rect 346216 273828 346268 273834
rect 346216 273770 346268 273776
rect 346228 266422 346256 273770
rect 347044 271992 347096 271998
rect 347044 271934 347096 271940
rect 346400 270496 346452 270502
rect 346400 270438 346452 270444
rect 346216 266416 346268 266422
rect 346216 266358 346268 266364
rect 345966 264302 346164 264330
rect 346412 264316 346440 270438
rect 347056 267646 347084 271934
rect 347240 270978 347268 277780
rect 347792 277766 348450 277794
rect 347688 273896 347740 273902
rect 347688 273838 347740 273844
rect 347228 270972 347280 270978
rect 347228 270914 347280 270920
rect 347044 267640 347096 267646
rect 347044 267582 347096 267588
rect 347320 266960 347372 266966
rect 347320 266902 347372 266908
rect 346860 266416 346912 266422
rect 346860 266358 346912 266364
rect 346872 264316 346900 266358
rect 347332 264316 347360 266902
rect 347700 266422 347728 273838
rect 347792 270366 347820 277766
rect 349068 276548 349120 276554
rect 349068 276490 349120 276496
rect 348976 276004 349028 276010
rect 348976 275946 349028 275952
rect 348516 274644 348568 274650
rect 348516 274586 348568 274592
rect 347780 270360 347832 270366
rect 347780 270302 347832 270308
rect 347688 266416 347740 266422
rect 347688 266358 347740 266364
rect 347780 266416 347832 266422
rect 347780 266358 347832 266364
rect 347792 264316 347820 266358
rect 348528 264330 348556 274586
rect 348988 264330 349016 275946
rect 349080 266422 349108 276490
rect 349632 274446 349660 277780
rect 350448 276616 350500 276622
rect 350448 276558 350500 276564
rect 350356 274576 350408 274582
rect 350356 274518 350408 274524
rect 349620 274440 349672 274446
rect 349620 274382 349672 274388
rect 349804 272060 349856 272066
rect 349804 272002 349856 272008
rect 349816 267578 349844 272002
rect 349988 267640 350040 267646
rect 349988 267582 350040 267588
rect 349804 267572 349856 267578
rect 349804 267514 349856 267520
rect 349068 266416 349120 266422
rect 349068 266358 349120 266364
rect 349528 266416 349580 266422
rect 349528 266358 349580 266364
rect 349068 265532 349120 265538
rect 349068 265474 349120 265480
rect 348266 264302 348556 264330
rect 348634 264302 349016 264330
rect 349080 264316 349108 265474
rect 349540 264316 349568 266358
rect 350000 264316 350028 267582
rect 350368 266422 350396 274518
rect 350356 266416 350408 266422
rect 350356 266358 350408 266364
rect 350460 264316 350488 276558
rect 350736 271726 350764 277780
rect 351828 275936 351880 275942
rect 351828 275878 351880 275884
rect 351736 274508 351788 274514
rect 351736 274450 351788 274456
rect 350724 271720 350776 271726
rect 350724 271662 350776 271668
rect 351748 266422 351776 274450
rect 350908 266416 350960 266422
rect 350908 266358 350960 266364
rect 351736 266416 351788 266422
rect 351736 266358 351788 266364
rect 350920 264316 350948 266358
rect 351840 265690 351868 275878
rect 351932 270298 351960 277780
rect 353024 274440 353076 274446
rect 353024 274382 353076 274388
rect 351920 270292 351972 270298
rect 351920 270234 351972 270240
rect 352656 267572 352708 267578
rect 352656 267514 352708 267520
rect 352196 266416 352248 266422
rect 352196 266358 352248 266364
rect 351656 265662 351868 265690
rect 351656 264330 351684 265662
rect 351736 265600 351788 265606
rect 351736 265542 351788 265548
rect 351302 264302 351684 264330
rect 351748 264316 351776 265542
rect 352208 264316 352236 266358
rect 352668 264316 352696 267514
rect 353036 266422 353064 274382
rect 353128 274310 353156 277780
rect 353208 277364 353260 277370
rect 353208 277306 353260 277312
rect 353116 274304 353168 274310
rect 353116 274246 353168 274252
rect 353024 266416 353076 266422
rect 353024 266358 353076 266364
rect 353220 264330 353248 277306
rect 354324 271046 354352 277780
rect 354692 277766 355534 277794
rect 356072 277766 356730 277794
rect 354404 275868 354456 275874
rect 354404 275810 354456 275816
rect 354312 271040 354364 271046
rect 354312 270982 354364 270988
rect 353300 269272 353352 269278
rect 353300 269214 353352 269220
rect 353312 267238 353340 269214
rect 354416 267734 354444 275810
rect 354692 270230 354720 277766
rect 355968 277296 356020 277302
rect 355968 277238 356020 277244
rect 354864 270428 354916 270434
rect 354864 270370 354916 270376
rect 354680 270224 354732 270230
rect 354680 270166 354732 270172
rect 354324 267706 354444 267734
rect 353300 267232 353352 267238
rect 353300 267174 353352 267180
rect 353852 264512 353904 264518
rect 353852 264454 353904 264460
rect 353864 264330 353892 264454
rect 354324 264330 354352 267706
rect 354404 266348 354456 266354
rect 354404 266290 354456 266296
rect 353142 264302 353248 264330
rect 353602 264302 353892 264330
rect 353970 264302 354352 264330
rect 354416 264316 354444 266290
rect 354876 264316 354904 270370
rect 355324 267504 355376 267510
rect 355324 267446 355376 267452
rect 355336 264316 355364 267446
rect 355980 264330 356008 277238
rect 356072 270162 356100 277766
rect 357348 275800 357400 275806
rect 357348 275742 357400 275748
rect 357256 274372 357308 274378
rect 357256 274314 357308 274320
rect 356060 270156 356112 270162
rect 356060 270098 356112 270104
rect 357268 267170 357296 274314
rect 356244 267164 356296 267170
rect 356244 267106 356296 267112
rect 357256 267164 357308 267170
rect 357256 267106 357308 267112
rect 355810 264302 356008 264330
rect 356256 264316 356284 267106
rect 357360 266422 357388 275742
rect 357912 273222 357940 277780
rect 358728 277228 358780 277234
rect 358728 277170 358780 277176
rect 357900 273216 357952 273222
rect 357900 273158 357952 273164
rect 358636 272468 358688 272474
rect 358636 272410 358688 272416
rect 357992 267436 358044 267442
rect 357992 267378 358044 267384
rect 356612 266416 356664 266422
rect 356612 266358 356664 266364
rect 357348 266416 357400 266422
rect 357348 266358 357400 266364
rect 357532 266416 357584 266422
rect 357532 266358 357584 266364
rect 356624 264316 356652 266358
rect 357072 266280 357124 266286
rect 357072 266222 357124 266228
rect 357084 264316 357112 266222
rect 357544 264316 357572 266358
rect 358004 264316 358032 267378
rect 358648 266422 358676 272410
rect 358636 266416 358688 266422
rect 358636 266358 358688 266364
rect 358740 264330 358768 277170
rect 359016 271658 359044 277780
rect 360108 277568 360160 277574
rect 360108 277510 360160 277516
rect 360016 271720 360068 271726
rect 360016 271662 360068 271668
rect 359004 271652 359056 271658
rect 359004 271594 359056 271600
rect 359924 270768 359976 270774
rect 359924 270710 359976 270716
rect 358912 267164 358964 267170
rect 358912 267106 358964 267112
rect 358478 264302 358768 264330
rect 358924 264316 358952 267106
rect 359372 266416 359424 266422
rect 359372 266358 359424 266364
rect 359384 264316 359412 266358
rect 359936 264330 359964 270710
rect 360028 266422 360056 271662
rect 360120 267170 360148 277510
rect 360212 274038 360240 277780
rect 360396 277766 361422 277794
rect 362328 277766 362618 277794
rect 362972 277766 363814 277794
rect 360200 274032 360252 274038
rect 360200 273974 360252 273980
rect 360200 270360 360252 270366
rect 360200 270302 360252 270308
rect 360108 267164 360160 267170
rect 360108 267106 360160 267112
rect 360016 266416 360068 266422
rect 360016 266358 360068 266364
rect 359766 264302 359964 264330
rect 360212 264316 360240 270302
rect 360396 269074 360424 277766
rect 362224 275732 362276 275738
rect 362224 275674 362276 275680
rect 360844 271924 360896 271930
rect 360844 271866 360896 271872
rect 360384 269068 360436 269074
rect 360384 269010 360436 269016
rect 360660 267368 360712 267374
rect 360660 267310 360712 267316
rect 360672 264316 360700 267310
rect 360856 267306 360884 271866
rect 362236 271726 362264 275674
rect 362224 271720 362276 271726
rect 362224 271662 362276 271668
rect 362328 271590 362356 277766
rect 362592 274304 362644 274310
rect 362592 274246 362644 274252
rect 362316 271584 362368 271590
rect 362316 271526 362368 271532
rect 361488 270836 361540 270842
rect 361488 270778 361540 270784
rect 360844 267300 360896 267306
rect 360844 267242 360896 267248
rect 361500 264330 361528 270778
rect 361580 269068 361632 269074
rect 361580 269010 361632 269016
rect 361146 264302 361528 264330
rect 361592 264316 361620 269010
rect 362040 267164 362092 267170
rect 362040 267106 362092 267112
rect 362052 264316 362080 267106
rect 362408 266416 362460 266422
rect 362408 266358 362460 266364
rect 362420 264316 362448 266358
rect 362604 264330 362632 274246
rect 362684 271584 362736 271590
rect 362684 271526 362736 271532
rect 362696 267170 362724 271526
rect 362776 270904 362828 270910
rect 362776 270846 362828 270852
rect 362684 267164 362736 267170
rect 362684 267106 362736 267112
rect 362788 266422 362816 270846
rect 362972 270026 363000 277766
rect 363512 275664 363564 275670
rect 363512 275606 363564 275612
rect 363524 271590 363552 275606
rect 364996 273154 365024 277780
rect 365628 274236 365680 274242
rect 365628 274178 365680 274184
rect 364984 273148 365036 273154
rect 364984 273090 365036 273096
rect 363604 272400 363656 272406
rect 363604 272342 363656 272348
rect 363512 271584 363564 271590
rect 363512 271526 363564 271532
rect 362960 270020 363012 270026
rect 362960 269962 363012 269968
rect 363328 267300 363380 267306
rect 363328 267242 363380 267248
rect 362776 266416 362828 266422
rect 362776 266358 362828 266364
rect 362604 264302 362894 264330
rect 363340 264316 363368 267242
rect 363616 267238 363644 272342
rect 365536 271652 365588 271658
rect 365536 271594 365588 271600
rect 365444 271040 365496 271046
rect 365444 270982 365496 270988
rect 364156 270972 364208 270978
rect 364156 270914 364208 270920
rect 363604 267232 363656 267238
rect 363604 267174 363656 267180
rect 364168 264330 364196 270914
rect 364248 270292 364300 270298
rect 364248 270234 364300 270240
rect 363814 264302 364196 264330
rect 364260 264316 364288 270234
rect 364708 266416 364760 266422
rect 364708 266358 364760 266364
rect 364720 264316 364748 266358
rect 365456 264330 365484 270982
rect 365548 266422 365576 271594
rect 365536 266416 365588 266422
rect 365536 266358 365588 266364
rect 365640 264330 365668 274178
rect 366100 271522 366128 277780
rect 367008 275596 367060 275602
rect 367008 275538 367060 275544
rect 366916 271856 366968 271862
rect 366916 271798 366968 271804
rect 366088 271516 366140 271522
rect 366088 271458 366140 271464
rect 365720 267776 365772 267782
rect 365720 267718 365772 267724
rect 365732 267238 365760 267718
rect 365720 267232 365772 267238
rect 365720 267174 365772 267180
rect 365996 267232 366048 267238
rect 365996 267174 366048 267180
rect 365102 264302 365484 264330
rect 365562 264302 365668 264330
rect 366008 264316 366036 267174
rect 366456 266416 366508 266422
rect 366456 266358 366508 266364
rect 366468 264316 366496 266358
rect 366928 264316 366956 271798
rect 367020 271658 367048 275538
rect 367296 273426 367324 277780
rect 368388 275528 368440 275534
rect 368388 275470 368440 275476
rect 367284 273420 367336 273426
rect 367284 273362 367336 273368
rect 368296 273216 368348 273222
rect 368296 273158 368348 273164
rect 368112 271788 368164 271794
rect 368112 271730 368164 271736
rect 367008 271652 367060 271658
rect 367008 271594 367060 271600
rect 367008 271108 367060 271114
rect 367008 271050 367060 271056
rect 367020 266422 367048 271050
rect 367008 266416 367060 266422
rect 367008 266358 367060 266364
rect 367376 266416 367428 266422
rect 367376 266358 367428 266364
rect 367388 264316 367416 266358
rect 368124 264330 368152 271730
rect 368308 264330 368336 273158
rect 368400 266422 368428 275470
rect 368492 268938 368520 277780
rect 369492 271720 369544 271726
rect 369492 271662 369544 271668
rect 368480 268932 368532 268938
rect 368480 268874 368532 268880
rect 368664 267164 368716 267170
rect 368664 267106 368716 267112
rect 368388 266416 368440 266422
rect 368388 266358 368440 266364
rect 367770 264302 368152 264330
rect 368230 264302 368336 264330
rect 368676 264316 368704 267106
rect 369504 264330 369532 271662
rect 369688 271454 369716 277780
rect 370780 271652 370832 271658
rect 370780 271594 370832 271600
rect 369676 271448 369728 271454
rect 369676 271390 369728 271396
rect 369584 270224 369636 270230
rect 369584 270166 369636 270172
rect 369150 264302 369532 264330
rect 369596 264316 369624 270166
rect 370044 266416 370096 266422
rect 370044 266358 370096 266364
rect 370056 264316 370084 266358
rect 370792 264330 370820 271594
rect 370884 271386 370912 277780
rect 371344 277766 372094 277794
rect 371238 275360 371294 275369
rect 371238 275295 371294 275304
rect 371252 271538 371280 275295
rect 371068 271510 371280 271538
rect 370872 271380 370924 271386
rect 370872 271322 370924 271328
rect 370872 268932 370924 268938
rect 370872 268874 370924 268880
rect 370530 264302 370820 264330
rect 370884 264316 370912 268874
rect 371068 266422 371096 271510
rect 371344 268326 371372 277766
rect 372528 274168 372580 274174
rect 372528 274110 372580 274116
rect 372160 271584 372212 271590
rect 372160 271526 372212 271532
rect 371332 268320 371384 268326
rect 371332 268262 371384 268268
rect 371884 267844 371936 267850
rect 371884 267786 371936 267792
rect 371332 267096 371384 267102
rect 371332 267038 371384 267044
rect 371056 266416 371108 266422
rect 371056 266358 371108 266364
rect 371344 264316 371372 267038
rect 371896 267034 371924 267786
rect 371884 267028 371936 267034
rect 371884 266970 371936 266976
rect 372172 264330 372200 271526
rect 372540 264330 372568 274110
rect 373276 271318 373304 277780
rect 374380 274106 374408 277780
rect 375392 277766 375590 277794
rect 375196 274984 375248 274990
rect 375196 274926 375248 274932
rect 374368 274100 374420 274106
rect 374368 274042 374420 274048
rect 373816 271516 373868 271522
rect 373816 271458 373868 271464
rect 373264 271312 373316 271318
rect 373264 271254 373316 271260
rect 372712 268320 372764 268326
rect 372712 268262 372764 268268
rect 371818 264302 372200 264330
rect 372278 264302 372568 264330
rect 372724 264316 372752 268262
rect 373172 266212 373224 266218
rect 373172 266154 373224 266160
rect 373184 264316 373212 266154
rect 373828 264330 373856 271458
rect 375208 270638 375236 274926
rect 375288 271448 375340 271454
rect 375288 271390 375340 271396
rect 375196 270632 375248 270638
rect 375196 270574 375248 270580
rect 374000 270156 374052 270162
rect 374000 270098 374052 270104
rect 373566 264302 373856 264330
rect 374012 264316 374040 270098
rect 374460 266144 374512 266150
rect 374460 266086 374512 266092
rect 374472 264316 374500 266086
rect 375300 264330 375328 271390
rect 375392 269006 375420 277766
rect 376668 274100 376720 274106
rect 376668 274042 376720 274048
rect 376576 271380 376628 271386
rect 376576 271322 376628 271328
rect 376482 270056 376538 270065
rect 376482 269991 376538 270000
rect 375380 269000 375432 269006
rect 375380 268942 375432 268948
rect 375380 267028 375432 267034
rect 375380 266970 375432 266976
rect 374946 264302 375328 264330
rect 375392 264316 375420 266970
rect 376496 266422 376524 269991
rect 376484 266416 376536 266422
rect 376484 266358 376536 266364
rect 375840 266076 375892 266082
rect 375840 266018 375892 266024
rect 375852 264316 375880 266018
rect 376588 264330 376616 271322
rect 376680 267034 376708 274042
rect 376772 271250 376800 277780
rect 376956 277766 377982 277794
rect 378152 277766 379178 277794
rect 376760 271244 376812 271250
rect 376760 271186 376812 271192
rect 376956 269958 376984 277766
rect 378048 274032 378100 274038
rect 378048 273974 378100 273980
rect 377956 271312 378008 271318
rect 377956 271254 378008 271260
rect 376944 269952 376996 269958
rect 376944 269894 376996 269900
rect 376668 267028 376720 267034
rect 376668 266970 376720 266976
rect 376668 266416 376720 266422
rect 376668 266358 376720 266364
rect 376234 264302 376616 264330
rect 376680 264316 376708 266358
rect 377128 266008 377180 266014
rect 377128 265950 377180 265956
rect 377140 264316 377168 265950
rect 377968 264330 377996 271254
rect 377614 264302 377996 264330
rect 378060 264316 378088 273974
rect 378152 268802 378180 277766
rect 379334 271280 379390 271289
rect 379334 271215 379390 271224
rect 379428 271244 379480 271250
rect 378140 268796 378192 268802
rect 378140 268738 378192 268744
rect 378876 266416 378928 266422
rect 378876 266358 378928 266364
rect 378508 265940 378560 265946
rect 378508 265882 378560 265888
rect 378520 264316 378548 265882
rect 378888 264316 378916 266358
rect 379348 264316 379376 271215
rect 379428 271186 379480 271192
rect 379440 266422 379468 271186
rect 380360 271182 380388 277780
rect 380912 277766 381570 277794
rect 382292 277766 382674 277794
rect 380808 277160 380860 277166
rect 380808 277102 380860 277108
rect 380348 271176 380400 271182
rect 380348 271118 380400 271124
rect 380716 269952 380768 269958
rect 380716 269894 380768 269900
rect 379428 266416 379480 266422
rect 379428 266358 379480 266364
rect 379796 266416 379848 266422
rect 379796 266358 379848 266364
rect 379808 264316 379836 266358
rect 380256 265872 380308 265878
rect 380256 265814 380308 265820
rect 380268 264316 380296 265814
rect 380728 264316 380756 269894
rect 380820 266422 380848 277102
rect 380912 269278 380940 277766
rect 382186 274136 382242 274145
rect 382186 274071 382242 274080
rect 381636 270020 381688 270026
rect 381636 269962 381688 269968
rect 380900 269272 380952 269278
rect 380900 269214 380952 269220
rect 380808 266416 380860 266422
rect 380808 266358 380860 266364
rect 381176 265804 381228 265810
rect 381176 265746 381228 265752
rect 381188 264316 381216 265746
rect 381648 264316 381676 269962
rect 382200 264330 382228 274071
rect 382292 268258 382320 277766
rect 383476 277092 383528 277098
rect 383476 277034 383528 277040
rect 383382 272776 383438 272785
rect 383382 272711 383438 272720
rect 382280 268252 382332 268258
rect 382280 268194 382332 268200
rect 382464 267028 382516 267034
rect 382464 266970 382516 266976
rect 382030 264302 382228 264330
rect 382476 264316 382504 266970
rect 382924 266416 382976 266422
rect 382924 266358 382976 266364
rect 382936 264316 382964 266358
rect 383396 264316 383424 272711
rect 383488 267034 383516 277034
rect 383568 277024 383620 277030
rect 383568 276966 383620 276972
rect 383476 267028 383528 267034
rect 383476 266970 383528 266976
rect 383580 266422 383608 276966
rect 383856 273086 383884 277780
rect 385052 273970 385080 277780
rect 385236 277766 386262 277794
rect 385040 273964 385092 273970
rect 385040 273906 385092 273912
rect 383844 273080 383896 273086
rect 383844 273022 383896 273028
rect 385236 268734 385264 277766
rect 387248 276956 387300 276962
rect 387248 276898 387300 276904
rect 385960 271176 386012 271182
rect 385960 271118 386012 271124
rect 385224 268728 385276 268734
rect 385224 268670 385276 268676
rect 385132 268048 385184 268054
rect 385132 267990 385184 267996
rect 383568 266416 383620 266422
rect 383568 266358 383620 266364
rect 384304 265736 384356 265742
rect 384304 265678 384356 265684
rect 383844 265668 383896 265674
rect 383844 265610 383896 265616
rect 383856 264316 383884 265610
rect 384316 264316 384344 265678
rect 384948 264444 385000 264450
rect 384948 264386 385000 264392
rect 384960 264330 384988 264386
rect 384698 264302 384988 264330
rect 385144 264316 385172 267990
rect 385972 264330 386000 271118
rect 386050 269920 386106 269929
rect 386050 269855 386106 269864
rect 385618 264302 386000 264330
rect 386064 264316 386092 269855
rect 386512 268184 386564 268190
rect 386512 268126 386564 268132
rect 386524 264316 386552 268126
rect 387260 264330 387288 276898
rect 387444 273018 387472 277780
rect 387812 277766 388654 277794
rect 389192 277766 389758 277794
rect 387432 273012 387484 273018
rect 387432 272954 387484 272960
rect 387812 267782 387840 277766
rect 388168 275324 388220 275330
rect 388168 275266 388220 275272
rect 388180 269822 388208 275266
rect 388168 269816 388220 269822
rect 388168 269758 388220 269764
rect 388720 269816 388772 269822
rect 388720 269758 388772 269764
rect 388168 268252 388220 268258
rect 388168 268194 388220 268200
rect 387800 267776 387852 267782
rect 387800 267718 387852 267724
rect 387616 264376 387668 264382
rect 386998 264302 387288 264330
rect 387366 264324 387616 264330
rect 388180 264330 388208 268194
rect 388258 265840 388314 265849
rect 388258 265775 388314 265784
rect 387366 264318 387668 264324
rect 387366 264302 387656 264318
rect 387826 264302 388208 264330
rect 388272 264316 388300 265775
rect 388732 264316 388760 269758
rect 389192 268666 389220 277766
rect 389916 276888 389968 276894
rect 389916 276830 389968 276836
rect 389180 268660 389232 268666
rect 389180 268602 389232 268608
rect 389178 267064 389234 267073
rect 389178 266999 389234 267008
rect 389192 264316 389220 266999
rect 389928 264330 389956 276830
rect 390376 273964 390428 273970
rect 390376 273906 390428 273912
rect 390388 264330 390416 273906
rect 390940 272950 390968 277780
rect 391664 277500 391716 277506
rect 391664 277442 391716 277448
rect 390928 272944 390980 272950
rect 390928 272886 390980 272892
rect 390468 267776 390520 267782
rect 390468 267718 390520 267724
rect 389666 264302 389956 264330
rect 390034 264302 390416 264330
rect 390480 264316 390508 267718
rect 390928 266416 390980 266422
rect 390928 266358 390980 266364
rect 390940 264316 390968 266358
rect 391676 264330 391704 277442
rect 391938 275496 391994 275505
rect 391938 275431 391994 275440
rect 391756 272332 391808 272338
rect 391756 272274 391808 272280
rect 391768 266422 391796 272274
rect 391848 269000 391900 269006
rect 391848 268942 391900 268948
rect 391756 266416 391808 266422
rect 391756 266358 391808 266364
rect 391414 264302 391704 264330
rect 391860 264316 391888 268942
rect 391952 268326 391980 275431
rect 392136 272406 392164 277780
rect 392124 272400 392176 272406
rect 392124 272342 392176 272348
rect 393136 272400 393188 272406
rect 393136 272342 393188 272348
rect 391940 268320 391992 268326
rect 391940 268262 391992 268268
rect 393148 266422 393176 272342
rect 393228 268796 393280 268802
rect 393228 268738 393280 268744
rect 392308 266416 392360 266422
rect 392308 266358 392360 266364
rect 393136 266416 393188 266422
rect 393136 266358 393188 266364
rect 392320 264316 392348 266358
rect 393240 264330 393268 268738
rect 393332 268598 393360 277780
rect 394424 273148 394476 273154
rect 394424 273090 394476 273096
rect 394056 268728 394108 268734
rect 394056 268670 394108 268676
rect 393320 268592 393372 268598
rect 393320 268534 393372 268540
rect 393596 266416 393648 266422
rect 393596 266358 393648 266364
rect 392794 264314 393084 264330
rect 392794 264308 393096 264314
rect 392794 264302 393044 264308
rect 393162 264302 393268 264330
rect 393608 264316 393636 266358
rect 394068 264316 394096 268670
rect 394436 266422 394464 273090
rect 394528 272882 394556 277780
rect 394712 277766 395738 277794
rect 396092 277766 396934 277794
rect 394516 272876 394568 272882
rect 394516 272818 394568 272824
rect 394516 268660 394568 268666
rect 394516 268602 394568 268608
rect 394424 266416 394476 266422
rect 394424 266358 394476 266364
rect 394528 264316 394556 268602
rect 394712 267850 394740 277766
rect 395710 271144 395766 271153
rect 395710 271079 395766 271088
rect 394974 269784 395030 269793
rect 394974 269719 395030 269728
rect 394700 267844 394752 267850
rect 394700 267786 394752 267792
rect 394988 264316 395016 269719
rect 395724 264330 395752 271079
rect 395804 268592 395856 268598
rect 395804 268534 395856 268540
rect 395462 264302 395752 264330
rect 395816 264316 395844 268534
rect 396092 268530 396120 277766
rect 397276 273080 397328 273086
rect 397276 273022 397328 273028
rect 396080 268524 396132 268530
rect 396080 268466 396132 268472
rect 397184 268524 397236 268530
rect 397184 268466 397236 268472
rect 396264 266416 396316 266422
rect 396264 266358 396316 266364
rect 396276 264316 396304 266358
rect 397196 264316 397224 268466
rect 397288 266422 397316 273022
rect 398024 272814 398052 277780
rect 398748 277432 398800 277438
rect 398748 277374 398800 277380
rect 398656 272944 398708 272950
rect 398656 272886 398708 272892
rect 398012 272808 398064 272814
rect 398012 272750 398064 272756
rect 398470 268696 398526 268705
rect 398470 268631 398526 268640
rect 397644 267028 397696 267034
rect 397644 266970 397696 266976
rect 397276 266416 397328 266422
rect 397276 266358 397328 266364
rect 397656 264316 397684 266970
rect 398104 266416 398156 266422
rect 398104 266358 398156 266364
rect 398116 264316 398144 266358
rect 398484 264316 398512 268631
rect 398668 267034 398696 272886
rect 398656 267028 398708 267034
rect 398656 266970 398708 266976
rect 398760 266422 398788 277374
rect 398840 274712 398892 274718
rect 398840 274654 398892 274660
rect 398852 268462 398880 274654
rect 398932 273012 398984 273018
rect 398932 272954 398984 272960
rect 398840 268456 398892 268462
rect 398840 268398 398892 268404
rect 398748 266416 398800 266422
rect 398748 266358 398800 266364
rect 398944 264316 398972 272954
rect 399220 271930 399248 277780
rect 400232 277766 400430 277794
rect 401626 277766 401732 277794
rect 399208 271924 399260 271930
rect 399208 271866 399260 271872
rect 399852 268456 399904 268462
rect 399852 268398 399904 268404
rect 399024 267028 399076 267034
rect 399024 266970 399076 266976
rect 399036 266558 399064 266970
rect 399024 266552 399076 266558
rect 399024 266494 399076 266500
rect 399864 264316 399892 268398
rect 400232 268394 400260 277766
rect 401600 274780 401652 274786
rect 401600 274722 401652 274728
rect 401046 274000 401102 274009
rect 401046 273935 401102 273944
rect 400312 272876 400364 272882
rect 400312 272818 400364 272824
rect 400220 268388 400272 268394
rect 400220 268330 400272 268336
rect 400324 264316 400352 272818
rect 401060 264330 401088 273935
rect 401612 272746 401640 274722
rect 401600 272740 401652 272746
rect 401600 272682 401652 272688
rect 401704 272678 401732 277766
rect 402808 275330 402836 277780
rect 403900 276820 403952 276826
rect 403900 276762 403952 276768
rect 402796 275324 402848 275330
rect 402796 275266 402848 275272
rect 401784 274916 401836 274922
rect 401784 274858 401836 274864
rect 401692 272672 401744 272678
rect 401692 272614 401744 272620
rect 401796 268870 401824 274858
rect 401968 272808 402020 272814
rect 401968 272750 402020 272756
rect 401784 268864 401836 268870
rect 401784 268806 401836 268812
rect 401140 268388 401192 268394
rect 401140 268330 401192 268336
rect 400798 264302 401088 264330
rect 401152 264316 401180 268330
rect 401980 264330 402008 272750
rect 402980 272740 403032 272746
rect 402980 272682 403032 272688
rect 402518 268424 402574 268433
rect 402518 268359 402574 268368
rect 402058 266520 402114 266529
rect 402058 266455 402114 266464
rect 401626 264302 402008 264330
rect 402072 264316 402100 266455
rect 402532 264316 402560 268359
rect 402992 264316 403020 272682
rect 403440 271924 403492 271930
rect 403440 271866 403492 271872
rect 403452 264316 403480 271866
rect 403912 264316 403940 276762
rect 404004 274718 404032 277780
rect 403992 274712 404044 274718
rect 403992 274654 404044 274660
rect 404268 274712 404320 274718
rect 404268 274654 404320 274660
rect 404174 272640 404230 272649
rect 404174 272575 404230 272584
rect 404188 264330 404216 272575
rect 404280 272134 404308 274654
rect 405200 272610 405228 277780
rect 406304 274786 406332 277780
rect 406660 276752 406712 276758
rect 406660 276694 406712 276700
rect 406292 274780 406344 274786
rect 406292 274722 406344 274728
rect 405648 272672 405700 272678
rect 405648 272614 405700 272620
rect 405188 272604 405240 272610
rect 405188 272546 405240 272552
rect 404268 272128 404320 272134
rect 404268 272070 404320 272076
rect 404360 272128 404412 272134
rect 404360 272070 404412 272076
rect 404372 271930 404400 272070
rect 404360 271924 404412 271930
rect 404360 271866 404412 271872
rect 404360 268864 404412 268870
rect 404360 268806 404412 268812
rect 404372 267073 404400 268806
rect 404358 267064 404414 267073
rect 404358 266999 404414 267008
rect 404726 266384 404782 266393
rect 404726 266319 404782 266328
rect 404188 264302 404294 264330
rect 404740 264316 404768 266319
rect 405186 265704 405242 265713
rect 405186 265639 405242 265648
rect 405200 264316 405228 265639
rect 405660 264316 405688 272614
rect 406106 271416 406162 271425
rect 406106 271351 406162 271360
rect 405738 268560 405794 268569
rect 405738 268495 405794 268504
rect 405752 266529 405780 268495
rect 405738 266520 405794 266529
rect 405738 266455 405794 266464
rect 406120 264316 406148 271351
rect 406672 264330 406700 276694
rect 407500 274922 407528 277780
rect 408512 277766 408710 277794
rect 407488 274916 407540 274922
rect 407488 274858 407540 274864
rect 407028 274848 407080 274854
rect 407028 274790 407080 274796
rect 406934 272504 406990 272513
rect 406934 272439 406990 272448
rect 406594 264302 406700 264330
rect 406948 264316 406976 272439
rect 407040 267986 407068 274790
rect 408512 274666 408540 277766
rect 409788 276684 409840 276690
rect 409788 276626 409840 276632
rect 409694 275224 409750 275233
rect 409694 275159 409750 275168
rect 408592 274780 408644 274786
rect 408592 274722 408644 274728
rect 408420 274638 408540 274666
rect 408316 272604 408368 272610
rect 408316 272546 408368 272552
rect 407028 267980 407080 267986
rect 407028 267922 407080 267928
rect 407394 267336 407450 267345
rect 407394 267271 407450 267280
rect 407408 264316 407436 267271
rect 407854 265568 407910 265577
rect 407854 265503 407910 265512
rect 407868 264316 407896 265503
rect 408328 264316 408356 272546
rect 408420 272542 408448 274638
rect 408408 272536 408460 272542
rect 408408 272478 408460 272484
rect 408604 272270 408632 274722
rect 409604 272536 409656 272542
rect 409604 272478 409656 272484
rect 408592 272264 408644 272270
rect 408592 272206 408644 272212
rect 408776 266484 408828 266490
rect 408776 266426 408828 266432
rect 408788 264316 408816 266426
rect 409236 266416 409288 266422
rect 409236 266358 409288 266364
rect 409248 264316 409276 266358
rect 409616 264316 409644 272478
rect 409708 266490 409736 275159
rect 409696 266484 409748 266490
rect 409696 266426 409748 266432
rect 409800 266422 409828 276626
rect 409892 274718 409920 277780
rect 409972 274916 410024 274922
rect 409972 274858 410024 274864
rect 409880 274712 409932 274718
rect 409880 274654 409932 274660
rect 409984 272202 410012 274858
rect 411088 274854 411116 277780
rect 411076 274848 411128 274854
rect 411076 274790 411128 274796
rect 412284 274786 412312 277780
rect 412652 277766 413402 277794
rect 412548 275324 412600 275330
rect 412548 275266 412600 275272
rect 412272 274780 412324 274786
rect 412272 274722 412324 274728
rect 411902 273864 411958 273873
rect 411902 273799 411958 273808
rect 410432 272264 410484 272270
rect 410432 272206 410484 272212
rect 409972 272196 410024 272202
rect 409972 272138 410024 272144
rect 409880 267844 409932 267850
rect 409880 267786 409932 267792
rect 409892 267034 409920 267786
rect 409880 267028 409932 267034
rect 409880 266970 409932 266976
rect 410064 266552 410116 266558
rect 410064 266494 410116 266500
rect 409788 266416 409840 266422
rect 409788 266358 409840 266364
rect 410076 264316 410104 266494
rect 410444 266490 410472 272206
rect 410982 267200 411038 267209
rect 410982 267135 411038 267144
rect 410432 266484 410484 266490
rect 410432 266426 410484 266432
rect 410524 266416 410576 266422
rect 410524 266358 410576 266364
rect 410536 264316 410564 266358
rect 410996 264316 411024 267135
rect 411444 266484 411496 266490
rect 411444 266426 411496 266432
rect 411456 264316 411484 266426
rect 411916 266393 411944 273799
rect 412270 267064 412326 267073
rect 412270 266999 412326 267008
rect 411902 266384 411958 266393
rect 411902 266319 411958 266328
rect 412284 264330 412312 266999
rect 412560 266490 412588 275266
rect 412652 267850 412680 277766
rect 414584 276282 414612 277780
rect 414572 276276 414624 276282
rect 414572 276218 414624 276224
rect 415780 271998 415808 277780
rect 416976 273562 417004 277780
rect 416964 273556 417016 273562
rect 416964 273498 417016 273504
rect 415768 271992 415820 271998
rect 415768 271934 415820 271940
rect 412640 267844 412692 267850
rect 412640 267786 412692 267792
rect 417424 267028 417476 267034
rect 417424 266970 417476 266976
rect 417436 266558 417464 266970
rect 417424 266552 417476 266558
rect 417424 266494 417476 266500
rect 412548 266484 412600 266490
rect 412548 266426 412600 266432
rect 418172 265198 418200 277780
rect 419368 274922 419396 277780
rect 419552 277766 420578 277794
rect 419356 274916 419408 274922
rect 419356 274858 419408 274864
rect 419552 268122 419580 277766
rect 421668 276350 421696 277780
rect 421656 276344 421708 276350
rect 421656 276286 421708 276292
rect 422864 272066 422892 277780
rect 422944 272264 422996 272270
rect 422944 272206 422996 272212
rect 422852 272060 422904 272066
rect 422852 272002 422904 272008
rect 419540 268116 419592 268122
rect 419540 268058 419592 268064
rect 422956 266626 422984 272206
rect 424060 272202 424088 277780
rect 425072 277766 425270 277794
rect 424048 272196 424100 272202
rect 424048 272138 424100 272144
rect 422944 266620 422996 266626
rect 422944 266562 422996 266568
rect 425072 265266 425100 277766
rect 426452 267918 426480 277780
rect 427648 275058 427676 277780
rect 428844 276418 428872 277780
rect 428832 276412 428884 276418
rect 428832 276354 428884 276360
rect 427636 275052 427688 275058
rect 427636 274994 427688 275000
rect 427728 275052 427780 275058
rect 427728 274994 427780 275000
rect 427740 273494 427768 274994
rect 427728 273488 427780 273494
rect 427728 273430 427780 273436
rect 429948 270706 429976 277780
rect 431144 272270 431172 277780
rect 431972 277766 432354 277794
rect 433352 277766 433550 277794
rect 431132 272264 431184 272270
rect 431132 272206 431184 272212
rect 431224 272264 431276 272270
rect 431224 272206 431276 272212
rect 429936 270700 429988 270706
rect 429936 270642 429988 270648
rect 426440 267912 426492 267918
rect 426440 267854 426492 267860
rect 431236 266694 431264 272206
rect 431224 266688 431276 266694
rect 431224 266630 431276 266636
rect 431972 265334 432000 277766
rect 433352 265402 433380 277766
rect 434732 274990 434760 277780
rect 435928 276486 435956 277780
rect 435916 276480 435968 276486
rect 435916 276422 435968 276428
rect 434720 274984 434772 274990
rect 434720 274926 434772 274932
rect 438228 272270 438256 277780
rect 438872 277766 439438 277794
rect 443880 277788 444222 277794
rect 443828 277782 444222 277788
rect 438216 272264 438268 272270
rect 438216 272206 438268 272212
rect 438872 265470 438900 277766
rect 441816 275126 441844 277780
rect 441804 275120 441856 275126
rect 441804 275062 441856 275068
rect 443012 269346 443040 277780
rect 443840 277766 444222 277782
rect 444392 277766 445326 277794
rect 445772 277766 446522 277794
rect 447336 277778 447718 277794
rect 447324 277772 447718 277778
rect 443000 269340 443052 269346
rect 443000 269282 443052 269288
rect 444392 266762 444420 277766
rect 445772 269414 445800 277766
rect 447376 277766 447718 277772
rect 447324 277714 447376 277720
rect 448900 275398 448928 277780
rect 449912 277766 450110 277794
rect 448888 275392 448940 275398
rect 448888 275334 448940 275340
rect 448980 275392 449032 275398
rect 448980 275334 449032 275340
rect 448992 271425 449020 275334
rect 448978 271416 449034 271425
rect 448978 271351 449034 271360
rect 449912 269890 449940 277766
rect 449900 269884 449952 269890
rect 449900 269826 449952 269832
rect 445760 269408 445812 269414
rect 445760 269350 445812 269356
rect 444380 266756 444432 266762
rect 444380 266698 444432 266704
rect 438860 265464 438912 265470
rect 438860 265406 438912 265412
rect 433340 265396 433392 265402
rect 433340 265338 433392 265344
rect 431960 265328 432012 265334
rect 431960 265270 432012 265276
rect 425060 265260 425112 265266
rect 425060 265202 425112 265208
rect 418160 265192 418212 265198
rect 418160 265134 418212 265140
rect 451292 264586 451320 277780
rect 452488 277710 452516 277780
rect 452672 277766 453606 277794
rect 452476 277704 452528 277710
rect 452476 277646 452528 277652
rect 451372 269884 451424 269890
rect 451372 269826 451424 269832
rect 451384 266422 451412 269826
rect 452672 269482 452700 277766
rect 454788 277642 454816 277780
rect 455432 277766 455998 277794
rect 456812 277766 457194 277794
rect 454776 277636 454828 277642
rect 454776 277578 454828 277584
rect 452660 269476 452712 269482
rect 452660 269418 452712 269424
rect 455432 266830 455460 277766
rect 456812 270094 456840 277766
rect 458376 275058 458404 277780
rect 459572 275466 459600 277780
rect 459756 277766 460690 277794
rect 459560 275460 459612 275466
rect 459560 275402 459612 275408
rect 459652 275460 459704 275466
rect 459652 275402 459704 275408
rect 458364 275052 458416 275058
rect 458364 274994 458416 275000
rect 458180 274848 458232 274854
rect 458180 274790 458232 274796
rect 458192 273630 458220 274790
rect 458180 273624 458232 273630
rect 458180 273566 458232 273572
rect 459664 272134 459692 275402
rect 459652 272128 459704 272134
rect 459652 272070 459704 272076
rect 456800 270088 456852 270094
rect 456800 270030 456852 270036
rect 457996 270088 458048 270094
rect 457996 270030 458048 270036
rect 458008 267345 458036 270030
rect 459756 269550 459784 277766
rect 461872 274854 461900 277780
rect 462332 277766 463082 277794
rect 463712 277766 464278 277794
rect 461860 274848 461912 274854
rect 461860 274790 461912 274796
rect 459744 269544 459796 269550
rect 459744 269486 459796 269492
rect 457994 267336 458050 267345
rect 457994 267271 458050 267280
rect 462332 266898 462360 277766
rect 463712 269618 463740 277766
rect 465460 273698 465488 277780
rect 466656 275194 466684 277780
rect 466644 275188 466696 275194
rect 466644 275130 466696 275136
rect 466736 275188 466788 275194
rect 466736 275130 466788 275136
rect 465448 273692 465500 273698
rect 465448 273634 465500 273640
rect 466748 270774 466776 275130
rect 466736 270768 466788 270774
rect 466736 270710 466788 270716
rect 467852 269686 467880 277780
rect 468956 273766 468984 277780
rect 469232 277766 470166 277794
rect 470612 277766 471362 277794
rect 468944 273760 468996 273766
rect 468944 273702 468996 273708
rect 467840 269680 467892 269686
rect 467840 269622 467892 269628
rect 463700 269612 463752 269618
rect 463700 269554 463752 269560
rect 469232 267714 469260 277766
rect 470612 269754 470640 277766
rect 472544 273834 472572 277780
rect 473740 275262 473768 277780
rect 474752 277766 474950 277794
rect 473728 275256 473780 275262
rect 473728 275198 473780 275204
rect 474188 275256 474240 275262
rect 474188 275198 474240 275204
rect 472532 273828 472584 273834
rect 472532 273770 472584 273776
rect 470600 269748 470652 269754
rect 470600 269690 470652 269696
rect 470692 269748 470744 269754
rect 470692 269690 470744 269696
rect 469220 267708 469272 267714
rect 469220 267650 469272 267656
rect 470704 266966 470732 269690
rect 474200 268054 474228 275198
rect 474752 270502 474780 277766
rect 476132 273902 476160 277780
rect 476316 277766 477250 277794
rect 476120 273896 476172 273902
rect 476120 273838 476172 273844
rect 474740 270496 474792 270502
rect 474740 270438 474792 270444
rect 476316 269754 476344 277766
rect 478432 276554 478460 277780
rect 478420 276548 478472 276554
rect 478420 276490 478472 276496
rect 479628 274650 479656 277780
rect 480824 276010 480852 277780
rect 481652 277766 482034 277794
rect 480812 276004 480864 276010
rect 480812 275946 480864 275952
rect 479616 274644 479668 274650
rect 479616 274586 479668 274592
rect 476304 269748 476356 269754
rect 476304 269690 476356 269696
rect 474188 268048 474240 268054
rect 474188 267990 474240 267996
rect 470692 266960 470744 266966
rect 470692 266902 470744 266908
rect 462320 266892 462372 266898
rect 462320 266834 462372 266840
rect 455420 266824 455472 266830
rect 455420 266766 455472 266772
rect 451372 266416 451424 266422
rect 451372 266358 451424 266364
rect 481652 265538 481680 277766
rect 483216 274582 483244 277780
rect 483400 277766 484334 277794
rect 483204 274576 483256 274582
rect 483204 274518 483256 274524
rect 483400 267646 483428 277766
rect 485516 276622 485544 277780
rect 485504 276616 485556 276622
rect 485504 276558 485556 276564
rect 486712 274514 486740 277780
rect 487160 276004 487212 276010
rect 487160 275946 487212 275952
rect 486700 274508 486752 274514
rect 486700 274450 486752 274456
rect 487172 268190 487200 275946
rect 487908 275942 487936 277780
rect 488552 277766 489118 277794
rect 487896 275936 487948 275942
rect 487896 275878 487948 275884
rect 487160 268184 487212 268190
rect 487160 268126 487212 268132
rect 483388 267640 483440 267646
rect 483388 267582 483440 267588
rect 488552 265606 488580 277766
rect 490300 274446 490328 277780
rect 491496 277394 491524 277780
rect 491404 277366 491524 277394
rect 492600 277370 492628 277780
rect 492692 277766 493810 277794
rect 490288 274440 490340 274446
rect 490288 274382 490340 274388
rect 491404 267578 491432 277366
rect 492588 277364 492640 277370
rect 492588 277306 492640 277312
rect 491392 267572 491444 267578
rect 491392 267514 491444 267520
rect 488540 265600 488592 265606
rect 488540 265542 488592 265548
rect 481640 265532 481692 265538
rect 481640 265474 481692 265480
rect 451280 264580 451332 264586
rect 451280 264522 451332 264528
rect 492692 264518 492720 277766
rect 494992 275874 495020 277780
rect 495452 277766 496202 277794
rect 496832 277766 497398 277794
rect 498212 277766 498594 277794
rect 494980 275868 495032 275874
rect 494980 275810 495032 275816
rect 495452 266354 495480 277766
rect 496728 275868 496780 275874
rect 496728 275810 496780 275816
rect 496740 270842 496768 275810
rect 496728 270836 496780 270842
rect 496728 270778 496780 270784
rect 496832 270434 496860 277766
rect 496820 270428 496872 270434
rect 496820 270370 496872 270376
rect 498212 267510 498240 277766
rect 499776 277302 499804 277780
rect 499764 277296 499816 277302
rect 499764 277238 499816 277244
rect 500880 274378 500908 277780
rect 502076 275806 502104 277780
rect 502352 277766 503286 277794
rect 502064 275800 502116 275806
rect 502064 275742 502116 275748
rect 502248 275800 502300 275806
rect 502248 275742 502300 275748
rect 500868 274372 500920 274378
rect 500868 274314 500920 274320
rect 502260 268258 502288 275742
rect 502248 268252 502300 268258
rect 502248 268194 502300 268200
rect 498200 267504 498252 267510
rect 498200 267446 498252 267452
rect 495440 266348 495492 266354
rect 495440 266290 495492 266296
rect 502352 266286 502380 277766
rect 504468 272474 504496 277780
rect 505112 277766 505678 277794
rect 504456 272468 504508 272474
rect 504456 272410 504508 272416
rect 505112 267442 505140 277766
rect 506860 277234 506888 277780
rect 507964 277574 507992 277780
rect 507952 277568 508004 277574
rect 507952 277510 508004 277516
rect 506848 277228 506900 277234
rect 506848 277170 506900 277176
rect 509160 275738 509188 277780
rect 509148 275732 509200 275738
rect 509148 275674 509200 275680
rect 510356 275194 510384 277780
rect 510632 277766 511566 277794
rect 512012 277766 512762 277794
rect 510344 275188 510396 275194
rect 510344 275130 510396 275136
rect 510528 274712 510580 274718
rect 510528 274654 510580 274660
rect 510540 270910 510568 274654
rect 510528 270904 510580 270910
rect 510528 270846 510580 270852
rect 510632 270366 510660 277766
rect 510620 270360 510672 270366
rect 510620 270302 510672 270308
rect 505100 267436 505152 267442
rect 505100 267378 505152 267384
rect 512012 267374 512040 277766
rect 513944 275874 513972 277780
rect 514772 277766 515154 277794
rect 513932 275868 513984 275874
rect 513932 275810 513984 275816
rect 513472 275732 513524 275738
rect 513472 275674 513524 275680
rect 513484 272338 513512 275674
rect 513472 272332 513524 272338
rect 513472 272274 513524 272280
rect 514772 269074 514800 277766
rect 516244 275670 516272 277780
rect 516232 275664 516284 275670
rect 516232 275606 516284 275612
rect 516140 274780 516192 274786
rect 516140 274722 516192 274728
rect 516152 270978 516180 274722
rect 517440 274718 517468 277780
rect 517428 274712 517480 274718
rect 517428 274654 517480 274660
rect 518636 274310 518664 277780
rect 518912 277766 519846 277794
rect 518624 274304 518676 274310
rect 518624 274246 518676 274252
rect 516140 270972 516192 270978
rect 516140 270914 516192 270920
rect 514760 269068 514812 269074
rect 514760 269010 514812 269016
rect 512000 267368 512052 267374
rect 512000 267310 512052 267316
rect 518912 267306 518940 277766
rect 521028 274718 521056 277780
rect 521672 277766 522238 277794
rect 521568 275664 521620 275670
rect 521568 275606 521620 275612
rect 521016 274712 521068 274718
rect 521016 274654 521068 274660
rect 521580 272406 521608 275606
rect 521568 272400 521620 272406
rect 521568 272342 521620 272348
rect 521672 270298 521700 277766
rect 523420 275602 523448 277780
rect 523408 275596 523460 275602
rect 523408 275538 523460 275544
rect 523684 275596 523736 275602
rect 523684 275538 523736 275544
rect 521660 270292 521712 270298
rect 521660 270234 521712 270240
rect 523696 267782 523724 275538
rect 524524 271046 524552 277780
rect 525720 274242 525748 277780
rect 525812 277766 526930 277794
rect 525708 274236 525760 274242
rect 525708 274178 525760 274184
rect 524512 271040 524564 271046
rect 524512 270982 524564 270988
rect 523684 267776 523736 267782
rect 523684 267718 523736 267724
rect 518900 267300 518952 267306
rect 518900 267242 518952 267248
rect 525812 267238 525840 277766
rect 528112 271114 528140 277780
rect 529308 271862 529336 277780
rect 530504 275534 530532 277780
rect 530492 275528 530544 275534
rect 530492 275470 530544 275476
rect 529296 271856 529348 271862
rect 529296 271798 529348 271804
rect 531608 271794 531636 277780
rect 532804 273222 532832 277780
rect 532896 277766 534014 277794
rect 532792 273216 532844 273222
rect 532792 273158 532844 273164
rect 531596 271788 531648 271794
rect 531596 271730 531648 271736
rect 528100 271108 528152 271114
rect 528100 271050 528152 271056
rect 525800 267232 525852 267238
rect 525800 267174 525852 267180
rect 532896 267170 532924 277766
rect 535196 271726 535224 277780
rect 535472 277766 536406 277794
rect 535184 271720 535236 271726
rect 535184 271662 535236 271668
rect 535472 270230 535500 277766
rect 537588 275369 537616 277780
rect 537574 275360 537630 275369
rect 537574 275295 537630 275304
rect 538784 271658 538812 277780
rect 539612 277766 539902 277794
rect 538772 271652 538824 271658
rect 538772 271594 538824 271600
rect 535460 270224 535512 270230
rect 535460 270166 535512 270172
rect 539612 268938 539640 277766
rect 541084 277394 541112 277780
rect 540992 277366 541112 277394
rect 539600 268932 539652 268938
rect 539600 268874 539652 268880
rect 532884 267164 532936 267170
rect 532884 267106 532936 267112
rect 540992 267102 541020 277366
rect 542280 271590 542308 277780
rect 543476 274174 543504 277780
rect 543740 275528 543792 275534
rect 544672 275505 544700 277780
rect 545132 277766 545882 277794
rect 543740 275470 543792 275476
rect 544658 275496 544714 275505
rect 543464 274168 543516 274174
rect 543464 274110 543516 274116
rect 542268 271584 542320 271590
rect 542268 271526 542320 271532
rect 543752 269006 543780 275470
rect 544658 275431 544714 275440
rect 543740 269000 543792 269006
rect 543740 268942 543792 268948
rect 540980 267096 541032 267102
rect 540980 267038 541032 267044
rect 502340 266280 502392 266286
rect 502340 266222 502392 266228
rect 545132 266218 545160 277766
rect 547064 271522 547092 277780
rect 547892 277766 548182 277794
rect 547052 271516 547104 271522
rect 547052 271458 547104 271464
rect 547892 270162 547920 277766
rect 549364 277394 549392 277780
rect 549272 277366 549392 277394
rect 547880 270156 547932 270162
rect 547880 270098 547932 270104
rect 545120 266212 545172 266218
rect 545120 266154 545172 266160
rect 549272 266150 549300 277366
rect 550560 271454 550588 277780
rect 551756 274106 551784 277780
rect 552032 277766 552966 277794
rect 551744 274100 551796 274106
rect 551744 274042 551796 274048
rect 550548 271448 550600 271454
rect 550548 271390 550600 271396
rect 549260 266144 549312 266150
rect 549260 266086 549312 266092
rect 552032 266082 552060 277766
rect 554148 271386 554176 277780
rect 554792 277766 555266 277794
rect 556172 277766 556462 277794
rect 554136 271380 554188 271386
rect 554136 271322 554188 271328
rect 554792 270065 554820 277766
rect 554778 270056 554834 270065
rect 554778 269991 554834 270000
rect 552020 266076 552072 266082
rect 552020 266018 552072 266024
rect 556172 266014 556200 277766
rect 557644 271318 557672 277780
rect 558840 274038 558868 277780
rect 558932 277766 560050 277794
rect 558828 274032 558880 274038
rect 558828 273974 558880 273980
rect 557632 271312 557684 271318
rect 557632 271254 557684 271260
rect 556160 266008 556212 266014
rect 556160 265950 556212 265956
rect 558932 265946 558960 277766
rect 561232 271250 561260 277780
rect 562428 271289 562456 277780
rect 563532 277166 563560 277780
rect 564452 277766 564742 277794
rect 563520 277160 563572 277166
rect 563520 277102 563572 277108
rect 562414 271280 562470 271289
rect 561220 271244 561272 271250
rect 562414 271215 562470 271224
rect 561220 271186 561272 271192
rect 558920 265940 558972 265946
rect 558920 265882 558972 265888
rect 564452 265878 564480 277766
rect 565924 269958 565952 277780
rect 566016 277766 567134 277794
rect 567212 277766 568330 277794
rect 565912 269952 565964 269958
rect 565912 269894 565964 269900
rect 564440 265872 564492 265878
rect 564440 265814 564492 265820
rect 566016 265810 566044 277766
rect 567212 270026 567240 277766
rect 569512 274145 569540 277780
rect 570708 277098 570736 277780
rect 570696 277092 570748 277098
rect 570696 277034 570748 277040
rect 571812 277030 571840 277780
rect 571800 277024 571852 277030
rect 571800 276966 571852 276972
rect 569498 274136 569554 274145
rect 569498 274071 569554 274080
rect 573008 272785 573036 277780
rect 574204 277394 574232 277780
rect 574112 277366 574232 277394
rect 574296 277766 575414 277794
rect 575492 277766 576610 277794
rect 572994 272776 573050 272785
rect 572994 272711 573050 272720
rect 567200 270020 567252 270026
rect 567200 269962 567252 269968
rect 566004 265804 566056 265810
rect 566004 265746 566056 265752
rect 574112 265674 574140 277366
rect 574296 265742 574324 277766
rect 574284 265736 574336 265742
rect 574284 265678 574336 265684
rect 574100 265668 574152 265674
rect 574100 265610 574152 265616
rect 492680 264512 492732 264518
rect 492680 264454 492732 264460
rect 575492 264450 575520 277766
rect 577792 275262 577820 277780
rect 577780 275256 577832 275262
rect 577780 275198 577832 275204
rect 578896 271182 578924 277780
rect 579632 277766 580106 277794
rect 578884 271176 578936 271182
rect 578884 271118 578936 271124
rect 579632 269929 579660 277766
rect 581288 275942 581316 277780
rect 582484 276962 582512 277780
rect 582576 277766 583694 277794
rect 582472 276956 582524 276962
rect 582472 276898 582524 276904
rect 581276 275936 581328 275942
rect 581276 275878 581328 275884
rect 581644 275868 581696 275874
rect 581644 275810 581696 275816
rect 579618 269920 579674 269929
rect 579618 269855 579674 269864
rect 581656 268802 581684 275810
rect 581644 268796 581696 268802
rect 581644 268738 581696 268744
rect 575480 264444 575532 264450
rect 575480 264386 575532 264392
rect 582576 264382 582604 277766
rect 583760 276004 583812 276010
rect 583760 275946 583812 275952
rect 583772 273154 583800 275946
rect 584876 275806 584904 277780
rect 585152 277766 586086 277794
rect 586532 277766 587190 277794
rect 587912 277766 588386 277794
rect 584864 275800 584916 275806
rect 584864 275742 584916 275748
rect 583760 273148 583812 273154
rect 583760 273090 583812 273096
rect 585152 265849 585180 277766
rect 586532 269822 586560 277766
rect 586520 269816 586572 269822
rect 586520 269758 586572 269764
rect 587912 268870 587940 277766
rect 589568 276894 589596 277780
rect 589556 276888 589608 276894
rect 589556 276830 589608 276836
rect 590764 273970 590792 277780
rect 591960 275602 591988 277780
rect 593156 275738 593184 277780
rect 594352 277506 594380 277780
rect 594340 277500 594392 277506
rect 594340 277442 594392 277448
rect 593144 275732 593196 275738
rect 593144 275674 593196 275680
rect 591948 275596 592000 275602
rect 591948 275538 592000 275544
rect 593420 275596 593472 275602
rect 593420 275538 593472 275544
rect 590752 273964 590804 273970
rect 590752 273906 590804 273912
rect 593432 273086 593460 275538
rect 595456 275534 595484 277780
rect 596652 275670 596680 277780
rect 597572 277766 597862 277794
rect 596640 275664 596692 275670
rect 596640 275606 596692 275612
rect 595444 275528 595496 275534
rect 595444 275470 595496 275476
rect 593420 273080 593472 273086
rect 593420 273022 593472 273028
rect 587900 268864 587952 268870
rect 587900 268806 587952 268812
rect 585138 265840 585194 265849
rect 585138 265775 585194 265784
rect 411930 264302 412312 264330
rect 582564 264376 582616 264382
rect 582564 264318 582616 264324
rect 597572 264314 597600 277766
rect 599044 275874 599072 277780
rect 600240 276010 600268 277780
rect 600332 277766 601450 277794
rect 601712 277766 602554 277794
rect 603092 277766 603750 277794
rect 600228 276004 600280 276010
rect 600228 275946 600280 275952
rect 599032 275868 599084 275874
rect 599032 275810 599084 275816
rect 597836 275664 597888 275670
rect 597836 275606 597888 275612
rect 597848 272950 597876 275606
rect 600044 275528 600096 275534
rect 600044 275470 600096 275476
rect 600056 273018 600084 275470
rect 600044 273012 600096 273018
rect 600044 272954 600096 272960
rect 597836 272944 597888 272950
rect 597836 272886 597888 272892
rect 600332 268734 600360 277766
rect 600320 268728 600372 268734
rect 600320 268670 600372 268676
rect 601712 268666 601740 277766
rect 603092 269793 603120 277766
rect 604932 271153 604960 277780
rect 605852 277766 606142 277794
rect 604918 271144 604974 271153
rect 604918 271079 604974 271088
rect 603078 269784 603134 269793
rect 603078 269719 603134 269728
rect 601700 268660 601752 268666
rect 601700 268602 601752 268608
rect 605852 268598 605880 277766
rect 607324 275602 607352 277780
rect 607416 277766 608534 277794
rect 608612 277766 609730 277794
rect 607312 275596 607364 275602
rect 607312 275538 607364 275544
rect 605840 268592 605892 268598
rect 605840 268534 605892 268540
rect 597560 264308 597612 264314
rect 393044 264250 393096 264256
rect 597560 264250 597612 264256
rect 396998 264208 397054 264217
rect 194626 264166 194916 264194
rect 396750 264166 396998 264194
rect 401230 264208 401286 264217
rect 399418 264178 399800 264194
rect 399418 264172 399812 264178
rect 399418 264166 399760 264172
rect 396998 264143 397054 264152
rect 607416 264178 607444 277766
rect 608612 268530 608640 277766
rect 610820 275670 610848 277780
rect 612016 277438 612044 277780
rect 612752 277766 613226 277794
rect 612004 277432 612056 277438
rect 612004 277374 612056 277380
rect 610808 275664 610860 275670
rect 610808 275606 610860 275612
rect 612752 268705 612780 277766
rect 614408 275534 614436 277780
rect 615604 277394 615632 277780
rect 615512 277366 615632 277394
rect 615696 277766 616814 277794
rect 614396 275528 614448 275534
rect 614396 275470 614448 275476
rect 612738 268696 612794 268705
rect 612738 268631 612794 268640
rect 608600 268524 608652 268530
rect 608600 268466 608652 268472
rect 401230 264143 401232 264152
rect 399760 264114 399812 264120
rect 401284 264143 401286 264152
rect 607404 264172 607456 264178
rect 401232 264114 401284 264120
rect 607404 264114 607456 264120
rect 615512 264110 615540 277366
rect 615696 268462 615724 277766
rect 617996 272882 618024 277780
rect 619100 274009 619128 277780
rect 619652 277766 620310 277794
rect 619086 274000 619142 274009
rect 619086 273935 619142 273944
rect 617984 272876 618036 272882
rect 617984 272818 618036 272824
rect 615684 268456 615736 268462
rect 615684 268398 615736 268404
rect 619652 268394 619680 277766
rect 621492 272814 621520 277780
rect 622412 277766 622702 277794
rect 621480 272808 621532 272814
rect 621480 272750 621532 272756
rect 622412 268569 622440 277766
rect 623884 277394 623912 277780
rect 623792 277366 623912 277394
rect 622398 268560 622454 268569
rect 622398 268495 622454 268504
rect 623792 268433 623820 277366
rect 625080 272746 625108 277780
rect 626184 275466 626212 277780
rect 627380 276826 627408 277780
rect 627368 276820 627420 276826
rect 627368 276762 627420 276768
rect 626172 275460 626224 275466
rect 626172 275402 626224 275408
rect 625068 272740 625120 272746
rect 625068 272682 625120 272688
rect 628576 272649 628604 277780
rect 629772 273873 629800 277780
rect 630692 277766 630982 277794
rect 629758 273864 629814 273873
rect 629758 273799 629814 273808
rect 628562 272640 628618 272649
rect 628562 272575 628618 272584
rect 623778 268424 623834 268433
rect 619640 268388 619692 268394
rect 623778 268359 623834 268368
rect 619640 268330 619692 268336
rect 630692 265713 630720 277766
rect 632164 272678 632192 277780
rect 633360 275398 633388 277780
rect 634464 276758 634492 277780
rect 634452 276752 634504 276758
rect 634452 276694 634504 276700
rect 633348 275392 633400 275398
rect 633348 275334 633400 275340
rect 632152 272672 632204 272678
rect 632152 272614 632204 272620
rect 635660 272513 635688 277780
rect 636212 277766 636870 277794
rect 637592 277766 638066 277794
rect 635646 272504 635702 272513
rect 635646 272439 635702 272448
rect 636212 270094 636240 277766
rect 636200 270088 636252 270094
rect 636200 270030 636252 270036
rect 630678 265704 630734 265713
rect 630678 265639 630734 265648
rect 637592 265577 637620 277766
rect 639248 272610 639276 277780
rect 640444 275233 640472 277780
rect 641640 276690 641668 277780
rect 641628 276684 641680 276690
rect 641628 276626 641680 276632
rect 640430 275224 640486 275233
rect 640430 275159 640486 275168
rect 639236 272604 639288 272610
rect 639236 272546 639288 272552
rect 642744 272542 642772 277780
rect 643112 277766 643954 277794
rect 644492 277766 645150 277794
rect 642732 272536 642784 272542
rect 642732 272478 642784 272484
rect 643112 267034 643140 277766
rect 644492 269890 644520 277766
rect 644480 269884 644532 269890
rect 644480 269826 644532 269832
rect 645872 267209 645900 278310
rect 646044 278248 646096 278254
rect 646044 278190 646096 278196
rect 645858 267200 645914 267209
rect 645858 267135 645914 267144
rect 643100 267028 643152 267034
rect 643100 266970 643152 266976
rect 637578 265568 637634 265577
rect 637578 265503 637634 265512
rect 615500 264104 615552 264110
rect 615500 264046 615552 264052
rect 415306 262304 415362 262313
rect 415306 262239 415308 262248
rect 415360 262239 415362 262248
rect 572720 262268 572772 262274
rect 415308 262210 415360 262216
rect 572720 262210 572772 262216
rect 414202 259176 414258 259185
rect 414202 259111 414258 259120
rect 189078 258632 189134 258641
rect 189078 258567 189134 258576
rect 189092 258398 189120 258567
rect 185216 258392 185268 258398
rect 185216 258334 185268 258340
rect 189080 258392 189132 258398
rect 189080 258334 189132 258340
rect 185228 253201 185256 258334
rect 414216 258126 414244 259111
rect 414204 258120 414256 258126
rect 414204 258062 414256 258068
rect 571524 258120 571576 258126
rect 571524 258062 571576 258068
rect 415306 255912 415362 255921
rect 415306 255847 415362 255856
rect 415320 255338 415348 255847
rect 415308 255332 415360 255338
rect 415308 255274 415360 255280
rect 571432 255332 571484 255338
rect 571432 255274 571484 255280
rect 185214 253192 185270 253201
rect 185214 253127 185270 253136
rect 414386 252784 414442 252793
rect 414386 252719 414442 252728
rect 414400 252618 414428 252719
rect 414388 252612 414440 252618
rect 414388 252554 414440 252560
rect 414202 249520 414258 249529
rect 414202 249455 414258 249464
rect 414216 248470 414244 249455
rect 414204 248464 414256 248470
rect 414204 248406 414256 248412
rect 438216 248464 438268 248470
rect 438216 248406 438268 248412
rect 190366 248024 190422 248033
rect 190366 247959 190422 247968
rect 189722 247208 189778 247217
rect 189722 247143 189778 247152
rect 117964 245676 118016 245682
rect 117964 245618 118016 245624
rect 65156 231600 65208 231606
rect 65156 231542 65208 231548
rect 64144 231464 64196 231470
rect 64144 231406 64196 231412
rect 54484 231396 54536 231402
rect 54484 231338 54536 231344
rect 53104 231192 53156 231198
rect 53104 231134 53156 231140
rect 64142 229936 64198 229945
rect 64142 229871 64198 229880
rect 57886 229800 57942 229809
rect 57886 229735 57942 229744
rect 56324 228472 56376 228478
rect 56324 228414 56376 228420
rect 53656 228404 53708 228410
rect 53656 228346 53708 228352
rect 52736 225616 52788 225622
rect 52736 225558 52788 225564
rect 52276 219428 52328 219434
rect 52276 219370 52328 219376
rect 52184 215960 52236 215966
rect 52184 215902 52236 215908
rect 46204 214600 46256 214606
rect 46204 214542 46256 214548
rect 50344 214396 50396 214402
rect 50344 214338 50396 214344
rect 50068 214328 50120 214334
rect 50068 214270 50120 214276
rect 47216 214260 47268 214266
rect 47216 214202 47268 214208
rect 47228 212537 47256 214202
rect 47214 212528 47270 212537
rect 47214 212463 47270 212472
rect 44730 211304 44786 211313
rect 44730 211239 44786 211248
rect 50080 210633 50108 214270
rect 50066 210624 50122 210633
rect 50066 210559 50122 210568
rect 42798 209264 42854 209273
rect 42798 209199 42854 209208
rect 39302 208584 39358 208593
rect 39302 208519 39358 208528
rect 31298 204912 31354 204921
rect 31298 204847 31354 204856
rect 31114 204504 31170 204513
rect 31114 204439 31170 204448
rect 35806 203280 35862 203289
rect 35806 203215 35862 203224
rect 35820 202910 35848 203215
rect 35808 202904 35860 202910
rect 35808 202846 35860 202852
rect 31022 199336 31078 199345
rect 31022 199271 31078 199280
rect 39316 197713 39344 208519
rect 39302 197704 39358 197713
rect 39302 197639 39358 197648
rect 41878 197160 41934 197169
rect 41878 197095 41934 197104
rect 41892 196656 41920 197095
rect 41786 195256 41842 195265
rect 41786 195191 41842 195200
rect 41800 194820 41828 195191
rect 42064 193180 42116 193186
rect 42064 193122 42116 193128
rect 42076 192984 42104 193122
rect 42168 191690 42196 191760
rect 42156 191684 42208 191690
rect 42156 191626 42208 191632
rect 42064 191480 42116 191486
rect 42064 191422 42116 191428
rect 42076 191148 42104 191422
rect 42156 190868 42208 190874
rect 42156 190810 42208 190816
rect 42168 190468 42196 190810
rect 41786 190224 41842 190233
rect 41786 190159 41842 190168
rect 41800 189924 41828 190159
rect 42156 187672 42208 187678
rect 42156 187614 42208 187620
rect 42168 187445 42196 187614
rect 42154 187368 42210 187377
rect 42154 187303 42210 187312
rect 42168 186796 42196 187303
rect 42064 186312 42116 186318
rect 42064 186254 42116 186260
rect 42076 186184 42104 186254
rect 42812 185910 42840 209199
rect 44178 208040 44234 208049
rect 44178 207975 44234 207984
rect 42890 207632 42946 207641
rect 42890 207567 42946 207576
rect 42904 186318 42932 207567
rect 43350 206816 43406 206825
rect 43350 206751 43406 206760
rect 43166 206408 43222 206417
rect 43166 206343 43222 206352
rect 42982 206000 43038 206009
rect 42982 205935 43038 205944
rect 42996 187678 43024 205935
rect 43180 191486 43208 206343
rect 43258 205184 43314 205193
rect 43258 205119 43314 205128
rect 43272 191690 43300 205119
rect 43364 193186 43392 206751
rect 43442 205592 43498 205601
rect 43442 205527 43498 205536
rect 43352 193180 43404 193186
rect 43352 193122 43404 193128
rect 43260 191684 43312 191690
rect 43260 191626 43312 191632
rect 43168 191480 43220 191486
rect 43168 191422 43220 191428
rect 43456 190874 43484 205527
rect 43444 190868 43496 190874
rect 43444 190810 43496 190816
rect 42984 187672 43036 187678
rect 42984 187614 43036 187620
rect 42892 186312 42944 186318
rect 42892 186254 42944 186260
rect 42156 185904 42208 185910
rect 42156 185846 42208 185852
rect 42800 185904 42852 185910
rect 42800 185846 42852 185852
rect 42168 185605 42196 185846
rect 41878 184240 41934 184249
rect 41878 184175 41934 184184
rect 41892 183765 41920 184175
rect 44192 183462 44220 207975
rect 50356 202910 50384 214338
rect 50344 202904 50396 202910
rect 50344 202846 50396 202852
rect 42156 183456 42208 183462
rect 42156 183398 42208 183404
rect 44180 183456 44232 183462
rect 44180 183398 44232 183404
rect 42168 183124 42196 183398
rect 41786 183016 41842 183025
rect 41786 182951 41842 182960
rect 41800 182477 41828 182951
rect 52196 52465 52224 215902
rect 52288 52494 52316 219370
rect 52748 217410 52776 225558
rect 53668 217410 53696 228346
rect 56048 225684 56100 225690
rect 56048 225626 56100 225632
rect 55126 222864 55182 222873
rect 55126 222799 55182 222808
rect 54392 219496 54444 219502
rect 54392 219438 54444 219444
rect 54404 217410 54432 219438
rect 55140 217410 55168 222799
rect 56060 217410 56088 225626
rect 56336 219502 56364 228414
rect 56600 223576 56652 223582
rect 56600 223518 56652 223524
rect 56612 219502 56640 223518
rect 56874 221504 56930 221513
rect 56874 221439 56930 221448
rect 56324 219496 56376 219502
rect 56324 219438 56376 219444
rect 56600 219496 56652 219502
rect 56600 219438 56652 219444
rect 56888 217410 56916 221439
rect 57900 219434 57928 229735
rect 62120 229152 62172 229158
rect 62120 229094 62172 229100
rect 59266 226944 59322 226953
rect 59266 226879 59322 226888
rect 58622 223000 58678 223009
rect 58622 222935 58678 222944
rect 57808 219406 57928 219434
rect 57808 217410 57836 219406
rect 58636 217410 58664 222935
rect 59280 217410 59308 226879
rect 62132 226386 62160 229094
rect 62762 227080 62818 227089
rect 62762 227015 62818 227024
rect 62040 226358 62160 226386
rect 61934 224224 61990 224233
rect 61934 224159 61990 224168
rect 60280 221468 60332 221474
rect 60280 221410 60332 221416
rect 60292 217410 60320 221410
rect 61108 220788 61160 220794
rect 61108 220730 61160 220736
rect 61120 217410 61148 220730
rect 61948 219434 61976 224159
rect 62040 223650 62068 226358
rect 62028 223644 62080 223650
rect 62028 223586 62080 223592
rect 61948 219406 62068 219434
rect 62040 217410 62068 219406
rect 62776 217410 62804 227015
rect 63408 221536 63460 221542
rect 63408 221478 63460 221484
rect 63420 217410 63448 221478
rect 64156 220794 64184 229871
rect 65168 229158 65196 231542
rect 91744 229900 91796 229906
rect 91744 229842 91796 229848
rect 82820 229832 82872 229838
rect 82820 229774 82872 229780
rect 73804 229764 73856 229770
rect 73804 229706 73856 229712
rect 65156 229152 65208 229158
rect 65156 229094 65208 229100
rect 72974 227216 73030 227225
rect 72974 227151 73030 227160
rect 72054 224496 72110 224505
rect 72054 224431 72110 224440
rect 69478 224360 69534 224369
rect 69478 224295 69534 224304
rect 69020 223032 69072 223038
rect 69020 222974 69072 222980
rect 68744 222964 68796 222970
rect 68744 222906 68796 222912
rect 65340 222896 65392 222902
rect 65340 222838 65392 222844
rect 64144 220788 64196 220794
rect 64144 220730 64196 220736
rect 64512 220108 64564 220114
rect 64512 220050 64564 220056
rect 64524 217410 64552 220050
rect 65352 217410 65380 222838
rect 66994 221640 67050 221649
rect 66994 221575 67050 221584
rect 66076 220244 66128 220250
rect 66076 220186 66128 220192
rect 66088 217410 66116 220186
rect 67008 217410 67036 221575
rect 67546 220144 67602 220153
rect 67546 220079 67602 220088
rect 67560 217410 67588 220079
rect 68756 217410 68784 222906
rect 69032 220250 69060 222974
rect 69020 220244 69072 220250
rect 69020 220186 69072 220192
rect 69492 217410 69520 224295
rect 70214 221776 70270 221785
rect 70214 221711 70270 221720
rect 70228 217410 70256 221711
rect 71228 220788 71280 220794
rect 71228 220730 71280 220736
rect 71240 217410 71268 220730
rect 72068 217410 72096 224431
rect 72988 217410 73016 227151
rect 73710 221912 73766 221921
rect 73710 221847 73766 221856
rect 73724 217410 73752 221847
rect 73816 220794 73844 229706
rect 82832 227798 82860 229774
rect 90546 228440 90602 228449
rect 90546 228375 90602 228384
rect 86866 228304 86922 228313
rect 86866 228239 86922 228248
rect 77944 227792 77996 227798
rect 77944 227734 77996 227740
rect 82820 227792 82872 227798
rect 82820 227734 82872 227740
rect 84660 227792 84712 227798
rect 84660 227734 84712 227740
rect 76288 225752 76340 225758
rect 76288 225694 76340 225700
rect 75368 223100 75420 223106
rect 75368 223042 75420 223048
rect 73804 220788 73856 220794
rect 73804 220730 73856 220736
rect 74446 220280 74502 220289
rect 74446 220215 74502 220224
rect 74460 217410 74488 220215
rect 75380 217410 75408 223042
rect 76300 217410 76328 225694
rect 77024 221604 77076 221610
rect 77024 221546 77076 221552
rect 77036 217410 77064 221546
rect 77956 217410 77984 227734
rect 82728 227180 82780 227186
rect 82728 227122 82780 227128
rect 78494 224632 78550 224641
rect 78494 224567 78550 224576
rect 78508 217410 78536 224567
rect 82176 223168 82228 223174
rect 82176 223110 82228 223116
rect 80428 221672 80480 221678
rect 80428 221614 80480 221620
rect 79600 220312 79652 220318
rect 79600 220254 79652 220260
rect 79612 217410 79640 220254
rect 80440 217410 80468 221614
rect 81256 220176 81308 220182
rect 81256 220118 81308 220124
rect 81268 217410 81296 220118
rect 82188 217410 82216 223110
rect 82740 217410 82768 227122
rect 83832 221740 83884 221746
rect 83832 221682 83884 221688
rect 83844 217410 83872 221682
rect 84672 217410 84700 227734
rect 86316 225820 86368 225826
rect 86316 225762 86368 225768
rect 85488 221808 85540 221814
rect 85488 221750 85540 221756
rect 85500 217410 85528 221750
rect 86328 217410 86356 225762
rect 86880 217410 86908 228239
rect 89534 225584 89590 225593
rect 89534 225519 89590 225528
rect 88156 224256 88208 224262
rect 88156 224198 88208 224204
rect 88168 217410 88196 224198
rect 88892 221876 88944 221882
rect 88892 221818 88944 221824
rect 88904 217410 88932 221818
rect 89548 217410 89576 225519
rect 90560 217410 90588 228375
rect 91756 227798 91784 229842
rect 117228 229016 117280 229022
rect 117228 228958 117280 228964
rect 114192 228948 114244 228954
rect 114192 228890 114244 228896
rect 110696 228880 110748 228886
rect 110696 228822 110748 228828
rect 107476 228812 107528 228818
rect 107476 228754 107528 228760
rect 103980 228744 104032 228750
rect 103980 228686 104032 228692
rect 100668 228676 100720 228682
rect 100668 228618 100720 228624
rect 97264 228608 97316 228614
rect 97264 228550 97316 228556
rect 93768 228540 93820 228546
rect 93768 228482 93820 228488
rect 91744 227792 91796 227798
rect 91744 227734 91796 227740
rect 91376 227384 91428 227390
rect 91376 227326 91428 227332
rect 91388 217410 91416 227326
rect 93030 225720 93086 225729
rect 93030 225655 93086 225664
rect 92294 223136 92350 223145
rect 92294 223071 92350 223080
rect 92308 217410 92336 223071
rect 93044 217410 93072 225655
rect 93780 217410 93808 228482
rect 96528 225888 96580 225894
rect 96528 225830 96580 225836
rect 95608 223236 95660 223242
rect 95608 223178 95660 223184
rect 94780 220244 94832 220250
rect 94780 220186 94832 220192
rect 94792 217410 94820 220186
rect 95620 217410 95648 223178
rect 96540 217410 96568 225830
rect 97276 217410 97304 228550
rect 99840 225956 99892 225962
rect 99840 225898 99892 225904
rect 99010 223272 99066 223281
rect 99010 223207 99066 223216
rect 97816 219564 97868 219570
rect 97816 219506 97868 219512
rect 97828 217410 97856 219506
rect 99024 217410 99052 223207
rect 99852 217410 99880 225898
rect 100680 217410 100708 228618
rect 103244 226024 103296 226030
rect 103244 225966 103296 225972
rect 101496 224324 101548 224330
rect 101496 224266 101548 224272
rect 100760 222012 100812 222018
rect 100760 221954 100812 221960
rect 100772 220318 100800 221954
rect 100760 220312 100812 220318
rect 100760 220254 100812 220260
rect 101508 217410 101536 224266
rect 101956 223304 102008 223310
rect 101956 223246 102008 223252
rect 52440 217382 52776 217410
rect 53268 217382 53696 217410
rect 54096 217382 54432 217410
rect 54924 217382 55168 217410
rect 55752 217382 56088 217410
rect 56580 217382 56916 217410
rect 57408 217382 57836 217410
rect 58328 217382 58664 217410
rect 59156 217382 59308 217410
rect 59984 217382 60320 217410
rect 60812 217382 61148 217410
rect 61640 217382 62068 217410
rect 62468 217382 62804 217410
rect 63296 217382 63448 217410
rect 64216 217382 64552 217410
rect 65044 217382 65380 217410
rect 65872 217382 66116 217410
rect 66700 217382 67036 217410
rect 67528 217382 67588 217410
rect 68356 217382 68784 217410
rect 69184 217382 69520 217410
rect 70104 217382 70256 217410
rect 70932 217382 71268 217410
rect 71760 217382 72096 217410
rect 72588 217382 73016 217410
rect 73416 217382 73752 217410
rect 74244 217382 74488 217410
rect 75072 217382 75408 217410
rect 75992 217382 76328 217410
rect 76820 217382 77064 217410
rect 77648 217382 77984 217410
rect 78476 217382 78536 217410
rect 79304 217382 79640 217410
rect 80132 217382 80468 217410
rect 80960 217382 81296 217410
rect 81880 217382 82216 217410
rect 82708 217382 82768 217410
rect 83536 217382 83872 217410
rect 84364 217382 84700 217410
rect 85192 217382 85528 217410
rect 86020 217382 86356 217410
rect 86848 217382 86908 217410
rect 87768 217382 88196 217410
rect 88596 217382 88932 217410
rect 89424 217382 89576 217410
rect 90252 217382 90588 217410
rect 91080 217382 91416 217410
rect 91908 217382 92336 217410
rect 92736 217382 93072 217410
rect 93656 217382 93808 217410
rect 94484 217382 94820 217410
rect 95312 217382 95648 217410
rect 96140 217382 96568 217410
rect 96968 217382 97304 217410
rect 97796 217382 97856 217410
rect 98624 217382 99052 217410
rect 99544 217382 99880 217410
rect 100372 217382 100708 217410
rect 101200 217382 101536 217410
rect 101968 217410 101996 223246
rect 103256 217410 103284 225966
rect 103992 217410 104020 228686
rect 106556 226092 106608 226098
rect 106556 226034 106608 226040
rect 105728 223372 105780 223378
rect 105728 223314 105780 223320
rect 104716 220312 104768 220318
rect 104716 220254 104768 220260
rect 104728 217410 104756 220254
rect 105740 217410 105768 223314
rect 106568 217410 106596 226034
rect 107488 217410 107516 228754
rect 108212 227520 108264 227526
rect 108212 227462 108264 227468
rect 108224 217410 108252 227462
rect 109868 226160 109920 226166
rect 109868 226102 109920 226108
rect 108856 223440 108908 223446
rect 108856 223382 108908 223388
rect 108868 217410 108896 223382
rect 109880 217410 109908 226102
rect 110708 217410 110736 228822
rect 112996 226228 113048 226234
rect 112996 226170 113048 226176
rect 112444 221944 112496 221950
rect 112444 221886 112496 221892
rect 111616 220448 111668 220454
rect 111616 220390 111668 220396
rect 111628 217410 111656 220390
rect 112456 217410 112484 221886
rect 113008 217410 113036 226170
rect 114204 217410 114232 228890
rect 116584 226296 116636 226302
rect 116584 226238 116636 226244
rect 114928 224732 114980 224738
rect 114928 224674 114980 224680
rect 114940 217410 114968 224674
rect 115756 223508 115808 223514
rect 115756 223450 115808 223456
rect 115768 217410 115796 223450
rect 116596 217410 116624 226238
rect 117240 217410 117268 228958
rect 117976 218657 118004 245618
rect 175002 241632 175058 241641
rect 175002 241567 175004 241576
rect 175056 241567 175058 241576
rect 175004 241538 175056 241544
rect 155868 240848 155920 240854
rect 155868 240790 155920 240796
rect 155880 236026 155908 240790
rect 184940 237448 184992 237454
rect 189080 237448 189132 237454
rect 184940 237390 184992 237396
rect 189078 237416 189080 237425
rect 189132 237416 189134 237425
rect 153108 236020 153160 236026
rect 153108 235962 153160 235968
rect 155868 236020 155920 236026
rect 155868 235962 155920 235968
rect 153120 233918 153148 235962
rect 184952 234682 184980 237390
rect 189078 237351 189134 237360
rect 184860 234654 184980 234682
rect 130384 233912 130436 233918
rect 130384 233854 130436 233860
rect 153108 233912 153160 233918
rect 153108 233854 153160 233860
rect 120816 229084 120868 229090
rect 120816 229026 120868 229032
rect 119896 225548 119948 225554
rect 119896 225490 119948 225496
rect 119160 222080 119212 222086
rect 119160 222022 119212 222028
rect 118332 220584 118384 220590
rect 118332 220526 118384 220532
rect 117962 218648 118018 218657
rect 117962 218583 118018 218592
rect 118344 217410 118372 220526
rect 118700 218068 118752 218074
rect 118700 218010 118752 218016
rect 101968 217382 102028 217410
rect 102856 217382 103284 217410
rect 103684 217382 104020 217410
rect 104512 217382 104756 217410
rect 105432 217382 105768 217410
rect 106260 217382 106596 217410
rect 107088 217382 107516 217410
rect 107916 217382 108252 217410
rect 108744 217382 108896 217410
rect 109572 217382 109908 217410
rect 110400 217382 110736 217410
rect 111320 217382 111656 217410
rect 112148 217382 112484 217410
rect 112976 217382 113036 217410
rect 113804 217382 114232 217410
rect 114632 217382 114968 217410
rect 115460 217382 115796 217410
rect 116288 217382 116624 217410
rect 117208 217382 117268 217410
rect 118036 217382 118372 217410
rect 118712 216442 118740 218010
rect 119172 217410 119200 222022
rect 119908 217410 119936 225490
rect 120828 217410 120856 229026
rect 127532 228336 127584 228342
rect 127532 228278 127584 228284
rect 124128 227044 124180 227050
rect 124128 226986 124180 226992
rect 123392 225480 123444 225486
rect 123392 225422 123444 225428
rect 122472 222148 122524 222154
rect 122472 222090 122524 222096
rect 121276 220516 121328 220522
rect 121276 220458 121328 220464
rect 118864 217382 119200 217410
rect 119692 217382 119936 217410
rect 120520 217382 120856 217410
rect 121288 217410 121316 220458
rect 122484 217410 122512 222090
rect 123404 217410 123432 225422
rect 124140 217410 124168 226986
rect 125048 226976 125100 226982
rect 125048 226918 125100 226924
rect 124864 226364 124916 226370
rect 124864 226306 124916 226312
rect 124876 218074 124904 226306
rect 124864 218068 124916 218074
rect 124864 218010 124916 218016
rect 125060 217410 125088 226918
rect 126796 225412 126848 225418
rect 126796 225354 126848 225360
rect 125876 223576 125928 223582
rect 125876 223518 125928 223524
rect 125888 217410 125916 223518
rect 126808 217410 126836 225354
rect 127544 217410 127572 228278
rect 130396 226370 130424 233854
rect 184860 232558 184888 234654
rect 177120 232552 177172 232558
rect 177120 232494 177172 232500
rect 184848 232552 184900 232558
rect 184848 232494 184900 232500
rect 177132 231606 177160 232494
rect 189736 231606 189764 247143
rect 190380 231742 190408 247959
rect 191102 247344 191158 247353
rect 191102 247279 191158 247288
rect 190368 231736 190420 231742
rect 190368 231678 190420 231684
rect 191116 231674 191144 247279
rect 415306 246392 415362 246401
rect 415306 246327 415362 246336
rect 415320 245682 415348 246327
rect 415308 245676 415360 245682
rect 415308 245618 415360 245624
rect 438124 245676 438176 245682
rect 438124 245618 438176 245624
rect 414386 243128 414442 243137
rect 414386 243063 414442 243072
rect 414400 242962 414428 243063
rect 414388 242956 414440 242962
rect 414388 242898 414440 242904
rect 414938 240000 414994 240009
rect 414938 239935 414994 239944
rect 414952 238814 414980 239935
rect 414940 238808 414992 238814
rect 414940 238750 414992 238756
rect 428464 238808 428516 238814
rect 428464 238750 428516 238756
rect 414202 236736 414258 236745
rect 414202 236671 414258 236680
rect 414216 232558 414244 236671
rect 415306 233608 415362 233617
rect 415306 233543 415362 233552
rect 415320 233306 415348 233543
rect 415308 233300 415360 233306
rect 415308 233242 415360 233248
rect 427084 233300 427136 233306
rect 427084 233242 427136 233248
rect 414204 232552 414256 232558
rect 414204 232494 414256 232500
rect 427096 232490 427124 233242
rect 427084 232484 427136 232490
rect 427084 232426 427136 232432
rect 263704 231798 263902 231826
rect 428476 231810 428504 238750
rect 438136 233918 438164 245618
rect 438228 238066 438256 248406
rect 438216 238060 438268 238066
rect 438216 238002 438268 238008
rect 438124 233912 438176 233918
rect 438124 233854 438176 233860
rect 428464 231804 428516 231810
rect 191104 231668 191156 231674
rect 191104 231610 191156 231616
rect 177120 231600 177172 231606
rect 177120 231542 177172 231548
rect 189724 231600 189776 231606
rect 189724 231542 189776 231548
rect 179328 230444 179380 230450
rect 179328 230386 179380 230392
rect 175188 230376 175240 230382
rect 175188 230318 175240 230324
rect 169668 230308 169720 230314
rect 169668 230250 169720 230256
rect 136364 230240 136416 230246
rect 136364 230182 136416 230188
rect 132408 229968 132460 229974
rect 132408 229910 132460 229916
rect 131028 228268 131080 228274
rect 131028 228210 131080 228216
rect 130384 226364 130436 226370
rect 130384 226306 130436 226312
rect 130108 225344 130160 225350
rect 130108 225286 130160 225292
rect 129280 221400 129332 221406
rect 129280 221342 129332 221348
rect 128176 220652 128228 220658
rect 128176 220594 128228 220600
rect 128188 217410 128216 220594
rect 129292 217410 129320 221342
rect 130120 217410 130148 225286
rect 131040 217410 131068 228210
rect 132316 222828 132368 222834
rect 132316 222770 132368 222776
rect 131764 220788 131816 220794
rect 131764 220730 131816 220736
rect 131776 217410 131804 220730
rect 132328 217410 132356 222770
rect 132420 220794 132448 229910
rect 134248 227112 134300 227118
rect 134248 227054 134300 227060
rect 133512 225276 133564 225282
rect 133512 225218 133564 225224
rect 132408 220788 132460 220794
rect 132408 220730 132460 220736
rect 133524 217410 133552 225218
rect 134260 217410 134288 227054
rect 135996 224392 136048 224398
rect 135996 224334 136048 224340
rect 134984 220720 135036 220726
rect 134984 220662 135036 220668
rect 134996 217410 135024 220662
rect 136008 217410 136036 224334
rect 136376 224330 136404 230182
rect 155868 230172 155920 230178
rect 155868 230114 155920 230120
rect 146208 230104 146260 230110
rect 146208 230046 146260 230052
rect 139308 230036 139360 230042
rect 139308 229978 139360 229984
rect 137744 228200 137796 228206
rect 137744 228142 137796 228148
rect 136364 224324 136416 224330
rect 136364 224266 136416 224272
rect 136548 224324 136600 224330
rect 136548 224266 136600 224272
rect 136560 217410 136588 224266
rect 137756 217410 137784 228142
rect 139216 224460 139268 224466
rect 139216 224402 139268 224408
rect 138480 220788 138532 220794
rect 138480 220730 138532 220736
rect 138492 217410 138520 220730
rect 139228 217410 139256 224402
rect 139320 220794 139348 229978
rect 140044 229696 140096 229702
rect 140044 229638 140096 229644
rect 140056 227186 140084 229638
rect 144368 228132 144420 228138
rect 144368 228074 144420 228080
rect 143448 227316 143500 227322
rect 143448 227258 143500 227264
rect 141056 227248 141108 227254
rect 141056 227190 141108 227196
rect 140044 227180 140096 227186
rect 140044 227122 140096 227128
rect 140136 227180 140188 227186
rect 140136 227122 140188 227128
rect 139308 220788 139360 220794
rect 139308 220730 139360 220736
rect 140148 217410 140176 227122
rect 141068 217410 141096 227190
rect 142712 224528 142764 224534
rect 142712 224470 142764 224476
rect 141884 220788 141936 220794
rect 141884 220730 141936 220736
rect 141896 217410 141924 220730
rect 142724 217410 142752 224470
rect 143460 217410 143488 227258
rect 144380 217410 144408 228074
rect 146116 224596 146168 224602
rect 146116 224538 146168 224544
rect 145196 220380 145248 220386
rect 145196 220322 145248 220328
rect 145208 217410 145236 220322
rect 146128 217410 146156 224538
rect 146220 220386 146248 230046
rect 151820 229628 151872 229634
rect 151820 229570 151872 229576
rect 149704 229560 149756 229566
rect 149704 229502 149756 229508
rect 146392 229492 146444 229498
rect 146392 229434 146444 229440
rect 146404 227390 146432 229434
rect 149716 227526 149744 229502
rect 149704 227520 149756 227526
rect 149704 227462 149756 227468
rect 150348 227520 150400 227526
rect 150348 227462 150400 227468
rect 147588 227452 147640 227458
rect 147588 227394 147640 227400
rect 146392 227384 146444 227390
rect 146392 227326 146444 227332
rect 146944 227384 146996 227390
rect 146944 227326 146996 227332
rect 146208 220380 146260 220386
rect 146208 220322 146260 220328
rect 146956 217410 146984 227326
rect 147600 217410 147628 227394
rect 149428 224664 149480 224670
rect 149428 224606 149480 224612
rect 148600 220040 148652 220046
rect 148600 219982 148652 219988
rect 148612 217410 148640 219982
rect 149440 217410 149468 224606
rect 150360 217410 150388 227462
rect 151832 224738 151860 229570
rect 154488 228064 154540 228070
rect 154488 228006 154540 228012
rect 153660 227588 153712 227594
rect 153660 227530 153712 227536
rect 151820 224732 151872 224738
rect 151820 224674 151872 224680
rect 152924 224732 152976 224738
rect 152924 224674 152976 224680
rect 151084 221332 151136 221338
rect 151084 221274 151136 221280
rect 151096 217410 151124 221274
rect 151728 219972 151780 219978
rect 151728 219914 151780 219920
rect 151740 217410 151768 219914
rect 152936 217410 152964 224674
rect 153672 217410 153700 227530
rect 154500 217410 154528 228006
rect 155776 224800 155828 224806
rect 155776 224742 155828 224748
rect 155316 220380 155368 220386
rect 155316 220322 155368 220328
rect 155328 217410 155356 220322
rect 121288 217382 121348 217410
rect 122176 217382 122512 217410
rect 123096 217382 123432 217410
rect 123924 217382 124168 217410
rect 124752 217382 125088 217410
rect 125580 217382 125916 217410
rect 126408 217382 126836 217410
rect 127236 217382 127572 217410
rect 128064 217382 128216 217410
rect 128984 217382 129320 217410
rect 129812 217382 130148 217410
rect 130640 217382 131068 217410
rect 131468 217382 131804 217410
rect 132296 217382 132356 217410
rect 133124 217382 133552 217410
rect 133952 217382 134288 217410
rect 134872 217382 135024 217410
rect 135700 217382 136036 217410
rect 136528 217382 136588 217410
rect 137356 217382 137784 217410
rect 138184 217382 138520 217410
rect 139012 217382 139256 217410
rect 139840 217382 140176 217410
rect 140760 217382 141096 217410
rect 141588 217382 141924 217410
rect 142416 217382 142752 217410
rect 143244 217382 143488 217410
rect 144072 217382 144408 217410
rect 144900 217382 145236 217410
rect 145728 217382 146156 217410
rect 146648 217382 146984 217410
rect 147476 217382 147628 217410
rect 148304 217382 148640 217410
rect 149132 217382 149468 217410
rect 149960 217382 150388 217410
rect 150788 217382 151124 217410
rect 151616 217382 151768 217410
rect 152536 217382 152964 217410
rect 153364 217382 153700 217410
rect 154192 217382 154528 217410
rect 155020 217382 155356 217410
rect 155788 217410 155816 224742
rect 155880 220386 155908 230114
rect 162860 229356 162912 229362
rect 162860 229298 162912 229304
rect 161296 227996 161348 228002
rect 161296 227938 161348 227944
rect 160376 227724 160428 227730
rect 160376 227666 160428 227672
rect 157064 227656 157116 227662
rect 157064 227598 157116 227604
rect 155868 220380 155920 220386
rect 155868 220322 155920 220328
rect 157076 217410 157104 227598
rect 159548 224868 159600 224874
rect 159548 224810 159600 224816
rect 157800 221264 157852 221270
rect 157800 221206 157852 221212
rect 157812 217410 157840 221206
rect 158628 219904 158680 219910
rect 158628 219846 158680 219852
rect 158640 217410 158668 219846
rect 159560 217410 159588 224810
rect 160388 217410 160416 227666
rect 161308 217410 161336 227938
rect 162872 226982 162900 229298
rect 162860 226976 162912 226982
rect 162860 226918 162912 226924
rect 163688 226976 163740 226982
rect 163688 226918 163740 226924
rect 162768 224936 162820 224942
rect 162768 224878 162820 224884
rect 162032 222692 162084 222698
rect 162032 222634 162084 222640
rect 162044 217410 162072 222634
rect 162780 217410 162808 224878
rect 163700 217410 163728 226918
rect 166908 226908 166960 226914
rect 166908 226850 166960 226856
rect 164608 226840 164660 226846
rect 164608 226782 164660 226788
rect 164620 217410 164648 226782
rect 166264 224188 166316 224194
rect 166264 224130 166316 224136
rect 165436 219836 165488 219842
rect 165436 219778 165488 219784
rect 165448 217410 165476 219778
rect 166276 217410 166304 224130
rect 166920 217410 166948 226850
rect 169576 224120 169628 224126
rect 169576 224062 169628 224068
rect 167920 221196 167972 221202
rect 167920 221138 167972 221144
rect 167932 217410 167960 221138
rect 168748 220380 168800 220386
rect 168748 220322 168800 220328
rect 168760 217410 168788 220322
rect 169588 217410 169616 224062
rect 169680 220386 169708 230250
rect 171048 227928 171100 227934
rect 171048 227870 171100 227876
rect 170496 225208 170548 225214
rect 170496 225150 170548 225156
rect 169668 220380 169720 220386
rect 169668 220322 169720 220328
rect 170508 217410 170536 225150
rect 171060 217410 171088 227870
rect 173808 226772 173860 226778
rect 173808 226714 173860 226720
rect 172980 224052 173032 224058
rect 172980 223994 173032 224000
rect 172152 219768 172204 219774
rect 172152 219710 172204 219716
rect 172164 217410 172192 219710
rect 172992 217410 173020 223994
rect 173820 217410 173848 226714
rect 174636 226704 174688 226710
rect 174636 226646 174688 226652
rect 174648 217410 174676 226646
rect 175200 217410 175228 230318
rect 177212 226636 177264 226642
rect 177212 226578 177264 226584
rect 176476 223984 176528 223990
rect 176476 223926 176528 223932
rect 176488 217410 176516 223926
rect 177224 217410 177252 226578
rect 177856 222760 177908 222766
rect 177856 222702 177908 222708
rect 177868 217410 177896 222702
rect 179340 220386 179368 230386
rect 186964 229424 187016 229430
rect 186964 229366 187016 229372
rect 180800 229288 180852 229294
rect 180800 229230 180852 229236
rect 180616 225140 180668 225146
rect 180616 225082 180668 225088
rect 179696 223916 179748 223922
rect 179696 223858 179748 223864
rect 178868 220380 178920 220386
rect 178868 220322 178920 220328
rect 179328 220380 179380 220386
rect 179328 220322 179380 220328
rect 178880 217410 178908 220322
rect 179708 217410 179736 223858
rect 180628 217410 180656 225082
rect 180812 222698 180840 229230
rect 183192 223848 183244 223854
rect 183192 223790 183244 223796
rect 180800 222692 180852 222698
rect 180800 222634 180852 222640
rect 181352 222692 181404 222698
rect 181352 222634 181404 222640
rect 181364 217410 181392 222634
rect 181996 219632 182048 219638
rect 181996 219574 182048 219580
rect 182008 217410 182036 219574
rect 183204 217410 183232 223790
rect 186228 223780 186280 223786
rect 186228 223722 186280 223728
rect 184756 222556 184808 222562
rect 184756 222498 184808 222504
rect 183928 221128 183980 221134
rect 183928 221070 183980 221076
rect 183940 217410 183968 221070
rect 184768 217410 184796 222498
rect 185584 219700 185636 219706
rect 185584 219642 185636 219648
rect 185596 217410 185624 219642
rect 186240 217410 186268 223722
rect 186976 219706 187004 229366
rect 192312 228410 192340 231676
rect 192404 231662 192602 231690
rect 192680 231662 192970 231690
rect 192300 228404 192352 228410
rect 192300 228346 192352 228352
rect 190276 226568 190328 226574
rect 190276 226510 190328 226516
rect 187332 222624 187384 222630
rect 187332 222566 187384 222572
rect 186964 219700 187016 219706
rect 186964 219642 187016 219648
rect 187344 217410 187372 222566
rect 188160 222488 188212 222494
rect 188160 222430 188212 222436
rect 188172 217410 188200 222430
rect 189816 221060 189868 221066
rect 189816 221002 189868 221008
rect 188896 219632 188948 219638
rect 188896 219574 188948 219580
rect 188908 217410 188936 219574
rect 189828 217410 189856 221002
rect 155788 217382 155848 217410
rect 156676 217382 157104 217410
rect 157504 217382 157840 217410
rect 158424 217382 158668 217410
rect 159252 217382 159588 217410
rect 160080 217382 160416 217410
rect 160908 217382 161336 217410
rect 161736 217382 162072 217410
rect 162564 217382 162808 217410
rect 163392 217382 163728 217410
rect 164312 217382 164648 217410
rect 165140 217382 165476 217410
rect 165968 217382 166304 217410
rect 166796 217382 166948 217410
rect 167624 217382 167960 217410
rect 168452 217382 168788 217410
rect 169280 217382 169616 217410
rect 170200 217382 170536 217410
rect 171028 217382 171088 217410
rect 171856 217382 172192 217410
rect 172684 217382 173020 217410
rect 173512 217382 173848 217410
rect 174340 217382 174676 217410
rect 175168 217382 175228 217410
rect 176088 217382 176516 217410
rect 176916 217382 177252 217410
rect 177744 217382 177896 217410
rect 178572 217382 178908 217410
rect 179400 217382 179736 217410
rect 180228 217382 180656 217410
rect 181056 217382 181392 217410
rect 181976 217382 182036 217410
rect 182804 217382 183232 217410
rect 183632 217382 183968 217410
rect 184460 217382 184796 217410
rect 185288 217382 185624 217410
rect 186116 217382 186268 217410
rect 186944 217382 187372 217410
rect 187864 217382 188200 217410
rect 188692 217382 188936 217410
rect 189520 217382 189856 217410
rect 190288 217410 190316 226510
rect 192404 222873 192432 231662
rect 192680 225622 192708 231662
rect 193324 228478 193352 231676
rect 193416 231662 193706 231690
rect 193312 228472 193364 228478
rect 193312 228414 193364 228420
rect 192668 225616 192720 225622
rect 192668 225558 192720 225564
rect 192852 225004 192904 225010
rect 192852 224946 192904 224952
rect 192390 222864 192446 222873
rect 192390 222799 192446 222808
rect 191564 222420 191616 222426
rect 191564 222362 191616 222368
rect 191576 217410 191604 222362
rect 192300 220380 192352 220386
rect 192300 220322 192352 220328
rect 192312 217410 192340 220322
rect 192864 220114 192892 224946
rect 193416 221513 193444 231662
rect 194060 223009 194088 231676
rect 194140 228404 194192 228410
rect 194140 228346 194192 228352
rect 194046 223000 194102 223009
rect 193956 222964 194008 222970
rect 194046 222935 194102 222944
rect 193956 222906 194008 222912
rect 193968 222290 193996 222906
rect 193956 222284 194008 222290
rect 193956 222226 194008 222232
rect 193402 221504 193458 221513
rect 193402 221439 193458 221448
rect 192944 220992 192996 220998
rect 192944 220934 192996 220940
rect 192852 220108 192904 220114
rect 192852 220050 192904 220056
rect 192956 217410 192984 220934
rect 194152 219434 194180 228346
rect 194428 225690 194456 231676
rect 194796 229809 194824 231676
rect 194888 231662 195178 231690
rect 194782 229800 194838 229809
rect 194782 229735 194838 229744
rect 194416 225684 194468 225690
rect 194416 225626 194468 225632
rect 194888 221474 194916 231662
rect 194968 228472 195020 228478
rect 194968 228414 195020 228420
rect 194876 221468 194928 221474
rect 194876 221410 194928 221416
rect 194980 219434 195008 228414
rect 195440 224233 195468 231676
rect 195808 226953 195836 231676
rect 196176 229945 196204 231676
rect 196268 231662 196558 231690
rect 196162 229936 196218 229945
rect 196162 229871 196218 229880
rect 195794 226944 195850 226953
rect 195794 226879 195850 226888
rect 195426 224224 195482 224233
rect 195426 224159 195482 224168
rect 196268 221542 196296 231662
rect 196622 230344 196678 230353
rect 196622 230279 196678 230288
rect 196532 222352 196584 222358
rect 196532 222294 196584 222300
rect 196256 221536 196308 221542
rect 196256 221478 196308 221484
rect 195152 220924 195204 220930
rect 195152 220866 195204 220872
rect 195164 219502 195192 220866
rect 195704 219564 195756 219570
rect 195704 219506 195756 219512
rect 195152 219496 195204 219502
rect 195152 219438 195204 219444
rect 194060 219406 194180 219434
rect 194888 219406 195008 219434
rect 194060 217410 194088 219406
rect 194888 217410 194916 219406
rect 195716 217410 195744 219506
rect 196544 217410 196572 222294
rect 196636 220153 196664 230279
rect 196912 222902 196940 231676
rect 197280 227089 197308 231676
rect 197266 227080 197322 227089
rect 197266 227015 197322 227024
rect 197648 225010 197676 231676
rect 197740 231662 198030 231690
rect 197636 225004 197688 225010
rect 197636 224946 197688 224952
rect 196900 222896 196952 222902
rect 196900 222838 196952 222844
rect 197740 221649 197768 231662
rect 198188 223032 198240 223038
rect 198188 222974 198240 222980
rect 197726 221640 197782 221649
rect 197726 221575 197782 221584
rect 197268 221536 197320 221542
rect 197268 221478 197320 221484
rect 196622 220144 196678 220153
rect 196622 220079 196678 220088
rect 197280 217410 197308 221478
rect 198200 217410 198228 222974
rect 198292 222290 198320 231676
rect 198384 231662 198674 231690
rect 198384 222970 198412 231662
rect 199028 230353 199056 231676
rect 199120 231662 199410 231690
rect 199014 230344 199070 230353
rect 199014 230279 199070 230288
rect 199016 225684 199068 225690
rect 199016 225626 199068 225632
rect 198372 222964 198424 222970
rect 198372 222906 198424 222912
rect 198280 222284 198332 222290
rect 198280 222226 198332 222232
rect 199028 217410 199056 225626
rect 199120 221785 199148 231662
rect 199764 224505 199792 231676
rect 199750 224496 199806 224505
rect 199750 224431 199806 224440
rect 200132 224369 200160 231676
rect 200500 229770 200528 231676
rect 200592 231662 200882 231690
rect 200488 229764 200540 229770
rect 200488 229706 200540 229712
rect 200118 224360 200174 224369
rect 200118 224295 200174 224304
rect 199936 222964 199988 222970
rect 199936 222906 199988 222912
rect 199106 221776 199162 221785
rect 199106 221711 199162 221720
rect 199948 217410 199976 222906
rect 200592 221921 200620 231662
rect 200672 229764 200724 229770
rect 200672 229706 200724 229712
rect 200684 225690 200712 229706
rect 200672 225684 200724 225690
rect 200672 225626 200724 225632
rect 201144 223106 201172 231676
rect 201512 227225 201540 231676
rect 201604 231662 201894 231690
rect 201972 231662 202262 231690
rect 201498 227216 201554 227225
rect 201498 227151 201554 227160
rect 201408 225616 201460 225622
rect 201408 225558 201460 225564
rect 201132 223100 201184 223106
rect 201132 223042 201184 223048
rect 200764 222896 200816 222902
rect 200764 222838 200816 222844
rect 200578 221912 200634 221921
rect 200578 221847 200634 221856
rect 200776 217410 200804 222838
rect 201420 217410 201448 225558
rect 201604 220289 201632 231662
rect 201972 221610 202000 231662
rect 202616 224641 202644 231676
rect 202984 225758 203012 231676
rect 203352 229838 203380 231676
rect 203444 231662 203734 231690
rect 203340 229832 203392 229838
rect 203340 229774 203392 229780
rect 202972 225752 203024 225758
rect 202972 225694 203024 225700
rect 203248 225684 203300 225690
rect 203248 225626 203300 225632
rect 202602 224632 202658 224641
rect 202602 224567 202658 224576
rect 201960 221604 202012 221610
rect 201960 221546 202012 221552
rect 202420 221604 202472 221610
rect 202420 221546 202472 221552
rect 201590 220280 201646 220289
rect 202432 220250 202460 221546
rect 201590 220215 201646 220224
rect 202420 220244 202472 220250
rect 202420 220186 202472 220192
rect 202420 219496 202472 219502
rect 202420 219438 202472 219444
rect 202432 217410 202460 219438
rect 203260 217410 203288 225626
rect 203444 221678 203472 231662
rect 203524 229832 203576 229838
rect 203524 229774 203576 229780
rect 203432 221672 203484 221678
rect 203432 221614 203484 221620
rect 203536 220182 203564 229774
rect 203996 223174 204024 231676
rect 203984 223168 204036 223174
rect 203984 223110 204036 223116
rect 204364 222018 204392 231676
rect 204732 229838 204760 231676
rect 204824 231662 205114 231690
rect 205192 231662 205482 231690
rect 204720 229832 204772 229838
rect 204720 229774 204772 229780
rect 204352 222012 204404 222018
rect 204352 221954 204404 221960
rect 204824 221746 204852 231662
rect 204904 223100 204956 223106
rect 204904 223042 204956 223048
rect 204812 221740 204864 221746
rect 204812 221682 204864 221688
rect 204168 221672 204220 221678
rect 204168 221614 204220 221620
rect 204180 220318 204208 221614
rect 204168 220312 204220 220318
rect 204168 220254 204220 220260
rect 203524 220176 203576 220182
rect 203524 220118 203576 220124
rect 204076 220176 204128 220182
rect 204076 220118 204128 220124
rect 204088 217410 204116 220118
rect 204916 217410 204944 223042
rect 205192 221814 205220 231662
rect 205836 229702 205864 231676
rect 206204 229906 206232 231676
rect 206192 229900 206244 229906
rect 206192 229842 206244 229848
rect 205824 229696 205876 229702
rect 205824 229638 205876 229644
rect 206572 228313 206600 231676
rect 206664 231662 206862 231690
rect 206558 228304 206614 228313
rect 206558 228239 206614 228248
rect 205548 221876 205600 221882
rect 205548 221818 205600 221824
rect 205180 221808 205232 221814
rect 205180 221750 205232 221756
rect 205560 217410 205588 221818
rect 206664 221746 206692 231662
rect 206744 229832 206796 229838
rect 206744 229774 206796 229780
rect 206756 221882 206784 229774
rect 207216 225826 207244 231676
rect 207204 225820 207256 225826
rect 207204 225762 207256 225768
rect 206836 225752 206888 225758
rect 206836 225694 206888 225700
rect 206744 221876 206796 221882
rect 206744 221818 206796 221824
rect 206652 221740 206704 221746
rect 206652 221682 206704 221688
rect 206192 220516 206244 220522
rect 206192 220458 206244 220464
rect 206204 220250 206232 220458
rect 206192 220244 206244 220250
rect 206192 220186 206244 220192
rect 206848 217410 206876 225694
rect 207584 224262 207612 231676
rect 207952 228449 207980 231676
rect 208044 231662 208334 231690
rect 207938 228440 207994 228449
rect 207938 228375 207994 228384
rect 207572 224256 207624 224262
rect 207572 224198 207624 224204
rect 208044 223145 208072 231662
rect 208308 225820 208360 225826
rect 208308 225762 208360 225768
rect 208030 223136 208086 223145
rect 208030 223071 208086 223080
rect 206928 221808 206980 221814
rect 206928 221750 206980 221756
rect 206940 220454 206968 221750
rect 208216 221740 208268 221746
rect 208216 221682 208268 221688
rect 208228 220522 208256 221682
rect 208216 220516 208268 220522
rect 208216 220458 208268 220464
rect 206928 220448 206980 220454
rect 206928 220390 206980 220396
rect 207480 220312 207532 220318
rect 207480 220254 207532 220260
rect 207492 217410 207520 220254
rect 208320 217410 208348 225762
rect 208688 225593 208716 231676
rect 209056 229498 209084 231676
rect 209044 229492 209096 229498
rect 209044 229434 209096 229440
rect 209424 228546 209452 231676
rect 209412 228540 209464 228546
rect 209412 228482 209464 228488
rect 208674 225584 208730 225593
rect 208674 225519 208730 225528
rect 209596 223372 209648 223378
rect 209596 223314 209648 223320
rect 209608 223174 209636 223314
rect 209700 223242 209728 231676
rect 209872 228540 209924 228546
rect 209872 228482 209924 228488
rect 209688 223236 209740 223242
rect 209688 223178 209740 223184
rect 209596 223168 209648 223174
rect 209596 223110 209648 223116
rect 209688 221468 209740 221474
rect 209688 221410 209740 221416
rect 209136 220108 209188 220114
rect 209136 220050 209188 220056
rect 209148 217410 209176 220050
rect 209700 217410 209728 221410
rect 209884 220182 209912 228482
rect 210068 225729 210096 231676
rect 210160 231662 210450 231690
rect 210054 225720 210110 225729
rect 210054 225655 210110 225664
rect 210160 221610 210188 231662
rect 210804 228614 210832 231676
rect 210792 228608 210844 228614
rect 210792 228550 210844 228556
rect 211172 223281 211200 231676
rect 211540 225894 211568 231676
rect 211632 231662 211922 231690
rect 211528 225888 211580 225894
rect 211528 225830 211580 225836
rect 211158 223272 211214 223281
rect 211158 223207 211214 223216
rect 210148 221604 210200 221610
rect 210148 221546 210200 221552
rect 211632 220930 211660 231662
rect 212276 228682 212304 231676
rect 212448 229900 212500 229906
rect 212448 229842 212500 229848
rect 212264 228676 212316 228682
rect 212264 228618 212316 228624
rect 211712 225888 211764 225894
rect 211712 225830 211764 225836
rect 211620 220924 211672 220930
rect 211620 220866 211672 220872
rect 209872 220176 209924 220182
rect 209872 220118 209924 220124
rect 210792 220176 210844 220182
rect 210792 220118 210844 220124
rect 210804 217410 210832 220118
rect 211724 217410 211752 225830
rect 212460 217410 212488 229842
rect 212552 223242 212580 231676
rect 212920 225962 212948 231676
rect 213288 230246 213316 231676
rect 213276 230240 213328 230246
rect 213276 230182 213328 230188
rect 213656 228750 213684 231676
rect 213644 228744 213696 228750
rect 213644 228686 213696 228692
rect 213828 228608 213880 228614
rect 213828 228550 213880 228556
rect 212908 225956 212960 225962
rect 212908 225898 212960 225904
rect 212540 223236 212592 223242
rect 212540 223178 212592 223184
rect 213368 221604 213420 221610
rect 213368 221546 213420 221552
rect 213380 217410 213408 221546
rect 213840 220318 213868 228550
rect 213920 223508 213972 223514
rect 213920 223450 213972 223456
rect 213828 220312 213880 220318
rect 213828 220254 213880 220260
rect 213932 220250 213960 223450
rect 214024 223174 214052 231676
rect 214392 226030 214420 231676
rect 214484 231662 214774 231690
rect 214380 226024 214432 226030
rect 214380 225966 214432 225972
rect 214012 223168 214064 223174
rect 214012 223110 214064 223116
rect 214484 221678 214512 231662
rect 215128 228818 215156 231676
rect 215116 228812 215168 228818
rect 215116 228754 215168 228760
rect 215116 228676 215168 228682
rect 215116 228618 215168 228624
rect 214472 221672 214524 221678
rect 214472 221614 214524 221620
rect 214196 220720 214248 220726
rect 214196 220662 214248 220668
rect 213920 220244 213972 220250
rect 213920 220186 213972 220192
rect 214208 217410 214236 220662
rect 215128 217410 215156 228618
rect 215300 225956 215352 225962
rect 215300 225898 215352 225904
rect 215312 220726 215340 225898
rect 215404 223310 215432 231676
rect 215772 226098 215800 231676
rect 216140 229566 216168 231676
rect 216128 229560 216180 229566
rect 216128 229502 216180 229508
rect 216508 228886 216536 231676
rect 216496 228880 216548 228886
rect 216496 228822 216548 228828
rect 216680 228812 216732 228818
rect 216680 228754 216732 228760
rect 215760 226092 215812 226098
rect 215760 226034 215812 226040
rect 215392 223304 215444 223310
rect 215392 223246 215444 223252
rect 216588 221672 216640 221678
rect 216588 221614 216640 221620
rect 215300 220720 215352 220726
rect 215300 220662 215352 220668
rect 215852 220244 215904 220250
rect 215852 220186 215904 220192
rect 215864 217410 215892 220186
rect 216600 217410 216628 221614
rect 216692 220590 216720 228754
rect 216876 221950 216904 231676
rect 217244 226166 217272 231676
rect 217336 231662 217626 231690
rect 217232 226160 217284 226166
rect 217232 226102 217284 226108
rect 216864 221944 216916 221950
rect 216864 221886 216916 221892
rect 217336 221814 217364 231662
rect 217980 228954 218008 231676
rect 217968 228948 218020 228954
rect 217968 228890 218020 228896
rect 218060 226160 218112 226166
rect 218060 226102 218112 226108
rect 217324 221808 217376 221814
rect 217324 221750 217376 221756
rect 218072 220658 218100 226102
rect 218256 223378 218284 231676
rect 218624 226234 218652 231676
rect 218992 229634 219020 231676
rect 219256 230240 219308 230246
rect 219256 230182 219308 230188
rect 218980 229628 219032 229634
rect 218980 229570 219032 229576
rect 218612 226228 218664 226234
rect 218612 226170 218664 226176
rect 218244 223372 218296 223378
rect 218244 223314 218296 223320
rect 218428 221808 218480 221814
rect 218428 221750 218480 221756
rect 218060 220652 218112 220658
rect 218060 220594 218112 220600
rect 216680 220584 216732 220590
rect 216680 220526 216732 220532
rect 217600 220312 217652 220318
rect 217600 220254 217652 220260
rect 217612 217410 217640 220254
rect 218440 217410 218468 221750
rect 219268 217410 219296 230182
rect 219360 229022 219388 231676
rect 219636 231662 219742 231690
rect 219348 229016 219400 229022
rect 219348 228958 219400 228964
rect 219636 222086 219664 231662
rect 220096 226302 220124 231676
rect 220188 231662 220478 231690
rect 220084 226296 220136 226302
rect 220084 226238 220136 226244
rect 219624 222080 219676 222086
rect 219624 222022 219676 222028
rect 220084 221876 220136 221882
rect 220084 221818 220136 221824
rect 220096 217410 220124 221818
rect 220188 221746 220216 231662
rect 220832 229090 220860 231676
rect 221016 231662 221122 231690
rect 221200 231662 221490 231690
rect 220820 229084 220872 229090
rect 220820 229026 220872 229032
rect 220636 226024 220688 226030
rect 220636 225966 220688 225972
rect 220176 221740 220228 221746
rect 220176 221682 220228 221688
rect 220648 217410 220676 225966
rect 221016 222154 221044 231662
rect 221200 225554 221228 231662
rect 221188 225548 221240 225554
rect 221188 225490 221240 225496
rect 221844 223514 221872 231676
rect 222108 228744 222160 228750
rect 222108 228686 222160 228692
rect 221832 223508 221884 223514
rect 221832 223450 221884 223456
rect 221004 222148 221056 222154
rect 221004 222090 221056 222096
rect 221740 221740 221792 221746
rect 221740 221682 221792 221688
rect 221752 217410 221780 221682
rect 222120 220794 222148 228686
rect 222212 227050 222240 231676
rect 222200 227044 222252 227050
rect 222200 226986 222252 226992
rect 222580 223582 222608 231676
rect 222948 225486 222976 231676
rect 223316 229362 223344 231676
rect 223304 229356 223356 229362
rect 223304 229298 223356 229304
rect 223684 228342 223712 231676
rect 223776 231662 223974 231690
rect 223672 228336 223724 228342
rect 223672 228278 223724 228284
rect 223120 226228 223172 226234
rect 223120 226170 223172 226176
rect 222936 225480 222988 225486
rect 222936 225422 222988 225428
rect 222568 223576 222620 223582
rect 222568 223518 222620 223524
rect 222108 220788 222160 220794
rect 222108 220730 222160 220736
rect 222568 220448 222620 220454
rect 222568 220390 222620 220396
rect 222580 217410 222608 220390
rect 223132 220046 223160 226170
rect 223488 222012 223540 222018
rect 223488 221954 223540 221960
rect 223120 220040 223172 220046
rect 223120 219982 223172 219988
rect 223500 217410 223528 221954
rect 223776 221406 223804 231662
rect 224040 228948 224092 228954
rect 224040 228890 224092 228896
rect 223764 221400 223816 221406
rect 223764 221342 223816 221348
rect 224052 219978 224080 228890
rect 224328 225418 224356 231676
rect 224696 228818 224724 231676
rect 224684 228812 224736 228818
rect 224684 228754 224736 228760
rect 225064 228274 225092 231676
rect 225052 228268 225104 228274
rect 225052 228210 225104 228216
rect 224960 226092 225012 226098
rect 224960 226034 225012 226040
rect 224316 225412 224368 225418
rect 224316 225354 224368 225360
rect 224868 221944 224920 221950
rect 224868 221886 224920 221892
rect 224316 220380 224368 220386
rect 224316 220322 224368 220328
rect 224040 219972 224092 219978
rect 224040 219914 224092 219920
rect 224328 217410 224356 220322
rect 224880 217410 224908 221886
rect 224972 220522 225000 226034
rect 225432 222834 225460 231676
rect 225800 225350 225828 231676
rect 226168 229974 226196 231676
rect 226156 229968 226208 229974
rect 226156 229910 226208 229916
rect 226248 229968 226300 229974
rect 226248 229910 226300 229916
rect 225788 225344 225840 225350
rect 225788 225286 225840 225292
rect 225420 222828 225472 222834
rect 225420 222770 225472 222776
rect 224960 220516 225012 220522
rect 224960 220458 225012 220464
rect 226260 219434 226288 229910
rect 226536 227118 226564 231676
rect 226524 227112 226576 227118
rect 226524 227054 226576 227060
rect 226812 224398 226840 231676
rect 227180 225282 227208 231676
rect 227272 231662 227562 231690
rect 227272 226166 227300 231662
rect 227536 229696 227588 229702
rect 227536 229638 227588 229644
rect 227260 226160 227312 226166
rect 227260 226102 227312 226108
rect 227352 226160 227404 226166
rect 227352 226102 227404 226108
rect 227168 225276 227220 225282
rect 227168 225218 227220 225224
rect 226800 224392 226852 224398
rect 226800 224334 226852 224340
rect 226800 222080 226852 222086
rect 226800 222022 226852 222028
rect 226076 219406 226288 219434
rect 226076 217410 226104 219406
rect 226812 217410 226840 222022
rect 227364 219910 227392 226102
rect 227352 219904 227404 219910
rect 227352 219846 227404 219852
rect 227548 217410 227576 229638
rect 227720 228880 227772 228886
rect 227720 228822 227772 228828
rect 227732 219842 227760 228822
rect 227916 228206 227944 231676
rect 227904 228200 227956 228206
rect 227904 228142 227956 228148
rect 228284 224466 228312 231676
rect 228272 224460 228324 224466
rect 228272 224402 228324 224408
rect 228652 224330 228680 231676
rect 229020 230042 229048 231676
rect 229008 230036 229060 230042
rect 229008 229978 229060 229984
rect 229388 227254 229416 231676
rect 229376 227248 229428 227254
rect 229376 227190 229428 227196
rect 229664 224534 229692 231676
rect 230032 227186 230060 231676
rect 230296 228812 230348 228818
rect 230296 228754 230348 228760
rect 230020 227180 230072 227186
rect 230020 227122 230072 227128
rect 229652 224528 229704 224534
rect 229652 224470 229704 224476
rect 228640 224324 228692 224330
rect 228640 224266 228692 224272
rect 228456 222148 228508 222154
rect 228456 222090 228508 222096
rect 227720 219836 227772 219842
rect 227720 219778 227772 219784
rect 228468 217410 228496 222090
rect 229376 220584 229428 220590
rect 229376 220526 229428 220532
rect 229388 217410 229416 220526
rect 230308 217410 230336 228754
rect 230400 228750 230428 231676
rect 230388 228744 230440 228750
rect 230388 228686 230440 228692
rect 230768 228138 230796 231676
rect 230756 228132 230808 228138
rect 230756 228074 230808 228080
rect 231136 224602 231164 231676
rect 231504 227322 231532 231676
rect 231872 230110 231900 231676
rect 231860 230104 231912 230110
rect 231860 230046 231912 230052
rect 232240 227458 232268 231676
rect 232332 231662 232530 231690
rect 232228 227452 232280 227458
rect 232228 227394 232280 227400
rect 231492 227316 231544 227322
rect 231492 227258 231544 227264
rect 232332 224670 232360 231662
rect 232884 227390 232912 231676
rect 233148 230104 233200 230110
rect 233148 230046 233200 230052
rect 232872 227384 232924 227390
rect 232872 227326 232924 227332
rect 232780 227248 232832 227254
rect 232780 227190 232832 227196
rect 232320 224664 232372 224670
rect 232320 224606 232372 224612
rect 231124 224596 231176 224602
rect 231124 224538 231176 224544
rect 232412 224324 232464 224330
rect 232412 224266 232464 224272
rect 231676 221400 231728 221406
rect 231676 221342 231728 221348
rect 231032 220516 231084 220522
rect 231032 220458 231084 220464
rect 231044 217410 231072 220458
rect 231688 217410 231716 221342
rect 232424 219774 232452 224266
rect 232688 220788 232740 220794
rect 232688 220730 232740 220736
rect 232412 219768 232464 219774
rect 232412 219710 232464 219716
rect 232700 217410 232728 220730
rect 232792 219706 232820 227190
rect 233160 220794 233188 230046
rect 233252 226234 233280 231676
rect 233528 231662 233634 231690
rect 233528 229094 233556 231662
rect 233436 229066 233556 229094
rect 233240 226228 233292 226234
rect 233240 226170 233292 226176
rect 233436 221338 233464 229066
rect 233516 228812 233568 228818
rect 233516 228754 233568 228760
rect 233424 221332 233476 221338
rect 233424 221274 233476 221280
rect 233148 220788 233200 220794
rect 233148 220730 233200 220736
rect 232780 219700 232832 219706
rect 232780 219642 232832 219648
rect 233528 217410 233556 228754
rect 233988 224738 234016 231676
rect 234356 227526 234384 231676
rect 234528 230036 234580 230042
rect 234528 229978 234580 229984
rect 234344 227520 234396 227526
rect 234344 227462 234396 227468
rect 233976 224732 234028 224738
rect 233976 224674 234028 224680
rect 234540 219434 234568 229978
rect 234724 228954 234752 231676
rect 234712 228948 234764 228954
rect 234712 228890 234764 228896
rect 235092 228070 235120 231676
rect 235080 228064 235132 228070
rect 235080 228006 235132 228012
rect 234712 227112 234764 227118
rect 234712 227054 234764 227060
rect 234620 224460 234672 224466
rect 234620 224402 234672 224408
rect 234632 219638 234660 224402
rect 234620 219632 234672 219638
rect 234620 219574 234672 219580
rect 234724 219570 234752 227054
rect 235368 224806 235396 231676
rect 235736 227594 235764 231676
rect 236104 230178 236132 231676
rect 236196 231662 236486 231690
rect 236092 230172 236144 230178
rect 236092 230114 236144 230120
rect 235724 227588 235776 227594
rect 235724 227530 235776 227536
rect 235356 224800 235408 224806
rect 235356 224742 235408 224748
rect 235264 221332 235316 221338
rect 235264 221274 235316 221280
rect 234712 219564 234764 219570
rect 234712 219506 234764 219512
rect 234448 219406 234568 219434
rect 234448 217410 234476 219406
rect 235276 217410 235304 221274
rect 236196 221270 236224 231662
rect 236840 224874 236868 231676
rect 237208 227662 237236 231676
rect 237196 227656 237248 227662
rect 237196 227598 237248 227604
rect 237380 227180 237432 227186
rect 237380 227122 237432 227128
rect 237012 227044 237064 227050
rect 237012 226986 237064 226992
rect 236828 224868 236880 224874
rect 236828 224810 236880 224816
rect 236184 221264 236236 221270
rect 236184 221206 236236 221212
rect 235908 220652 235960 220658
rect 235908 220594 235960 220600
rect 235920 217410 235948 220594
rect 237024 217410 237052 226986
rect 237392 219502 237420 227122
rect 237576 226166 237604 231676
rect 237944 228002 237972 231676
rect 237932 227996 237984 228002
rect 237932 227938 237984 227944
rect 237564 226160 237616 226166
rect 237564 226102 237616 226108
rect 238220 224942 238248 231676
rect 238588 227730 238616 231676
rect 238956 229294 238984 231676
rect 238944 229288 238996 229294
rect 238944 229230 238996 229236
rect 238576 227724 238628 227730
rect 238576 227666 238628 227672
rect 239324 226846 239352 231676
rect 239312 226840 239364 226846
rect 239312 226782 239364 226788
rect 238208 224936 238260 224942
rect 238208 224878 238260 224884
rect 239692 224194 239720 231676
rect 239784 231662 240074 231690
rect 239784 226982 239812 231662
rect 240048 230172 240100 230178
rect 240048 230114 240100 230120
rect 239772 226976 239824 226982
rect 239772 226918 239824 226924
rect 239956 224256 240008 224262
rect 239956 224198 240008 224204
rect 239680 224188 239732 224194
rect 239680 224130 239732 224136
rect 238576 221264 238628 221270
rect 238576 221206 238628 221212
rect 237748 220720 237800 220726
rect 237748 220662 237800 220668
rect 237380 219496 237432 219502
rect 237380 219438 237432 219444
rect 237760 217410 237788 220662
rect 238588 217410 238616 221206
rect 239404 220788 239456 220794
rect 239404 220730 239456 220736
rect 239416 217410 239444 220730
rect 239968 217410 239996 224198
rect 240060 220794 240088 230114
rect 240428 228886 240456 231676
rect 240520 231662 240810 231690
rect 240416 228880 240468 228886
rect 240416 228822 240468 228828
rect 240520 221202 240548 231662
rect 241072 224126 241100 231676
rect 241440 226914 241468 231676
rect 241808 230314 241836 231676
rect 241796 230308 241848 230314
rect 241796 230250 241848 230256
rect 242176 227934 242204 231676
rect 242164 227928 242216 227934
rect 242164 227870 242216 227876
rect 241428 226908 241480 226914
rect 241428 226850 241480 226856
rect 241060 224120 241112 224126
rect 241060 224062 241112 224068
rect 242544 224058 242572 231676
rect 242912 225214 242940 231676
rect 242900 225208 242952 225214
rect 242900 225150 242952 225156
rect 243280 224330 243308 231676
rect 243648 226710 243676 231676
rect 243636 226704 243688 226710
rect 243636 226646 243688 226652
rect 243268 224324 243320 224330
rect 243268 224266 243320 224272
rect 243636 224324 243688 224330
rect 243636 224266 243688 224272
rect 242532 224052 242584 224058
rect 242532 223994 242584 224000
rect 240508 221196 240560 221202
rect 240508 221138 240560 221144
rect 241980 221196 242032 221202
rect 241980 221138 242032 221144
rect 240048 220788 240100 220794
rect 240048 220730 240100 220736
rect 241152 220788 241204 220794
rect 241152 220730 241204 220736
rect 241164 217410 241192 220730
rect 241992 217410 242020 221138
rect 242808 219904 242860 219910
rect 242808 219846 242860 219852
rect 242820 217410 242848 219846
rect 243648 217410 243676 224266
rect 243924 223990 243952 231676
rect 244188 230308 244240 230314
rect 244188 230250 244240 230256
rect 243912 223984 243964 223990
rect 243912 223926 243964 223932
rect 244200 217410 244228 230250
rect 244292 226778 244320 231676
rect 244660 230382 244688 231676
rect 244648 230376 244700 230382
rect 244648 230318 244700 230324
rect 244924 229560 244976 229566
rect 244924 229502 244976 229508
rect 244280 226772 244332 226778
rect 244280 226714 244332 226720
rect 244936 221542 244964 229502
rect 245028 222766 245056 231676
rect 245396 223922 245424 231676
rect 245764 226642 245792 231676
rect 246132 230450 246160 231676
rect 246120 230444 246172 230450
rect 246120 230386 246172 230392
rect 245752 226636 245804 226642
rect 245752 226578 245804 226584
rect 245384 223916 245436 223922
rect 245384 223858 245436 223864
rect 245016 222760 245068 222766
rect 245016 222702 245068 222708
rect 246500 222698 246528 231676
rect 246776 223854 246804 231676
rect 246948 230376 247000 230382
rect 246948 230318 247000 230324
rect 246856 224392 246908 224398
rect 246856 224334 246908 224340
rect 246764 223848 246816 223854
rect 246764 223790 246816 223796
rect 246488 222692 246540 222698
rect 246488 222634 246540 222640
rect 244924 221536 244976 221542
rect 244924 221478 244976 221484
rect 245292 221536 245344 221542
rect 245292 221478 245344 221484
rect 245304 217410 245332 221478
rect 246120 219972 246172 219978
rect 246120 219914 246172 219920
rect 246132 217410 246160 219914
rect 246868 217410 246896 224334
rect 246960 219978 246988 230318
rect 247144 225146 247172 231676
rect 247512 227254 247540 231676
rect 247500 227248 247552 227254
rect 247500 227190 247552 227196
rect 247132 225140 247184 225146
rect 247132 225082 247184 225088
rect 247880 222562 247908 231676
rect 248248 223786 248276 231676
rect 248630 231662 248736 231690
rect 248328 229628 248380 229634
rect 248328 229570 248380 229576
rect 248236 223780 248288 223786
rect 248236 223722 248288 223728
rect 247868 222556 247920 222562
rect 247868 222498 247920 222504
rect 248340 220046 248368 229570
rect 248708 229094 248736 231662
rect 248984 229430 249012 231676
rect 248972 229424 249024 229430
rect 248972 229366 249024 229372
rect 248616 229066 248736 229094
rect 248616 221134 248644 229066
rect 249352 222494 249380 231676
rect 249444 231662 249642 231690
rect 249340 222488 249392 222494
rect 249340 222430 249392 222436
rect 248604 221128 248656 221134
rect 248604 221070 248656 221076
rect 248696 221128 248748 221134
rect 248696 221070 248748 221076
rect 247868 220040 247920 220046
rect 247868 219982 247920 219988
rect 248328 220040 248380 220046
rect 248328 219982 248380 219988
rect 246948 219972 247000 219978
rect 246948 219914 247000 219920
rect 247880 217410 247908 219982
rect 248708 217410 248736 221070
rect 249444 221066 249472 231662
rect 249996 222630 250024 231676
rect 250364 224466 250392 231676
rect 250352 224460 250404 224466
rect 250352 224402 250404 224408
rect 250352 223168 250404 223174
rect 250352 223110 250404 223116
rect 249984 222624 250036 222630
rect 249984 222566 250036 222572
rect 249432 221060 249484 221066
rect 249432 221002 249484 221008
rect 249524 219904 249576 219910
rect 249524 219846 249576 219852
rect 249536 217410 249564 219846
rect 250364 217410 250392 223110
rect 250732 222426 250760 231676
rect 250824 231662 251114 231690
rect 250720 222420 250772 222426
rect 250720 222362 250772 222368
rect 250824 220998 250852 231662
rect 251468 226574 251496 231676
rect 251456 226568 251508 226574
rect 251456 226510 251508 226516
rect 251836 226098 251864 231676
rect 252204 228478 252232 231676
rect 252296 231662 252494 231690
rect 252192 228472 252244 228478
rect 252192 228414 252244 228420
rect 252008 228336 252060 228342
rect 252008 228278 252060 228284
rect 251824 226092 251876 226098
rect 251824 226034 251876 226040
rect 250812 220992 250864 220998
rect 250812 220934 250864 220940
rect 250996 219768 251048 219774
rect 250996 219710 251048 219716
rect 251008 217410 251036 219710
rect 252020 217410 252048 228278
rect 252296 222358 252324 231662
rect 252848 228410 252876 231676
rect 252836 228404 252888 228410
rect 252836 228346 252888 228352
rect 253216 227118 253244 231676
rect 253204 227112 253256 227118
rect 253204 227054 253256 227060
rect 253584 223038 253612 231676
rect 253848 226092 253900 226098
rect 253848 226034 253900 226040
rect 253572 223032 253624 223038
rect 253572 222974 253624 222980
rect 252284 222352 252336 222358
rect 252284 222294 252336 222300
rect 252100 220108 252152 220114
rect 252100 220050 252152 220056
rect 252112 219706 252140 220050
rect 252928 219904 252980 219910
rect 252928 219846 252980 219852
rect 252100 219700 252152 219706
rect 252100 219642 252152 219648
rect 252940 217410 252968 219846
rect 253860 217410 253888 226034
rect 253952 222970 253980 231676
rect 254320 229566 254348 231676
rect 254688 229770 254716 231676
rect 254676 229764 254728 229770
rect 254676 229706 254728 229712
rect 254308 229560 254360 229566
rect 254308 229502 254360 229508
rect 255056 225622 255084 231676
rect 255228 229764 255280 229770
rect 255228 229706 255280 229712
rect 255136 227112 255188 227118
rect 255136 227054 255188 227060
rect 255044 225616 255096 225622
rect 255044 225558 255096 225564
rect 253940 222964 253992 222970
rect 253940 222906 253992 222912
rect 254584 220176 254636 220182
rect 254584 220118 254636 220124
rect 254596 217410 254624 220118
rect 255148 217410 255176 227054
rect 255240 220182 255268 229706
rect 255332 225690 255360 231676
rect 255320 225684 255372 225690
rect 255320 225626 255372 225632
rect 255700 222902 255728 231676
rect 255964 229220 256016 229226
rect 255964 229162 256016 229168
rect 255688 222896 255740 222902
rect 255688 222838 255740 222844
rect 255228 220176 255280 220182
rect 255228 220118 255280 220124
rect 255976 220114 256004 229162
rect 256068 227186 256096 231676
rect 256056 227180 256108 227186
rect 256056 227122 256108 227128
rect 256436 223106 256464 231676
rect 256804 225758 256832 231676
rect 257172 228546 257200 231676
rect 257540 229838 257568 231676
rect 257528 229832 257580 229838
rect 257528 229774 257580 229780
rect 257344 229152 257396 229158
rect 257344 229094 257396 229100
rect 257160 228540 257212 228546
rect 257160 228482 257212 228488
rect 256792 225752 256844 225758
rect 256792 225694 256844 225700
rect 257068 225616 257120 225622
rect 257068 225558 257120 225564
rect 256424 223100 256476 223106
rect 256424 223042 256476 223048
rect 255964 220108 256016 220114
rect 255964 220050 256016 220056
rect 256240 219836 256292 219842
rect 256240 219778 256292 219784
rect 256252 217410 256280 219778
rect 257080 217410 257108 225558
rect 257356 219706 257384 229094
rect 257908 225826 257936 231676
rect 258198 231662 258304 231690
rect 257896 225820 257948 225826
rect 257896 225762 257948 225768
rect 258276 221474 258304 231662
rect 258552 228614 258580 231676
rect 258920 229158 258948 231676
rect 259012 231662 259302 231690
rect 258908 229152 258960 229158
rect 258908 229094 258960 229100
rect 258540 228608 258592 228614
rect 258540 228550 258592 228556
rect 258816 227180 258868 227186
rect 258816 227122 258868 227128
rect 258264 221468 258316 221474
rect 258264 221410 258316 221416
rect 257896 220176 257948 220182
rect 257896 220118 257948 220124
rect 257344 219700 257396 219706
rect 257344 219642 257396 219648
rect 257908 217410 257936 220118
rect 258828 217410 258856 227122
rect 259012 225894 259040 231662
rect 259368 229832 259420 229838
rect 259368 229774 259420 229780
rect 259000 225888 259052 225894
rect 259000 225830 259052 225836
rect 259380 217410 259408 229774
rect 259656 221610 259684 231676
rect 259920 229968 259972 229974
rect 259920 229910 259972 229916
rect 259932 229702 259960 229910
rect 259920 229696 259972 229702
rect 259920 229638 259972 229644
rect 260024 229226 260052 231676
rect 260104 229968 260156 229974
rect 260104 229910 260156 229916
rect 260012 229220 260064 229226
rect 260012 229162 260064 229168
rect 259644 221604 259696 221610
rect 259644 221546 259696 221552
rect 260116 220318 260144 229910
rect 260392 229906 260420 231676
rect 260380 229900 260432 229906
rect 260380 229842 260432 229848
rect 260760 228682 260788 231676
rect 260748 228676 260800 228682
rect 260748 228618 260800 228624
rect 260564 228404 260616 228410
rect 260564 228346 260616 228352
rect 260104 220312 260156 220318
rect 260104 220254 260156 220260
rect 260576 217410 260604 228346
rect 261036 221678 261064 231676
rect 261404 225962 261432 231676
rect 261496 231662 261786 231690
rect 261864 231662 262154 231690
rect 262324 231662 262522 231690
rect 261392 225956 261444 225962
rect 261392 225898 261444 225904
rect 261024 221672 261076 221678
rect 261024 221614 261076 221620
rect 261496 220250 261524 231662
rect 261864 221814 261892 231662
rect 262220 230444 262272 230450
rect 262220 230386 262272 230392
rect 262232 230246 262260 230386
rect 262220 230240 262272 230246
rect 262220 230182 262272 230188
rect 262128 222896 262180 222902
rect 262128 222838 262180 222844
rect 261852 221808 261904 221814
rect 261852 221750 261904 221756
rect 261484 220244 261536 220250
rect 261484 220186 261536 220192
rect 261300 219700 261352 219706
rect 261300 219642 261352 219648
rect 261312 217410 261340 219642
rect 262140 217410 262168 222838
rect 262324 221882 262352 231662
rect 262772 230240 262824 230246
rect 262772 230182 262824 230188
rect 262784 230042 262812 230182
rect 262772 230036 262824 230042
rect 262772 229978 262824 229984
rect 262876 229974 262904 231676
rect 263244 230450 263272 231676
rect 263612 230450 263640 231676
rect 263232 230444 263284 230450
rect 263232 230386 263284 230392
rect 263600 230444 263652 230450
rect 263600 230386 263652 230392
rect 262864 229968 262916 229974
rect 262864 229910 262916 229916
rect 263508 229900 263560 229906
rect 263508 229842 263560 229848
rect 263416 225684 263468 225690
rect 263416 225626 263468 225632
rect 262312 221876 262364 221882
rect 262312 221818 262364 221824
rect 262588 220584 262640 220590
rect 262588 220526 262640 220532
rect 262956 220584 263008 220590
rect 262956 220526 263008 220532
rect 262600 220250 262628 220526
rect 262588 220244 262640 220250
rect 262588 220186 262640 220192
rect 262968 217410 262996 220526
rect 190288 217382 190348 217410
rect 191176 217382 191604 217410
rect 192004 217382 192340 217410
rect 192832 217382 192984 217410
rect 193752 217382 194088 217410
rect 194580 217382 194916 217410
rect 195408 217382 195744 217410
rect 196236 217382 196572 217410
rect 197064 217382 197308 217410
rect 197892 217382 198228 217410
rect 198720 217382 199056 217410
rect 199640 217382 199976 217410
rect 200468 217382 200804 217410
rect 201296 217382 201448 217410
rect 202124 217382 202460 217410
rect 202952 217382 203288 217410
rect 203780 217382 204116 217410
rect 204608 217382 204944 217410
rect 205528 217382 205588 217410
rect 206356 217382 206876 217410
rect 207184 217382 207520 217410
rect 208012 217382 208348 217410
rect 208840 217382 209176 217410
rect 209668 217382 209728 217410
rect 210496 217382 210832 217410
rect 211416 217382 211752 217410
rect 212244 217382 212488 217410
rect 213072 217382 213408 217410
rect 213900 217382 214236 217410
rect 214728 217382 215156 217410
rect 215556 217382 215892 217410
rect 216384 217382 216628 217410
rect 217304 217382 217640 217410
rect 218132 217382 218468 217410
rect 218960 217382 219296 217410
rect 219788 217382 220124 217410
rect 220616 217382 220676 217410
rect 221444 217382 221780 217410
rect 222272 217382 222608 217410
rect 223192 217382 223528 217410
rect 224020 217382 224356 217410
rect 224848 217382 224908 217410
rect 225676 217382 226104 217410
rect 226504 217382 226840 217410
rect 227332 217382 227576 217410
rect 228160 217382 228496 217410
rect 229080 217382 229416 217410
rect 229908 217382 230336 217410
rect 230736 217382 231072 217410
rect 231564 217382 231716 217410
rect 232392 217382 232728 217410
rect 233220 217382 233556 217410
rect 234048 217382 234476 217410
rect 234968 217382 235304 217410
rect 235796 217382 235948 217410
rect 236624 217382 237052 217410
rect 237452 217382 237788 217410
rect 238280 217382 238616 217410
rect 239108 217382 239444 217410
rect 239936 217382 239996 217410
rect 240856 217382 241192 217410
rect 241684 217382 242020 217410
rect 242512 217382 242848 217410
rect 243340 217382 243676 217410
rect 244168 217382 244228 217410
rect 244996 217382 245332 217410
rect 245824 217382 246160 217410
rect 246744 217382 246896 217410
rect 247572 217382 247908 217410
rect 248400 217382 248736 217410
rect 249228 217382 249564 217410
rect 250056 217382 250392 217410
rect 250884 217382 251036 217410
rect 251712 217382 252048 217410
rect 252632 217382 252968 217410
rect 253460 217382 253888 217410
rect 254288 217382 254624 217410
rect 255116 217382 255176 217410
rect 255944 217382 256280 217410
rect 256772 217382 257108 217410
rect 257600 217382 257936 217410
rect 258520 217382 258856 217410
rect 259348 217382 259408 217410
rect 260176 217382 260604 217410
rect 261004 217382 261340 217410
rect 261832 217382 262168 217410
rect 262660 217382 262996 217410
rect 263428 217410 263456 225626
rect 263520 220590 263548 229842
rect 263704 222018 263732 231798
rect 428464 231746 428516 231752
rect 263784 230444 263836 230450
rect 263784 230386 263836 230392
rect 263692 222012 263744 222018
rect 263692 221954 263744 221960
rect 263796 221746 263824 230386
rect 264256 226030 264284 231676
rect 264348 231662 264638 231690
rect 265006 231662 265204 231690
rect 264244 226024 264296 226030
rect 264244 225966 264296 225972
rect 263784 221740 263836 221746
rect 263784 221682 263836 221688
rect 263508 220584 263560 220590
rect 263508 220526 263560 220532
rect 264348 220454 264376 231662
rect 265176 221950 265204 231662
rect 265268 231662 265374 231690
rect 265452 231662 265742 231690
rect 265268 222086 265296 231662
rect 265256 222080 265308 222086
rect 265256 222022 265308 222028
rect 265164 221944 265216 221950
rect 265164 221886 265216 221892
rect 264336 220448 264388 220454
rect 264336 220390 264388 220396
rect 265452 220386 265480 231662
rect 266096 229702 266124 231676
rect 266084 229696 266136 229702
rect 266084 229638 266136 229644
rect 265532 222964 265584 222970
rect 265532 222906 265584 222912
rect 265440 220380 265492 220386
rect 265440 220322 265492 220328
rect 264704 220312 264756 220318
rect 264704 220254 264756 220260
rect 264716 217410 264744 220254
rect 265544 217410 265572 222906
rect 266464 222154 266492 231676
rect 266740 228750 266768 231676
rect 267108 229566 267136 231676
rect 267200 231662 267490 231690
rect 267096 229560 267148 229566
rect 267096 229502 267148 229508
rect 266728 228744 266780 228750
rect 266728 228686 266780 228692
rect 266452 222148 266504 222154
rect 266452 222090 266504 222096
rect 267200 220250 267228 231662
rect 267844 221406 267872 231676
rect 268212 228818 268240 231676
rect 268304 231662 268594 231690
rect 268200 228812 268252 228818
rect 268200 228754 268252 228760
rect 267832 221400 267884 221406
rect 267832 221342 267884 221348
rect 268304 220522 268332 231662
rect 268948 230042 268976 231676
rect 269224 231662 269330 231690
rect 268936 230036 268988 230042
rect 268936 229978 268988 229984
rect 268384 229696 268436 229702
rect 268384 229638 268436 229644
rect 268292 220516 268344 220522
rect 268292 220458 268344 220464
rect 268016 220380 268068 220386
rect 268016 220322 268068 220328
rect 267188 220244 267240 220250
rect 267188 220186 267240 220192
rect 266176 220108 266228 220114
rect 266176 220050 266228 220056
rect 266188 217410 266216 220050
rect 267188 219496 267240 219502
rect 267188 219438 267240 219444
rect 267200 217410 267228 219438
rect 268028 217410 268056 220322
rect 268396 219502 268424 229638
rect 268936 224460 268988 224466
rect 268936 224402 268988 224408
rect 268384 219496 268436 219502
rect 268384 219438 268436 219444
rect 268948 217410 268976 224402
rect 269224 221338 269252 231662
rect 269592 227050 269620 231676
rect 269960 230246 269988 231676
rect 270052 231662 270342 231690
rect 269948 230240 270000 230246
rect 269948 230182 270000 230188
rect 269580 227044 269632 227050
rect 269580 226986 269632 226992
rect 269212 221332 269264 221338
rect 269212 221274 269264 221280
rect 269672 220788 269724 220794
rect 269672 220730 269724 220736
rect 269684 217410 269712 220730
rect 270052 220658 270080 231662
rect 270408 230036 270460 230042
rect 270408 229978 270460 229984
rect 270316 229968 270368 229974
rect 270316 229910 270368 229916
rect 270132 229560 270184 229566
rect 270132 229502 270184 229508
rect 270144 220726 270172 229502
rect 270328 220794 270356 229910
rect 270316 220788 270368 220794
rect 270316 220730 270368 220736
rect 270132 220720 270184 220726
rect 270132 220662 270184 220668
rect 270040 220652 270092 220658
rect 270040 220594 270092 220600
rect 270420 217410 270448 229978
rect 270696 221270 270724 231676
rect 271064 224262 271092 231676
rect 271328 230376 271380 230382
rect 271328 230318 271380 230324
rect 271144 230104 271196 230110
rect 271144 230046 271196 230052
rect 271052 224256 271104 224262
rect 271052 224198 271104 224204
rect 270684 221264 270736 221270
rect 270684 221206 270736 221212
rect 271156 219774 271184 230046
rect 271236 229288 271288 229294
rect 271236 229230 271288 229236
rect 271248 220182 271276 229230
rect 271340 220794 271368 230318
rect 271432 229566 271460 231676
rect 271800 230178 271828 231676
rect 271984 231662 272182 231690
rect 272260 231662 272458 231690
rect 271788 230172 271840 230178
rect 271788 230114 271840 230120
rect 271420 229560 271472 229566
rect 271420 229502 271472 229508
rect 271984 221202 272012 231662
rect 272260 224330 272288 231662
rect 272812 230382 272840 231676
rect 272904 231662 273194 231690
rect 273456 231662 273562 231690
rect 273640 231662 273930 231690
rect 272800 230376 272852 230382
rect 272800 230318 272852 230324
rect 272248 224324 272300 224330
rect 272248 224266 272300 224272
rect 272248 221468 272300 221474
rect 272248 221410 272300 221416
rect 271972 221196 272024 221202
rect 271972 221138 272024 221144
rect 271328 220788 271380 220794
rect 271328 220730 271380 220736
rect 271420 220244 271472 220250
rect 271420 220186 271472 220192
rect 271236 220176 271288 220182
rect 271236 220118 271288 220124
rect 271144 219768 271196 219774
rect 271144 219710 271196 219716
rect 271432 217410 271460 220186
rect 272260 217410 272288 221410
rect 272904 220046 272932 231662
rect 272984 229560 273036 229566
rect 272984 229502 273036 229508
rect 272892 220040 272944 220046
rect 272892 219982 272944 219988
rect 272996 219706 273024 229502
rect 273456 221542 273484 231662
rect 273640 224398 273668 231662
rect 274284 230314 274312 231676
rect 274652 230450 274680 231676
rect 274836 231662 275034 231690
rect 275112 231662 275310 231690
rect 274640 230444 274692 230450
rect 274640 230386 274692 230392
rect 274272 230308 274324 230314
rect 274272 230250 274324 230256
rect 274548 230308 274600 230314
rect 274548 230250 274600 230256
rect 273904 229492 273956 229498
rect 273904 229434 273956 229440
rect 273916 229094 273944 229434
rect 273824 229066 273944 229094
rect 273628 224392 273680 224398
rect 273628 224334 273680 224340
rect 273444 221536 273496 221542
rect 273444 221478 273496 221484
rect 273076 220652 273128 220658
rect 273076 220594 273128 220600
rect 272984 219700 273036 219706
rect 272984 219642 273036 219648
rect 273088 217410 273116 220594
rect 273824 220318 273852 229066
rect 274560 220794 274588 230250
rect 274836 221134 274864 231662
rect 275112 223174 275140 231662
rect 275284 230172 275336 230178
rect 275284 230114 275336 230120
rect 275100 223168 275152 223174
rect 275100 223110 275152 223116
rect 274824 221128 274876 221134
rect 274824 221070 274876 221076
rect 273904 220788 273956 220794
rect 273904 220730 273956 220736
rect 274548 220788 274600 220794
rect 274548 220730 274600 220736
rect 273812 220312 273864 220318
rect 273812 220254 273864 220260
rect 273916 217410 273944 220730
rect 274456 220720 274508 220726
rect 274456 220662 274508 220668
rect 274468 217410 274496 220662
rect 275296 220250 275324 230114
rect 275664 229634 275692 231676
rect 276046 231662 276244 231690
rect 275652 229628 275704 229634
rect 275652 229570 275704 229576
rect 275376 229424 275428 229430
rect 275376 229366 275428 229372
rect 275388 220386 275416 229366
rect 275560 221536 275612 221542
rect 275560 221478 275612 221484
rect 275376 220380 275428 220386
rect 275376 220322 275428 220328
rect 275284 220244 275336 220250
rect 275284 220186 275336 220192
rect 275572 217410 275600 221478
rect 276216 219978 276244 231662
rect 276400 228478 276428 231676
rect 276492 231662 276782 231690
rect 276388 228472 276440 228478
rect 276388 228414 276440 228420
rect 276492 226098 276520 231662
rect 276756 230444 276808 230450
rect 276756 230386 276808 230392
rect 276664 230240 276716 230246
rect 276664 230182 276716 230188
rect 276480 226092 276532 226098
rect 276480 226034 276532 226040
rect 276676 220726 276704 230182
rect 276664 220720 276716 220726
rect 276664 220662 276716 220668
rect 276768 220658 276796 230386
rect 277136 230110 277164 231676
rect 277518 231662 277624 231690
rect 277124 230104 277176 230110
rect 277124 230046 277176 230052
rect 277216 230104 277268 230110
rect 277216 230046 277268 230052
rect 277228 229702 277256 230046
rect 277216 229696 277268 229702
rect 277216 229638 277268 229644
rect 277308 229628 277360 229634
rect 277308 229570 277360 229576
rect 277492 229628 277544 229634
rect 277492 229570 277544 229576
rect 276756 220652 276808 220658
rect 276756 220594 276808 220600
rect 276204 219972 276256 219978
rect 276204 219914 276256 219920
rect 276480 219496 276532 219502
rect 276480 219438 276532 219444
rect 276492 217410 276520 219438
rect 277320 217410 277348 229570
rect 277504 229362 277532 229570
rect 277492 229356 277544 229362
rect 277492 229298 277544 229304
rect 277596 219910 277624 231662
rect 277768 230444 277820 230450
rect 277768 230386 277820 230392
rect 277780 230178 277808 230386
rect 277676 230172 277728 230178
rect 277676 230114 277728 230120
rect 277768 230172 277820 230178
rect 277768 230114 277820 230120
rect 277688 229634 277716 230114
rect 277676 229628 277728 229634
rect 277676 229570 277728 229576
rect 277872 227118 277900 231676
rect 278044 230308 278096 230314
rect 278044 230250 278096 230256
rect 277860 227112 277912 227118
rect 277860 227054 277912 227060
rect 277584 219904 277636 219910
rect 277584 219846 277636 219852
rect 278056 219502 278084 230250
rect 278148 225622 278176 231676
rect 278516 229770 278544 231676
rect 278898 231662 279004 231690
rect 278504 229764 278556 229770
rect 278504 229706 278556 229712
rect 278688 229764 278740 229770
rect 278688 229706 278740 229712
rect 278136 225616 278188 225622
rect 278136 225558 278188 225564
rect 278700 220794 278728 229706
rect 278136 220788 278188 220794
rect 278136 220730 278188 220736
rect 278688 220788 278740 220794
rect 278688 220730 278740 220736
rect 278044 219496 278096 219502
rect 278044 219438 278096 219444
rect 278148 217410 278176 220730
rect 278596 220108 278648 220114
rect 278596 220050 278648 220056
rect 263428 217382 263488 217410
rect 264408 217382 264744 217410
rect 265236 217382 265572 217410
rect 266064 217382 266216 217410
rect 266892 217382 267228 217410
rect 267720 217382 268056 217410
rect 268548 217382 268976 217410
rect 269376 217382 269712 217410
rect 270296 217382 270448 217410
rect 271124 217382 271460 217410
rect 271952 217382 272288 217410
rect 272780 217382 273116 217410
rect 273608 217382 273944 217410
rect 274436 217382 274496 217410
rect 275264 217382 275600 217410
rect 276184 217382 276520 217410
rect 277012 217382 277348 217410
rect 277840 217382 278176 217410
rect 278608 217410 278636 220050
rect 278976 219842 279004 231662
rect 279252 227186 279280 231676
rect 279424 230376 279476 230382
rect 279424 230318 279476 230324
rect 279240 227180 279292 227186
rect 279240 227122 279292 227128
rect 279436 220182 279464 230318
rect 279620 228410 279648 231676
rect 279988 229294 280016 231676
rect 280356 229838 280384 231676
rect 280344 229832 280396 229838
rect 280344 229774 280396 229780
rect 280068 229696 280120 229702
rect 280068 229638 280120 229644
rect 279976 229288 280028 229294
rect 279976 229230 280028 229236
rect 279608 228404 279660 228410
rect 279608 228346 279660 228352
rect 279424 220176 279476 220182
rect 279424 220118 279476 220124
rect 278964 219836 279016 219842
rect 278964 219778 279016 219784
rect 280080 219434 280108 229638
rect 280724 222902 280752 231676
rect 281000 225690 281028 231676
rect 281092 231662 281382 231690
rect 281092 229566 281120 231662
rect 281736 229906 281764 231676
rect 281724 229900 281776 229906
rect 281724 229842 281776 229848
rect 281356 229832 281408 229838
rect 281356 229774 281408 229780
rect 281080 229560 281132 229566
rect 281080 229502 281132 229508
rect 280988 225684 281040 225690
rect 280988 225626 281040 225632
rect 280712 222896 280764 222902
rect 280712 222838 280764 222844
rect 280620 220176 280672 220182
rect 280620 220118 280672 220124
rect 279896 219406 280108 219434
rect 279896 217410 279924 219406
rect 280632 217410 280660 220118
rect 281368 217410 281396 229774
rect 281448 229288 281500 229294
rect 281448 229230 281500 229236
rect 281460 220182 281488 229230
rect 282104 222970 282132 231676
rect 282472 230110 282500 231676
rect 282460 230104 282512 230110
rect 282460 230046 282512 230052
rect 282840 229498 282868 231676
rect 283208 230382 283236 231676
rect 283196 230376 283248 230382
rect 283196 230318 283248 230324
rect 282828 229492 282880 229498
rect 282828 229434 282880 229440
rect 282828 229220 282880 229226
rect 282828 229162 282880 229168
rect 282092 222964 282144 222970
rect 282092 222906 282144 222912
rect 282840 220794 282868 229162
rect 283576 224466 283604 231676
rect 283852 230042 283880 231676
rect 283840 230036 283892 230042
rect 283840 229978 283892 229984
rect 284116 229900 284168 229906
rect 284116 229842 284168 229848
rect 283564 224460 283616 224466
rect 283564 224402 283616 224408
rect 284128 220794 284156 229842
rect 284220 229430 284248 231676
rect 284588 229974 284616 231676
rect 284680 231662 284970 231690
rect 284576 229968 284628 229974
rect 284576 229910 284628 229916
rect 284208 229424 284260 229430
rect 284208 229366 284260 229372
rect 284208 229152 284260 229158
rect 284208 229094 284260 229100
rect 282368 220788 282420 220794
rect 282368 220730 282420 220736
rect 282828 220788 282880 220794
rect 282828 220730 282880 220736
rect 283196 220788 283248 220794
rect 283196 220730 283248 220736
rect 284116 220788 284168 220794
rect 284116 220730 284168 220736
rect 281448 220176 281500 220182
rect 281448 220118 281500 220124
rect 282380 217410 282408 220730
rect 283208 217410 283236 220730
rect 284220 219434 284248 229094
rect 284680 221474 284708 231662
rect 285324 230450 285352 231676
rect 285312 230444 285364 230450
rect 285312 230386 285364 230392
rect 285496 230036 285548 230042
rect 285496 229978 285548 229984
rect 284668 221468 284720 221474
rect 284668 221410 284720 221416
rect 284852 219972 284904 219978
rect 284852 219914 284904 219920
rect 284128 219406 284248 219434
rect 284128 217410 284156 219406
rect 284864 217410 284892 219914
rect 285508 217410 285536 229978
rect 285588 229968 285640 229974
rect 285588 229910 285640 229916
rect 285600 219978 285628 229910
rect 285692 229634 285720 231676
rect 286060 230178 286088 231676
rect 286152 231662 286442 231690
rect 286048 230172 286100 230178
rect 286048 230114 286100 230120
rect 285680 229628 285732 229634
rect 285680 229570 285732 229576
rect 286152 221542 286180 231662
rect 286704 229362 286732 231676
rect 286968 230308 287020 230314
rect 286968 230250 287020 230256
rect 286692 229356 286744 229362
rect 286692 229298 286744 229304
rect 286140 221536 286192 221542
rect 286140 221478 286192 221484
rect 286980 220794 287008 230250
rect 287072 230246 287100 231676
rect 287440 230382 287468 231676
rect 287532 231662 287822 231690
rect 287428 230376 287480 230382
rect 287428 230318 287480 230324
rect 287060 230240 287112 230246
rect 287060 230182 287112 230188
rect 286508 220788 286560 220794
rect 286508 220730 286560 220736
rect 286968 220788 287020 220794
rect 286968 220730 287020 220736
rect 287336 220788 287388 220794
rect 287336 220730 287388 220736
rect 285588 219972 285640 219978
rect 285588 219914 285640 219920
rect 286520 217410 286548 220730
rect 287348 217410 287376 220730
rect 287532 220182 287560 231662
rect 288176 229294 288204 231676
rect 288348 230444 288400 230450
rect 288348 230386 288400 230392
rect 288164 229288 288216 229294
rect 288164 229230 288216 229236
rect 287520 220176 287572 220182
rect 287520 220118 287572 220124
rect 288360 217410 288388 230386
rect 288544 229770 288572 231676
rect 288532 229764 288584 229770
rect 288532 229706 288584 229712
rect 288912 229702 288940 231676
rect 288900 229696 288952 229702
rect 288900 229638 288952 229644
rect 289280 229226 289308 231676
rect 289268 229220 289320 229226
rect 289268 229162 289320 229168
rect 289556 229158 289584 231676
rect 289924 229838 289952 231676
rect 290292 229906 290320 231676
rect 290660 230042 290688 231676
rect 290752 231662 291042 231690
rect 290648 230036 290700 230042
rect 290648 229978 290700 229984
rect 290280 229900 290332 229906
rect 290280 229842 290332 229848
rect 289912 229832 289964 229838
rect 289912 229774 289964 229780
rect 289544 229152 289596 229158
rect 289544 229094 289596 229100
rect 290752 229094 290780 231662
rect 291396 229974 291424 231676
rect 291764 230314 291792 231676
rect 291856 231662 292146 231690
rect 292224 231662 292422 231690
rect 291752 230308 291804 230314
rect 291752 230250 291804 230256
rect 291384 229968 291436 229974
rect 291384 229910 291436 229916
rect 290660 229066 290780 229094
rect 290660 220794 290688 229066
rect 290648 220788 290700 220794
rect 290648 220730 290700 220736
rect 290740 220788 290792 220794
rect 290740 220730 290792 220736
rect 289084 220720 289136 220726
rect 289084 220662 289136 220668
rect 289096 217410 289124 220662
rect 289636 220040 289688 220046
rect 289636 219982 289688 219988
rect 289648 217410 289676 219982
rect 290752 217410 290780 220730
rect 291856 220726 291884 231662
rect 292224 220794 292252 231662
rect 292776 230450 292804 231676
rect 292868 231662 293158 231690
rect 293236 231662 293526 231690
rect 292764 230444 292816 230450
rect 292764 230386 292816 230392
rect 292580 229152 292632 229158
rect 292580 229094 292632 229100
rect 292592 224262 292620 229094
rect 292580 224256 292632 224262
rect 292580 224198 292632 224204
rect 292212 220788 292264 220794
rect 292212 220730 292264 220736
rect 292488 220788 292540 220794
rect 292488 220730 292540 220736
rect 291844 220720 291896 220726
rect 291844 220662 291896 220668
rect 291476 220652 291528 220658
rect 291476 220594 291528 220600
rect 291488 217410 291516 220594
rect 292500 217410 292528 220730
rect 292868 220046 292896 231662
rect 293236 220794 293264 231662
rect 293880 229158 293908 231676
rect 293868 229152 293920 229158
rect 293868 229094 293920 229100
rect 294248 228410 294276 231676
rect 294236 228404 294288 228410
rect 294236 228346 294288 228352
rect 294052 228200 294104 228206
rect 294052 228142 294104 228148
rect 293960 226976 294012 226982
rect 293960 226918 294012 226924
rect 293500 224256 293552 224262
rect 293500 224198 293552 224204
rect 293224 220788 293276 220794
rect 293224 220730 293276 220736
rect 292856 220040 292908 220046
rect 292856 219982 292908 219988
rect 293224 219836 293276 219842
rect 293224 219778 293276 219784
rect 293236 217410 293264 219778
rect 278608 217382 278668 217410
rect 279496 217382 279924 217410
rect 280324 217382 280660 217410
rect 281152 217382 281396 217410
rect 282072 217382 282408 217410
rect 282900 217382 283236 217410
rect 283728 217382 284156 217410
rect 284556 217382 284892 217410
rect 285384 217382 285536 217410
rect 286212 217382 286548 217410
rect 287040 217382 287376 217410
rect 287960 217382 288388 217410
rect 288788 217382 289124 217410
rect 289616 217382 289676 217410
rect 290444 217382 290780 217410
rect 291272 217382 291516 217410
rect 292100 217382 292528 217410
rect 292928 217382 293264 217410
rect 293512 217410 293540 224198
rect 293972 219842 294000 226918
rect 294064 220658 294092 228142
rect 294616 226982 294644 231676
rect 294998 231662 295196 231690
rect 295168 229106 295196 231662
rect 295260 229226 295288 231676
rect 295536 231662 295642 231690
rect 295904 231662 296010 231690
rect 295248 229220 295300 229226
rect 295248 229162 295300 229168
rect 295168 229078 295380 229106
rect 294604 226976 294656 226982
rect 294604 226918 294656 226924
rect 294972 220788 295024 220794
rect 294972 220730 295024 220736
rect 294052 220652 294104 220658
rect 294052 220594 294104 220600
rect 293960 219836 294012 219842
rect 293960 219778 294012 219784
rect 294984 217410 295012 220730
rect 293512 217382 293848 217410
rect 294676 217382 295012 217410
rect 295352 217410 295380 229078
rect 295536 220794 295564 231662
rect 295524 220788 295576 220794
rect 295524 220730 295576 220736
rect 295904 217410 295932 231662
rect 296364 229294 296392 231676
rect 296732 229362 296760 231676
rect 296824 231662 297114 231690
rect 296720 229356 296772 229362
rect 296720 229298 296772 229304
rect 296352 229288 296404 229294
rect 296352 229230 296404 229236
rect 296824 217870 296852 231662
rect 297468 229226 297496 231676
rect 297850 231662 298048 231690
rect 296904 229220 296956 229226
rect 296904 229162 296956 229168
rect 297456 229220 297508 229226
rect 297456 229162 297508 229168
rect 296812 217864 296864 217870
rect 296812 217806 296864 217812
rect 296916 217410 296944 229162
rect 298020 220794 298048 231662
rect 298112 229158 298140 231676
rect 298480 229430 298508 231676
rect 298848 229838 298876 231676
rect 299230 231662 299336 231690
rect 298836 229832 298888 229838
rect 298836 229774 298888 229780
rect 298468 229424 298520 229430
rect 298468 229366 298520 229372
rect 298468 229288 298520 229294
rect 298468 229230 298520 229236
rect 298100 229152 298152 229158
rect 298100 229094 298152 229100
rect 298008 220788 298060 220794
rect 298008 220730 298060 220736
rect 297640 217864 297692 217870
rect 297640 217806 297692 217812
rect 297652 217410 297680 217806
rect 298480 217410 298508 229230
rect 299308 220522 299336 231662
rect 299480 229220 299532 229226
rect 299480 229162 299532 229168
rect 299388 229152 299440 229158
rect 299388 229094 299440 229100
rect 299400 220590 299428 229094
rect 299492 224954 299520 229162
rect 299584 229158 299612 231676
rect 299952 230450 299980 231676
rect 300334 231662 300624 231690
rect 299940 230444 299992 230450
rect 299940 230386 299992 230392
rect 300124 229356 300176 229362
rect 300124 229298 300176 229304
rect 299572 229152 299624 229158
rect 299572 229094 299624 229100
rect 299492 224926 299612 224954
rect 299388 220584 299440 220590
rect 299388 220526 299440 220532
rect 299296 220516 299348 220522
rect 299296 220458 299348 220464
rect 299584 217410 299612 224926
rect 300136 217410 300164 229298
rect 300492 229152 300544 229158
rect 300492 229094 300544 229100
rect 300504 219638 300532 229094
rect 300492 219632 300544 219638
rect 300492 219574 300544 219580
rect 300596 219502 300624 231662
rect 300688 229566 300716 231676
rect 300978 231662 301268 231690
rect 301346 231662 301636 231690
rect 301714 231662 302004 231690
rect 300676 229560 300728 229566
rect 300676 229502 300728 229508
rect 301136 229424 301188 229430
rect 301136 229366 301188 229372
rect 300584 219496 300636 219502
rect 300584 219438 300636 219444
rect 301148 219434 301176 229366
rect 301240 221474 301268 231662
rect 301228 221468 301280 221474
rect 301228 221410 301280 221416
rect 301608 219570 301636 231662
rect 301976 220114 302004 231662
rect 302068 229770 302096 231676
rect 302056 229764 302108 229770
rect 302056 229706 302108 229712
rect 302436 225690 302464 231676
rect 302818 231662 303108 231690
rect 303186 231662 303476 231690
rect 302516 229832 302568 229838
rect 302516 229774 302568 229780
rect 302528 229094 302556 229774
rect 302528 229066 302648 229094
rect 302424 225684 302476 225690
rect 302424 225626 302476 225632
rect 302240 220788 302292 220794
rect 302240 220730 302292 220736
rect 301964 220108 302016 220114
rect 301964 220050 302016 220056
rect 301596 219564 301648 219570
rect 301596 219506 301648 219512
rect 301148 219406 301268 219434
rect 301240 217410 301268 219406
rect 302252 217410 302280 220730
rect 295352 217382 295504 217410
rect 295904 217382 296332 217410
rect 296916 217382 297160 217410
rect 297652 217382 297988 217410
rect 298480 217382 298816 217410
rect 299584 217382 299736 217410
rect 300136 217382 300564 217410
rect 301240 217382 301392 217410
rect 302220 217382 302280 217410
rect 302620 217410 302648 229066
rect 303080 220726 303108 231662
rect 303068 220720 303120 220726
rect 303068 220662 303120 220668
rect 303448 220658 303476 231662
rect 303540 229838 303568 231676
rect 303528 229832 303580 229838
rect 303528 229774 303580 229780
rect 303816 225758 303844 231676
rect 304198 231662 304488 231690
rect 304566 231662 304856 231690
rect 303988 230444 304040 230450
rect 303988 230386 304040 230392
rect 304000 229094 304028 230386
rect 304000 229066 304304 229094
rect 303804 225752 303856 225758
rect 303804 225694 303856 225700
rect 303436 220652 303488 220658
rect 303436 220594 303488 220600
rect 303620 220584 303672 220590
rect 303620 220526 303672 220532
rect 303632 217410 303660 220526
rect 304276 217410 304304 229066
rect 304460 220182 304488 231662
rect 304828 220590 304856 231662
rect 304920 229906 304948 231676
rect 304908 229900 304960 229906
rect 304908 229842 304960 229848
rect 305288 227050 305316 231676
rect 305656 230382 305684 231676
rect 306038 231662 306144 231690
rect 305644 230376 305696 230382
rect 305644 230318 305696 230324
rect 305552 229560 305604 229566
rect 305552 229502 305604 229508
rect 305276 227044 305328 227050
rect 305276 226986 305328 226992
rect 305564 220862 305592 229502
rect 305552 220856 305604 220862
rect 305552 220798 305604 220804
rect 304816 220584 304868 220590
rect 304816 220526 304868 220532
rect 305276 220516 305328 220522
rect 305276 220458 305328 220464
rect 304448 220176 304500 220182
rect 304448 220118 304500 220124
rect 305288 217410 305316 220458
rect 306116 220454 306144 231662
rect 306196 230376 306248 230382
rect 306196 230318 306248 230324
rect 306208 220522 306236 230318
rect 306392 223038 306420 231676
rect 306668 228546 306696 231676
rect 307036 230382 307064 231676
rect 307024 230376 307076 230382
rect 307024 230318 307076 230324
rect 306656 228540 306708 228546
rect 306656 228482 306708 228488
rect 306380 223032 306432 223038
rect 306380 222974 306432 222980
rect 306196 220516 306248 220522
rect 306196 220458 306248 220464
rect 306104 220448 306156 220454
rect 306104 220390 306156 220396
rect 307404 220318 307432 231676
rect 307576 230376 307628 230382
rect 307576 230318 307628 230324
rect 307588 220386 307616 230318
rect 307772 224398 307800 231676
rect 308140 228410 308168 231676
rect 308128 228404 308180 228410
rect 308128 228346 308180 228352
rect 307760 224392 307812 224398
rect 307760 224334 307812 224340
rect 308508 222902 308536 231676
rect 308784 231662 308890 231690
rect 308496 222896 308548 222902
rect 308496 222838 308548 222844
rect 308588 220856 308640 220862
rect 308588 220798 308640 220804
rect 307576 220380 307628 220386
rect 307576 220322 307628 220328
rect 307392 220312 307444 220318
rect 307392 220254 307444 220260
rect 306932 219632 306984 219638
rect 306932 219574 306984 219580
rect 306380 219496 306432 219502
rect 306380 219438 306432 219444
rect 306392 217410 306420 219438
rect 306944 217410 306972 219574
rect 307760 219564 307812 219570
rect 307760 219506 307812 219512
rect 307772 217410 307800 219506
rect 308600 217410 308628 220798
rect 308784 220250 308812 231662
rect 309244 224330 309272 231676
rect 309520 227458 309548 231676
rect 309888 228478 309916 231676
rect 309876 228472 309928 228478
rect 309876 228414 309928 228420
rect 309508 227452 309560 227458
rect 309508 227394 309560 227400
rect 309232 224324 309284 224330
rect 309232 224266 309284 224272
rect 308772 220244 308824 220250
rect 308772 220186 308824 220192
rect 310256 220114 310284 231676
rect 310624 229430 310652 231676
rect 310612 229424 310664 229430
rect 310612 229366 310664 229372
rect 310992 225622 311020 231676
rect 311164 229764 311216 229770
rect 311164 229706 311216 229712
rect 310980 225616 311032 225622
rect 310980 225558 311032 225564
rect 311176 222154 311204 229706
rect 311360 224262 311388 231676
rect 311728 230246 311756 231676
rect 312096 230382 312124 231676
rect 312084 230376 312136 230382
rect 312084 230318 312136 230324
rect 311716 230240 311768 230246
rect 311716 230182 311768 230188
rect 312372 230042 312400 231676
rect 312360 230036 312412 230042
rect 312360 229978 312412 229984
rect 311624 229900 311676 229906
rect 311624 229842 311676 229848
rect 311348 224256 311400 224262
rect 311348 224198 311400 224204
rect 311636 223174 311664 229842
rect 312544 229832 312596 229838
rect 312544 229774 312596 229780
rect 311624 223168 311676 223174
rect 311624 223110 311676 223116
rect 312556 222154 312584 229774
rect 312740 227322 312768 231676
rect 313108 229294 313136 231676
rect 313188 230376 313240 230382
rect 313188 230318 313240 230324
rect 313096 229288 313148 229294
rect 313096 229230 313148 229236
rect 312728 227316 312780 227322
rect 312728 227258 312780 227264
rect 311164 222148 311216 222154
rect 311164 222090 311216 222096
rect 311992 222148 312044 222154
rect 311992 222090 312044 222096
rect 312544 222148 312596 222154
rect 312544 222090 312596 222096
rect 310520 221468 310572 221474
rect 310520 221410 310572 221416
rect 309416 220108 309468 220114
rect 309416 220050 309468 220056
rect 310244 220108 310296 220114
rect 310244 220050 310296 220056
rect 309428 217410 309456 220050
rect 310532 217410 310560 221410
rect 311164 220720 311216 220726
rect 311164 220662 311216 220668
rect 311176 217410 311204 220662
rect 312004 217410 312032 222090
rect 313200 221202 313228 230318
rect 313476 229634 313504 231676
rect 313844 229974 313872 231676
rect 313832 229968 313884 229974
rect 313832 229910 313884 229916
rect 313464 229628 313516 229634
rect 313464 229570 313516 229576
rect 313556 225684 313608 225690
rect 313556 225626 313608 225632
rect 313188 221196 313240 221202
rect 313188 221138 313240 221144
rect 312820 220652 312872 220658
rect 312820 220594 312872 220600
rect 312832 217410 312860 220594
rect 313568 217410 313596 225626
rect 314212 223106 314240 231676
rect 314580 230382 314608 231676
rect 314948 230450 314976 231676
rect 314936 230444 314988 230450
rect 314936 230386 314988 230392
rect 314568 230376 314620 230382
rect 314568 230318 314620 230324
rect 314568 229628 314620 229634
rect 314568 229570 314620 229576
rect 314476 229424 314528 229430
rect 314476 229366 314528 229372
rect 314488 225690 314516 229366
rect 314476 225684 314528 225690
rect 314476 225626 314528 225632
rect 314200 223100 314252 223106
rect 314200 223042 314252 223048
rect 314580 221270 314608 229570
rect 315224 229362 315252 231676
rect 315304 230240 315356 230246
rect 315304 230182 315356 230188
rect 315212 229356 315264 229362
rect 315212 229298 315264 229304
rect 315316 229094 315344 230182
rect 315316 229066 315436 229094
rect 315304 222148 315356 222154
rect 315304 222090 315356 222096
rect 314568 221264 314620 221270
rect 314568 221206 314620 221212
rect 314660 220176 314712 220182
rect 314660 220118 314712 220124
rect 314672 217410 314700 220118
rect 315316 217410 315344 222090
rect 315408 220182 315436 229066
rect 315592 227390 315620 231676
rect 315868 231662 315974 231690
rect 315868 230110 315896 231662
rect 315948 230444 316000 230450
rect 315948 230386 316000 230392
rect 315856 230104 315908 230110
rect 315856 230046 315908 230052
rect 315580 227384 315632 227390
rect 315580 227326 315632 227332
rect 315960 221338 315988 230386
rect 316328 230382 316356 231676
rect 316316 230376 316368 230382
rect 316316 230318 316368 230324
rect 316696 229906 316724 231676
rect 316684 229900 316736 229906
rect 316684 229842 316736 229848
rect 317064 222970 317092 231676
rect 317328 230376 317380 230382
rect 317328 230318 317380 230324
rect 317052 222964 317104 222970
rect 317052 222906 317104 222912
rect 317340 221406 317368 230318
rect 317432 230178 317460 231676
rect 317800 230382 317828 231676
rect 317788 230376 317840 230382
rect 317788 230318 317840 230324
rect 317420 230172 317472 230178
rect 317420 230114 317472 230120
rect 318076 229838 318104 231676
rect 318064 229832 318116 229838
rect 318064 229774 318116 229780
rect 318064 229288 318116 229294
rect 318064 229230 318116 229236
rect 317420 225752 317472 225758
rect 317420 225694 317472 225700
rect 317328 221400 317380 221406
rect 317328 221342 317380 221348
rect 315948 221332 316000 221338
rect 315948 221274 316000 221280
rect 316132 220584 316184 220590
rect 316132 220526 316184 220532
rect 315396 220176 315448 220182
rect 315396 220118 315448 220124
rect 316144 217410 316172 220526
rect 317432 217410 317460 225694
rect 317880 220516 317932 220522
rect 317880 220458 317932 220464
rect 302620 217382 303048 217410
rect 303632 217382 303876 217410
rect 304276 217382 304704 217410
rect 305288 217382 305624 217410
rect 306392 217382 306452 217410
rect 306944 217382 307280 217410
rect 307772 217382 308108 217410
rect 308600 217382 308936 217410
rect 309428 217382 309764 217410
rect 310532 217382 310592 217410
rect 311176 217382 311512 217410
rect 312004 217382 312340 217410
rect 312832 217382 313168 217410
rect 313568 217382 313996 217410
rect 314672 217382 314824 217410
rect 315316 217382 315652 217410
rect 316144 217382 316480 217410
rect 317400 217382 317460 217410
rect 317892 217410 317920 220458
rect 318076 220046 318104 229230
rect 318444 227254 318472 231676
rect 318812 230450 318840 231676
rect 319194 231662 319484 231690
rect 319562 231662 319852 231690
rect 318800 230444 318852 230450
rect 318800 230386 318852 230392
rect 318708 230376 318760 230382
rect 318708 230318 318760 230324
rect 319260 230376 319312 230382
rect 319260 230318 319312 230324
rect 318432 227248 318484 227254
rect 318432 227190 318484 227196
rect 318720 222154 318748 230318
rect 319272 223242 319300 230318
rect 319352 230308 319404 230314
rect 319352 230250 319404 230256
rect 319260 223236 319312 223242
rect 319260 223178 319312 223184
rect 318892 223168 318944 223174
rect 318892 223110 318944 223116
rect 318708 222148 318760 222154
rect 318708 222090 318760 222096
rect 318064 220040 318116 220046
rect 318064 219982 318116 219988
rect 318904 217410 318932 223110
rect 319364 220522 319392 230250
rect 319456 221542 319484 231662
rect 319444 221536 319496 221542
rect 319444 221478 319496 221484
rect 319824 221474 319852 231662
rect 319916 230382 319944 231676
rect 319904 230376 319956 230382
rect 319904 230318 319956 230324
rect 320284 230246 320312 231676
rect 320652 230382 320680 231676
rect 320942 231662 321232 231690
rect 320640 230376 320692 230382
rect 320640 230318 320692 230324
rect 320272 230240 320324 230246
rect 320272 230182 320324 230188
rect 320272 227044 320324 227050
rect 320272 226986 320324 226992
rect 319812 221468 319864 221474
rect 319812 221410 319864 221416
rect 319352 220516 319404 220522
rect 319352 220458 319404 220464
rect 319536 220448 319588 220454
rect 319536 220390 319588 220396
rect 319548 217410 319576 220390
rect 320284 217410 320312 226986
rect 321204 222018 321232 231662
rect 321296 227186 321324 231676
rect 321664 230382 321692 231676
rect 322046 231662 322336 231690
rect 322414 231662 322704 231690
rect 321376 230376 321428 230382
rect 321376 230318 321428 230324
rect 321652 230376 321704 230382
rect 321652 230318 321704 230324
rect 321284 227180 321336 227186
rect 321284 227122 321336 227128
rect 321388 222086 321416 230318
rect 322204 230104 322256 230110
rect 322204 230046 322256 230052
rect 321928 223032 321980 223038
rect 321928 222974 321980 222980
rect 321376 222080 321428 222086
rect 321376 222022 321428 222028
rect 321192 222012 321244 222018
rect 321192 221954 321244 221960
rect 321560 220380 321612 220386
rect 321560 220322 321612 220328
rect 321572 217410 321600 220322
rect 317892 217382 318228 217410
rect 318904 217382 319056 217410
rect 319548 217382 319884 217410
rect 320284 217382 320712 217410
rect 321540 217382 321600 217410
rect 321940 217410 321968 222974
rect 322216 219910 322244 230046
rect 322308 221950 322336 231662
rect 322296 221944 322348 221950
rect 322296 221886 322348 221892
rect 322676 221882 322704 231662
rect 322768 226030 322796 231676
rect 323136 229702 323164 231676
rect 323124 229696 323176 229702
rect 323124 229638 323176 229644
rect 323504 229158 323532 231676
rect 323780 230110 323808 231676
rect 323768 230104 323820 230110
rect 323768 230046 323820 230052
rect 323492 229152 323544 229158
rect 323492 229094 323544 229100
rect 323676 228540 323728 228546
rect 323676 228482 323728 228488
rect 322756 226024 322808 226030
rect 322756 225966 322808 225972
rect 322664 221876 322716 221882
rect 322664 221818 322716 221824
rect 322940 220312 322992 220318
rect 322940 220254 322992 220260
rect 322204 219904 322256 219910
rect 322204 219846 322256 219852
rect 322952 217410 322980 220254
rect 323688 217410 323716 228482
rect 324148 225826 324176 231676
rect 324516 229158 324544 231676
rect 324884 229226 324912 231676
rect 325266 231662 325464 231690
rect 324872 229220 324924 229226
rect 324872 229162 324924 229168
rect 324228 229152 324280 229158
rect 324228 229094 324280 229100
rect 324504 229152 324556 229158
rect 324504 229094 324556 229100
rect 325332 229152 325384 229158
rect 325332 229094 325384 229100
rect 324136 225820 324188 225826
rect 324136 225762 324188 225768
rect 324240 221814 324268 229094
rect 324504 222896 324556 222902
rect 324504 222838 324556 222844
rect 324228 221808 324280 221814
rect 324228 221750 324280 221756
rect 324516 217410 324544 222838
rect 325344 220794 325372 229094
rect 325436 221610 325464 231662
rect 325516 229220 325568 229226
rect 325516 229162 325568 229168
rect 325528 221746 325556 229162
rect 325620 227050 325648 231676
rect 326002 231662 326292 231690
rect 326370 231662 326568 231690
rect 325608 227044 325660 227050
rect 325608 226986 325660 226992
rect 325700 224392 325752 224398
rect 325700 224334 325752 224340
rect 325516 221740 325568 221746
rect 325516 221682 325568 221688
rect 325424 221604 325476 221610
rect 325424 221546 325476 221552
rect 325332 220788 325384 220794
rect 325332 220730 325384 220736
rect 325712 217410 325740 224334
rect 326264 220726 326292 231662
rect 326344 230444 326396 230450
rect 326344 230386 326396 230392
rect 326356 229770 326384 230386
rect 326344 229764 326396 229770
rect 326344 229706 326396 229712
rect 326540 221678 326568 231662
rect 326632 223038 326660 231676
rect 327000 225962 327028 231676
rect 327368 229566 327396 231676
rect 327356 229560 327408 229566
rect 327356 229502 327408 229508
rect 327736 228886 327764 231676
rect 327724 228880 327776 228886
rect 327724 228822 327776 228828
rect 328104 228750 328132 231676
rect 328472 229226 328500 231676
rect 328460 229220 328512 229226
rect 328460 229162 328512 229168
rect 328840 229158 328868 231676
rect 328828 229152 328880 229158
rect 328828 229094 328880 229100
rect 329208 228954 329236 231676
rect 329196 228948 329248 228954
rect 329196 228890 329248 228896
rect 328092 228744 328144 228750
rect 328092 228686 328144 228692
rect 327816 228472 327868 228478
rect 327816 228414 327868 228420
rect 327080 228404 327132 228410
rect 327080 228346 327132 228352
rect 326988 225956 327040 225962
rect 326988 225898 327040 225904
rect 326620 223032 326672 223038
rect 326620 222974 326672 222980
rect 326528 221672 326580 221678
rect 326528 221614 326580 221620
rect 326252 220720 326304 220726
rect 326252 220662 326304 220668
rect 326252 220244 326304 220250
rect 326252 220186 326304 220192
rect 326264 217410 326292 220186
rect 327092 217410 327120 228346
rect 327828 217410 327856 228414
rect 329484 227118 329512 231676
rect 329564 229220 329616 229226
rect 329564 229162 329616 229168
rect 329472 227112 329524 227118
rect 329472 227054 329524 227060
rect 328736 224324 328788 224330
rect 328736 224266 328788 224272
rect 328748 217410 328776 224266
rect 329576 220658 329604 229162
rect 329852 229158 329880 231676
rect 330234 231662 330524 231690
rect 329656 229152 329708 229158
rect 329656 229094 329708 229100
rect 329840 229152 329892 229158
rect 329840 229094 329892 229100
rect 329564 220652 329616 220658
rect 329564 220594 329616 220600
rect 329668 220590 329696 229094
rect 330392 227452 330444 227458
rect 330392 227394 330444 227400
rect 329656 220584 329708 220590
rect 329656 220526 329708 220532
rect 329840 220108 329892 220114
rect 329840 220050 329892 220056
rect 329852 217410 329880 220050
rect 330404 217410 330432 227394
rect 330496 220386 330524 231662
rect 330588 228818 330616 231676
rect 330576 228812 330628 228818
rect 330576 228754 330628 228760
rect 330956 223174 330984 231676
rect 331324 230450 331352 231676
rect 331312 230444 331364 230450
rect 331312 230386 331364 230392
rect 331692 229634 331720 231676
rect 331680 229628 331732 229634
rect 331680 229570 331732 229576
rect 331036 229152 331088 229158
rect 331036 229094 331088 229100
rect 330944 223168 330996 223174
rect 330944 223110 330996 223116
rect 331048 220454 331076 229094
rect 332060 229022 332088 231676
rect 332232 230444 332284 230450
rect 332232 230386 332284 230392
rect 332048 229016 332100 229022
rect 332048 228958 332100 228964
rect 331220 225684 331272 225690
rect 331220 225626 331272 225632
rect 331036 220448 331088 220454
rect 331036 220390 331088 220396
rect 330484 220380 330536 220386
rect 330484 220322 330536 220328
rect 331232 217870 331260 225626
rect 331312 224256 331364 224262
rect 331312 224198 331364 224204
rect 331220 217864 331272 217870
rect 331220 217806 331272 217812
rect 331324 217410 331352 224198
rect 332244 220318 332272 230386
rect 332336 224534 332364 231676
rect 332416 229628 332468 229634
rect 332416 229570 332468 229576
rect 332324 224528 332376 224534
rect 332324 224470 332376 224476
rect 332232 220312 332284 220318
rect 332232 220254 332284 220260
rect 332428 220250 332456 229570
rect 332704 229566 332732 231676
rect 333072 230450 333100 231676
rect 333454 231662 333652 231690
rect 333624 230518 333652 231662
rect 333716 231662 333822 231690
rect 333612 230512 333664 230518
rect 333612 230454 333664 230460
rect 333060 230444 333112 230450
rect 333060 230386 333112 230392
rect 332692 229560 332744 229566
rect 332692 229502 332744 229508
rect 333716 224466 333744 231662
rect 333888 230444 333940 230450
rect 333888 230386 333940 230392
rect 333796 229560 333848 229566
rect 333796 229502 333848 229508
rect 333704 224460 333756 224466
rect 333704 224402 333756 224408
rect 332416 220244 332468 220250
rect 332416 220186 332468 220192
rect 333808 220182 333836 229502
rect 332968 220176 333020 220182
rect 332968 220118 333020 220124
rect 333796 220176 333848 220182
rect 333796 220118 333848 220124
rect 332140 217864 332192 217870
rect 332140 217806 332192 217812
rect 332152 217410 332180 217806
rect 332980 217410 333008 220118
rect 333900 220114 333928 230386
rect 334176 228138 334204 231676
rect 334544 229430 334572 231676
rect 334624 230172 334676 230178
rect 334624 230114 334676 230120
rect 334532 229424 334584 229430
rect 334532 229366 334584 229372
rect 334164 228132 334216 228138
rect 334164 228074 334216 228080
rect 333980 227316 334032 227322
rect 333980 227258 334032 227264
rect 333888 220108 333940 220114
rect 333888 220050 333940 220056
rect 333992 217870 334020 227258
rect 334072 225616 334124 225622
rect 334072 225558 334124 225564
rect 333980 217864 334032 217870
rect 333980 217806 334032 217812
rect 334084 217410 334112 225558
rect 334636 219638 334664 230114
rect 334716 229764 334768 229770
rect 334716 229706 334768 229712
rect 334728 219706 334756 229706
rect 334912 228682 334940 231676
rect 334900 228676 334952 228682
rect 334900 228618 334952 228624
rect 335188 227322 335216 231676
rect 335176 227316 335228 227322
rect 335176 227258 335228 227264
rect 335556 224602 335584 231676
rect 335924 226098 335952 231676
rect 336292 228614 336320 231676
rect 336660 230178 336688 231676
rect 337042 231662 337332 231690
rect 337410 231662 337700 231690
rect 336648 230172 336700 230178
rect 336648 230114 336700 230120
rect 337016 230036 337068 230042
rect 337016 229978 337068 229984
rect 337028 229094 337056 229978
rect 337028 229066 337148 229094
rect 336280 228608 336332 228614
rect 336280 228550 336332 228556
rect 335912 226092 335964 226098
rect 335912 226034 335964 226040
rect 335544 224596 335596 224602
rect 335544 224538 335596 224544
rect 335544 221196 335596 221202
rect 335544 221138 335596 221144
rect 334716 219700 334768 219706
rect 334716 219642 334768 219648
rect 334624 219632 334676 219638
rect 334624 219574 334676 219580
rect 334716 217864 334768 217870
rect 334716 217806 334768 217812
rect 334728 217410 334756 217806
rect 335556 217410 335584 221138
rect 336740 220040 336792 220046
rect 336740 219982 336792 219988
rect 336752 217410 336780 219982
rect 321940 217382 322368 217410
rect 322952 217382 323288 217410
rect 323688 217382 324116 217410
rect 324516 217382 324944 217410
rect 325712 217382 325772 217410
rect 326264 217382 326600 217410
rect 327092 217382 327428 217410
rect 327828 217382 328256 217410
rect 328748 217382 329176 217410
rect 329852 217382 330004 217410
rect 330404 217382 330832 217410
rect 331324 217382 331660 217410
rect 332152 217382 332488 217410
rect 332980 217382 333316 217410
rect 334084 217382 334144 217410
rect 334728 217382 335064 217410
rect 335556 217382 335892 217410
rect 336720 217382 336780 217410
rect 337120 217410 337148 229066
rect 337304 223718 337332 231662
rect 337384 230240 337436 230246
rect 337384 230182 337436 230188
rect 337292 223712 337344 223718
rect 337292 223654 337344 223660
rect 337396 219774 337424 230182
rect 337672 222902 337700 231662
rect 337764 228546 337792 231676
rect 338040 229566 338068 231676
rect 338028 229560 338080 229566
rect 338028 229502 338080 229508
rect 337752 228540 337804 228546
rect 337752 228482 337804 228488
rect 338408 224126 338436 231676
rect 338790 231662 339080 231690
rect 338764 230376 338816 230382
rect 338764 230318 338816 230324
rect 338396 224120 338448 224126
rect 338396 224062 338448 224068
rect 338120 223100 338172 223106
rect 338120 223042 338172 223048
rect 337660 222896 337712 222902
rect 337660 222838 337712 222844
rect 337384 219768 337436 219774
rect 337384 219710 337436 219716
rect 338132 217410 338160 223042
rect 338776 219842 338804 230318
rect 339052 225214 339080 231662
rect 339144 230314 339172 231676
rect 339132 230308 339184 230314
rect 339132 230250 339184 230256
rect 339512 229498 339540 231676
rect 339500 229492 339552 229498
rect 339500 229434 339552 229440
rect 339040 225208 339092 225214
rect 339040 225150 339092 225156
rect 339880 224398 339908 231676
rect 340144 229696 340196 229702
rect 340144 229638 340196 229644
rect 339868 224392 339920 224398
rect 339868 224334 339920 224340
rect 338856 221264 338908 221270
rect 338856 221206 338908 221212
rect 338764 219836 338816 219842
rect 338764 219778 338816 219784
rect 338868 217410 338896 221206
rect 339684 220516 339736 220522
rect 339684 220458 339736 220464
rect 339696 217410 339724 220458
rect 340156 219978 340184 229638
rect 340248 225146 340276 231676
rect 340616 228206 340644 231676
rect 340892 229702 340920 231676
rect 341274 231662 341472 231690
rect 341248 229968 341300 229974
rect 341248 229910 341300 229916
rect 340880 229696 340932 229702
rect 340880 229638 340932 229644
rect 340604 228200 340656 228206
rect 340604 228142 340656 228148
rect 340236 225140 340288 225146
rect 340236 225082 340288 225088
rect 340144 219972 340196 219978
rect 340144 219914 340196 219920
rect 341260 217410 341288 229910
rect 341340 227384 341392 227390
rect 341340 227326 341392 227332
rect 337120 217382 337548 217410
rect 338132 217382 338376 217410
rect 338868 217382 339204 217410
rect 339696 217382 340032 217410
rect 340952 217382 341288 217410
rect 341352 217410 341380 227326
rect 341444 224330 341472 231662
rect 341524 229628 341576 229634
rect 341524 229570 341576 229576
rect 341432 224324 341484 224330
rect 341432 224266 341484 224272
rect 341536 220046 341564 229570
rect 341628 225690 341656 231676
rect 341996 230382 342024 231676
rect 341984 230376 342036 230382
rect 341984 230318 342036 230324
rect 342364 229362 342392 231676
rect 342352 229356 342404 229362
rect 342352 229298 342404 229304
rect 341616 225684 341668 225690
rect 341616 225626 341668 225632
rect 342732 224194 342760 231676
rect 342904 229424 342956 229430
rect 342904 229366 342956 229372
rect 342720 224188 342772 224194
rect 342720 224130 342772 224136
rect 342260 221332 342312 221338
rect 342260 221274 342312 221280
rect 341524 220040 341576 220046
rect 341524 219982 341576 219988
rect 342272 217410 342300 221274
rect 342916 220522 342944 229366
rect 343100 225758 343128 231676
rect 343272 229356 343324 229362
rect 343272 229298 343324 229304
rect 343088 225752 343140 225758
rect 343088 225694 343140 225700
rect 343284 221066 343312 229298
rect 343468 228070 343496 231676
rect 343744 230042 343772 231676
rect 343732 230036 343784 230042
rect 343732 229978 343784 229984
rect 343824 229288 343876 229294
rect 343824 229230 343876 229236
rect 343456 228064 343508 228070
rect 343456 228006 343508 228012
rect 343272 221060 343324 221066
rect 343272 221002 343324 221008
rect 342904 220516 342956 220522
rect 342904 220458 342956 220464
rect 343088 219904 343140 219910
rect 343088 219846 343140 219852
rect 343100 217410 343128 219846
rect 343836 217410 343864 229230
rect 344112 224262 344140 231676
rect 344480 225622 344508 231676
rect 344848 229770 344876 231676
rect 344836 229764 344888 229770
rect 344836 229706 344888 229712
rect 345216 228478 345244 231676
rect 345584 229974 345612 231676
rect 345572 229968 345624 229974
rect 345572 229910 345624 229916
rect 345204 228472 345256 228478
rect 345204 228414 345256 228420
rect 344468 225616 344520 225622
rect 344468 225558 344520 225564
rect 345952 225282 345980 231676
rect 346320 228410 346348 231676
rect 346492 229900 346544 229906
rect 346492 229842 346544 229848
rect 346308 228404 346360 228410
rect 346308 228346 346360 228352
rect 345940 225276 345992 225282
rect 345940 225218 345992 225224
rect 344100 224256 344152 224262
rect 344100 224198 344152 224204
rect 346504 224210 346532 229842
rect 346596 229094 346624 231676
rect 346596 229066 346716 229094
rect 346504 224182 346624 224210
rect 345020 222964 345072 222970
rect 345020 222906 345072 222912
rect 345032 217410 345060 222906
rect 345572 221400 345624 221406
rect 345572 221342 345624 221348
rect 345584 217410 345612 221342
rect 346492 219632 346544 219638
rect 346492 219574 346544 219580
rect 346504 217410 346532 219574
rect 346596 219434 346624 224182
rect 346688 222970 346716 229066
rect 346964 223854 346992 231676
rect 347332 223990 347360 231676
rect 347700 230246 347728 231676
rect 347688 230240 347740 230246
rect 347688 230182 347740 230188
rect 348068 229094 348096 231676
rect 348068 229066 348188 229094
rect 348056 227248 348108 227254
rect 348056 227190 348108 227196
rect 347320 223984 347372 223990
rect 347320 223926 347372 223932
rect 346952 223848 347004 223854
rect 346952 223790 347004 223796
rect 346676 222964 346728 222970
rect 346676 222906 346728 222912
rect 346596 219406 347268 219434
rect 347240 217410 347268 219406
rect 348068 217410 348096 227190
rect 348160 223106 348188 229066
rect 348436 223922 348464 231676
rect 348804 225350 348832 231676
rect 349172 228274 349200 231676
rect 349160 228268 349212 228274
rect 349160 228210 349212 228216
rect 348792 225344 348844 225350
rect 348792 225286 348844 225292
rect 348424 223916 348476 223922
rect 348424 223858 348476 223864
rect 348148 223100 348200 223106
rect 348148 223042 348200 223048
rect 349448 222426 349476 231676
rect 349816 224058 349844 231676
rect 349804 224052 349856 224058
rect 349804 223994 349856 224000
rect 349436 222420 349488 222426
rect 349436 222362 349488 222368
rect 349160 222148 349212 222154
rect 349160 222090 349212 222096
rect 349172 217410 349200 222090
rect 349804 219700 349856 219706
rect 349804 219642 349856 219648
rect 349816 217410 349844 219642
rect 350184 219434 350212 231676
rect 350552 229634 350580 231676
rect 350934 231662 351224 231690
rect 351302 231662 351592 231690
rect 350908 229832 350960 229838
rect 350908 229774 350960 229780
rect 350540 229628 350592 229634
rect 350540 229570 350592 229576
rect 350632 223236 350684 223242
rect 350632 223178 350684 223184
rect 350172 219428 350224 219434
rect 350172 219370 350224 219376
rect 350644 217870 350672 223178
rect 350632 217864 350684 217870
rect 350632 217806 350684 217812
rect 350920 217410 350948 229774
rect 351196 222494 351224 231662
rect 351184 222488 351236 222494
rect 351184 222430 351236 222436
rect 351564 221202 351592 231662
rect 351656 226574 351684 231676
rect 352024 229906 352052 231676
rect 352012 229900 352064 229906
rect 352012 229842 352064 229848
rect 351644 226568 351696 226574
rect 351644 226510 351696 226516
rect 352300 223446 352328 231676
rect 352564 229560 352616 229566
rect 352564 229502 352616 229508
rect 352288 223440 352340 223446
rect 352288 223382 352340 223388
rect 352576 221542 352604 229502
rect 352668 222562 352696 231676
rect 353050 231662 353248 231690
rect 352656 222556 352708 222562
rect 352656 222498 352708 222504
rect 352380 221536 352432 221542
rect 352380 221478 352432 221484
rect 352564 221536 352616 221542
rect 352564 221478 352616 221484
rect 351552 221196 351604 221202
rect 351552 221138 351604 221144
rect 351460 217864 351512 217870
rect 351460 217806 351512 217812
rect 351472 217410 351500 217806
rect 352392 217410 352420 221478
rect 353220 219298 353248 231662
rect 353404 228342 353432 231676
rect 353392 228336 353444 228342
rect 353392 228278 353444 228284
rect 353772 222630 353800 231676
rect 354154 231662 354444 231690
rect 353944 229492 353996 229498
rect 353944 229434 353996 229440
rect 353760 222624 353812 222630
rect 353760 222566 353812 222572
rect 353956 221338 353984 229434
rect 354036 221468 354088 221474
rect 354036 221410 354088 221416
rect 353944 221332 353996 221338
rect 353944 221274 353996 221280
rect 353300 219768 353352 219774
rect 353300 219710 353352 219716
rect 353208 219292 353260 219298
rect 353208 219234 353260 219240
rect 353312 217410 353340 219710
rect 354048 217410 354076 221410
rect 354416 219366 354444 231662
rect 354508 226642 354536 231676
rect 354772 229968 354824 229974
rect 354772 229910 354824 229916
rect 354784 229094 354812 229910
rect 354876 229566 354904 231676
rect 354864 229560 354916 229566
rect 354864 229502 354916 229508
rect 354784 229066 354904 229094
rect 354772 227180 354824 227186
rect 354772 227122 354824 227128
rect 354496 226636 354548 226642
rect 354496 226578 354548 226584
rect 354404 219360 354456 219366
rect 354404 219302 354456 219308
rect 354784 217410 354812 227122
rect 354876 223786 354904 229066
rect 354864 223780 354916 223786
rect 354864 223722 354916 223728
rect 355152 222698 355180 231676
rect 355520 229498 355548 231676
rect 355508 229492 355560 229498
rect 355508 229434 355560 229440
rect 355888 226710 355916 231676
rect 356256 229974 356284 231676
rect 356244 229968 356296 229974
rect 356244 229910 356296 229916
rect 355876 226704 355928 226710
rect 355876 226646 355928 226652
rect 356624 222766 356652 231676
rect 356992 225894 357020 231676
rect 357072 229968 357124 229974
rect 357072 229910 357124 229916
rect 356980 225888 357032 225894
rect 356980 225830 357032 225836
rect 356612 222760 356664 222766
rect 356612 222702 356664 222708
rect 355140 222692 355192 222698
rect 355140 222634 355192 222640
rect 356060 222080 356112 222086
rect 356060 222022 356112 222028
rect 356072 217410 356100 222022
rect 357084 221270 357112 229910
rect 357360 226778 357388 231676
rect 357728 229294 357756 231676
rect 357716 229288 357768 229294
rect 357716 229230 357768 229236
rect 357348 226772 357400 226778
rect 357348 226714 357400 226720
rect 358004 222834 358032 231676
rect 358176 226024 358228 226030
rect 358176 225966 358228 225972
rect 357992 222828 358044 222834
rect 357992 222770 358044 222776
rect 357532 222012 357584 222018
rect 357532 221954 357584 221960
rect 357072 221264 357124 221270
rect 357072 221206 357124 221212
rect 356520 219836 356572 219842
rect 356520 219778 356572 219784
rect 341352 217382 341780 217410
rect 342272 217382 342608 217410
rect 343100 217382 343436 217410
rect 343836 217382 344264 217410
rect 345032 217382 345092 217410
rect 345584 217382 345920 217410
rect 346504 217382 346840 217410
rect 347240 217382 347668 217410
rect 348068 217382 348496 217410
rect 349172 217382 349324 217410
rect 349816 217382 350152 217410
rect 350920 217382 350980 217410
rect 351472 217382 351808 217410
rect 352392 217382 352728 217410
rect 353312 217382 353556 217410
rect 354048 217382 354384 217410
rect 354784 217382 355212 217410
rect 356040 217382 356100 217410
rect 356532 217410 356560 219778
rect 357544 217410 357572 221954
rect 358188 217410 358216 225966
rect 358372 225418 358400 231676
rect 358740 227662 358768 231676
rect 359108 229974 359136 231676
rect 359096 229968 359148 229974
rect 359096 229910 359148 229916
rect 358728 227656 358780 227662
rect 358728 227598 358780 227604
rect 358360 225412 358412 225418
rect 358360 225354 358412 225360
rect 359476 223582 359504 231676
rect 359844 225486 359872 231676
rect 360108 229968 360160 229974
rect 360108 229910 360160 229916
rect 359832 225480 359884 225486
rect 359832 225422 359884 225428
rect 359464 223576 359516 223582
rect 359464 223518 359516 223524
rect 359096 221944 359148 221950
rect 359096 221886 359148 221892
rect 359108 217410 359136 221886
rect 360120 221338 360148 229910
rect 360212 226846 360240 231676
rect 360580 229974 360608 231676
rect 360870 231662 361160 231690
rect 360568 229968 360620 229974
rect 360568 229910 360620 229916
rect 360292 227044 360344 227050
rect 360292 226986 360344 226992
rect 360200 226840 360252 226846
rect 360200 226782 360252 226788
rect 360108 221332 360160 221338
rect 360108 221274 360160 221280
rect 360200 219972 360252 219978
rect 360200 219914 360252 219920
rect 360212 217410 360240 219914
rect 360304 219502 360332 226986
rect 361132 223514 361160 231662
rect 361224 229430 361252 231676
rect 361304 229968 361356 229974
rect 361304 229910 361356 229916
rect 361212 229424 361264 229430
rect 361212 229366 361264 229372
rect 361120 223508 361172 223514
rect 361120 223450 361172 223456
rect 360752 221876 360804 221882
rect 360752 221818 360804 221824
rect 360292 219496 360344 219502
rect 360292 219438 360344 219444
rect 360764 217410 360792 221818
rect 361316 221406 361344 229910
rect 361592 226914 361620 231676
rect 361960 229974 361988 231676
rect 361948 229968 362000 229974
rect 361948 229910 362000 229916
rect 362328 229838 362356 231676
rect 362710 231662 362908 231690
rect 362684 229968 362736 229974
rect 362684 229910 362736 229916
rect 362316 229832 362368 229838
rect 362316 229774 362368 229780
rect 361580 226908 361632 226914
rect 361580 226850 361632 226856
rect 361580 225820 361632 225826
rect 361580 225762 361632 225768
rect 361304 221400 361356 221406
rect 361304 221342 361356 221348
rect 361592 217410 361620 225762
rect 362696 222154 362724 229910
rect 362880 225554 362908 231662
rect 363064 226982 363092 231676
rect 363432 229362 363460 231676
rect 363722 231662 364012 231690
rect 363420 229356 363472 229362
rect 363420 229298 363472 229304
rect 363144 227316 363196 227322
rect 363144 227258 363196 227264
rect 363052 226976 363104 226982
rect 363052 226918 363104 226924
rect 362960 225956 363012 225962
rect 362960 225898 363012 225904
rect 362868 225548 362920 225554
rect 362868 225490 362920 225496
rect 362684 222148 362736 222154
rect 362684 222090 362736 222096
rect 362408 221808 362460 221814
rect 362408 221750 362460 221756
rect 362420 217410 362448 221750
rect 362972 219842 363000 225898
rect 363156 219910 363184 227258
rect 363984 222018 364012 231662
rect 364076 226302 364104 231676
rect 364248 229968 364300 229974
rect 364168 229916 364248 229922
rect 364168 229910 364300 229916
rect 364168 229894 364288 229910
rect 364168 229838 364196 229894
rect 364156 229832 364208 229838
rect 364156 229774 364208 229780
rect 364248 229832 364300 229838
rect 364248 229774 364300 229780
rect 364260 229566 364288 229774
rect 364248 229560 364300 229566
rect 364248 229502 364300 229508
rect 364156 229356 364208 229362
rect 364156 229298 364208 229304
rect 364064 226296 364116 226302
rect 364064 226238 364116 226244
rect 364168 222086 364196 229298
rect 364444 227730 364472 231676
rect 364826 231662 365116 231690
rect 364524 230104 364576 230110
rect 364524 230046 364576 230052
rect 364432 227724 364484 227730
rect 364432 227666 364484 227672
rect 364156 222080 364208 222086
rect 364156 222022 364208 222028
rect 363972 222012 364024 222018
rect 363972 221954 364024 221960
rect 363236 220788 363288 220794
rect 363236 220730 363288 220736
rect 363144 219904 363196 219910
rect 363144 219846 363196 219852
rect 362960 219836 363012 219842
rect 362960 219778 363012 219784
rect 363248 217410 363276 220730
rect 364536 217410 364564 230046
rect 365088 221950 365116 231662
rect 365180 229090 365208 231676
rect 365168 229084 365220 229090
rect 365168 229026 365220 229032
rect 365260 227112 365312 227118
rect 365260 227054 365312 227060
rect 365076 221944 365128 221950
rect 365076 221886 365128 221892
rect 365272 219978 365300 227054
rect 365548 226234 365576 231676
rect 365916 227594 365944 231676
rect 366298 231662 366496 231690
rect 365904 227588 365956 227594
rect 365904 227530 365956 227536
rect 365536 226228 365588 226234
rect 365536 226170 365588 226176
rect 366468 221882 366496 231662
rect 366560 229566 366588 231676
rect 366548 229560 366600 229566
rect 366548 229502 366600 229508
rect 366928 226166 366956 231676
rect 367296 227526 367324 231676
rect 367678 231662 367968 231690
rect 367284 227520 367336 227526
rect 367284 227462 367336 227468
rect 366916 226160 366968 226166
rect 366916 226102 366968 226108
rect 367652 226092 367704 226098
rect 367652 226034 367704 226040
rect 367008 223168 367060 223174
rect 367008 223110 367060 223116
rect 366456 221876 366508 221882
rect 366456 221818 366508 221824
rect 365812 221740 365864 221746
rect 365812 221682 365864 221688
rect 365260 219972 365312 219978
rect 365260 219914 365312 219920
rect 364984 219496 365036 219502
rect 364984 219438 365036 219444
rect 356532 217382 356868 217410
rect 357544 217382 357696 217410
rect 358188 217382 358616 217410
rect 359108 217382 359444 217410
rect 360212 217382 360272 217410
rect 360764 217382 361100 217410
rect 361592 217382 361928 217410
rect 362420 217382 362756 217410
rect 363248 217382 363584 217410
rect 364504 217382 364564 217410
rect 364996 217410 365024 219438
rect 365824 217410 365852 221682
rect 367020 220794 367048 223110
rect 367468 221604 367520 221610
rect 367468 221546 367520 221552
rect 367008 220788 367060 220794
rect 367008 220730 367060 220736
rect 366640 220720 366692 220726
rect 366640 220662 366692 220668
rect 366652 217410 366680 220662
rect 367480 217410 367508 221546
rect 367664 220726 367692 226034
rect 367940 221814 367968 231662
rect 368032 224942 368060 231676
rect 368400 226098 368428 231676
rect 368768 227458 368796 231676
rect 369150 231662 369348 231690
rect 368756 227452 368808 227458
rect 368756 227394 368808 227400
rect 368388 226092 368440 226098
rect 368388 226034 368440 226040
rect 368020 224936 368072 224942
rect 368020 224878 368072 224884
rect 367928 221808 367980 221814
rect 367928 221750 367980 221756
rect 369320 221746 369348 231662
rect 369412 229226 369440 231676
rect 369400 229220 369452 229226
rect 369400 229162 369452 229168
rect 369780 226030 369808 231676
rect 370148 227390 370176 231676
rect 370530 231662 370820 231690
rect 370228 229016 370280 229022
rect 370228 228958 370280 228964
rect 370136 227384 370188 227390
rect 370136 227326 370188 227332
rect 369768 226024 369820 226030
rect 369768 225966 369820 225972
rect 369308 221740 369360 221746
rect 369308 221682 369360 221688
rect 369124 221672 369176 221678
rect 369124 221614 369176 221620
rect 367652 220720 367704 220726
rect 367652 220662 367704 220668
rect 368480 219836 368532 219842
rect 368480 219778 368532 219784
rect 368492 217410 368520 219778
rect 369136 217410 369164 221614
rect 370240 220046 370268 228958
rect 370792 221678 370820 231662
rect 370884 224806 370912 231676
rect 371252 225962 371280 231676
rect 371332 228948 371384 228954
rect 371332 228890 371384 228896
rect 371240 225956 371292 225962
rect 371240 225898 371292 225904
rect 370872 224800 370924 224806
rect 370872 224742 370924 224748
rect 371240 223032 371292 223038
rect 371240 222974 371292 222980
rect 370780 221672 370832 221678
rect 370780 221614 370832 221620
rect 370044 220040 370096 220046
rect 370044 219982 370096 219988
rect 370228 220040 370280 220046
rect 370228 219982 370280 219988
rect 370056 217410 370084 219982
rect 371252 217410 371280 222974
rect 371344 219502 371372 228890
rect 371620 227322 371648 231676
rect 371884 230444 371936 230450
rect 371884 230386 371936 230392
rect 371608 227316 371660 227322
rect 371608 227258 371660 227264
rect 371896 220658 371924 230386
rect 371988 229362 372016 231676
rect 371976 229356 372028 229362
rect 371976 229298 372028 229304
rect 372264 224738 372292 231676
rect 372632 225826 372660 231676
rect 372712 228880 372764 228886
rect 372712 228822 372764 228828
rect 372620 225820 372672 225826
rect 372620 225762 372672 225768
rect 372252 224732 372304 224738
rect 372252 224674 372304 224680
rect 372620 224528 372672 224534
rect 372620 224470 372672 224476
rect 371700 220652 371752 220658
rect 371700 220594 371752 220600
rect 371884 220652 371936 220658
rect 371884 220594 371936 220600
rect 371332 219496 371384 219502
rect 371332 219438 371384 219444
rect 364996 217382 365332 217410
rect 365824 217382 366160 217410
rect 366652 217382 366988 217410
rect 367480 217382 367816 217410
rect 368492 217382 368644 217410
rect 369136 217382 369472 217410
rect 370056 217382 370392 217410
rect 371220 217382 371280 217410
rect 371712 217410 371740 220594
rect 372632 219774 372660 224470
rect 372620 219768 372672 219774
rect 372620 219710 372672 219716
rect 372724 217410 372752 228822
rect 373000 227254 373028 231676
rect 373368 229022 373396 231676
rect 373356 229016 373408 229022
rect 373356 228958 373408 228964
rect 372988 227248 373040 227254
rect 372988 227190 373040 227196
rect 373736 224670 373764 231676
rect 374104 230382 374132 231676
rect 374092 230376 374144 230382
rect 374092 230318 374144 230324
rect 374092 228744 374144 228750
rect 374092 228686 374144 228692
rect 373724 224664 373776 224670
rect 373724 224606 373776 224612
rect 373356 220584 373408 220590
rect 373356 220526 373408 220532
rect 373368 217410 373396 220526
rect 374104 217410 374132 228686
rect 374472 227186 374500 231676
rect 374460 227180 374512 227186
rect 374460 227122 374512 227128
rect 374840 227118 374868 231676
rect 375116 228954 375144 231676
rect 375104 228948 375156 228954
rect 375104 228890 375156 228896
rect 375288 228812 375340 228818
rect 375288 228754 375340 228760
rect 374828 227112 374880 227118
rect 374828 227054 374880 227060
rect 375300 219842 375328 228754
rect 375484 227866 375512 231676
rect 375852 230081 375880 231676
rect 376024 230172 376076 230178
rect 376024 230114 376076 230120
rect 375838 230072 375894 230081
rect 375838 230007 375894 230016
rect 375472 227860 375524 227866
rect 375472 227802 375524 227808
rect 376036 220454 376064 230114
rect 376116 229288 376168 229294
rect 376116 229230 376168 229236
rect 376128 221134 376156 229230
rect 376220 223281 376248 231676
rect 376588 228886 376616 231676
rect 376956 230353 376984 231676
rect 376942 230344 376998 230353
rect 376942 230279 376998 230288
rect 376576 228880 376628 228886
rect 376576 228822 376628 228828
rect 377324 227798 377352 231676
rect 377404 230376 377456 230382
rect 377404 230318 377456 230324
rect 377312 227792 377364 227798
rect 377312 227734 377364 227740
rect 377416 224874 377444 230318
rect 377404 224868 377456 224874
rect 377404 224810 377456 224816
rect 377692 224777 377720 231676
rect 377968 228818 377996 231676
rect 378232 230308 378284 230314
rect 378232 230250 378284 230256
rect 377956 228812 378008 228818
rect 377956 228754 378008 228760
rect 378244 227934 378272 230250
rect 378336 230178 378364 231676
rect 378324 230172 378376 230178
rect 378324 230114 378376 230120
rect 378704 229945 378732 231676
rect 378690 229936 378746 229945
rect 378690 229871 378746 229880
rect 378508 228132 378560 228138
rect 378508 228074 378560 228080
rect 378232 227928 378284 227934
rect 378232 227870 378284 227876
rect 377678 224768 377734 224777
rect 377678 224703 377734 224712
rect 377312 224596 377364 224602
rect 377312 224538 377364 224544
rect 376206 223272 376262 223281
rect 376206 223207 376262 223216
rect 376116 221128 376168 221134
rect 376116 221070 376168 221076
rect 375380 220448 375432 220454
rect 375380 220390 375432 220396
rect 376024 220448 376076 220454
rect 376024 220390 376076 220396
rect 375288 219836 375340 219842
rect 375288 219778 375340 219784
rect 375392 217410 375420 220390
rect 376944 220380 376996 220386
rect 376944 220322 376996 220328
rect 375932 219496 375984 219502
rect 375932 219438 375984 219444
rect 371712 217382 372048 217410
rect 372724 217382 372876 217410
rect 373368 217382 373704 217410
rect 374104 217382 374532 217410
rect 375360 217382 375420 217410
rect 375944 217410 375972 219438
rect 376956 217410 376984 220322
rect 377324 219638 377352 224538
rect 378048 224460 378100 224466
rect 378048 224402 378100 224408
rect 378060 220386 378088 224402
rect 378048 220380 378100 220386
rect 378048 220322 378100 220328
rect 378416 220312 378468 220318
rect 378416 220254 378468 220260
rect 377588 219972 377640 219978
rect 377588 219914 377640 219920
rect 377312 219632 377364 219638
rect 377312 219574 377364 219580
rect 377600 217410 377628 219914
rect 378428 217410 378456 220254
rect 378520 219502 378548 228074
rect 378784 223712 378836 223718
rect 378784 223654 378836 223660
rect 378796 220318 378824 223654
rect 379072 223145 379100 231676
rect 379058 223136 379114 223145
rect 379058 223071 379114 223080
rect 378784 220312 378836 220318
rect 378784 220254 378836 220260
rect 378508 219496 378560 219502
rect 378508 219438 378560 219444
rect 379440 219230 379468 231676
rect 379520 229492 379572 229498
rect 379520 229434 379572 229440
rect 379532 229378 379560 229434
rect 379532 229350 379744 229378
rect 379716 229294 379744 229350
rect 379704 229288 379756 229294
rect 379704 229230 379756 229236
rect 379808 223038 379836 231676
rect 380176 229809 380204 231676
rect 380162 229800 380218 229809
rect 380162 229735 380218 229744
rect 380256 229696 380308 229702
rect 380256 229638 380308 229644
rect 379796 223032 379848 223038
rect 379796 222974 379848 222980
rect 380268 220930 380296 229638
rect 380348 227792 380400 227798
rect 380348 227734 380400 227740
rect 380256 220924 380308 220930
rect 380256 220866 380308 220872
rect 380360 220425 380388 227734
rect 380544 227361 380572 231676
rect 380716 230444 380768 230450
rect 380716 230386 380768 230392
rect 380728 228138 380756 230386
rect 380716 228132 380768 228138
rect 380716 228074 380768 228080
rect 380530 227352 380586 227361
rect 380530 227287 380586 227296
rect 380716 224120 380768 224126
rect 380716 224062 380768 224068
rect 380346 220416 380402 220425
rect 380346 220351 380402 220360
rect 380728 220250 380756 224062
rect 380072 220244 380124 220250
rect 380072 220186 380124 220192
rect 380716 220244 380768 220250
rect 380716 220186 380768 220192
rect 379520 219836 379572 219842
rect 379520 219778 379572 219784
rect 379428 219224 379480 219230
rect 379428 219166 379480 219172
rect 379532 217410 379560 219778
rect 380084 217410 380112 220186
rect 380820 219162 380848 231676
rect 381188 229158 381216 231676
rect 381556 230217 381584 231676
rect 381542 230208 381598 230217
rect 381542 230143 381598 230152
rect 381176 229152 381228 229158
rect 381176 229094 381228 229100
rect 380992 227860 381044 227866
rect 380992 227802 381044 227808
rect 380900 220788 380952 220794
rect 380900 220730 380952 220736
rect 380808 219156 380860 219162
rect 380808 219098 380860 219104
rect 380912 217410 380940 220730
rect 381004 219842 381032 227802
rect 381924 224641 381952 231676
rect 382096 229492 382148 229498
rect 382096 229434 382148 229440
rect 382108 229226 382136 229434
rect 382292 229226 382320 231676
rect 382464 229424 382516 229430
rect 382464 229366 382516 229372
rect 382096 229220 382148 229226
rect 382096 229162 382148 229168
rect 382280 229220 382332 229226
rect 382280 229162 382332 229168
rect 382188 229152 382240 229158
rect 382188 229094 382240 229100
rect 381910 224632 381966 224641
rect 381910 224567 381966 224576
rect 382200 220289 382228 229094
rect 382476 225214 382504 229366
rect 382660 229158 382688 231676
rect 382648 229152 382700 229158
rect 382648 229094 382700 229100
rect 383028 227225 383056 231676
rect 383410 231662 383608 231690
rect 383476 229220 383528 229226
rect 383476 229162 383528 229168
rect 383384 229152 383436 229158
rect 383384 229094 383436 229100
rect 383014 227216 383070 227225
rect 383014 227151 383070 227160
rect 382280 225208 382332 225214
rect 382280 225150 382332 225156
rect 382464 225208 382516 225214
rect 382464 225150 382516 225156
rect 382186 220280 382242 220289
rect 382186 220215 382242 220224
rect 382292 220182 382320 225150
rect 381820 220176 381872 220182
rect 381820 220118 381872 220124
rect 382280 220176 382332 220182
rect 382280 220118 382332 220124
rect 380992 219836 381044 219842
rect 380992 219778 381044 219784
rect 381832 217410 381860 220118
rect 383396 220046 383424 229094
rect 382648 220040 382700 220046
rect 382648 219982 382700 219988
rect 383384 220040 383436 220046
rect 383384 219982 383436 219988
rect 382660 217410 382688 219982
rect 383488 219094 383516 229162
rect 383476 219088 383528 219094
rect 383476 219030 383528 219036
rect 383580 219026 383608 231662
rect 383672 229158 383700 231676
rect 383660 229152 383712 229158
rect 383660 229094 383712 229100
rect 384040 224505 384068 231676
rect 384408 229294 384436 231676
rect 384790 231662 384896 231690
rect 384396 229288 384448 229294
rect 384396 229230 384448 229236
rect 384026 224496 384082 224505
rect 384026 224431 384082 224440
rect 384868 220153 384896 231662
rect 385144 230518 385172 231676
rect 385132 230512 385184 230518
rect 385132 230454 385184 230460
rect 385512 229158 385540 231676
rect 385684 230036 385736 230042
rect 385684 229978 385736 229984
rect 384948 229152 385000 229158
rect 384948 229094 385000 229100
rect 385500 229152 385552 229158
rect 385500 229094 385552 229100
rect 384854 220144 384910 220153
rect 383660 220108 383712 220114
rect 384854 220079 384910 220088
rect 383660 220050 383712 220056
rect 383568 219020 383620 219026
rect 383568 218962 383620 218968
rect 383672 217410 383700 220050
rect 384960 219978 384988 229094
rect 385500 225140 385552 225146
rect 385500 225082 385552 225088
rect 385512 220114 385540 225082
rect 385696 220998 385724 229978
rect 385880 223174 385908 231676
rect 386248 226001 386276 231676
rect 386420 230240 386472 230246
rect 386420 230182 386472 230188
rect 386328 229152 386380 229158
rect 386328 229094 386380 229100
rect 386234 225992 386290 226001
rect 386234 225927 386290 225936
rect 385868 223168 385920 223174
rect 385868 223110 385920 223116
rect 385684 220992 385736 220998
rect 385684 220934 385736 220940
rect 385960 220652 386012 220658
rect 385960 220594 386012 220600
rect 385500 220108 385552 220114
rect 385500 220050 385552 220056
rect 384948 219972 385000 219978
rect 384948 219914 385000 219920
rect 384304 219768 384356 219774
rect 384304 219710 384356 219716
rect 384316 217410 384344 219710
rect 385132 219496 385184 219502
rect 385132 219438 385184 219444
rect 385144 217410 385172 219438
rect 385972 217410 386000 220594
rect 386340 218958 386368 229094
rect 386432 228002 386460 230182
rect 386524 229158 386552 231676
rect 386892 229226 386920 231676
rect 386604 229220 386656 229226
rect 386604 229162 386656 229168
rect 386880 229220 386932 229226
rect 386880 229162 386932 229168
rect 386512 229152 386564 229158
rect 386512 229094 386564 229100
rect 386420 227996 386472 228002
rect 386420 227938 386472 227944
rect 386616 225146 386644 229162
rect 387260 228721 387288 231676
rect 387628 230042 387656 231676
rect 387996 230110 388024 231676
rect 387984 230104 388036 230110
rect 387984 230046 388036 230052
rect 387616 230036 387668 230042
rect 387616 229978 387668 229984
rect 387800 229628 387852 229634
rect 387800 229570 387852 229576
rect 387708 229152 387760 229158
rect 387708 229094 387760 229100
rect 387246 228712 387302 228721
rect 387246 228647 387302 228656
rect 387156 228064 387208 228070
rect 387156 228006 387208 228012
rect 386604 225140 386656 225146
rect 386604 225082 386656 225088
rect 386420 224392 386472 224398
rect 386420 224334 386472 224340
rect 386432 219706 386460 224334
rect 386788 220516 386840 220522
rect 386788 220458 386840 220464
rect 386420 219700 386472 219706
rect 386420 219642 386472 219648
rect 386328 218952 386380 218958
rect 386328 218894 386380 218900
rect 386800 217410 386828 220458
rect 387168 219774 387196 228006
rect 387156 219768 387208 219774
rect 387156 219710 387208 219716
rect 387720 218890 387748 229094
rect 387812 228070 387840 229570
rect 387800 228064 387852 228070
rect 387800 228006 387852 228012
rect 388364 227089 388392 231676
rect 388444 229220 388496 229226
rect 388444 229162 388496 229168
rect 388350 227080 388406 227089
rect 388350 227015 388406 227024
rect 387800 223168 387852 223174
rect 387800 223110 387852 223116
rect 387812 220794 387840 223110
rect 387800 220788 387852 220794
rect 387800 220730 387852 220736
rect 388456 220658 388484 229162
rect 388732 224602 388760 231676
rect 388720 224596 388772 224602
rect 388720 224538 388772 224544
rect 389100 223378 389128 231676
rect 389272 228676 389324 228682
rect 389272 228618 389324 228624
rect 389088 223372 389140 223378
rect 389088 223314 389140 223320
rect 389180 223032 389232 223038
rect 389180 222974 389232 222980
rect 388444 220652 388496 220658
rect 388444 220594 388496 220600
rect 389192 220561 389220 222974
rect 389178 220552 389234 220561
rect 389178 220487 389234 220496
rect 387800 220380 387852 220386
rect 387800 220322 387852 220328
rect 387708 218884 387760 218890
rect 387708 218826 387760 218832
rect 387812 217410 387840 220322
rect 388536 219632 388588 219638
rect 388536 219574 388588 219580
rect 388548 217410 388576 219574
rect 389284 217410 389312 228618
rect 389376 223009 389404 231676
rect 389744 224534 389772 231676
rect 390112 229226 390140 231676
rect 390100 229220 390152 229226
rect 390100 229162 390152 229168
rect 389732 224528 389784 224534
rect 389732 224470 389784 224476
rect 389362 223000 389418 223009
rect 389362 222935 389418 222944
rect 390480 222873 390508 231676
rect 390848 230382 390876 231676
rect 391230 231662 391520 231690
rect 390836 230376 390888 230382
rect 390836 230318 390888 230324
rect 390652 222896 390704 222902
rect 390466 222864 390522 222873
rect 390652 222838 390704 222844
rect 390466 222799 390522 222808
rect 390560 220720 390612 220726
rect 390560 220662 390612 220668
rect 390572 217410 390600 220662
rect 390664 219502 390692 222838
rect 391492 220522 391520 231662
rect 391584 223242 391612 231676
rect 391848 230376 391900 230382
rect 391848 230318 391900 230324
rect 391572 223236 391624 223242
rect 391572 223178 391624 223184
rect 391480 220516 391532 220522
rect 391480 220458 391532 220464
rect 391020 219904 391072 219910
rect 391020 219846 391072 219852
rect 390652 219496 390704 219502
rect 390652 219438 390704 219444
rect 375944 217382 376280 217410
rect 376956 217382 377108 217410
rect 377600 217382 377936 217410
rect 378428 217382 378764 217410
rect 379532 217382 379592 217410
rect 380084 217382 380420 217410
rect 380912 217382 381248 217410
rect 381832 217382 382168 217410
rect 382660 217382 382996 217410
rect 383672 217382 383824 217410
rect 384316 217382 384652 217410
rect 385144 217382 385480 217410
rect 385972 217382 386308 217410
rect 386800 217382 387136 217410
rect 387812 217382 388056 217410
rect 388548 217382 388884 217410
rect 389284 217382 389712 217410
rect 390540 217382 390600 217410
rect 391032 217410 391060 219846
rect 391860 218822 391888 230318
rect 391952 228750 391980 231676
rect 392228 229430 392256 231676
rect 392610 231662 392900 231690
rect 392216 229424 392268 229430
rect 392216 229366 392268 229372
rect 391940 228744 391992 228750
rect 391940 228686 391992 228692
rect 392584 228608 392636 228614
rect 392584 228550 392636 228556
rect 391940 220312 391992 220318
rect 391940 220254 391992 220260
rect 391848 218816 391900 218822
rect 391848 218758 391900 218764
rect 391952 217410 391980 220254
rect 392596 217410 392624 228550
rect 392872 221785 392900 231662
rect 392964 228682 392992 231676
rect 393332 230382 393360 231676
rect 393700 230450 393728 231676
rect 393688 230444 393740 230450
rect 393688 230386 393740 230392
rect 393320 230376 393372 230382
rect 393320 230318 393372 230324
rect 393412 229492 393464 229498
rect 393412 229434 393464 229440
rect 392952 228676 393004 228682
rect 392952 228618 393004 228624
rect 393424 224126 393452 229434
rect 394068 225865 394096 231676
rect 394450 231662 394556 231690
rect 394054 225856 394110 225865
rect 394054 225791 394110 225800
rect 393412 224120 393464 224126
rect 393412 224062 393464 224068
rect 392858 221776 392914 221785
rect 392858 221711 392914 221720
rect 394528 220386 394556 231662
rect 394608 230376 394660 230382
rect 394608 230318 394660 230324
rect 394620 220454 394648 230318
rect 394804 223038 394832 231676
rect 395094 231662 395384 231690
rect 395356 229378 395384 231662
rect 395448 230314 395476 231676
rect 395436 230308 395488 230314
rect 395436 230250 395488 230256
rect 395356 229350 395476 229378
rect 395448 229226 395476 229350
rect 395344 229220 395396 229226
rect 395344 229162 395396 229168
rect 395436 229220 395488 229226
rect 395436 229162 395488 229168
rect 394792 223032 394844 223038
rect 394792 222974 394844 222980
rect 395356 220590 395384 229162
rect 395816 229094 395844 231676
rect 396198 231662 396488 231690
rect 396566 231662 396856 231690
rect 396934 231662 397224 231690
rect 395816 229066 396028 229094
rect 395712 223372 395764 223378
rect 395712 223314 395764 223320
rect 395724 220726 395752 223314
rect 396000 223242 396028 229066
rect 396172 228540 396224 228546
rect 396172 228482 396224 228488
rect 395988 223236 396040 223242
rect 395988 223178 396040 223184
rect 395712 220720 395764 220726
rect 395712 220662 395764 220668
rect 394700 220584 394752 220590
rect 394700 220526 394752 220532
rect 395344 220584 395396 220590
rect 395344 220526 395396 220532
rect 394608 220448 394660 220454
rect 394608 220390 394660 220396
rect 394516 220380 394568 220386
rect 394516 220322 394568 220328
rect 393596 219496 393648 219502
rect 393596 219438 393648 219444
rect 393608 217410 393636 219438
rect 394712 217410 394740 220526
rect 395252 220244 395304 220250
rect 395252 220186 395304 220192
rect 395264 217410 395292 220186
rect 396184 217410 396212 228482
rect 396460 225729 396488 231662
rect 396724 230308 396776 230314
rect 396724 230250 396776 230256
rect 396446 225720 396502 225729
rect 396446 225655 396502 225664
rect 396736 220318 396764 230250
rect 396724 220312 396776 220318
rect 396724 220254 396776 220260
rect 396828 220250 396856 231662
rect 397196 221649 397224 231662
rect 397288 228614 397316 231676
rect 397656 230382 397684 231676
rect 397644 230376 397696 230382
rect 397644 230318 397696 230324
rect 397276 228608 397328 228614
rect 397276 228550 397328 228556
rect 397932 223174 397960 231676
rect 398104 230240 398156 230246
rect 398104 230182 398156 230188
rect 398116 229906 398144 230182
rect 398104 229900 398156 229906
rect 398104 229842 398156 229848
rect 398104 229628 398156 229634
rect 398104 229570 398156 229576
rect 398116 229362 398144 229570
rect 398104 229356 398156 229362
rect 398104 229298 398156 229304
rect 398300 228546 398328 231676
rect 398564 230376 398616 230382
rect 398564 230318 398616 230324
rect 398288 228540 398340 228546
rect 398288 228482 398340 228488
rect 398288 223304 398340 223310
rect 398288 223246 398340 223252
rect 397920 223168 397972 223174
rect 397920 223110 397972 223116
rect 398300 223038 398328 223246
rect 398288 223032 398340 223038
rect 398288 222974 398340 222980
rect 397182 221640 397238 221649
rect 397182 221575 397238 221584
rect 397736 221536 397788 221542
rect 397736 221478 397788 221484
rect 396816 220244 396868 220250
rect 396816 220186 396868 220192
rect 396908 220176 396960 220182
rect 396908 220118 396960 220124
rect 396920 217410 396948 220118
rect 397748 217410 397776 221478
rect 398576 220182 398604 230318
rect 398668 230314 398696 231676
rect 399036 230382 399064 231676
rect 399024 230376 399076 230382
rect 399024 230318 399076 230324
rect 398656 230308 398708 230314
rect 398656 230250 398708 230256
rect 399404 228585 399432 231676
rect 399484 230036 399536 230042
rect 399484 229978 399536 229984
rect 399390 228576 399446 228585
rect 399390 228511 399446 228520
rect 399392 227928 399444 227934
rect 399392 227870 399444 227876
rect 398564 220176 398616 220182
rect 398564 220118 398616 220124
rect 398840 219700 398892 219706
rect 398840 219642 398892 219648
rect 398852 217410 398880 219642
rect 399404 217410 399432 227870
rect 399496 219910 399524 229978
rect 399772 229906 399800 231676
rect 400048 231662 400154 231690
rect 399760 229900 399812 229906
rect 399760 229842 399812 229848
rect 400048 224466 400076 231662
rect 400128 230376 400180 230382
rect 400128 230318 400180 230324
rect 400036 224460 400088 224466
rect 400036 224402 400088 224408
rect 400140 221610 400168 230318
rect 400508 225593 400536 231676
rect 400680 230444 400732 230450
rect 400680 230386 400732 230392
rect 400494 225584 400550 225593
rect 400494 225519 400550 225528
rect 400692 221921 400720 230386
rect 400784 229702 400812 231676
rect 400864 230308 400916 230314
rect 400864 230250 400916 230256
rect 400876 230042 400904 230250
rect 400864 230036 400916 230042
rect 400864 229978 400916 229984
rect 400772 229696 400824 229702
rect 400772 229638 400824 229644
rect 401152 224369 401180 231676
rect 401520 229498 401548 231676
rect 401888 230450 401916 231676
rect 401876 230444 401928 230450
rect 401876 230386 401928 230392
rect 401508 229492 401560 229498
rect 401508 229434 401560 229440
rect 402256 224398 402284 231676
rect 402624 228449 402652 231676
rect 402992 230314 403020 231676
rect 403360 230382 403388 231676
rect 403348 230376 403400 230382
rect 403348 230318 403400 230324
rect 402980 230308 403032 230314
rect 402980 230250 403032 230256
rect 403072 230240 403124 230246
rect 403072 230182 403124 230188
rect 402610 228440 402666 228449
rect 402610 228375 402666 228384
rect 402980 228200 403032 228206
rect 402980 228142 403032 228148
rect 402244 224392 402296 224398
rect 401138 224360 401194 224369
rect 402244 224334 402296 224340
rect 401138 224295 401194 224304
rect 401876 224324 401928 224330
rect 401876 224266 401928 224272
rect 400678 221912 400734 221921
rect 400678 221847 400734 221856
rect 400128 221604 400180 221610
rect 400128 221546 400180 221552
rect 401140 221468 401192 221474
rect 401140 221410 401192 221416
rect 400312 220108 400364 220114
rect 400312 220050 400364 220056
rect 399484 219904 399536 219910
rect 399484 219846 399536 219852
rect 400324 217410 400352 220050
rect 401152 217410 401180 221410
rect 401888 217410 401916 224266
rect 402992 217410 403020 228142
rect 403084 227934 403112 230182
rect 403072 227928 403124 227934
rect 403072 227870 403124 227876
rect 403636 225690 403664 231676
rect 404018 231662 404308 231690
rect 404386 231662 404676 231690
rect 404280 230466 404308 231662
rect 404280 230438 404400 230466
rect 404372 230382 404400 230438
rect 404176 230376 404228 230382
rect 404176 230318 404228 230324
rect 404360 230376 404412 230382
rect 404360 230318 404412 230324
rect 403532 225684 403584 225690
rect 403532 225626 403584 225632
rect 403624 225684 403676 225690
rect 403624 225626 403676 225632
rect 403544 217410 403572 225626
rect 404188 221542 404216 230318
rect 404268 230308 404320 230314
rect 404268 230250 404320 230256
rect 404176 221536 404228 221542
rect 404176 221478 404228 221484
rect 404280 220114 404308 230250
rect 404360 229628 404412 229634
rect 404360 229570 404412 229576
rect 404372 228206 404400 229570
rect 404360 228200 404412 228206
rect 404360 228142 404412 228148
rect 404648 223038 404676 231662
rect 404740 230314 404768 231676
rect 404728 230308 404780 230314
rect 404728 230250 404780 230256
rect 405004 229492 405056 229498
rect 405004 229434 405056 229440
rect 404636 223032 404688 223038
rect 404636 222974 404688 222980
rect 405016 221513 405044 229434
rect 405108 229158 405136 231676
rect 405096 229152 405148 229158
rect 405096 229094 405148 229100
rect 405476 224330 405504 231676
rect 405858 231662 406148 231690
rect 406016 228132 406068 228138
rect 406016 228074 406068 228080
rect 405464 224324 405516 224330
rect 405464 224266 405516 224272
rect 405832 224188 405884 224194
rect 405832 224130 405884 224136
rect 405002 221504 405058 221513
rect 405002 221439 405058 221448
rect 404452 220924 404504 220930
rect 404452 220866 404504 220872
rect 404268 220108 404320 220114
rect 404268 220050 404320 220056
rect 404464 217410 404492 220866
rect 405844 217410 405872 224130
rect 406028 219434 406056 228074
rect 406120 224233 406148 231662
rect 406212 230246 406240 231676
rect 406502 231662 406792 231690
rect 406660 230376 406712 230382
rect 406660 230318 406712 230324
rect 406200 230240 406252 230246
rect 406200 230182 406252 230188
rect 406672 229770 406700 230318
rect 406384 229764 406436 229770
rect 406384 229706 406436 229712
rect 406660 229764 406712 229770
rect 406660 229706 406712 229712
rect 406106 224224 406162 224233
rect 406106 224159 406162 224168
rect 406396 219570 406424 229706
rect 406764 221474 406792 231662
rect 406856 230382 406884 231676
rect 406844 230376 406896 230382
rect 406844 230318 406896 230324
rect 407028 229968 407080 229974
rect 407028 229910 407080 229916
rect 407040 228138 407068 229910
rect 407224 229362 407252 231676
rect 407396 229832 407448 229838
rect 407396 229774 407448 229780
rect 407212 229356 407264 229362
rect 407212 229298 407264 229304
rect 407408 229226 407436 229774
rect 407304 229220 407356 229226
rect 407304 229162 407356 229168
rect 407396 229220 407448 229226
rect 407396 229162 407448 229168
rect 407028 228132 407080 228138
rect 407028 228074 407080 228080
rect 407316 225758 407344 229162
rect 407120 225752 407172 225758
rect 407120 225694 407172 225700
rect 407304 225752 407356 225758
rect 407304 225694 407356 225700
rect 406752 221468 406804 221474
rect 406752 221410 406804 221416
rect 406384 219564 406436 219570
rect 406384 219506 406436 219512
rect 406028 219406 406148 219434
rect 391032 217382 391368 217410
rect 391952 217382 392196 217410
rect 392596 217382 393024 217410
rect 393608 217382 393944 217410
rect 394712 217382 394772 217410
rect 395264 217382 395600 217410
rect 396184 217382 396428 217410
rect 396920 217382 397256 217410
rect 397748 217382 398084 217410
rect 398852 217382 398912 217410
rect 399404 217382 399832 217410
rect 400324 217382 400660 217410
rect 401152 217382 401488 217410
rect 401888 217382 402316 217410
rect 402992 217382 403144 217410
rect 403544 217382 403972 217410
rect 404464 217382 404800 217410
rect 405720 217382 405872 217410
rect 406120 217410 406148 219406
rect 407132 217410 407160 225694
rect 407592 222902 407620 231676
rect 407764 230036 407816 230042
rect 407764 229978 407816 229984
rect 407776 229498 407804 229978
rect 407856 229900 407908 229906
rect 407856 229842 407908 229848
rect 407868 229634 407896 229842
rect 407856 229628 407908 229634
rect 407856 229570 407908 229576
rect 407764 229492 407816 229498
rect 407764 229434 407816 229440
rect 407764 229220 407816 229226
rect 407764 229162 407816 229168
rect 407776 225026 407804 229162
rect 407960 226953 407988 231676
rect 408328 230042 408356 231676
rect 408316 230036 408368 230042
rect 408316 229978 408368 229984
rect 408500 228472 408552 228478
rect 408500 228414 408552 228420
rect 407946 226944 408002 226953
rect 407946 226879 408002 226888
rect 407776 224998 407988 225026
rect 407580 222896 407632 222902
rect 407580 222838 407632 222844
rect 407960 221066 407988 224998
rect 407856 221060 407908 221066
rect 407856 221002 407908 221008
rect 407948 221060 408000 221066
rect 407948 221002 408000 221008
rect 407868 217410 407896 221002
rect 408512 219502 408540 228414
rect 408696 224262 408724 231676
rect 409064 229838 409092 231676
rect 409340 229974 409368 231676
rect 409328 229968 409380 229974
rect 409328 229910 409380 229916
rect 409052 229832 409104 229838
rect 409052 229774 409104 229780
rect 409708 227050 409736 231676
rect 409788 230308 409840 230314
rect 409788 230250 409840 230256
rect 409800 228478 409828 230250
rect 409972 230240 410024 230246
rect 409972 230182 410024 230188
rect 409880 229560 409932 229566
rect 409880 229502 409932 229508
rect 409788 228472 409840 228478
rect 409788 228414 409840 228420
rect 409696 227044 409748 227050
rect 409696 226986 409748 226992
rect 408592 224256 408644 224262
rect 408592 224198 408644 224204
rect 408684 224256 408736 224262
rect 408684 224198 408736 224204
rect 408500 219496 408552 219502
rect 408500 219438 408552 219444
rect 408604 217410 408632 224198
rect 409892 223718 409920 229502
rect 409984 229158 410012 230182
rect 410076 229226 410104 231676
rect 410444 229906 410472 231676
rect 410432 229900 410484 229906
rect 410432 229842 410484 229848
rect 410064 229220 410116 229226
rect 410064 229162 410116 229168
rect 409972 229152 410024 229158
rect 409972 229094 410024 229100
rect 410812 228410 410840 231676
rect 410904 231662 411194 231690
rect 410904 229158 410932 231662
rect 410984 230376 411036 230382
rect 410984 230318 411036 230324
rect 411168 230376 411220 230382
rect 411168 230318 411220 230324
rect 410892 229152 410944 229158
rect 410892 229094 410944 229100
rect 409972 228404 410024 228410
rect 409972 228346 410024 228352
rect 410800 228404 410852 228410
rect 410800 228346 410852 228352
rect 409880 223712 409932 223718
rect 409880 223654 409932 223660
rect 409984 219774 410012 228346
rect 410996 225622 411024 230318
rect 411076 229832 411128 229838
rect 411076 229774 411128 229780
rect 411088 228313 411116 229774
rect 411180 229770 411208 230318
rect 411548 229770 411576 231676
rect 411168 229764 411220 229770
rect 411168 229706 411220 229712
rect 411536 229764 411588 229770
rect 411536 229706 411588 229712
rect 411916 229566 411944 231676
rect 507952 230512 508004 230518
rect 507952 230454 508004 230460
rect 456156 230444 456208 230450
rect 456156 230386 456208 230392
rect 428646 230344 428702 230353
rect 428646 230279 428702 230288
rect 411996 230036 412048 230042
rect 411996 229978 412048 229984
rect 411904 229560 411956 229566
rect 411904 229502 411956 229508
rect 412008 229362 412036 229978
rect 422300 229560 422352 229566
rect 422300 229502 422352 229508
rect 411996 229356 412048 229362
rect 411996 229298 412048 229304
rect 411260 229288 411312 229294
rect 411260 229230 411312 229236
rect 411074 228304 411130 228313
rect 411074 228239 411130 228248
rect 410248 225616 410300 225622
rect 410248 225558 410300 225564
rect 410984 225616 411036 225622
rect 410984 225558 411036 225564
rect 409880 219768 409932 219774
rect 409880 219710 409932 219716
rect 409972 219768 410024 219774
rect 409972 219710 410024 219716
rect 409892 217410 409920 219710
rect 406120 217382 406548 217410
rect 407132 217382 407376 217410
rect 407868 217382 408204 217410
rect 408604 217382 409032 217410
rect 409860 217382 409920 217410
rect 410260 217410 410288 225558
rect 411272 224194 411300 229230
rect 416228 229220 416280 229226
rect 416228 229162 416280 229168
rect 414020 225276 414072 225282
rect 414020 225218 414072 225224
rect 411260 224188 411312 224194
rect 411260 224130 411312 224136
rect 411996 223780 412048 223786
rect 411996 223722 412048 223728
rect 411260 220992 411312 220998
rect 411260 220934 411312 220940
rect 411272 217410 411300 220934
rect 412008 217410 412036 223722
rect 412916 219564 412968 219570
rect 412916 219506 412968 219512
rect 412928 217410 412956 219506
rect 414032 217410 414060 225218
rect 415492 223848 415544 223854
rect 415492 223790 415544 223796
rect 415308 222964 415360 222970
rect 415308 222906 415360 222912
rect 415320 219706 415348 222906
rect 415308 219700 415360 219706
rect 415308 219642 415360 219648
rect 414572 219496 414624 219502
rect 414572 219438 414624 219444
rect 414584 217410 414612 219438
rect 415504 217410 415532 223790
rect 416240 222970 416268 229162
rect 421012 229152 421064 229158
rect 421012 229094 421064 229100
rect 421024 229066 421328 229094
rect 419540 227996 419592 228002
rect 419540 227938 419592 227944
rect 417056 223984 417108 223990
rect 417056 223926 417108 223932
rect 416228 222964 416280 222970
rect 416228 222906 416280 222912
rect 416228 219768 416280 219774
rect 416228 219710 416280 219716
rect 416240 217410 416268 219710
rect 417068 217410 417096 223926
rect 418712 223916 418764 223922
rect 418712 223858 418764 223864
rect 418160 219700 418212 219706
rect 418160 219642 418212 219648
rect 418172 217410 418200 219642
rect 418724 217410 418752 223858
rect 419552 217410 419580 227938
rect 420368 225344 420420 225350
rect 420368 225286 420420 225292
rect 420380 217410 420408 225286
rect 421300 223106 421328 229066
rect 422312 228274 422340 229502
rect 422208 228268 422260 228274
rect 422208 228210 422260 228216
rect 422300 228268 422352 228274
rect 422300 228210 422352 228216
rect 422220 228154 422248 228210
rect 422220 228126 422340 228154
rect 421196 223100 421248 223106
rect 421196 223042 421248 223048
rect 421288 223100 421340 223106
rect 421288 223042 421340 223048
rect 421208 217410 421236 223042
rect 422312 217870 422340 228126
rect 426440 228064 426492 228070
rect 426440 228006 426492 228012
rect 422392 224052 422444 224058
rect 422392 223994 422444 224000
rect 422300 217864 422352 217870
rect 422300 217806 422352 217812
rect 422404 217410 422432 223994
rect 425060 222420 425112 222426
rect 425060 222362 425112 222368
rect 423864 219428 423916 219434
rect 423864 219370 423916 219376
rect 423036 217864 423088 217870
rect 423036 217806 423088 217812
rect 423048 217410 423076 217806
rect 423876 217410 423904 219370
rect 425072 217410 425100 222362
rect 425520 221196 425572 221202
rect 425520 221138 425572 221144
rect 410260 217382 410688 217410
rect 411272 217382 411608 217410
rect 412008 217382 412436 217410
rect 412928 217382 413264 217410
rect 414032 217382 414092 217410
rect 414584 217382 414920 217410
rect 415504 217382 415748 217410
rect 416240 217382 416576 217410
rect 417068 217382 417496 217410
rect 418172 217382 418324 217410
rect 418724 217382 419152 217410
rect 419552 217382 419980 217410
rect 420380 217382 420808 217410
rect 421208 217382 421636 217410
rect 422404 217382 422464 217410
rect 423048 217382 423384 217410
rect 423876 217382 424212 217410
rect 425040 217382 425100 217410
rect 425532 217410 425560 221138
rect 426452 217410 426480 228006
rect 427084 226568 427136 226574
rect 427084 226510 427136 226516
rect 427096 217410 427124 226510
rect 428660 222494 428688 230279
rect 443644 230172 443696 230178
rect 443644 230114 443696 230120
rect 438952 229492 439004 229498
rect 438952 229434 439004 229440
rect 431960 229424 432012 229430
rect 431960 229366 432012 229372
rect 429660 227928 429712 227934
rect 429660 227870 429712 227876
rect 429292 222556 429344 222562
rect 429292 222498 429344 222504
rect 427912 222488 427964 222494
rect 427912 222430 427964 222436
rect 428648 222488 428700 222494
rect 428648 222430 428700 222436
rect 427924 217410 427952 222430
rect 429304 217410 429332 222498
rect 425532 217382 425868 217410
rect 426452 217382 426696 217410
rect 427096 217382 427524 217410
rect 427924 217382 428352 217410
rect 429272 217382 429332 217410
rect 429672 217410 429700 227870
rect 431972 223446 432000 229366
rect 433340 228336 433392 228342
rect 433340 228278 433392 228284
rect 431316 223440 431368 223446
rect 431316 223382 431368 223388
rect 431960 223440 432012 223446
rect 431960 223382 432012 223388
rect 430580 219292 430632 219298
rect 430580 219234 430632 219240
rect 430592 217410 430620 219234
rect 431328 217410 431356 223382
rect 432236 219360 432288 219366
rect 432236 219302 432288 219308
rect 432248 217410 432276 219302
rect 433352 217410 433380 228278
rect 437480 226704 437532 226710
rect 437480 226646 437532 226652
rect 433800 226636 433852 226642
rect 433800 226578 433852 226584
rect 433812 217410 433840 226578
rect 434720 225140 434772 225146
rect 434720 225082 434772 225088
rect 434732 217870 434760 225082
rect 434812 222624 434864 222630
rect 434812 222566 434864 222572
rect 434720 217864 434772 217870
rect 434720 217806 434772 217812
rect 434824 217410 434852 222566
rect 436468 221060 436520 221066
rect 436468 221002 436520 221008
rect 435640 217864 435692 217870
rect 435640 217806 435692 217812
rect 435652 217410 435680 217806
rect 436480 217410 436508 221002
rect 437492 217410 437520 226646
rect 438964 225894 438992 229434
rect 440608 226772 440660 226778
rect 440608 226714 440660 226720
rect 438860 225888 438912 225894
rect 438860 225830 438912 225836
rect 438952 225888 439004 225894
rect 438952 225830 439004 225836
rect 438032 222692 438084 222698
rect 438032 222634 438084 222640
rect 438044 217410 438072 222634
rect 438872 217410 438900 225830
rect 439780 221264 439832 221270
rect 439780 221206 439832 221212
rect 439792 217410 439820 221206
rect 440620 217410 440648 226714
rect 441620 225412 441672 225418
rect 441620 225354 441672 225360
rect 441632 217870 441660 225354
rect 441712 222760 441764 222766
rect 441712 222702 441764 222708
rect 441620 217864 441672 217870
rect 441620 217806 441672 217812
rect 441724 217410 441752 222702
rect 443656 221270 443684 230114
rect 453304 229696 453356 229702
rect 453304 229638 453356 229644
rect 449164 229628 449216 229634
rect 449164 229570 449216 229576
rect 449176 227662 449204 229570
rect 444380 227656 444432 227662
rect 444380 227598 444432 227604
rect 449164 227656 449216 227662
rect 449164 227598 449216 227604
rect 443644 221264 443696 221270
rect 443644 221206 443696 221212
rect 443184 221128 443236 221134
rect 443184 221070 443236 221076
rect 442356 217864 442408 217870
rect 442356 217806 442408 217812
rect 442368 217410 442396 217806
rect 443196 217410 443224 221070
rect 444392 217410 444420 227598
rect 450636 226908 450688 226914
rect 450636 226850 450688 226856
rect 447324 226840 447376 226846
rect 447324 226782 447376 226788
rect 445760 225480 445812 225486
rect 445760 225422 445812 225428
rect 444748 222828 444800 222834
rect 444748 222770 444800 222776
rect 429672 217382 430100 217410
rect 430592 217382 430928 217410
rect 431328 217382 431756 217410
rect 432248 217382 432584 217410
rect 433352 217382 433412 217410
rect 433812 217382 434240 217410
rect 434824 217382 435160 217410
rect 435652 217382 435988 217410
rect 436480 217382 436816 217410
rect 437492 217382 437644 217410
rect 438044 217382 438472 217410
rect 438872 217382 439300 217410
rect 439792 217382 440128 217410
rect 440620 217382 441048 217410
rect 441724 217382 441876 217410
rect 442368 217382 442704 217410
rect 443196 217382 443532 217410
rect 444360 217382 444420 217410
rect 444760 217410 444788 222770
rect 445772 217410 445800 225422
rect 446588 221332 446640 221338
rect 446588 221274 446640 221280
rect 446600 217410 446628 221274
rect 447336 217410 447364 226782
rect 448980 225208 449032 225214
rect 448980 225150 449032 225156
rect 448612 223576 448664 223582
rect 448612 223518 448664 223524
rect 448624 217410 448652 223518
rect 444760 217382 445188 217410
rect 445772 217382 446016 217410
rect 446600 217382 446936 217410
rect 447336 217382 447764 217410
rect 448592 217382 448652 217410
rect 448992 217410 449020 225150
rect 449900 221400 449952 221406
rect 449900 221342 449952 221348
rect 449912 217410 449940 221342
rect 450648 217410 450676 226850
rect 452660 225548 452712 225554
rect 452660 225490 452712 225496
rect 451464 223508 451516 223514
rect 451464 223450 451516 223456
rect 451476 217410 451504 223450
rect 452672 217410 452700 225490
rect 453316 222154 453344 229638
rect 454040 228132 454092 228138
rect 454040 228074 454092 228080
rect 453212 222148 453264 222154
rect 453212 222090 453264 222096
rect 453304 222148 453356 222154
rect 453304 222090 453356 222096
rect 453224 217410 453252 222090
rect 454052 217870 454080 228074
rect 454132 226976 454184 226982
rect 454132 226918 454184 226924
rect 454040 217864 454092 217870
rect 454040 217806 454092 217812
rect 454144 217410 454172 226918
rect 456168 226302 456196 230386
rect 461584 230376 461636 230382
rect 461584 230318 461636 230324
rect 460940 229084 460992 229090
rect 460940 229026 460992 229032
rect 457352 227724 457404 227730
rect 457352 227666 457404 227672
rect 455696 226296 455748 226302
rect 455696 226238 455748 226244
rect 456156 226296 456208 226302
rect 456156 226238 456208 226244
rect 454960 217864 455012 217870
rect 454960 217806 455012 217812
rect 454972 217410 455000 217806
rect 455708 217410 455736 226238
rect 456800 222080 456852 222086
rect 456800 222022 456852 222028
rect 456812 217410 456840 222022
rect 457364 217410 457392 227666
rect 459560 226228 459612 226234
rect 459560 226170 459612 226176
rect 458364 222012 458416 222018
rect 458364 221954 458416 221960
rect 458376 217410 458404 221954
rect 459572 217410 459600 226170
rect 460020 221944 460072 221950
rect 460020 221886 460072 221892
rect 448992 217382 449420 217410
rect 449912 217382 450248 217410
rect 450648 217382 451076 217410
rect 451476 217382 451904 217410
rect 452672 217382 452824 217410
rect 453224 217382 453652 217410
rect 454144 217382 454480 217410
rect 454972 217382 455308 217410
rect 455708 217382 456136 217410
rect 456812 217382 456964 217410
rect 457364 217382 457792 217410
rect 458376 217382 458712 217410
rect 459540 217382 459600 217410
rect 460032 217410 460060 221886
rect 460952 217870 460980 229026
rect 461596 227594 461624 230318
rect 467104 230308 467156 230314
rect 467104 230250 467156 230256
rect 461216 227588 461268 227594
rect 461216 227530 461268 227536
rect 461584 227588 461636 227594
rect 461584 227530 461636 227536
rect 461228 219434 461256 227530
rect 464160 227520 464212 227526
rect 464160 227462 464212 227468
rect 462412 226160 462464 226166
rect 462412 226102 462464 226108
rect 461044 219406 461256 219434
rect 460940 217864 460992 217870
rect 460940 217806 460992 217812
rect 461044 217410 461072 219406
rect 461676 217864 461728 217870
rect 461676 217806 461728 217812
rect 461688 217410 461716 217806
rect 462424 217410 462452 226102
rect 463700 221876 463752 221882
rect 463700 221818 463752 221824
rect 463712 217410 463740 221818
rect 460032 217382 460368 217410
rect 461044 217382 461196 217410
rect 461688 217382 462024 217410
rect 462424 217382 462852 217410
rect 463680 217382 463740 217410
rect 464172 217410 464200 227462
rect 465080 226092 465132 226098
rect 465080 226034 465132 226040
rect 465092 217870 465120 226034
rect 465172 223712 465224 223718
rect 465172 223654 465224 223660
rect 465080 217864 465132 217870
rect 465080 217806 465132 217812
rect 465184 217410 465212 223654
rect 467116 221814 467144 230250
rect 469220 230240 469272 230246
rect 469220 230182 469272 230188
rect 478142 230208 478198 230217
rect 469232 227458 469260 230182
rect 478142 230143 478198 230152
rect 476120 228200 476172 228206
rect 476120 228142 476172 228148
rect 467840 227452 467892 227458
rect 467840 227394 467892 227400
rect 469220 227452 469272 227458
rect 469220 227394 469272 227400
rect 466736 221808 466788 221814
rect 466736 221750 466788 221756
rect 467104 221808 467156 221814
rect 467104 221750 467156 221756
rect 465908 217864 465960 217870
rect 465908 217806 465960 217812
rect 465920 217410 465948 217806
rect 466748 217410 466776 221750
rect 467852 217410 467880 227394
rect 470876 227384 470928 227390
rect 470876 227326 470928 227332
rect 469220 226024 469272 226030
rect 469220 225966 469272 225972
rect 468300 224936 468352 224942
rect 468300 224878 468352 224884
rect 468312 217410 468340 224878
rect 469232 217410 469260 225966
rect 470140 221740 470192 221746
rect 470140 221682 470192 221688
rect 470152 217410 470180 221682
rect 470888 217410 470916 227326
rect 474188 227316 474240 227322
rect 474188 227258 474240 227264
rect 471980 225956 472032 225962
rect 471980 225898 472032 225904
rect 471992 217870 472020 225898
rect 472072 224120 472124 224126
rect 472072 224062 472124 224068
rect 471980 217864 472032 217870
rect 471980 217806 472032 217812
rect 472084 217410 472112 224062
rect 473544 221672 473596 221678
rect 473544 221614 473596 221620
rect 472624 217864 472676 217870
rect 472624 217806 472676 217812
rect 472636 217410 472664 217806
rect 473556 217410 473584 221614
rect 474200 217410 474228 227258
rect 475016 224800 475068 224806
rect 475016 224742 475068 224748
rect 475028 217410 475056 224742
rect 476132 217870 476160 228142
rect 478156 227254 478184 230143
rect 486422 230072 486478 230081
rect 486422 230007 486478 230016
rect 480260 229016 480312 229022
rect 480260 228958 480312 228964
rect 477592 227248 477644 227254
rect 477592 227190 477644 227196
rect 478144 227248 478196 227254
rect 478144 227190 478196 227196
rect 476212 225820 476264 225826
rect 476212 225762 476264 225768
rect 476120 217864 476172 217870
rect 476120 217806 476172 217812
rect 476224 217410 476252 225762
rect 476856 217864 476908 217870
rect 476856 217806 476908 217812
rect 476868 217410 476896 217806
rect 477604 217410 477632 227190
rect 479248 224868 479300 224874
rect 479248 224810 479300 224816
rect 478972 224732 479024 224738
rect 478972 224674 479024 224680
rect 478984 217410 479012 224674
rect 464172 217382 464600 217410
rect 465184 217382 465428 217410
rect 465920 217382 466256 217410
rect 466748 217382 467084 217410
rect 467852 217382 467912 217410
rect 468312 217382 468740 217410
rect 469232 217382 469568 217410
rect 470152 217382 470488 217410
rect 470888 217382 471316 217410
rect 472084 217382 472144 217410
rect 472636 217382 472972 217410
rect 473556 217382 473800 217410
rect 474200 217382 474628 217410
rect 475028 217382 475456 217410
rect 476224 217382 476376 217410
rect 476868 217382 477204 217410
rect 477604 217382 478032 217410
rect 478860 217382 479012 217410
rect 479260 217410 479288 224810
rect 480272 217410 480300 228958
rect 483480 228948 483532 228954
rect 483480 228890 483532 228896
rect 480904 227180 480956 227186
rect 480904 227122 480956 227128
rect 480916 217410 480944 227122
rect 483112 227112 483164 227118
rect 483112 227054 483164 227060
rect 481824 224664 481876 224670
rect 481824 224606 481876 224612
rect 481836 217410 481864 224606
rect 483124 217410 483152 227054
rect 479260 217382 479688 217410
rect 480272 217382 480516 217410
rect 480916 217382 481344 217410
rect 481836 217382 482264 217410
rect 483092 217382 483152 217410
rect 483492 217410 483520 228890
rect 485136 228268 485188 228274
rect 485136 228210 485188 228216
rect 484400 219836 484452 219842
rect 484400 219778 484452 219784
rect 484412 217410 484440 219778
rect 485148 217410 485176 228210
rect 486436 218142 486464 230007
rect 493322 229936 493378 229945
rect 493322 229871 493378 229880
rect 493336 229094 493364 229871
rect 496082 229800 496138 229809
rect 496082 229735 496138 229744
rect 493336 229066 493456 229094
rect 487712 228880 487764 228886
rect 487712 228822 487764 228828
rect 486424 218136 486476 218142
rect 486424 218078 486476 218084
rect 486436 217410 486464 218078
rect 487528 218068 487580 218074
rect 487528 218010 487580 218016
rect 487540 217410 487568 218010
rect 483492 217382 483920 217410
rect 484412 217382 484748 217410
rect 485148 217382 485576 217410
rect 486404 217382 486464 217410
rect 487232 217382 487568 217410
rect 487724 217410 487752 228822
rect 491300 228812 491352 228818
rect 491300 228754 491352 228760
rect 490194 224768 490250 224777
rect 490194 224703 490250 224712
rect 487802 223272 487858 223281
rect 487802 223207 487858 223216
rect 487816 218482 487844 223207
rect 488540 222488 488592 222494
rect 488540 222430 488592 222436
rect 487804 218476 487856 218482
rect 487804 218418 487856 218424
rect 487816 218074 487844 218418
rect 487804 218068 487856 218074
rect 487804 218010 487856 218016
rect 488552 217410 488580 222430
rect 489458 220416 489514 220425
rect 489458 220351 489514 220360
rect 489472 218142 489500 220351
rect 489460 218136 489512 218142
rect 489460 218078 489512 218084
rect 489472 217410 489500 218078
rect 490208 217410 490236 224703
rect 490932 217728 490984 217734
rect 490932 217670 490984 217676
rect 490944 217410 490972 217670
rect 487724 217382 488152 217410
rect 488552 217396 488980 217410
rect 488552 217382 488994 217396
rect 489472 217382 489808 217410
rect 490208 217382 490972 217410
rect 491312 217410 491340 228754
rect 491944 221264 491996 221270
rect 491944 221206 491996 221212
rect 491312 217382 491464 217410
rect 488966 216730 488994 217382
rect 491956 216866 491984 221206
rect 493428 218210 493456 229066
rect 494150 223136 494206 223145
rect 494150 223071 494206 223080
rect 493416 218204 493468 218210
rect 493416 218146 493468 218152
rect 493428 217410 493456 218146
rect 494164 217410 494192 223071
rect 495622 220552 495678 220561
rect 495622 220487 495678 220496
rect 494520 219224 494572 219230
rect 494520 219166 494572 219172
rect 494532 217410 494560 219166
rect 495636 218414 495664 220487
rect 495624 218408 495676 218414
rect 495624 218350 495676 218356
rect 495992 218408 496044 218414
rect 495992 218350 496044 218356
rect 496004 217410 496032 218350
rect 496096 218278 496124 229735
rect 496910 227352 496966 227361
rect 496910 227287 496966 227296
rect 496084 218272 496136 218278
rect 496084 218214 496136 218220
rect 493120 217382 493456 217410
rect 494040 217394 494376 217410
rect 494040 217388 494388 217394
rect 494040 217382 494336 217388
rect 494532 217382 494868 217410
rect 495696 217382 496032 217410
rect 496096 217410 496124 218214
rect 496924 217410 496952 227287
rect 500224 227248 500276 227254
rect 500224 227190 500276 227196
rect 502522 227216 502578 227225
rect 499578 224632 499634 224641
rect 499578 224567 499634 224576
rect 498658 220280 498714 220289
rect 498658 220215 498714 220224
rect 498672 219638 498700 220215
rect 498660 219632 498712 219638
rect 498660 219574 498712 219580
rect 498200 219156 498252 219162
rect 498200 219098 498252 219104
rect 497648 217796 497700 217802
rect 497648 217738 497700 217744
rect 497660 217410 497688 217738
rect 498212 217410 498240 219098
rect 496096 217382 496524 217410
rect 496924 217382 497688 217410
rect 498180 217382 498240 217410
rect 498672 217410 498700 219574
rect 499592 217870 499620 224567
rect 500236 218346 500264 227190
rect 502522 227151 502578 227160
rect 502432 220040 502484 220046
rect 502432 219982 502484 219988
rect 502444 219570 502472 219982
rect 502432 219564 502484 219570
rect 502432 219506 502484 219512
rect 501236 219088 501288 219094
rect 501236 219030 501288 219036
rect 500224 218340 500276 218346
rect 500224 218282 500276 218288
rect 499580 217864 499632 217870
rect 499580 217806 499632 217812
rect 500236 217410 500264 218282
rect 500868 217864 500920 217870
rect 500868 217806 500920 217812
rect 500880 217410 500908 217806
rect 498672 217382 499008 217410
rect 499928 217382 500264 217410
rect 500756 217382 500908 217410
rect 501248 217410 501276 219030
rect 502444 217410 502472 219506
rect 501248 217382 501584 217410
rect 502412 217382 502472 217410
rect 494336 217330 494388 217336
rect 502536 216918 502564 227151
rect 505374 224496 505430 224505
rect 505374 224431 505430 224440
rect 504916 219972 504968 219978
rect 504916 219914 504968 219920
rect 504928 219502 504956 219914
rect 505008 219632 505060 219638
rect 505008 219574 505060 219580
rect 504916 219496 504968 219502
rect 504916 219438 504968 219444
rect 503720 219020 503772 219026
rect 503720 218962 503772 218968
rect 503732 217410 503760 218962
rect 504928 217410 504956 219438
rect 505020 219026 505048 219574
rect 505008 219020 505060 219026
rect 505008 218962 505060 218968
rect 503732 217382 504068 217410
rect 504896 217382 504956 217410
rect 505388 217410 505416 224431
rect 506480 224188 506532 224194
rect 506480 224130 506532 224136
rect 506492 217410 506520 224130
rect 507214 220144 507270 220153
rect 507214 220079 507270 220088
rect 507228 219473 507256 220079
rect 507214 219464 507270 219473
rect 507214 219399 507270 219408
rect 507228 217410 507256 219399
rect 507964 217410 507992 230454
rect 515404 230104 515456 230110
rect 515404 230046 515456 230052
rect 513378 228712 513434 228721
rect 513378 228647 513434 228656
rect 510710 225992 510766 226001
rect 510710 225927 510766 225936
rect 509884 220788 509936 220794
rect 509884 220730 509936 220736
rect 509896 219638 509924 220730
rect 509884 219632 509936 219638
rect 509884 219574 509936 219580
rect 508780 218952 508832 218958
rect 508780 218894 508832 218900
rect 508792 217410 508820 218894
rect 509896 217410 509924 219574
rect 510724 217682 510752 225927
rect 512828 220652 512880 220658
rect 512828 220594 512880 220600
rect 512840 219706 512868 220594
rect 512828 219700 512880 219706
rect 512828 219642 512880 219648
rect 511356 218884 511408 218890
rect 511356 218826 511408 218832
rect 510724 217654 510798 217682
rect 510770 217410 510798 217654
rect 511368 217410 511396 218826
rect 512840 217410 512868 219642
rect 505388 217382 506152 217410
rect 506492 217382 506644 217410
rect 507228 217382 507472 217410
rect 507964 217382 508544 217410
rect 508792 217382 509128 217410
rect 509896 217382 509956 217410
rect 510770 217396 510844 217410
rect 510784 217382 510844 217396
rect 511368 217382 511704 217410
rect 512532 217382 512868 217410
rect 506124 216986 506152 217382
rect 508516 217054 508544 217382
rect 508504 217048 508556 217054
rect 510816 217002 510844 217382
rect 513392 217138 513420 228647
rect 513840 219904 513892 219910
rect 513840 219846 513892 219852
rect 513852 217410 513880 219846
rect 515416 219774 515444 230046
rect 539600 230036 539652 230042
rect 539600 229978 539652 229984
rect 523040 228744 523092 228750
rect 523040 228686 523092 228692
rect 515494 227080 515550 227089
rect 515494 227015 515550 227024
rect 515404 219768 515456 219774
rect 515404 219710 515456 219716
rect 515416 217410 515444 219710
rect 515508 218618 515536 227015
rect 516232 224596 516284 224602
rect 516232 224538 516284 224544
rect 515496 218612 515548 218618
rect 515496 218554 515548 218560
rect 513852 217382 514188 217410
rect 515016 217382 515444 217410
rect 515508 217410 515536 218554
rect 516244 217410 516272 224538
rect 518900 224528 518952 224534
rect 518900 224470 518952 224476
rect 517978 223000 518034 223009
rect 517978 222935 518034 222944
rect 517520 220720 517572 220726
rect 517520 220662 517572 220668
rect 517532 217410 517560 220662
rect 517992 217410 518020 222935
rect 518912 217410 518940 224470
rect 520462 222864 520518 222873
rect 520462 222799 520518 222808
rect 520004 220584 520056 220590
rect 520004 220526 520056 220532
rect 520016 217410 520044 220526
rect 515508 217382 515844 217410
rect 516244 217382 516672 217410
rect 517532 217382 517592 217410
rect 517992 217382 518756 217410
rect 518912 217382 519248 217410
rect 520016 217382 520076 217410
rect 513656 217184 513708 217190
rect 513360 217132 513656 217138
rect 513360 217126 513708 217132
rect 511080 217116 511132 217122
rect 513360 217110 513696 217126
rect 511080 217058 511132 217064
rect 511092 217002 511120 217058
rect 508504 216990 508556 216996
rect 506112 216980 506164 216986
rect 510784 216974 511120 217002
rect 506112 216922 506164 216928
rect 502524 216912 502576 216918
rect 492586 216880 492642 216889
rect 491956 216838 492586 216866
rect 503536 216912 503588 216918
rect 502524 216854 502576 216860
rect 503240 216860 503536 216866
rect 503240 216854 503588 216860
rect 503240 216838 503576 216854
rect 492586 216815 492642 216824
rect 489090 216744 489146 216753
rect 488966 216716 489090 216730
rect 488980 216702 489090 216716
rect 489090 216679 489146 216688
rect 518728 216442 518756 217382
rect 520476 216458 520504 222799
rect 522580 220720 522632 220726
rect 522580 220662 522632 220668
rect 522592 220522 522620 220662
rect 522580 220516 522632 220522
rect 522580 220458 522632 220464
rect 521660 218816 521712 218822
rect 521660 218758 521712 218764
rect 521672 217410 521700 218758
rect 522592 217410 522620 220458
rect 523052 217938 523080 228686
rect 526352 228676 526404 228682
rect 526352 228618 526404 228624
rect 525064 223440 525116 223446
rect 525064 223382 525116 223388
rect 523132 223372 523184 223378
rect 523132 223314 523184 223320
rect 523040 217932 523092 217938
rect 523040 217874 523092 217880
rect 521672 217382 521732 217410
rect 522560 217382 522620 217410
rect 523144 216458 523172 223314
rect 525076 220522 525104 223382
rect 525890 221776 525946 221785
rect 525890 221711 525946 221720
rect 525064 220516 525116 220522
rect 525064 220458 525116 220464
rect 523960 217932 524012 217938
rect 523960 217874 524012 217880
rect 523972 217410 524000 217874
rect 525076 217410 525104 220458
rect 525904 217546 525932 221711
rect 525904 217518 525978 217546
rect 523972 217382 524308 217410
rect 525076 217382 525136 217410
rect 525950 216594 525978 217518
rect 526364 217410 526392 228618
rect 536840 228608 536892 228614
rect 536840 228550 536892 228556
rect 528926 225856 528982 225865
rect 528926 225791 528982 225800
rect 528098 221912 528154 221921
rect 528098 221847 528154 221856
rect 527272 220448 527324 220454
rect 527272 220390 527324 220396
rect 527284 217410 527312 220390
rect 528112 217410 528140 221847
rect 528940 217410 528968 225791
rect 531412 225752 531464 225758
rect 531412 225694 531464 225700
rect 534078 225720 534134 225729
rect 530584 223304 530636 223310
rect 530584 223246 530636 223252
rect 530124 220380 530176 220386
rect 530124 220322 530176 220328
rect 530136 217410 530164 220322
rect 526364 217382 526792 217410
rect 527284 217382 527620 217410
rect 528112 217396 528448 217410
rect 528112 217382 528462 217396
rect 528940 217382 529368 217410
rect 530136 217382 530196 217410
rect 525950 216580 526300 216594
rect 525964 216566 526300 216580
rect 520476 216442 521240 216458
rect 523144 216442 523816 216458
rect 526272 216442 526300 216566
rect 528434 216458 528462 217382
rect 530596 216458 530624 223246
rect 531424 217410 531452 225694
rect 534078 225655 534134 225664
rect 533068 223236 533120 223242
rect 533068 223178 533120 223184
rect 532700 220312 532752 220318
rect 532700 220254 532752 220260
rect 531424 217382 531852 217410
rect 532712 217002 532740 220254
rect 532974 217016 533030 217025
rect 532680 216974 532974 217002
rect 532974 216951 533030 216960
rect 533080 216458 533108 223178
rect 534092 217410 534120 225655
rect 536010 221640 536066 221649
rect 536010 221575 536066 221584
rect 535368 220244 535420 220250
rect 535368 220186 535420 220192
rect 535380 219842 535408 220186
rect 535368 219836 535420 219842
rect 535368 219778 535420 219784
rect 535380 217410 535408 219778
rect 534092 217382 534336 217410
rect 535256 217382 535408 217410
rect 536024 217410 536052 221575
rect 536852 217410 536880 228550
rect 538220 228540 538272 228546
rect 538220 228482 538272 228488
rect 537392 220176 537444 220182
rect 537392 220118 537444 220124
rect 537404 217410 537432 220118
rect 538232 217938 538260 228482
rect 539612 225758 539640 229978
rect 547144 229968 547196 229974
rect 547144 229910 547196 229916
rect 541530 228576 541586 228585
rect 541530 228511 541586 228520
rect 540428 225888 540480 225894
rect 540428 225830 540480 225836
rect 539600 225752 539652 225758
rect 539600 225694 539652 225700
rect 538312 223168 538364 223174
rect 538312 223110 538364 223116
rect 538220 217932 538272 217938
rect 538220 217874 538272 217880
rect 536024 217382 536420 217410
rect 536852 217382 536912 217410
rect 537404 217382 537984 217410
rect 528434 216444 528600 216458
rect 528448 216442 528600 216444
rect 530596 216442 531268 216458
rect 533080 216442 533844 216458
rect 536392 216442 536420 217382
rect 537956 217258 537984 217382
rect 537944 217252 537996 217258
rect 537944 217194 537996 217200
rect 538324 216458 538352 223110
rect 540440 219910 540468 225830
rect 541072 221604 541124 221610
rect 541072 221546 541124 221552
rect 540428 219904 540480 219910
rect 540428 219846 540480 219852
rect 539048 217932 539100 217938
rect 539048 217874 539100 217880
rect 539060 217410 539088 217874
rect 540440 217410 540468 219846
rect 541084 217546 541112 221546
rect 541084 217518 541158 217546
rect 539060 217382 539396 217410
rect 540224 217382 540468 217410
rect 541130 216594 541158 217518
rect 541544 217410 541572 228511
rect 543004 227656 543056 227662
rect 543004 227598 543056 227604
rect 543016 220114 543044 227598
rect 544014 225584 544070 225593
rect 544014 225519 544070 225528
rect 543188 224460 543240 224466
rect 543188 224402 543240 224408
rect 543004 220108 543056 220114
rect 543004 220050 543056 220056
rect 543016 217410 543044 220050
rect 543200 218550 543228 224402
rect 543188 218544 543240 218550
rect 543188 218486 543240 218492
rect 543648 218544 543700 218550
rect 543648 218486 543700 218492
rect 543660 217410 543688 218486
rect 541544 217382 541972 217410
rect 542800 217382 543044 217410
rect 543628 217382 543688 217410
rect 544028 217410 544056 225519
rect 545762 224360 545818 224369
rect 545762 224295 545818 224304
rect 545212 222148 545264 222154
rect 545212 222090 545264 222096
rect 545224 217410 545252 222090
rect 545776 220658 545804 224295
rect 547156 221610 547184 229910
rect 551284 229900 551336 229906
rect 551284 229842 551336 229848
rect 549258 228440 549314 228449
rect 549258 228375 549314 228384
rect 548156 226296 548208 226302
rect 548156 226238 548208 226244
rect 547144 221604 547196 221610
rect 547144 221546 547196 221552
rect 546682 221504 546738 221513
rect 546682 221439 546738 221448
rect 545764 220652 545816 220658
rect 545764 220594 545816 220600
rect 545776 217410 545804 220594
rect 546696 217410 546724 221439
rect 548168 220182 548196 226238
rect 548524 224392 548576 224398
rect 548524 224334 548576 224340
rect 548156 220176 548208 220182
rect 548156 220118 548208 220124
rect 548168 217410 548196 220118
rect 548536 219094 548564 224334
rect 548524 219088 548576 219094
rect 548524 219030 548576 219036
rect 544028 217382 544456 217410
rect 545224 217382 545620 217410
rect 545776 217382 546112 217410
rect 546696 217382 547032 217410
rect 547860 217382 548196 217410
rect 548536 217410 548564 219030
rect 549272 217410 549300 228375
rect 551296 221542 551324 229842
rect 563704 229832 563756 229838
rect 563704 229774 563756 229780
rect 553400 228472 553452 228478
rect 553400 228414 553452 228420
rect 552664 227588 552716 227594
rect 552664 227530 552716 227536
rect 552020 225684 552072 225690
rect 552020 225626 552072 225632
rect 550824 221536 550876 221542
rect 550824 221478 550876 221484
rect 551284 221536 551336 221542
rect 551284 221478 551336 221484
rect 549628 220040 549680 220046
rect 549628 219982 549680 219988
rect 549640 217462 549668 219982
rect 549628 217456 549680 217462
rect 548536 217382 548688 217410
rect 549272 217382 549516 217410
rect 550548 217456 550600 217462
rect 549628 217398 549680 217404
rect 550344 217404 550548 217410
rect 550344 217398 550600 217404
rect 550344 217382 550588 217398
rect 545592 217326 545620 217382
rect 545580 217320 545632 217326
rect 545580 217262 545632 217268
rect 541130 216580 541480 216594
rect 541144 216566 541480 216580
rect 538324 216442 538904 216458
rect 541452 216442 541480 216566
rect 550836 216458 550864 221478
rect 552032 217410 552060 225626
rect 552000 217382 552060 217410
rect 552676 220130 552704 227530
rect 553412 224954 553440 228414
rect 555424 227452 555476 227458
rect 555424 227394 555476 227400
rect 553412 224926 554176 224954
rect 553676 223032 553728 223038
rect 553676 222974 553728 222980
rect 552676 220114 552888 220130
rect 552676 220108 552900 220114
rect 552676 220102 552848 220108
rect 552676 217410 552704 220102
rect 552848 220050 552900 220056
rect 553688 217682 553716 222974
rect 553688 217666 553762 217682
rect 553688 217660 553774 217666
rect 553688 217654 553722 217660
rect 553722 217602 553774 217608
rect 552676 217382 552920 217410
rect 553734 217396 553762 217602
rect 554148 217410 554176 224926
rect 555436 219162 555464 227394
rect 561678 226944 561734 226953
rect 561678 226879 561734 226888
rect 560852 225752 560904 225758
rect 560852 225694 560904 225700
rect 559196 225616 559248 225622
rect 559196 225558 559248 225564
rect 556160 224324 556212 224330
rect 556160 224266 556212 224272
rect 555424 219156 555476 219162
rect 555424 219098 555476 219104
rect 555436 217410 555464 219098
rect 556172 217530 556200 224266
rect 556710 224224 556766 224233
rect 556710 224159 556766 224168
rect 556160 217524 556212 217530
rect 556160 217466 556212 217472
rect 554148 217382 554576 217410
rect 555404 217382 555464 217410
rect 556172 217410 556200 217466
rect 556724 217410 556752 224159
rect 557816 221808 557868 221814
rect 557816 221750 557868 221756
rect 557828 218958 557856 221750
rect 558460 221468 558512 221474
rect 558460 221410 558512 221416
rect 557816 218952 557868 218958
rect 557816 218894 557868 218900
rect 557828 217410 557856 218894
rect 558472 217410 558500 221410
rect 559208 217410 559236 225558
rect 560864 224954 560892 225694
rect 560772 224926 560892 224954
rect 560772 220182 560800 224926
rect 560944 222896 560996 222902
rect 560944 222838 560996 222844
rect 560760 220176 560812 220182
rect 560760 220118 560812 220124
rect 560772 217410 560800 220118
rect 556172 217382 556232 217410
rect 556724 217382 557060 217410
rect 557828 217382 557888 217410
rect 558472 217382 558868 217410
rect 559208 217382 559636 217410
rect 560464 217382 560800 217410
rect 560956 217410 560984 222838
rect 561692 217410 561720 226879
rect 563612 224256 563664 224262
rect 563612 224198 563664 224204
rect 561772 221604 561824 221610
rect 561772 221546 561824 221552
rect 561784 218890 561812 221546
rect 561772 218884 561824 218890
rect 561772 218826 561824 218832
rect 562876 218884 562928 218890
rect 562876 218826 562928 218832
rect 562888 217410 562916 218826
rect 563624 217410 563652 224198
rect 563716 220862 563744 229774
rect 570604 229764 570656 229770
rect 570604 229706 570656 229712
rect 568580 228404 568632 228410
rect 568580 228346 568632 228352
rect 564438 228304 564494 228313
rect 564438 228239 564494 228248
rect 563704 220856 563756 220862
rect 563704 220798 563756 220804
rect 564452 217410 564480 228239
rect 565912 227044 565964 227050
rect 565912 226986 565964 226992
rect 565452 221536 565504 221542
rect 565452 221478 565504 221484
rect 565464 218822 565492 221478
rect 565452 218816 565504 218822
rect 565452 218758 565504 218764
rect 565464 217410 565492 218758
rect 565924 217410 565952 226986
rect 567200 222964 567252 222970
rect 567200 222906 567252 222912
rect 567212 217410 567240 222906
rect 567936 220856 567988 220862
rect 567936 220798 567988 220804
rect 567948 218686 567976 220798
rect 567936 218680 567988 218686
rect 567936 218622 567988 218628
rect 560956 217382 561444 217410
rect 561692 217382 562120 217410
rect 562888 217382 562948 217410
rect 563624 217382 564112 217410
rect 564452 217382 564696 217410
rect 565464 217382 565524 217410
rect 565924 217382 566504 217410
rect 567180 217382 567240 217410
rect 567948 217410 567976 218622
rect 568592 217410 568620 228346
rect 569316 223100 569368 223106
rect 569316 223042 569368 223048
rect 568810 217592 568862 217598
rect 568810 217534 568862 217540
rect 568822 217410 568850 217534
rect 567948 217382 568008 217410
rect 568592 217396 568850 217410
rect 569328 217410 569356 223042
rect 570616 219230 570644 229706
rect 570604 219224 570656 219230
rect 570604 219166 570656 219172
rect 570616 217410 570644 219166
rect 571444 217410 571472 255274
rect 571536 229094 571564 258062
rect 571536 229066 571840 229094
rect 568592 217382 568836 217396
rect 569328 217382 569664 217410
rect 570584 217382 570644 217410
rect 571412 217382 571472 217410
rect 571812 217410 571840 229066
rect 572732 217410 572760 262210
rect 574744 252612 574796 252618
rect 574744 252554 574796 252560
rect 574100 238060 574152 238066
rect 574100 238002 574152 238008
rect 572812 233912 572864 233918
rect 572812 233854 572864 233860
rect 572824 229094 572852 233854
rect 574112 229094 574140 238002
rect 572824 229066 573496 229094
rect 574112 229066 574324 229094
rect 573468 217410 573496 229066
rect 574296 217410 574324 229066
rect 574756 222154 574784 252554
rect 646056 248414 646084 278190
rect 647528 275330 647556 277780
rect 648724 277394 648752 277780
rect 648632 277366 648752 277394
rect 647516 275324 647568 275330
rect 647516 275266 647568 275272
rect 648632 267073 648660 277366
rect 648618 267064 648674 267073
rect 648618 266999 648674 267008
rect 646056 248386 646176 248414
rect 621664 242956 621716 242962
rect 621664 242898 621716 242904
rect 604460 231736 604512 231742
rect 604460 231678 604512 231684
rect 604472 230518 604500 231678
rect 604460 230512 604512 230518
rect 604460 230454 604512 230460
rect 605748 230512 605800 230518
rect 605748 230454 605800 230460
rect 574744 222148 574796 222154
rect 574744 222090 574796 222096
rect 575480 222148 575532 222154
rect 575480 222090 575532 222096
rect 574928 220584 574980 220590
rect 574928 220526 574980 220532
rect 574836 220380 574888 220386
rect 574836 220322 574888 220328
rect 571812 217382 572240 217410
rect 572732 217382 573068 217410
rect 573468 217382 573896 217410
rect 574296 217382 574724 217410
rect 558840 216730 558868 217382
rect 561416 216782 561444 217382
rect 564084 216850 564112 217382
rect 564072 216844 564124 216850
rect 564072 216786 564124 216792
rect 561404 216776 561456 216782
rect 558840 216714 558960 216730
rect 561404 216718 561456 216724
rect 558840 216708 558972 216714
rect 558840 216702 558920 216708
rect 558920 216650 558972 216656
rect 550836 216442 551508 216458
rect 566476 216442 566504 217382
rect 574848 216442 574876 220322
rect 574940 216442 574968 220526
rect 575492 217410 575520 222090
rect 576400 220788 576452 220794
rect 576400 220730 576452 220736
rect 576308 220448 576360 220454
rect 576308 220390 576360 220396
rect 576216 219088 576268 219094
rect 576216 219030 576268 219036
rect 576032 218612 576084 218618
rect 576032 218554 576084 218560
rect 575940 218476 575992 218482
rect 575940 218418 575992 218424
rect 575848 217660 575900 217666
rect 575848 217602 575900 217608
rect 575492 217382 575552 217410
rect 575756 216776 575808 216782
rect 575756 216718 575808 216724
rect 575664 216708 575716 216714
rect 575664 216650 575716 216656
rect 118700 216436 118752 216442
rect 118700 216378 118752 216384
rect 518716 216436 518768 216442
rect 520476 216436 521252 216442
rect 520476 216430 521200 216436
rect 518716 216378 518768 216384
rect 523144 216436 523828 216442
rect 523144 216430 523776 216436
rect 521200 216378 521252 216384
rect 523776 216378 523828 216384
rect 526260 216436 526312 216442
rect 528448 216436 528612 216442
rect 528448 216430 528560 216436
rect 526260 216378 526312 216384
rect 530596 216436 531280 216442
rect 530596 216430 531228 216436
rect 528560 216378 528612 216384
rect 533080 216436 533856 216442
rect 533080 216430 533804 216436
rect 531228 216378 531280 216384
rect 533804 216378 533856 216384
rect 536380 216436 536432 216442
rect 538324 216436 538916 216442
rect 538324 216430 538864 216436
rect 536380 216378 536432 216384
rect 538864 216378 538916 216384
rect 541440 216436 541492 216442
rect 550836 216436 551520 216442
rect 550836 216430 551468 216436
rect 541440 216378 541492 216384
rect 551468 216378 551520 216384
rect 566464 216436 566516 216442
rect 566464 216378 566516 216384
rect 574836 216436 574888 216442
rect 574836 216378 574888 216384
rect 574928 216436 574980 216442
rect 574928 216378 574980 216384
rect 575676 213382 575704 216650
rect 575664 213376 575716 213382
rect 575664 213318 575716 213324
rect 575768 213314 575796 216718
rect 575860 213518 575888 217602
rect 575952 213926 575980 218418
rect 575940 213920 575992 213926
rect 575940 213862 575992 213868
rect 576044 213858 576072 218554
rect 576124 218544 576176 218550
rect 576124 218486 576176 218492
rect 576032 213852 576084 213858
rect 576032 213794 576084 213800
rect 576136 213722 576164 218486
rect 576124 213716 576176 213722
rect 576124 213658 576176 213664
rect 576228 213654 576256 219030
rect 576320 214606 576348 220390
rect 576412 214810 576440 220730
rect 577320 220720 577372 220726
rect 577320 220662 577372 220668
rect 576492 220652 576544 220658
rect 576492 220594 576544 220600
rect 576400 214804 576452 214810
rect 576400 214746 576452 214752
rect 576308 214600 576360 214606
rect 576308 214542 576360 214548
rect 576216 213648 576268 213654
rect 576216 213590 576268 213596
rect 576504 213586 576532 220594
rect 577136 220516 577188 220522
rect 577136 220458 577188 220464
rect 577044 216844 577096 216850
rect 577044 216786 577096 216792
rect 576492 213580 576544 213586
rect 576492 213522 576544 213528
rect 575848 213512 575900 213518
rect 575848 213454 575900 213460
rect 577056 213450 577084 216786
rect 577148 214742 577176 220458
rect 577136 214736 577188 214742
rect 577136 214678 577188 214684
rect 577332 214674 577360 220662
rect 577504 219156 577556 219162
rect 577504 219098 577556 219104
rect 577320 214668 577372 214674
rect 577320 214610 577372 214616
rect 577044 213444 577096 213450
rect 577044 213386 577096 213392
rect 575756 213308 575808 213314
rect 575756 213250 575808 213256
rect 577516 213246 577544 219098
rect 578148 217388 578200 217394
rect 578148 217330 578200 217336
rect 577872 216096 577924 216102
rect 577872 216038 577924 216044
rect 577884 213790 577912 216038
rect 577872 213784 577924 213790
rect 577872 213726 577924 213732
rect 577504 213240 577556 213246
rect 577504 213182 577556 213188
rect 578160 213178 578188 217330
rect 578882 216200 578938 216209
rect 578882 216135 578938 216144
rect 578148 213172 578200 213178
rect 578148 213114 578200 213120
rect 578422 211712 578478 211721
rect 578422 211647 578478 211656
rect 578436 206990 578464 211647
rect 578514 210216 578570 210225
rect 578514 210151 578570 210160
rect 578424 206984 578476 206990
rect 578424 206926 578476 206932
rect 578528 205630 578556 210151
rect 578896 209778 578924 216135
rect 579250 214704 579306 214713
rect 579250 214639 579306 214648
rect 578974 213208 579030 213217
rect 578974 213143 579030 213152
rect 578884 209772 578936 209778
rect 578884 209714 578936 209720
rect 578988 208350 579016 213143
rect 579264 209710 579292 214639
rect 583024 211200 583076 211206
rect 583024 211142 583076 211148
rect 579252 209704 579304 209710
rect 579252 209646 579304 209652
rect 579526 208720 579582 208729
rect 579526 208655 579582 208664
rect 578976 208344 579028 208350
rect 578976 208286 579028 208292
rect 578790 207224 578846 207233
rect 578790 207159 578846 207168
rect 578516 205624 578568 205630
rect 578516 205566 578568 205572
rect 578804 204270 578832 207159
rect 579434 205728 579490 205737
rect 579434 205663 579490 205672
rect 578792 204264 578844 204270
rect 578792 204206 578844 204212
rect 578882 204232 578938 204241
rect 578882 204167 578938 204176
rect 578896 201482 578924 204167
rect 579448 202842 579476 205663
rect 579540 205562 579568 208655
rect 579528 205556 579580 205562
rect 579528 205498 579580 205504
rect 579436 202836 579488 202842
rect 579436 202778 579488 202784
rect 579250 202736 579306 202745
rect 579250 202671 579306 202680
rect 578884 201476 578936 201482
rect 578884 201418 578936 201424
rect 579264 201414 579292 202671
rect 579252 201408 579304 201414
rect 579252 201350 579304 201356
rect 578238 201240 578294 201249
rect 578238 201175 578294 201184
rect 578252 200122 578280 201175
rect 578240 200116 578292 200122
rect 578240 200058 578292 200064
rect 578422 199744 578478 199753
rect 578422 199679 578478 199688
rect 578436 198694 578464 199679
rect 578424 198688 578476 198694
rect 578424 198630 578476 198636
rect 579066 198248 579122 198257
rect 579066 198183 579122 198192
rect 579080 197334 579108 198183
rect 579068 197328 579120 197334
rect 579068 197270 579120 197276
rect 579526 196752 579582 196761
rect 579526 196687 579582 196696
rect 579540 196654 579568 196687
rect 579528 196648 579580 196654
rect 579528 196590 579580 196596
rect 579528 195288 579580 195294
rect 579526 195256 579528 195265
rect 579580 195256 579582 195265
rect 579526 195191 579582 195200
rect 579528 193860 579580 193866
rect 579528 193802 579580 193808
rect 579540 193633 579568 193802
rect 579526 193624 579582 193633
rect 579526 193559 579582 193568
rect 579528 192500 579580 192506
rect 579528 192442 579580 192448
rect 579540 192137 579568 192442
rect 579526 192128 579582 192137
rect 579526 192063 579582 192072
rect 579252 191888 579304 191894
rect 579252 191830 579304 191836
rect 579264 190641 579292 191830
rect 579250 190632 579306 190641
rect 579250 190567 579306 190576
rect 578240 190528 578292 190534
rect 578240 190470 578292 190476
rect 578252 189145 578280 190470
rect 579528 189168 579580 189174
rect 578238 189136 578294 189145
rect 579528 189110 579580 189116
rect 578238 189071 578294 189080
rect 579252 189100 579304 189106
rect 579252 189042 579304 189048
rect 578884 187740 578936 187746
rect 578884 187682 578936 187688
rect 578896 184657 578924 187682
rect 579264 187649 579292 189042
rect 579250 187640 579306 187649
rect 579250 187575 579306 187584
rect 579436 186380 579488 186386
rect 579436 186322 579488 186328
rect 578976 184952 579028 184958
rect 578976 184894 579028 184900
rect 578882 184648 578938 184657
rect 578882 184583 578938 184592
rect 578240 182232 578292 182238
rect 578240 182174 578292 182180
rect 578252 177177 578280 182174
rect 578332 180940 578384 180946
rect 578332 180882 578384 180888
rect 578238 177168 578294 177177
rect 578238 177103 578294 177112
rect 578344 175681 578372 180882
rect 578424 180872 578476 180878
rect 578424 180814 578476 180820
rect 578330 175672 578386 175681
rect 578330 175607 578386 175616
rect 578436 174185 578464 180814
rect 578988 180794 579016 184894
rect 579344 183592 579396 183598
rect 579344 183534 579396 183540
rect 578896 180766 579016 180794
rect 578896 180169 578924 180766
rect 578882 180160 578938 180169
rect 578882 180095 578938 180104
rect 578792 179444 578844 179450
rect 578792 179386 578844 179392
rect 578700 178084 578752 178090
rect 578700 178026 578752 178032
rect 578422 174176 578478 174185
rect 578422 174111 578478 174120
rect 578712 171193 578740 178026
rect 578804 172689 578832 179386
rect 579356 178673 579384 183534
rect 579448 183161 579476 186322
rect 579540 186153 579568 189110
rect 579526 186144 579582 186153
rect 579526 186079 579582 186088
rect 579528 185020 579580 185026
rect 579528 184962 579580 184968
rect 579434 183152 579490 183161
rect 579434 183087 579490 183096
rect 579540 181665 579568 184962
rect 579526 181656 579582 181665
rect 579526 181591 579582 181600
rect 579342 178664 579398 178673
rect 579342 178599 579398 178608
rect 579436 176792 579488 176798
rect 579436 176734 579488 176740
rect 579344 176724 579396 176730
rect 579344 176666 579396 176672
rect 578790 172680 578846 172689
rect 578790 172615 578846 172624
rect 579160 172576 579212 172582
rect 579160 172518 579212 172524
rect 578698 171184 578754 171193
rect 578698 171119 578754 171128
rect 579068 169856 579120 169862
rect 579068 169798 579120 169804
rect 578884 169788 578936 169794
rect 578884 169730 578936 169736
rect 578608 167000 578660 167006
rect 578608 166942 578660 166948
rect 578620 166569 578648 166942
rect 578606 166560 578662 166569
rect 578606 166495 578662 166504
rect 578240 164484 578292 164490
rect 578240 164426 578292 164432
rect 578252 164393 578280 164426
rect 578238 164384 578294 164393
rect 578238 164319 578294 164328
rect 578896 157593 578924 169730
rect 578976 168428 579028 168434
rect 578976 168370 579028 168376
rect 578882 157584 578938 157593
rect 578882 157519 578938 157528
rect 578988 156097 579016 168370
rect 579080 159089 579108 169798
rect 579172 162081 579200 172518
rect 579252 171148 579304 171154
rect 579252 171090 579304 171096
rect 579158 162072 579214 162081
rect 579158 162007 579214 162016
rect 579264 160585 579292 171090
rect 579356 168065 579384 176666
rect 579448 169561 579476 176734
rect 580264 175296 580316 175302
rect 580264 175238 580316 175244
rect 579434 169552 579490 169561
rect 579434 169487 579490 169496
rect 579342 168056 579398 168065
rect 579342 167991 579398 168000
rect 580276 167006 580304 175238
rect 580356 173936 580408 173942
rect 580356 173878 580408 173884
rect 580264 167000 580316 167006
rect 580264 166942 580316 166948
rect 580368 164490 580396 173878
rect 581644 165640 581696 165646
rect 581644 165582 581696 165588
rect 580356 164484 580408 164490
rect 580356 164426 580408 164432
rect 579528 164212 579580 164218
rect 579528 164154 579580 164160
rect 579540 163577 579568 164154
rect 579526 163568 579582 163577
rect 579526 163503 579582 163512
rect 580264 162920 580316 162926
rect 580264 162862 580316 162868
rect 579250 160576 579306 160585
rect 579250 160511 579306 160520
rect 579160 160132 579212 160138
rect 579160 160074 579212 160080
rect 579066 159080 579122 159089
rect 579066 159015 579122 159024
rect 578974 156088 579030 156097
rect 578974 156023 579030 156032
rect 578332 154896 578384 154902
rect 578332 154838 578384 154844
rect 578344 154601 578372 154838
rect 578330 154592 578386 154601
rect 578330 154527 578386 154536
rect 579068 153332 579120 153338
rect 579068 153274 579120 153280
rect 578884 153264 578936 153270
rect 578884 153206 578936 153212
rect 578516 148640 578568 148646
rect 578514 148608 578516 148617
rect 578568 148608 578570 148617
rect 578514 148543 578570 148552
rect 578700 146192 578752 146198
rect 578700 146134 578752 146140
rect 578712 145489 578740 146134
rect 578698 145480 578754 145489
rect 578698 145415 578754 145424
rect 578700 143540 578752 143546
rect 578700 143482 578752 143488
rect 578712 142497 578740 143482
rect 578698 142488 578754 142497
rect 578698 142423 578754 142432
rect 578896 132025 578924 153206
rect 578976 150476 579028 150482
rect 578976 150418 579028 150424
rect 578882 132016 578938 132025
rect 578882 131951 578938 131960
rect 578332 130552 578384 130558
rect 578330 130520 578332 130529
rect 578384 130520 578386 130529
rect 578330 130455 578386 130464
rect 578988 129033 579016 150418
rect 579080 133521 579108 153274
rect 579172 139505 579200 160074
rect 579344 158772 579396 158778
rect 579344 158714 579396 158720
rect 579252 154624 579304 154630
rect 579252 154566 579304 154572
rect 579158 139496 579214 139505
rect 579158 139431 579214 139440
rect 579264 135017 579292 154566
rect 579356 141001 579384 158714
rect 579528 153196 579580 153202
rect 579528 153138 579580 153144
rect 579540 153105 579568 153138
rect 579526 153096 579582 153105
rect 579526 153031 579582 153040
rect 579436 151632 579488 151638
rect 579434 151600 579436 151609
rect 579488 151600 579490 151609
rect 579434 151535 579490 151544
rect 579436 150272 579488 150278
rect 579436 150214 579488 150220
rect 579448 150113 579476 150214
rect 579434 150104 579490 150113
rect 579434 150039 579490 150048
rect 580276 148646 580304 162862
rect 580356 151836 580408 151842
rect 580356 151778 580408 151784
rect 580264 148640 580316 148646
rect 580264 148582 580316 148588
rect 579528 147008 579580 147014
rect 579526 146976 579528 146985
rect 579580 146976 579582 146985
rect 579526 146911 579582 146920
rect 579620 146940 579672 146946
rect 579620 146882 579672 146888
rect 579526 143984 579582 143993
rect 579632 143970 579660 146882
rect 579582 143942 579660 143970
rect 579526 143919 579582 143928
rect 580264 143608 580316 143614
rect 580264 143550 580316 143556
rect 579342 140992 579398 141001
rect 579342 140927 579398 140936
rect 579526 138000 579582 138009
rect 579526 137935 579528 137944
rect 579580 137935 579582 137944
rect 579528 137906 579580 137912
rect 579528 136536 579580 136542
rect 579526 136504 579528 136513
rect 579580 136504 579582 136513
rect 579526 136439 579582 136448
rect 579250 135008 579306 135017
rect 579250 134943 579306 134952
rect 579066 133512 579122 133521
rect 579066 133447 579122 133456
rect 578974 129024 579030 129033
rect 578974 128959 579030 128968
rect 579528 128308 579580 128314
rect 579528 128250 579580 128256
rect 579540 127537 579568 128250
rect 579526 127528 579582 127537
rect 579526 127463 579582 127472
rect 578700 126064 578752 126070
rect 578698 126032 578700 126041
rect 578752 126032 578754 126041
rect 578698 125967 578754 125976
rect 578424 125588 578476 125594
rect 578424 125530 578476 125536
rect 578436 124545 578464 125530
rect 578422 124536 578478 124545
rect 578422 124471 578478 124480
rect 579252 124160 579304 124166
rect 579252 124102 579304 124108
rect 579264 122913 579292 124102
rect 579250 122904 579306 122913
rect 579250 122839 579306 122848
rect 579436 122120 579488 122126
rect 579436 122062 579488 122068
rect 579252 120080 579304 120086
rect 579252 120022 579304 120028
rect 579264 119921 579292 120022
rect 579250 119912 579306 119921
rect 579250 119847 579306 119856
rect 579160 118720 579212 118726
rect 579160 118662 579212 118668
rect 578516 118584 578568 118590
rect 578516 118526 578568 118532
rect 578528 118425 578556 118526
rect 578514 118416 578570 118425
rect 578514 118351 578570 118360
rect 579068 117360 579120 117366
rect 579068 117302 579120 117308
rect 578976 114572 579028 114578
rect 578976 114514 579028 114520
rect 578884 113212 578936 113218
rect 578884 113154 578936 113160
rect 578700 111784 578752 111790
rect 578700 111726 578752 111732
rect 578712 110945 578740 111726
rect 578698 110936 578754 110945
rect 578698 110871 578754 110880
rect 578792 108996 578844 109002
rect 578792 108938 578844 108944
rect 578804 107953 578832 108938
rect 578790 107944 578846 107953
rect 578790 107879 578846 107888
rect 578240 105188 578292 105194
rect 578240 105130 578292 105136
rect 578252 104961 578280 105130
rect 578238 104952 578294 104961
rect 578238 104887 578294 104896
rect 578332 102128 578384 102134
rect 578332 102070 578384 102076
rect 578344 101969 578372 102070
rect 578330 101960 578386 101969
rect 578330 101895 578386 101904
rect 578700 100360 578752 100366
rect 578698 100328 578700 100337
rect 578752 100328 578754 100337
rect 578698 100263 578754 100272
rect 578700 97640 578752 97646
rect 578700 97582 578752 97588
rect 578712 97345 578740 97582
rect 578698 97336 578754 97345
rect 578698 97271 578754 97280
rect 578516 96008 578568 96014
rect 578516 95950 578568 95956
rect 578528 95849 578556 95950
rect 578514 95840 578570 95849
rect 578514 95775 578570 95784
rect 578608 95192 578660 95198
rect 578608 95134 578660 95140
rect 578620 94353 578648 95134
rect 578606 94344 578662 94353
rect 578606 94279 578662 94288
rect 576124 77308 576176 77314
rect 576124 77250 576176 77256
rect 405096 53168 405148 53174
rect 405096 53110 405148 53116
rect 145380 53100 145432 53106
rect 145380 53042 145432 53048
rect 84824 52686 85160 52714
rect 52276 52488 52328 52494
rect 52182 52456 52238 52465
rect 52276 52430 52328 52436
rect 52182 52391 52238 52400
rect 85132 50289 85160 52686
rect 145392 50810 145420 53042
rect 150314 52465 150342 52700
rect 215832 52686 216168 52714
rect 281336 52686 281488 52714
rect 150300 52456 150356 52465
rect 150300 52391 150356 52400
rect 145084 50782 145420 50810
rect 216140 50425 216168 52686
rect 281460 50561 281488 52686
rect 346826 52494 346854 52700
rect 346814 52488 346866 52494
rect 346814 52430 346866 52436
rect 281446 50552 281502 50561
rect 281446 50487 281502 50496
rect 216126 50416 216182 50425
rect 216126 50351 216182 50360
rect 85118 50280 85174 50289
rect 85118 50215 85174 50224
rect 142356 44305 142384 46716
rect 194048 46232 194100 46238
rect 194048 46174 194100 46180
rect 142342 44296 142398 44305
rect 142342 44231 142398 44240
rect 187514 42120 187570 42129
rect 187358 42078 187514 42106
rect 194060 42092 194088 46174
rect 307298 43480 307354 43489
rect 307298 43415 307354 43424
rect 307312 42106 307340 43415
rect 310104 42392 310160 42401
rect 310104 42327 310160 42336
rect 307004 42078 307340 42106
rect 310118 42092 310146 42327
rect 361946 42120 362002 42129
rect 361790 42078 361946 42106
rect 187514 42055 187570 42064
rect 365074 42120 365130 42129
rect 364918 42078 365074 42106
rect 361946 42055 362002 42064
rect 405108 42106 405136 53110
rect 412344 52686 412496 52714
rect 477848 52686 478184 52714
rect 412468 46753 412496 52686
rect 478156 49774 478184 52686
rect 543016 52686 543352 52714
rect 543016 50289 543044 52686
rect 543002 50280 543058 50289
rect 543002 50215 543058 50224
rect 478144 49768 478196 49774
rect 478144 49710 478196 49716
rect 478788 49768 478840 49774
rect 478788 49710 478840 49716
rect 473174 47696 473230 47705
rect 473174 47631 473230 47640
rect 412454 46744 412510 46753
rect 412454 46679 412510 46688
rect 470138 46472 470194 46481
rect 470138 46407 470194 46416
rect 415122 46200 415178 46209
rect 415122 46135 415178 46144
rect 415136 42398 415164 46135
rect 419722 45248 419778 45257
rect 419722 45183 419778 45192
rect 419736 42772 419764 45183
rect 415124 42392 415176 42398
rect 415124 42334 415176 42340
rect 460570 42120 460626 42129
rect 405108 42078 405582 42106
rect 460368 42078 460570 42106
rect 365074 42055 365130 42064
rect 460570 42055 460626 42064
rect 416686 41848 416742 41857
rect 416622 41806 416686 41834
rect 470152 41820 470180 46407
rect 473188 42534 473216 47631
rect 473176 42528 473228 42534
rect 473176 42470 473228 42476
rect 471610 42120 471666 42129
rect 471408 42078 471610 42106
rect 471610 42055 471666 42064
rect 416686 41783 416742 41792
rect 478800 41585 478828 49710
rect 576136 47569 576164 77250
rect 578896 73273 578924 113154
rect 578988 76265 579016 114514
rect 579080 79393 579108 117302
rect 579172 82385 579200 118662
rect 579448 115433 579476 122062
rect 579528 121440 579580 121446
rect 579526 121408 579528 121417
rect 579580 121408 579582 121417
rect 579526 121343 579582 121352
rect 580276 118590 580304 143550
rect 580368 130558 580396 151778
rect 581656 151638 581684 165582
rect 581736 164280 581788 164286
rect 581736 164222 581788 164228
rect 581644 151632 581696 151638
rect 581644 151574 581696 151580
rect 581748 150278 581776 164222
rect 581736 150272 581788 150278
rect 581736 150214 581788 150220
rect 583036 147014 583064 211142
rect 603080 209772 603132 209778
rect 603080 209714 603132 209720
rect 603092 209545 603120 209714
rect 603172 209704 603224 209710
rect 603172 209646 603224 209652
rect 603078 209536 603134 209545
rect 603078 209471 603134 209480
rect 603184 208593 603212 209646
rect 603170 208584 603226 208593
rect 603170 208519 603226 208528
rect 603080 208344 603132 208350
rect 603080 208286 603132 208292
rect 603092 207505 603120 208286
rect 603078 207496 603134 207505
rect 603078 207431 603134 207440
rect 603080 206984 603132 206990
rect 603080 206926 603132 206932
rect 603092 206553 603120 206926
rect 603078 206544 603134 206553
rect 603078 206479 603134 206488
rect 603080 205624 603132 205630
rect 603080 205566 603132 205572
rect 603092 205465 603120 205566
rect 603172 205556 603224 205562
rect 603172 205498 603224 205504
rect 603078 205456 603134 205465
rect 603078 205391 603134 205400
rect 603184 204513 603212 205498
rect 603170 204504 603226 204513
rect 603170 204439 603226 204448
rect 603080 204264 603132 204270
rect 603080 204206 603132 204212
rect 603092 203425 603120 204206
rect 603078 203416 603134 203425
rect 603078 203351 603134 203360
rect 603080 202836 603132 202842
rect 603080 202778 603132 202784
rect 603092 202473 603120 202778
rect 603078 202464 603134 202473
rect 603078 202399 603134 202408
rect 603080 201476 603132 201482
rect 603080 201418 603132 201424
rect 603092 201385 603120 201418
rect 603172 201408 603224 201414
rect 603078 201376 603134 201385
rect 603172 201350 603224 201356
rect 603078 201311 603134 201320
rect 603184 200433 603212 201350
rect 603170 200424 603226 200433
rect 603170 200359 603226 200368
rect 603080 200116 603132 200122
rect 603080 200058 603132 200064
rect 603092 199345 603120 200058
rect 603078 199336 603134 199345
rect 603078 199271 603134 199280
rect 603080 198688 603132 198694
rect 603080 198630 603132 198636
rect 603092 198393 603120 198630
rect 603078 198384 603134 198393
rect 603078 198319 603134 198328
rect 603172 197328 603224 197334
rect 603078 197296 603134 197305
rect 603172 197270 603224 197276
rect 603078 197231 603134 197240
rect 603092 196654 603120 197231
rect 603080 196648 603132 196654
rect 603080 196590 603132 196596
rect 603184 196353 603212 197270
rect 603170 196344 603226 196353
rect 603170 196279 603226 196288
rect 603080 195288 603132 195294
rect 603078 195256 603080 195265
rect 603132 195256 603134 195265
rect 603078 195191 603134 195200
rect 603078 194304 603134 194313
rect 603078 194239 603134 194248
rect 603092 193866 603120 194239
rect 603080 193860 603132 193866
rect 603080 193802 603132 193808
rect 603078 193216 603134 193225
rect 603078 193151 603134 193160
rect 603092 192506 603120 193151
rect 603080 192500 603132 192506
rect 603080 192442 603132 192448
rect 603078 192264 603134 192273
rect 603078 192199 603134 192208
rect 603092 191894 603120 192199
rect 603080 191888 603132 191894
rect 603080 191830 603132 191836
rect 603078 191176 603134 191185
rect 603078 191111 603134 191120
rect 603092 190534 603120 191111
rect 603080 190528 603132 190534
rect 603080 190470 603132 190476
rect 603170 190224 603226 190233
rect 603170 190159 603226 190168
rect 603080 189168 603132 189174
rect 603078 189136 603080 189145
rect 603132 189136 603134 189145
rect 603184 189106 603212 190159
rect 603078 189071 603134 189080
rect 603172 189100 603224 189106
rect 603172 189042 603224 189048
rect 603078 188184 603134 188193
rect 603078 188119 603134 188128
rect 603092 187746 603120 188119
rect 603080 187740 603132 187746
rect 603080 187682 603132 187688
rect 603078 187096 603134 187105
rect 603078 187031 603134 187040
rect 603092 186386 603120 187031
rect 603080 186380 603132 186386
rect 603080 186322 603132 186328
rect 603170 186144 603226 186153
rect 603170 186079 603226 186088
rect 603078 185056 603134 185065
rect 603184 185026 603212 186079
rect 603078 184991 603134 185000
rect 603172 185020 603224 185026
rect 603092 184958 603120 184991
rect 603172 184962 603224 184968
rect 603080 184952 603132 184958
rect 603080 184894 603132 184900
rect 603078 184104 603134 184113
rect 603078 184039 603134 184048
rect 603092 183598 603120 184039
rect 603080 183592 603132 183598
rect 603080 183534 603132 183540
rect 603078 183016 603134 183025
rect 603078 182951 603134 182960
rect 603092 182238 603120 182951
rect 603080 182232 603132 182238
rect 603080 182174 603132 182180
rect 603170 182064 603226 182073
rect 603170 181999 603226 182008
rect 603078 180976 603134 180985
rect 603184 180946 603212 181999
rect 603078 180911 603134 180920
rect 603172 180940 603224 180946
rect 603092 180878 603120 180911
rect 603172 180882 603224 180888
rect 603080 180872 603132 180878
rect 603080 180814 603132 180820
rect 603078 180024 603134 180033
rect 603078 179959 603134 179968
rect 603092 179450 603120 179959
rect 603080 179444 603132 179450
rect 603080 179386 603132 179392
rect 603078 178936 603134 178945
rect 603078 178871 603134 178880
rect 603092 178090 603120 178871
rect 603080 178084 603132 178090
rect 603080 178026 603132 178032
rect 603170 177984 603226 177993
rect 603170 177919 603226 177928
rect 603078 176896 603134 176905
rect 603078 176831 603134 176840
rect 603092 176730 603120 176831
rect 603184 176798 603212 177919
rect 603172 176792 603224 176798
rect 603172 176734 603224 176740
rect 603080 176724 603132 176730
rect 603080 176666 603132 176672
rect 603078 175944 603134 175953
rect 603078 175879 603134 175888
rect 603092 175302 603120 175879
rect 603080 175296 603132 175302
rect 603080 175238 603132 175244
rect 603078 174856 603134 174865
rect 603078 174791 603134 174800
rect 603092 173942 603120 174791
rect 603080 173936 603132 173942
rect 603080 173878 603132 173884
rect 603722 173904 603778 173913
rect 603722 173839 603778 173848
rect 603078 172816 603134 172825
rect 603078 172751 603134 172760
rect 603092 172582 603120 172751
rect 603080 172576 603132 172582
rect 603080 172518 603132 172524
rect 603078 171864 603134 171873
rect 603078 171799 603134 171808
rect 603092 171154 603120 171799
rect 603080 171148 603132 171154
rect 603080 171090 603132 171096
rect 603170 170776 603226 170785
rect 603170 170711 603226 170720
rect 603184 169862 603212 170711
rect 603172 169856 603224 169862
rect 603078 169824 603134 169833
rect 603172 169798 603224 169804
rect 603078 169759 603080 169768
rect 603132 169759 603134 169768
rect 603080 169730 603132 169736
rect 603078 168736 603134 168745
rect 603078 168671 603134 168680
rect 603092 168434 603120 168671
rect 603080 168428 603132 168434
rect 603080 168370 603132 168376
rect 603078 167784 603134 167793
rect 603078 167719 603134 167728
rect 603092 167074 603120 167719
rect 583116 167068 583168 167074
rect 583116 167010 583168 167016
rect 603080 167068 603132 167074
rect 603080 167010 603132 167016
rect 583128 154902 583156 167010
rect 603078 165744 603134 165753
rect 603078 165679 603134 165688
rect 603092 165646 603120 165679
rect 603080 165640 603132 165646
rect 603080 165582 603132 165588
rect 603078 164656 603134 164665
rect 603078 164591 603134 164600
rect 603092 164286 603120 164591
rect 603080 164280 603132 164286
rect 603080 164222 603132 164228
rect 603736 164218 603764 173839
rect 603814 166696 603870 166705
rect 603814 166631 603870 166640
rect 603724 164212 603776 164218
rect 603724 164154 603776 164160
rect 603078 163704 603134 163713
rect 603078 163639 603134 163648
rect 603092 162926 603120 163639
rect 603080 162920 603132 162926
rect 603080 162862 603132 162868
rect 603078 162616 603134 162625
rect 603078 162551 603134 162560
rect 603092 161498 603120 162551
rect 603722 161664 603778 161673
rect 603722 161599 603778 161608
rect 584496 161492 584548 161498
rect 584496 161434 584548 161440
rect 603080 161492 603132 161498
rect 603080 161434 603132 161440
rect 584404 157412 584456 157418
rect 584404 157354 584456 157360
rect 583116 154896 583168 154902
rect 583116 154838 583168 154844
rect 583024 147008 583076 147014
rect 583024 146950 583076 146956
rect 583024 144968 583076 144974
rect 583024 144910 583076 144916
rect 581828 133952 581880 133958
rect 581828 133894 581880 133900
rect 581644 133204 581696 133210
rect 581644 133146 581696 133152
rect 580356 130552 580408 130558
rect 580356 130494 580408 130500
rect 580356 127016 580408 127022
rect 580356 126958 580408 126964
rect 580264 118584 580316 118590
rect 580264 118526 580316 118532
rect 579528 117292 579580 117298
rect 579528 117234 579580 117240
rect 579540 116929 579568 117234
rect 579526 116920 579582 116929
rect 579526 116855 579582 116864
rect 579434 115424 579490 115433
rect 579434 115359 579490 115368
rect 579252 114504 579304 114510
rect 579252 114446 579304 114452
rect 579264 113937 579292 114446
rect 579250 113928 579306 113937
rect 579250 113863 579306 113872
rect 579528 113144 579580 113150
rect 579528 113086 579580 113092
rect 579540 112441 579568 113086
rect 579526 112432 579582 112441
rect 579526 112367 579582 112376
rect 579528 110424 579580 110430
rect 579528 110366 579580 110372
rect 579540 109449 579568 110366
rect 579526 109440 579582 109449
rect 579526 109375 579582 109384
rect 579436 107092 579488 107098
rect 579436 107034 579488 107040
rect 579448 106457 579476 107034
rect 579434 106448 579490 106457
rect 579434 106383 579490 106392
rect 579344 103488 579396 103494
rect 579342 103456 579344 103465
rect 579396 103456 579398 103465
rect 579342 103391 579398 103400
rect 580264 100768 580316 100774
rect 580264 100710 580316 100716
rect 579528 99136 579580 99142
rect 579528 99078 579580 99084
rect 579540 98841 579568 99078
rect 579526 98832 579582 98841
rect 579526 98767 579582 98776
rect 579528 93832 579580 93838
rect 579528 93774 579580 93780
rect 579540 92857 579568 93774
rect 579526 92848 579582 92857
rect 579526 92783 579582 92792
rect 579528 92472 579580 92478
rect 579528 92414 579580 92420
rect 579540 91361 579568 92414
rect 579526 91352 579582 91361
rect 579526 91287 579582 91296
rect 579528 91044 579580 91050
rect 579528 90986 579580 90992
rect 579540 89865 579568 90986
rect 579526 89856 579582 89865
rect 579526 89791 579582 89800
rect 579528 89684 579580 89690
rect 579528 89626 579580 89632
rect 579540 88369 579568 89626
rect 579526 88360 579582 88369
rect 579526 88295 579582 88304
rect 579528 86964 579580 86970
rect 579528 86906 579580 86912
rect 579540 86873 579568 86906
rect 579526 86864 579582 86873
rect 579526 86799 579582 86808
rect 579528 85536 579580 85542
rect 579528 85478 579580 85484
rect 579540 85377 579568 85478
rect 579526 85368 579582 85377
rect 579526 85303 579582 85312
rect 579528 84176 579580 84182
rect 579528 84118 579580 84124
rect 579540 83881 579568 84118
rect 579526 83872 579582 83881
rect 579526 83807 579582 83816
rect 579158 82376 579214 82385
rect 579158 82311 579214 82320
rect 579528 80912 579580 80918
rect 579526 80880 579528 80889
rect 579580 80880 579582 80889
rect 579526 80815 579582 80824
rect 579066 79384 579122 79393
rect 579066 79319 579122 79328
rect 579528 78668 579580 78674
rect 579528 78610 579580 78616
rect 579540 77897 579568 78610
rect 579526 77888 579582 77897
rect 579526 77823 579582 77832
rect 579068 77376 579120 77382
rect 579068 77318 579120 77324
rect 578974 76256 579030 76265
rect 578974 76191 579030 76200
rect 578882 73264 578938 73273
rect 578882 73199 578938 73208
rect 578700 69012 578752 69018
rect 578700 68954 578752 68960
rect 578712 68785 578740 68954
rect 578698 68776 578754 68785
rect 578698 68711 578754 68720
rect 578700 64864 578752 64870
rect 578700 64806 578752 64812
rect 578712 64297 578740 64806
rect 578698 64288 578754 64297
rect 578698 64223 578754 64232
rect 578700 62076 578752 62082
rect 578700 62018 578752 62024
rect 578712 61305 578740 62018
rect 578698 61296 578754 61305
rect 578698 61231 578754 61240
rect 578884 60716 578936 60722
rect 578884 60658 578936 60664
rect 578896 59809 578924 60658
rect 578882 59800 578938 59809
rect 578882 59735 578938 59744
rect 578884 58812 578936 58818
rect 578884 58754 578936 58760
rect 578896 58313 578924 58754
rect 578882 58304 578938 58313
rect 578882 58239 578938 58248
rect 578884 57928 578936 57934
rect 578884 57870 578936 57876
rect 578332 57248 578384 57254
rect 578332 57190 578384 57196
rect 578240 55684 578292 55690
rect 578240 55626 578292 55632
rect 578252 55321 578280 55626
rect 578238 55312 578294 55321
rect 578238 55247 578294 55256
rect 578344 53825 578372 57190
rect 578896 56817 578924 57870
rect 578882 56808 578938 56817
rect 578882 56743 578938 56752
rect 578330 53816 578386 53825
rect 578330 53751 578386 53760
rect 579080 53106 579108 77318
rect 579528 75880 579580 75886
rect 579528 75822 579580 75828
rect 579540 74769 579568 75822
rect 579526 74760 579582 74769
rect 579526 74695 579582 74704
rect 579526 71768 579582 71777
rect 579526 71703 579528 71712
rect 579580 71703 579582 71712
rect 579528 71674 579580 71680
rect 579252 70304 579304 70310
rect 579250 70272 579252 70281
rect 579304 70272 579306 70281
rect 579250 70207 579306 70216
rect 579528 67584 579580 67590
rect 579528 67526 579580 67532
rect 579540 67289 579568 67526
rect 579526 67280 579582 67289
rect 579526 67215 579582 67224
rect 579528 65952 579580 65958
rect 579528 65894 579580 65900
rect 579540 65793 579568 65894
rect 579526 65784 579582 65793
rect 579526 65719 579582 65728
rect 579528 63504 579580 63510
rect 579528 63446 579580 63452
rect 579540 62801 579568 63446
rect 579526 62792 579582 62801
rect 579526 62727 579582 62736
rect 580276 55690 580304 100710
rect 580368 95198 580396 126958
rect 581656 120086 581684 133146
rect 581736 129804 581788 129810
rect 581736 129746 581788 129752
rect 581644 120080 581696 120086
rect 581644 120022 581696 120028
rect 581644 102196 581696 102202
rect 581644 102138 581696 102144
rect 580356 95192 580408 95198
rect 580356 95134 580408 95140
rect 581656 57934 581684 102138
rect 581748 97646 581776 129746
rect 581840 103494 581868 133894
rect 583036 121446 583064 144910
rect 584416 136542 584444 157354
rect 584508 146198 584536 161434
rect 603078 160576 603134 160585
rect 603078 160511 603134 160520
rect 603092 160138 603120 160511
rect 603080 160132 603132 160138
rect 603080 160074 603132 160080
rect 603078 159624 603134 159633
rect 603078 159559 603134 159568
rect 603092 158778 603120 159559
rect 603080 158772 603132 158778
rect 603080 158714 603132 158720
rect 603170 158536 603226 158545
rect 603170 158471 603226 158480
rect 603078 157584 603134 157593
rect 603078 157519 603134 157528
rect 592684 157480 592736 157486
rect 592684 157422 592736 157428
rect 585784 155984 585836 155990
rect 585784 155926 585836 155932
rect 584496 146192 584548 146198
rect 584496 146134 584548 146140
rect 584680 140072 584732 140078
rect 584680 140014 584732 140020
rect 584404 136536 584456 136542
rect 584404 136478 584456 136484
rect 584588 131164 584640 131170
rect 584588 131106 584640 131112
rect 583116 129872 583168 129878
rect 583116 129814 583168 129820
rect 583024 121440 583076 121446
rect 583024 121382 583076 121388
rect 581828 103488 581880 103494
rect 581828 103430 581880 103436
rect 583024 102264 583076 102270
rect 583024 102206 583076 102212
rect 581736 97640 581788 97646
rect 581736 97582 581788 97588
rect 581736 82136 581788 82142
rect 581736 82078 581788 82084
rect 581748 70310 581776 82078
rect 581736 70304 581788 70310
rect 581736 70246 581788 70252
rect 583036 58818 583064 102206
rect 583128 99142 583156 129814
rect 584496 128376 584548 128382
rect 584496 128318 584548 128324
rect 584404 103556 584456 103562
rect 584404 103498 584456 103504
rect 583116 99136 583168 99142
rect 583116 99078 583168 99084
rect 584416 60722 584444 103498
rect 584508 96014 584536 128318
rect 584600 100366 584628 131106
rect 584692 126070 584720 140014
rect 585796 137970 585824 155926
rect 589924 149116 589976 149122
rect 589924 149058 589976 149064
rect 587256 147688 587308 147694
rect 587256 147630 587308 147636
rect 587164 138032 587216 138038
rect 587164 137974 587216 137980
rect 585784 137964 585836 137970
rect 585784 137906 585836 137912
rect 585784 135312 585836 135318
rect 585784 135254 585836 135260
rect 584680 126064 584732 126070
rect 584680 126006 584732 126012
rect 585796 107098 585824 135254
rect 585968 134020 586020 134026
rect 585968 133962 586020 133968
rect 585876 107704 585928 107710
rect 585876 107646 585928 107652
rect 585784 107092 585836 107098
rect 585784 107034 585836 107040
rect 585784 104916 585836 104922
rect 585784 104858 585836 104864
rect 584588 100360 584640 100366
rect 584588 100302 584640 100308
rect 584496 96008 584548 96014
rect 584496 95950 584548 95956
rect 584496 87644 584548 87650
rect 584496 87586 584548 87592
rect 584508 80918 584536 87586
rect 584496 80912 584548 80918
rect 584496 80854 584548 80860
rect 585796 62082 585824 104858
rect 585888 65958 585916 107646
rect 585980 105194 586008 133962
rect 587176 111790 587204 137974
rect 587268 128314 587296 147630
rect 588636 140820 588688 140826
rect 588636 140762 588688 140768
rect 588544 136672 588596 136678
rect 588544 136614 588596 136620
rect 587256 128308 587308 128314
rect 587256 128250 587308 128256
rect 587256 125656 587308 125662
rect 587256 125598 587308 125604
rect 587164 111784 587216 111790
rect 587164 111726 587216 111732
rect 587164 106344 587216 106350
rect 587164 106286 587216 106292
rect 585968 105188 586020 105194
rect 585968 105130 586020 105136
rect 585876 65952 585928 65958
rect 585876 65894 585928 65900
rect 587176 63510 587204 106286
rect 587268 93838 587296 125598
rect 588556 109002 588584 136614
rect 588648 114510 588676 140762
rect 589936 125594 589964 149058
rect 591304 146328 591356 146334
rect 591304 146270 591356 146276
rect 590108 138100 590160 138106
rect 590108 138042 590160 138048
rect 589924 125588 589976 125594
rect 589924 125530 589976 125536
rect 590016 120148 590068 120154
rect 590016 120090 590068 120096
rect 588636 114504 588688 114510
rect 588636 114446 588688 114452
rect 589924 110492 589976 110498
rect 589924 110434 589976 110440
rect 588636 109064 588688 109070
rect 588636 109006 588688 109012
rect 588544 108996 588596 109002
rect 588544 108938 588596 108944
rect 588544 106412 588596 106418
rect 588544 106354 588596 106360
rect 587256 93832 587308 93838
rect 587256 93774 587308 93780
rect 588556 64870 588584 106354
rect 588648 67590 588676 109006
rect 589936 69018 589964 110434
rect 590028 84182 590056 120090
rect 590120 110430 590148 138042
rect 591316 124166 591344 146270
rect 592696 143546 592724 157422
rect 603092 157418 603120 157519
rect 603184 157486 603212 158471
rect 603172 157480 603224 157486
rect 603172 157422 603224 157428
rect 603080 157412 603132 157418
rect 603080 157354 603132 157360
rect 603078 156496 603134 156505
rect 603078 156431 603134 156440
rect 603092 155990 603120 156431
rect 603080 155984 603132 155990
rect 603080 155926 603132 155932
rect 603078 155544 603134 155553
rect 603078 155479 603134 155488
rect 603092 154630 603120 155479
rect 603080 154624 603132 154630
rect 603080 154566 603132 154572
rect 603170 154456 603226 154465
rect 603170 154391 603226 154400
rect 603078 153504 603134 153513
rect 603078 153439 603134 153448
rect 603092 153270 603120 153439
rect 603184 153338 603212 154391
rect 603172 153332 603224 153338
rect 603172 153274 603224 153280
rect 603080 153264 603132 153270
rect 603080 153206 603132 153212
rect 603078 152416 603134 152425
rect 603078 152351 603134 152360
rect 603092 151842 603120 152351
rect 603080 151836 603132 151842
rect 603080 151778 603132 151784
rect 603078 151464 603134 151473
rect 603078 151399 603134 151408
rect 603092 150482 603120 151399
rect 603080 150476 603132 150482
rect 603080 150418 603132 150424
rect 603078 150376 603134 150385
rect 603078 150311 603134 150320
rect 603092 149122 603120 150311
rect 603080 149116 603132 149122
rect 603080 149058 603132 149064
rect 603078 148336 603134 148345
rect 603078 148271 603134 148280
rect 603092 147694 603120 148271
rect 603080 147688 603132 147694
rect 603080 147630 603132 147636
rect 603078 147384 603134 147393
rect 603078 147319 603134 147328
rect 603092 146334 603120 147319
rect 603736 146946 603764 161599
rect 603828 153202 603856 166631
rect 603816 153196 603868 153202
rect 603816 153138 603868 153144
rect 603906 149424 603962 149433
rect 603906 149359 603962 149368
rect 603724 146940 603776 146946
rect 603724 146882 603776 146888
rect 603080 146328 603132 146334
rect 603080 146270 603132 146276
rect 603170 146296 603226 146305
rect 603170 146231 603226 146240
rect 603184 144974 603212 146231
rect 603722 145344 603778 145353
rect 603722 145279 603778 145288
rect 603172 144968 603224 144974
rect 603172 144910 603224 144916
rect 603078 144256 603134 144265
rect 603078 144191 603134 144200
rect 603092 143614 603120 144191
rect 603080 143608 603132 143614
rect 603080 143550 603132 143556
rect 592684 143540 592736 143546
rect 592684 143482 592736 143488
rect 603078 142216 603134 142225
rect 591488 142180 591540 142186
rect 603078 142151 603080 142160
rect 591488 142122 591540 142128
rect 603132 142151 603134 142160
rect 603080 142122 603132 142128
rect 591396 124228 591448 124234
rect 591396 124170 591448 124176
rect 591304 124160 591356 124166
rect 591304 124102 591356 124108
rect 591304 121508 591356 121514
rect 591304 121450 591356 121456
rect 590108 110424 590160 110430
rect 590108 110366 590160 110372
rect 591316 85542 591344 121450
rect 591408 91050 591436 124170
rect 591500 122126 591528 142122
rect 603078 141264 603134 141273
rect 603078 141199 603134 141208
rect 603092 140826 603120 141199
rect 603080 140820 603132 140826
rect 603080 140762 603132 140768
rect 603078 140176 603134 140185
rect 603078 140111 603134 140120
rect 603092 139466 603120 140111
rect 594156 139460 594208 139466
rect 594156 139402 594208 139408
rect 603080 139460 603132 139466
rect 603080 139402 603132 139408
rect 592776 132524 592828 132530
rect 592776 132466 592828 132472
rect 592684 122868 592736 122874
rect 592684 122810 592736 122816
rect 591488 122120 591540 122126
rect 591488 122062 591540 122068
rect 591396 91044 591448 91050
rect 591396 90986 591448 90992
rect 592696 89690 592724 122810
rect 592788 102134 592816 132466
rect 594064 125724 594116 125730
rect 594064 125666 594116 125672
rect 592776 102128 592828 102134
rect 592776 102070 592828 102076
rect 594076 92478 594104 125666
rect 594168 113150 594196 139402
rect 603170 139224 603226 139233
rect 603170 139159 603226 139168
rect 603078 138136 603134 138145
rect 603078 138071 603080 138080
rect 603132 138071 603134 138080
rect 603080 138042 603132 138048
rect 603184 138038 603212 139159
rect 603172 138032 603224 138038
rect 603172 137974 603224 137980
rect 603078 137184 603134 137193
rect 603078 137119 603134 137128
rect 603092 136678 603120 137119
rect 603080 136672 603132 136678
rect 603080 136614 603132 136620
rect 603078 136096 603134 136105
rect 603078 136031 603134 136040
rect 603092 135318 603120 136031
rect 603080 135312 603132 135318
rect 603080 135254 603132 135260
rect 603170 135144 603226 135153
rect 603170 135079 603226 135088
rect 603078 134056 603134 134065
rect 603184 134026 603212 135079
rect 603078 133991 603134 134000
rect 603172 134020 603224 134026
rect 603092 133958 603120 133991
rect 603172 133962 603224 133968
rect 603080 133952 603132 133958
rect 603080 133894 603132 133900
rect 603736 133210 603764 145279
rect 603814 143304 603870 143313
rect 603814 143239 603870 143248
rect 603724 133204 603776 133210
rect 603724 133146 603776 133152
rect 603078 133104 603134 133113
rect 603078 133039 603134 133048
rect 603092 132530 603120 133039
rect 603080 132524 603132 132530
rect 603080 132466 603132 132472
rect 603078 132016 603134 132025
rect 603078 131951 603134 131960
rect 603092 131170 603120 131951
rect 603080 131164 603132 131170
rect 603080 131106 603132 131112
rect 603170 131064 603226 131073
rect 603170 130999 603226 131008
rect 603078 129976 603134 129985
rect 603078 129911 603134 129920
rect 603092 129810 603120 129911
rect 603184 129878 603212 130999
rect 603172 129872 603224 129878
rect 603172 129814 603224 129820
rect 603080 129804 603132 129810
rect 603080 129746 603132 129752
rect 603078 129024 603134 129033
rect 603078 128959 603134 128968
rect 603092 128382 603120 128959
rect 603080 128376 603132 128382
rect 603080 128318 603132 128324
rect 603078 127936 603134 127945
rect 603078 127871 603134 127880
rect 603092 127022 603120 127871
rect 603080 127016 603132 127022
rect 603080 126958 603132 126964
rect 603170 126984 603226 126993
rect 603170 126919 603226 126928
rect 603078 125896 603134 125905
rect 603078 125831 603134 125840
rect 603092 125730 603120 125831
rect 603080 125724 603132 125730
rect 603080 125666 603132 125672
rect 603184 125662 603212 126919
rect 603172 125656 603224 125662
rect 603172 125598 603224 125604
rect 603078 124944 603134 124953
rect 603078 124879 603134 124888
rect 603092 124234 603120 124879
rect 603080 124228 603132 124234
rect 603080 124170 603132 124176
rect 603078 123856 603134 123865
rect 603078 123791 603134 123800
rect 598204 122936 598256 122942
rect 598204 122878 598256 122884
rect 596824 114640 596876 114646
rect 596824 114582 596876 114588
rect 594156 113144 594208 113150
rect 594156 113086 594208 113092
rect 595444 111852 595496 111858
rect 595444 111794 595496 111800
rect 594064 92472 594116 92478
rect 594064 92414 594116 92420
rect 592684 89684 592736 89690
rect 592684 89626 592736 89632
rect 591304 85536 591356 85542
rect 591304 85478 591356 85484
rect 590016 84176 590068 84182
rect 590016 84118 590068 84124
rect 595456 71738 595484 111794
rect 596836 75886 596864 114582
rect 598216 86970 598244 122878
rect 603092 122874 603120 123791
rect 603172 122936 603224 122942
rect 603170 122904 603172 122913
rect 603224 122904 603226 122913
rect 603080 122868 603132 122874
rect 603170 122839 603226 122848
rect 603080 122810 603132 122816
rect 603078 121816 603134 121825
rect 603078 121751 603134 121760
rect 603092 121514 603120 121751
rect 603080 121508 603132 121514
rect 603080 121450 603132 121456
rect 603078 120864 603134 120873
rect 603078 120799 603134 120808
rect 603092 120154 603120 120799
rect 603080 120148 603132 120154
rect 603080 120090 603132 120096
rect 603078 119776 603134 119785
rect 603078 119711 603134 119720
rect 603092 118726 603120 119711
rect 603722 118824 603778 118833
rect 603722 118759 603778 118768
rect 603080 118720 603132 118726
rect 603080 118662 603132 118668
rect 603078 117736 603134 117745
rect 603078 117671 603134 117680
rect 603092 117366 603120 117671
rect 603080 117360 603132 117366
rect 603080 117302 603132 117308
rect 602342 116784 602398 116793
rect 602342 116719 602398 116728
rect 600964 99408 601016 99414
rect 600964 99350 601016 99356
rect 598204 86964 598256 86970
rect 598204 86906 598256 86912
rect 596824 75880 596876 75886
rect 596824 75822 596876 75828
rect 595444 71732 595496 71738
rect 595444 71674 595496 71680
rect 589924 69012 589976 69018
rect 589924 68954 589976 68960
rect 588636 67584 588688 67590
rect 588636 67526 588688 67532
rect 588544 64864 588596 64870
rect 588544 64806 588596 64812
rect 587164 63504 587216 63510
rect 587164 63446 587216 63452
rect 585784 62076 585836 62082
rect 585784 62018 585836 62024
rect 584404 60716 584456 60722
rect 584404 60658 584456 60664
rect 583024 58812 583076 58818
rect 583024 58754 583076 58760
rect 581644 57928 581696 57934
rect 581644 57870 581696 57876
rect 600976 57254 601004 99350
rect 602356 78674 602384 116719
rect 603078 115696 603134 115705
rect 603078 115631 603134 115640
rect 603092 114578 603120 115631
rect 603170 114744 603226 114753
rect 603170 114679 603226 114688
rect 603184 114646 603212 114679
rect 603172 114640 603224 114646
rect 603172 114582 603224 114588
rect 603080 114572 603132 114578
rect 603080 114514 603132 114520
rect 603078 113656 603134 113665
rect 603078 113591 603134 113600
rect 603092 113218 603120 113591
rect 603080 113212 603132 113218
rect 603080 113154 603132 113160
rect 603078 112704 603134 112713
rect 603078 112639 603134 112648
rect 603092 111858 603120 112639
rect 603080 111852 603132 111858
rect 603080 111794 603132 111800
rect 603078 110664 603134 110673
rect 603078 110599 603134 110608
rect 603092 110498 603120 110599
rect 603080 110492 603132 110498
rect 603080 110434 603132 110440
rect 603078 109576 603134 109585
rect 603078 109511 603134 109520
rect 603092 109070 603120 109511
rect 603080 109064 603132 109070
rect 603080 109006 603132 109012
rect 603078 108624 603134 108633
rect 603078 108559 603134 108568
rect 603092 107710 603120 108559
rect 603080 107704 603132 107710
rect 603080 107646 603132 107652
rect 603170 107536 603226 107545
rect 603170 107471 603226 107480
rect 603078 106584 603134 106593
rect 603078 106519 603134 106528
rect 603092 106350 603120 106519
rect 603184 106418 603212 107471
rect 603172 106412 603224 106418
rect 603172 106354 603224 106360
rect 603080 106344 603132 106350
rect 603080 106286 603132 106292
rect 603078 105496 603134 105505
rect 603078 105431 603134 105440
rect 603092 104922 603120 105431
rect 603080 104916 603132 104922
rect 603080 104858 603132 104864
rect 603078 104544 603134 104553
rect 603078 104479 603134 104488
rect 603092 103562 603120 104479
rect 603080 103556 603132 103562
rect 603080 103498 603132 103504
rect 603170 103456 603226 103465
rect 603170 103391 603226 103400
rect 603078 102504 603134 102513
rect 603078 102439 603134 102448
rect 603092 102202 603120 102439
rect 603184 102270 603212 103391
rect 603172 102264 603224 102270
rect 603172 102206 603224 102212
rect 603080 102196 603132 102202
rect 603080 102138 603132 102144
rect 603078 101416 603134 101425
rect 603078 101351 603134 101360
rect 603092 100774 603120 101351
rect 603080 100768 603132 100774
rect 603080 100710 603132 100716
rect 603446 100464 603502 100473
rect 603446 100399 603502 100408
rect 603460 99414 603488 100399
rect 603448 99408 603500 99414
rect 603448 99350 603500 99356
rect 603736 87650 603764 118759
rect 603828 117298 603856 143239
rect 603920 140078 603948 149359
rect 603908 140072 603960 140078
rect 603908 140014 603960 140020
rect 603816 117292 603868 117298
rect 603816 117234 603868 117240
rect 603814 111616 603870 111625
rect 603814 111551 603870 111560
rect 603724 87644 603776 87650
rect 603724 87586 603776 87592
rect 603828 82142 603856 111551
rect 603816 82136 603868 82142
rect 603816 82078 603868 82084
rect 602344 78668 602396 78674
rect 602344 78610 602396 78616
rect 605760 77994 605788 230454
rect 617156 220176 617208 220182
rect 617156 220118 617208 220124
rect 609612 220108 609664 220114
rect 609612 220050 609664 220056
rect 607680 218952 607732 218958
rect 607680 218894 607732 218900
rect 607128 217728 607180 217734
rect 607128 217670 607180 217676
rect 606668 213920 606720 213926
rect 606668 213862 606720 213868
rect 606680 210202 606708 213862
rect 607140 210202 607168 217670
rect 607692 213926 607720 218894
rect 608508 217864 608560 217870
rect 608508 217806 608560 217812
rect 608048 217796 608100 217802
rect 608048 217738 608100 217744
rect 607680 213920 607732 213926
rect 607680 213862 607732 213868
rect 607588 213172 607640 213178
rect 607588 213114 607640 213120
rect 607600 210202 607628 213114
rect 608060 210202 608088 217738
rect 608520 210202 608548 217806
rect 609624 217394 609652 220050
rect 614120 220040 614172 220046
rect 614120 219982 614172 219988
rect 611728 219972 611780 219978
rect 611728 219914 611780 219920
rect 609888 219836 609940 219842
rect 609888 219778 609940 219784
rect 609900 217666 609928 219778
rect 609888 217660 609940 217666
rect 609888 217602 609940 217608
rect 609612 217388 609664 217394
rect 609612 217330 609664 217336
rect 610808 217184 610860 217190
rect 610808 217126 610860 217132
rect 610348 217116 610400 217122
rect 610348 217058 610400 217064
rect 609888 217048 609940 217054
rect 609888 216990 609940 216996
rect 609428 216980 609480 216986
rect 609428 216922 609480 216928
rect 608968 216912 609020 216918
rect 608968 216854 609020 216860
rect 608980 210202 609008 216854
rect 609440 210202 609468 216922
rect 609900 210202 609928 216990
rect 610360 210202 610388 217058
rect 610820 210202 610848 217126
rect 611740 216102 611768 219914
rect 613016 219904 613068 219910
rect 613016 219846 613068 219852
rect 613028 216374 613056 219846
rect 613016 216368 613068 216374
rect 613016 216310 613068 216316
rect 614132 216306 614160 219982
rect 616788 218884 616840 218890
rect 616788 218826 616840 218832
rect 614120 216300 614172 216306
rect 614120 216242 614172 216248
rect 611728 216096 611780 216102
rect 611728 216038 611780 216044
rect 615500 215892 615552 215898
rect 615500 215834 615552 215840
rect 615040 215824 615092 215830
rect 615040 215766 615092 215772
rect 614580 215756 614632 215762
rect 614580 215698 614632 215704
rect 614028 215688 614080 215694
rect 614028 215630 614080 215636
rect 613568 215620 613620 215626
rect 613568 215562 613620 215568
rect 613108 215552 613160 215558
rect 613108 215494 613160 215500
rect 612648 215484 612700 215490
rect 612648 215426 612700 215432
rect 612188 215416 612240 215422
rect 612188 215358 612240 215364
rect 611728 215348 611780 215354
rect 611728 215290 611780 215296
rect 611268 213852 611320 213858
rect 611268 213794 611320 213800
rect 611280 210202 611308 213794
rect 611740 210202 611768 215290
rect 612200 210202 612228 215358
rect 612660 210202 612688 215426
rect 613120 210202 613148 215494
rect 613580 210202 613608 215562
rect 614040 210202 614068 215630
rect 614592 210202 614620 215698
rect 615052 210202 615080 215766
rect 615512 210202 615540 215834
rect 615960 213784 616012 213790
rect 615960 213726 616012 213732
rect 615972 210202 616000 213726
rect 616800 213722 616828 218826
rect 617168 215966 617196 220118
rect 619548 218816 619600 218822
rect 619548 218758 619600 218764
rect 618352 217592 618404 217598
rect 618352 217534 618404 217540
rect 617156 215960 617208 215966
rect 617156 215902 617208 215908
rect 617800 215892 617852 215898
rect 617800 215834 617852 215840
rect 616420 213716 616472 213722
rect 616420 213658 616472 213664
rect 616788 213716 616840 213722
rect 616788 213658 616840 213664
rect 616432 210202 616460 213658
rect 617340 213648 617392 213654
rect 617340 213590 617392 213596
rect 616880 213580 616932 213586
rect 616880 213522 616932 213528
rect 616892 210202 616920 213522
rect 617352 210202 617380 213590
rect 617812 210202 617840 215834
rect 618260 213512 618312 213518
rect 618260 213454 618312 213460
rect 618272 210202 618300 213454
rect 618364 212566 618392 217534
rect 618720 217524 618772 217530
rect 618720 217466 618772 217472
rect 618352 212560 618404 212566
rect 618352 212502 618404 212508
rect 618732 210202 618760 217466
rect 619560 213382 619588 218758
rect 619732 218408 619784 218414
rect 619732 218350 619784 218356
rect 619744 213858 619772 218350
rect 620926 216744 620982 216753
rect 620926 216679 620982 216688
rect 620560 216028 620612 216034
rect 620560 215970 620612 215976
rect 619732 213852 619784 213858
rect 619732 213794 619784 213800
rect 620100 213444 620152 213450
rect 620100 213386 620152 213392
rect 619180 213376 619232 213382
rect 619180 213318 619232 213324
rect 619548 213376 619600 213382
rect 619548 213318 619600 213324
rect 619192 210202 619220 213318
rect 619640 213308 619692 213314
rect 619640 213250 619692 213256
rect 619652 210202 619680 213250
rect 620112 210202 620140 213386
rect 620572 210202 620600 215970
rect 620940 212650 620968 216679
rect 621676 213314 621704 242898
rect 639604 232552 639656 232558
rect 639604 232494 639656 232500
rect 639144 232484 639196 232490
rect 639144 232426 639196 232432
rect 639052 231804 639104 231810
rect 639052 231746 639104 231752
rect 636844 230512 636896 230518
rect 636844 230454 636896 230460
rect 625344 219768 625396 219774
rect 625344 219710 625396 219716
rect 625252 219700 625304 219706
rect 625252 219642 625304 219648
rect 623872 219632 623924 219638
rect 623872 219574 623924 219580
rect 623044 219564 623096 219570
rect 623044 219506 623096 219512
rect 622952 219020 623004 219026
rect 622952 218962 623004 218968
rect 622030 216880 622086 216889
rect 622030 216815 622086 216824
rect 621664 213308 621716 213314
rect 621664 213250 621716 213256
rect 620940 212622 621152 212650
rect 621020 212560 621072 212566
rect 621020 212502 621072 212508
rect 621032 210202 621060 212502
rect 606648 210174 606708 210202
rect 607108 210174 607168 210202
rect 607568 210174 607628 210202
rect 608028 210174 608088 210202
rect 608488 210174 608548 210202
rect 608948 210174 609008 210202
rect 609408 210174 609468 210202
rect 609868 210174 609928 210202
rect 610328 210174 610388 210202
rect 610788 210174 610848 210202
rect 611248 210174 611308 210202
rect 611708 210174 611768 210202
rect 612168 210174 612228 210202
rect 612628 210174 612688 210202
rect 613088 210174 613148 210202
rect 613548 210174 613608 210202
rect 614008 210174 614068 210202
rect 614560 210174 614620 210202
rect 615020 210174 615080 210202
rect 615480 210174 615540 210202
rect 615940 210174 616000 210202
rect 616400 210174 616460 210202
rect 616860 210174 616920 210202
rect 617320 210174 617380 210202
rect 617780 210174 617840 210202
rect 618240 210174 618300 210202
rect 618700 210174 618760 210202
rect 619160 210174 619220 210202
rect 619620 210174 619680 210202
rect 620080 210174 620140 210202
rect 620540 210174 620600 210202
rect 621000 210174 621060 210202
rect 621124 210066 621152 212622
rect 622044 210202 622072 216815
rect 622492 213852 622544 213858
rect 622492 213794 622544 213800
rect 622504 210202 622532 213794
rect 622964 210202 622992 218962
rect 622012 210174 622072 210202
rect 622472 210174 622532 210202
rect 622932 210174 622992 210202
rect 623056 210066 623084 219506
rect 623780 219496 623832 219502
rect 623780 219438 623832 219444
rect 623792 210338 623820 219438
rect 623884 214538 623912 219574
rect 623962 219464 624018 219473
rect 623962 219399 624018 219408
rect 623872 214532 623924 214538
rect 623872 214474 623924 214480
rect 623792 210310 623912 210338
rect 623884 210202 623912 210310
rect 623852 210174 623912 210202
rect 623976 210066 624004 219399
rect 624424 214532 624476 214538
rect 624424 214474 624476 214480
rect 624436 210066 624464 214474
rect 625264 210202 625292 219642
rect 625232 210174 625292 210202
rect 625356 210066 625384 219710
rect 635924 219224 635976 219230
rect 635924 219166 635976 219172
rect 627460 218680 627512 218686
rect 627460 218622 627512 218628
rect 626632 216232 626684 216238
rect 626632 216174 626684 216180
rect 626172 214804 626224 214810
rect 626172 214746 626224 214752
rect 626184 210202 626212 214746
rect 626644 210202 626672 216174
rect 627092 214668 627144 214674
rect 627092 214610 627144 214616
rect 627104 210202 627132 214610
rect 627472 213450 627500 218622
rect 633716 218136 633768 218142
rect 633716 218078 633768 218084
rect 629484 217660 629536 217666
rect 629484 217602 629536 217608
rect 628930 217016 628986 217025
rect 628930 216951 628986 216960
rect 628472 216164 628524 216170
rect 628472 216106 628524 216112
rect 627552 214736 627604 214742
rect 627552 214678 627604 214684
rect 627460 213444 627512 213450
rect 627460 213386 627512 213392
rect 627564 210202 627592 214678
rect 628012 214600 628064 214606
rect 628012 214542 628064 214548
rect 628024 210202 628052 214542
rect 628484 210202 628512 216106
rect 628944 210202 628972 216951
rect 629496 210202 629524 217602
rect 632244 217456 632296 217462
rect 632244 217398 632296 217404
rect 631324 217320 631376 217326
rect 631324 217262 631376 217268
rect 629944 217252 629996 217258
rect 629944 217194 629996 217200
rect 629956 210202 629984 217194
rect 630404 216368 630456 216374
rect 630404 216310 630456 216316
rect 630416 210202 630444 216310
rect 630864 216096 630916 216102
rect 630864 216038 630916 216044
rect 630876 210202 630904 216038
rect 631336 210202 631364 217262
rect 631784 216300 631836 216306
rect 631784 216242 631836 216248
rect 631796 210202 631824 216242
rect 632256 210202 632284 217398
rect 632704 217388 632756 217394
rect 632704 217330 632756 217336
rect 632716 210202 632744 217330
rect 633728 213926 633756 218078
rect 634084 215960 634136 215966
rect 634084 215902 634136 215908
rect 633624 213920 633676 213926
rect 633624 213862 633676 213868
rect 633716 213920 633768 213926
rect 633716 213862 633768 213868
rect 633164 213240 633216 213246
rect 633164 213182 633216 213188
rect 633176 210202 633204 213182
rect 633636 210202 633664 213862
rect 634096 210202 634124 215902
rect 634544 213716 634596 213722
rect 634544 213658 634596 213664
rect 634556 210202 634584 213658
rect 635464 213444 635516 213450
rect 635464 213386 635516 213392
rect 635004 213376 635056 213382
rect 635004 213318 635056 213324
rect 635016 210202 635044 213318
rect 635476 210202 635504 213386
rect 635936 210202 635964 219166
rect 636856 213926 636884 230454
rect 637856 218340 637908 218346
rect 637856 218282 637908 218288
rect 637396 218272 637448 218278
rect 637396 218214 637448 218220
rect 636936 218204 636988 218210
rect 636936 218146 636988 218152
rect 636384 213920 636436 213926
rect 636384 213862 636436 213868
rect 636844 213920 636896 213926
rect 636844 213862 636896 213868
rect 636396 210202 636424 213862
rect 636948 210202 636976 218146
rect 637408 210202 637436 218214
rect 637868 210202 637896 218282
rect 638316 218068 638368 218074
rect 638316 218010 638368 218016
rect 638328 210202 638356 218010
rect 638776 211200 638828 211206
rect 638776 211142 638828 211148
rect 638788 210202 638816 211142
rect 626152 210174 626212 210202
rect 626612 210174 626672 210202
rect 627072 210174 627132 210202
rect 627532 210174 627592 210202
rect 627992 210174 628052 210202
rect 628452 210174 628512 210202
rect 628912 210174 628972 210202
rect 629464 210174 629524 210202
rect 629924 210174 629984 210202
rect 630384 210174 630444 210202
rect 630844 210174 630904 210202
rect 631304 210174 631364 210202
rect 631764 210174 631824 210202
rect 632224 210174 632284 210202
rect 632684 210174 632744 210202
rect 633144 210174 633204 210202
rect 633604 210174 633664 210202
rect 634064 210174 634124 210202
rect 634524 210174 634584 210202
rect 634984 210174 635044 210202
rect 635444 210174 635504 210202
rect 635904 210174 635964 210202
rect 636364 210174 636424 210202
rect 636916 210174 636976 210202
rect 637376 210174 637436 210202
rect 637836 210174 637896 210202
rect 638296 210174 638356 210202
rect 638756 210174 638816 210202
rect 639064 210118 639092 231746
rect 639156 229094 639184 232426
rect 639156 229066 639368 229094
rect 639236 213920 639288 213926
rect 639236 213862 639288 213868
rect 639248 210202 639276 213862
rect 639216 210174 639276 210202
rect 639052 210112 639104 210118
rect 621124 210038 621460 210066
rect 623056 210038 623392 210066
rect 623976 210038 624312 210066
rect 624436 210038 624772 210066
rect 625356 210038 625692 210066
rect 639052 210054 639104 210060
rect 639340 210066 639368 229066
rect 639616 213926 639644 232494
rect 646148 229673 646176 248386
rect 649356 231532 649408 231538
rect 649356 231474 649408 231480
rect 646134 229664 646190 229673
rect 646134 229599 646190 229608
rect 649368 229094 649396 231474
rect 649368 229066 649580 229094
rect 639604 213920 639656 213926
rect 639604 213862 639656 213868
rect 640616 213920 640668 213926
rect 640616 213862 640668 213868
rect 640628 210202 640656 213862
rect 641076 213308 641128 213314
rect 641076 213250 641128 213256
rect 643836 213308 643888 213314
rect 643836 213250 643888 213256
rect 641088 210202 641116 213250
rect 642732 213240 642784 213246
rect 642732 213182 642784 213188
rect 641824 210310 642128 210338
rect 641824 210202 641852 210310
rect 640596 210174 640656 210202
rect 641056 210174 641116 210202
rect 641516 210174 641852 210202
rect 639788 210112 639840 210118
rect 639340 210038 639676 210066
rect 642100 210066 642128 210310
rect 642744 210202 642772 213182
rect 643204 210310 643508 210338
rect 643204 210202 643232 210310
rect 642436 210188 642772 210202
rect 642422 210174 642772 210188
rect 642896 210174 643232 210202
rect 642422 210066 642450 210174
rect 639840 210060 640136 210066
rect 639788 210054 640136 210060
rect 639800 210038 640136 210054
rect 642100 210052 642450 210066
rect 643480 210066 643508 210310
rect 643848 210202 643876 213250
rect 645584 213172 645636 213178
rect 645584 213114 645636 213120
rect 644492 210310 644980 210338
rect 644492 210202 644520 210310
rect 643816 210188 643876 210202
rect 643802 210174 643876 210188
rect 644368 210174 644520 210202
rect 643802 210066 643830 210174
rect 643480 210052 643830 210066
rect 644952 210066 644980 210310
rect 645596 210202 645624 213114
rect 647146 213072 647202 213081
rect 646964 213036 647016 213042
rect 647146 213007 647202 213016
rect 648526 213072 648582 213081
rect 648526 213007 648582 213016
rect 646964 212978 647016 212984
rect 646056 210310 646360 210338
rect 646056 210202 646084 210310
rect 645288 210188 645624 210202
rect 645274 210174 645624 210188
rect 645748 210174 646084 210202
rect 645274 210066 645302 210174
rect 644952 210052 645302 210066
rect 646332 210066 646360 210310
rect 646976 210202 647004 212978
rect 647160 210202 647188 213007
rect 647436 210310 647740 210338
rect 647436 210202 647464 210310
rect 646668 210188 647004 210202
rect 646654 210174 647004 210188
rect 647128 210174 647464 210202
rect 646654 210066 646682 210174
rect 646332 210052 646682 210066
rect 647712 210066 647740 210310
rect 648540 210202 648568 213007
rect 648816 210310 649120 210338
rect 648816 210202 648844 210310
rect 648508 210174 648844 210202
rect 649092 210066 649120 210310
rect 649552 210066 649580 229066
rect 650012 213178 650040 984642
rect 650104 213246 650132 984778
rect 651472 984768 651524 984774
rect 651472 984710 651524 984716
rect 651380 984632 651432 984638
rect 651380 984574 651432 984580
rect 650644 231328 650696 231334
rect 650644 231270 650696 231276
rect 650656 229094 650684 231270
rect 650656 229066 650960 229094
rect 650092 213240 650144 213246
rect 650092 213182 650144 213188
rect 650000 213172 650052 213178
rect 650000 213114 650052 213120
rect 650196 210310 650500 210338
rect 650196 210066 650224 210310
rect 642100 210038 642436 210052
rect 643480 210038 643816 210052
rect 644952 210038 645288 210052
rect 646332 210038 646668 210052
rect 647712 210038 648048 210066
rect 649092 210038 649428 210066
rect 649552 210038 650224 210066
rect 650472 210066 650500 210310
rect 650932 210066 650960 229066
rect 651392 213042 651420 984574
rect 651484 213314 651512 984710
rect 651654 975896 651710 975905
rect 651654 975831 651710 975840
rect 651668 975730 651696 975831
rect 651656 975724 651708 975730
rect 651656 975666 651708 975672
rect 652022 962568 652078 962577
rect 652022 962503 652078 962512
rect 651562 949376 651618 949385
rect 651562 949311 651618 949320
rect 651576 948122 651604 949311
rect 651564 948116 651616 948122
rect 651564 948058 651616 948064
rect 652036 939826 652064 962503
rect 652024 939820 652076 939826
rect 652024 939762 652076 939768
rect 658936 937242 658964 990218
rect 659016 957840 659068 957846
rect 659016 957782 659068 957788
rect 658924 937236 658976 937242
rect 658924 937178 658976 937184
rect 659028 937038 659056 957782
rect 651564 937032 651616 937038
rect 651564 936974 651616 936980
rect 659016 937032 659068 937038
rect 659016 936974 659068 936980
rect 651576 936193 651604 936974
rect 651562 936184 651618 936193
rect 651562 936119 651618 936128
rect 660316 935678 660344 991510
rect 661696 937378 661724 992938
rect 666744 992928 666796 992934
rect 666744 992870 666796 992876
rect 666560 991500 666612 991506
rect 666560 991442 666612 991448
rect 665456 984904 665508 984910
rect 665456 984846 665508 984852
rect 661684 937372 661736 937378
rect 661684 937314 661736 937320
rect 660304 935672 660356 935678
rect 660304 935614 660356 935620
rect 651562 922720 651618 922729
rect 651562 922655 651618 922664
rect 651576 921874 651604 922655
rect 651564 921868 651616 921874
rect 651564 921810 651616 921816
rect 664444 921868 664496 921874
rect 664444 921810 664496 921816
rect 651562 909528 651618 909537
rect 651562 909463 651564 909472
rect 651616 909463 651618 909472
rect 661684 909492 661736 909498
rect 651564 909434 651616 909440
rect 661684 909434 661736 909440
rect 651562 896200 651618 896209
rect 651562 896135 651618 896144
rect 651576 895694 651604 896135
rect 651564 895688 651616 895694
rect 651564 895630 651616 895636
rect 660304 895688 660356 895694
rect 660304 895630 660356 895636
rect 652022 882872 652078 882881
rect 652022 882807 652078 882816
rect 651562 869680 651618 869689
rect 651562 869615 651618 869624
rect 651576 869446 651604 869615
rect 651564 869440 651616 869446
rect 651564 869382 651616 869388
rect 652036 868698 652064 882807
rect 652024 868692 652076 868698
rect 652024 868634 652076 868640
rect 652574 856352 652630 856361
rect 652574 856287 652630 856296
rect 652588 855642 652616 856287
rect 652576 855636 652628 855642
rect 652576 855578 652628 855584
rect 651562 843024 651618 843033
rect 651562 842959 651618 842968
rect 651576 841838 651604 842959
rect 651564 841832 651616 841838
rect 651564 841774 651616 841780
rect 651562 829832 651618 829841
rect 651562 829767 651618 829776
rect 651576 829462 651604 829767
rect 651564 829456 651616 829462
rect 651564 829398 651616 829404
rect 659016 829456 659068 829462
rect 659016 829398 659068 829404
rect 651562 816504 651618 816513
rect 651562 816439 651618 816448
rect 651576 815658 651604 816439
rect 651564 815652 651616 815658
rect 651564 815594 651616 815600
rect 651562 803312 651618 803321
rect 651562 803247 651618 803256
rect 651576 803214 651604 803247
rect 651564 803208 651616 803214
rect 651564 803150 651616 803156
rect 658924 803208 658976 803214
rect 658924 803150 658976 803156
rect 651654 789984 651710 789993
rect 651654 789919 651710 789928
rect 651668 789410 651696 789919
rect 651656 789404 651708 789410
rect 651656 789346 651708 789352
rect 651562 776656 651618 776665
rect 651562 776591 651618 776600
rect 651576 775606 651604 776591
rect 651564 775600 651616 775606
rect 651564 775542 651616 775548
rect 651562 763328 651618 763337
rect 651562 763263 651618 763272
rect 651576 763230 651604 763263
rect 651564 763224 651616 763230
rect 651564 763166 651616 763172
rect 651562 750136 651618 750145
rect 651562 750071 651618 750080
rect 651576 749426 651604 750071
rect 651564 749420 651616 749426
rect 651564 749362 651616 749368
rect 651562 736808 651618 736817
rect 651562 736743 651618 736752
rect 651576 735622 651604 736743
rect 651564 735616 651616 735622
rect 651564 735558 651616 735564
rect 652022 723480 652078 723489
rect 652022 723415 652078 723424
rect 652036 723178 652064 723415
rect 652024 723172 652076 723178
rect 652024 723114 652076 723120
rect 651562 710288 651618 710297
rect 651562 710223 651618 710232
rect 651576 709374 651604 710223
rect 651564 709368 651616 709374
rect 651564 709310 651616 709316
rect 652022 696960 652078 696969
rect 652022 696895 652078 696904
rect 651838 683632 651894 683641
rect 651838 683567 651894 683576
rect 651852 683194 651880 683567
rect 651840 683188 651892 683194
rect 651840 683130 651892 683136
rect 651562 670440 651618 670449
rect 651562 670375 651618 670384
rect 651576 669390 651604 670375
rect 651564 669384 651616 669390
rect 651564 669326 651616 669332
rect 651562 657112 651618 657121
rect 651562 657047 651618 657056
rect 651576 656946 651604 657047
rect 651564 656940 651616 656946
rect 651564 656882 651616 656888
rect 651562 643784 651618 643793
rect 651562 643719 651618 643728
rect 651576 643142 651604 643719
rect 651564 643136 651616 643142
rect 651564 643078 651616 643084
rect 651562 630592 651618 630601
rect 651562 630527 651618 630536
rect 651576 629338 651604 630527
rect 651564 629332 651616 629338
rect 651564 629274 651616 629280
rect 651562 603936 651618 603945
rect 651562 603871 651618 603880
rect 651576 603158 651604 603871
rect 651564 603152 651616 603158
rect 651564 603094 651616 603100
rect 651562 590744 651618 590753
rect 651562 590679 651564 590688
rect 651616 590679 651618 590688
rect 651564 590650 651616 590656
rect 652036 581058 652064 696895
rect 658936 670818 658964 803150
rect 659028 779006 659056 829398
rect 659016 779000 659068 779006
rect 659016 778942 659068 778948
rect 659016 775600 659068 775606
rect 659016 775542 659068 775548
rect 659028 734874 659056 775542
rect 660316 760578 660344 895630
rect 661696 760714 661724 909434
rect 663064 841832 663116 841838
rect 663064 841774 663116 841780
rect 661776 789404 661828 789410
rect 661776 789346 661828 789352
rect 661684 760708 661736 760714
rect 661684 760650 661736 760656
rect 660304 760572 660356 760578
rect 660304 760514 660356 760520
rect 660304 735616 660356 735622
rect 660304 735558 660356 735564
rect 659016 734868 659068 734874
rect 659016 734810 659068 734816
rect 659016 683188 659068 683194
rect 659016 683130 659068 683136
rect 658924 670812 658976 670818
rect 658924 670754 658976 670760
rect 658924 669384 658976 669390
rect 658924 669326 658976 669332
rect 658936 643754 658964 669326
rect 658924 643748 658976 643754
rect 658924 643690 658976 643696
rect 652390 617264 652446 617273
rect 652390 617199 652446 617208
rect 652404 616894 652432 617199
rect 652392 616888 652444 616894
rect 652392 616830 652444 616836
rect 658924 616888 658976 616894
rect 658924 616830 658976 616836
rect 658936 599622 658964 616830
rect 658924 599616 658976 599622
rect 658924 599558 658976 599564
rect 652024 581052 652076 581058
rect 652024 580994 652076 581000
rect 659028 579834 659056 683130
rect 660316 625190 660344 735558
rect 661788 669458 661816 789346
rect 663076 715018 663104 841774
rect 664456 760850 664484 921810
rect 664536 763224 664588 763230
rect 664536 763166 664588 763172
rect 664444 760844 664496 760850
rect 664444 760786 664496 760792
rect 663064 715012 663116 715018
rect 663064 714954 663116 714960
rect 661776 669452 661828 669458
rect 661776 669394 661828 669400
rect 663064 656940 663116 656946
rect 663064 656882 663116 656888
rect 661684 629332 661736 629338
rect 661684 629274 661736 629280
rect 660304 625184 660356 625190
rect 660304 625126 660356 625132
rect 660304 603152 660356 603158
rect 660304 603094 660356 603100
rect 659016 579828 659068 579834
rect 659016 579770 659068 579776
rect 651562 577416 651618 577425
rect 651562 577351 651618 577360
rect 651576 576910 651604 577351
rect 651564 576904 651616 576910
rect 651564 576846 651616 576852
rect 659016 576904 659068 576910
rect 659016 576846 659068 576852
rect 652114 564088 652170 564097
rect 652114 564023 652170 564032
rect 652128 563106 652156 564023
rect 652116 563100 652168 563106
rect 652116 563042 652168 563048
rect 658924 563100 658976 563106
rect 658924 563042 658976 563048
rect 658936 554062 658964 563042
rect 658924 554056 658976 554062
rect 658924 553998 658976 554004
rect 651562 550896 651618 550905
rect 651562 550831 651618 550840
rect 651576 550662 651604 550831
rect 651564 550656 651616 550662
rect 651564 550598 651616 550604
rect 651562 537568 651618 537577
rect 651562 537503 651618 537512
rect 651576 536858 651604 537503
rect 651564 536852 651616 536858
rect 651564 536794 651616 536800
rect 651562 524240 651618 524249
rect 651562 524175 651618 524184
rect 651576 523054 651604 524175
rect 651564 523048 651616 523054
rect 651564 522990 651616 522996
rect 651562 511048 651618 511057
rect 651562 510983 651618 510992
rect 651576 510678 651604 510983
rect 651564 510672 651616 510678
rect 651564 510614 651616 510620
rect 651562 497720 651618 497729
rect 651562 497655 651618 497664
rect 651576 496874 651604 497655
rect 651564 496868 651616 496874
rect 651564 496810 651616 496816
rect 658924 496868 658976 496874
rect 658924 496810 658976 496816
rect 651562 484528 651618 484537
rect 651562 484463 651618 484472
rect 651576 484430 651604 484463
rect 651564 484424 651616 484430
rect 651564 484366 651616 484372
rect 651654 471200 651710 471209
rect 651654 471135 651710 471144
rect 651668 470626 651696 471135
rect 651656 470620 651708 470626
rect 651656 470562 651708 470568
rect 651562 457872 651618 457881
rect 651562 457807 651618 457816
rect 651576 456822 651604 457807
rect 651564 456816 651616 456822
rect 651564 456758 651616 456764
rect 651562 444544 651618 444553
rect 651562 444479 651618 444488
rect 651576 444446 651604 444479
rect 651564 444440 651616 444446
rect 651564 444382 651616 444388
rect 651562 431352 651618 431361
rect 651562 431287 651618 431296
rect 651576 430642 651604 431287
rect 651564 430636 651616 430642
rect 651564 430578 651616 430584
rect 651562 418024 651618 418033
rect 651562 417959 651618 417968
rect 651576 416838 651604 417959
rect 651564 416832 651616 416838
rect 651564 416774 651616 416780
rect 652022 404696 652078 404705
rect 652022 404631 652078 404640
rect 652036 404394 652064 404631
rect 652024 404388 652076 404394
rect 652024 404330 652076 404336
rect 651562 391504 651618 391513
rect 651562 391439 651618 391448
rect 651576 390590 651604 391439
rect 651564 390584 651616 390590
rect 651564 390526 651616 390532
rect 651564 378208 651616 378214
rect 651562 378176 651564 378185
rect 651616 378176 651618 378185
rect 651562 378111 651618 378120
rect 652022 364848 652078 364857
rect 652022 364783 652078 364792
rect 652036 364410 652064 364783
rect 652024 364404 652076 364410
rect 652024 364346 652076 364352
rect 658936 357610 658964 496810
rect 659028 491434 659056 576846
rect 660316 491570 660344 603094
rect 660396 536852 660448 536858
rect 660396 536794 660448 536800
rect 660304 491564 660356 491570
rect 660304 491506 660356 491512
rect 659016 491428 659068 491434
rect 659016 491370 659068 491376
rect 659016 444440 659068 444446
rect 659016 444382 659068 444388
rect 658924 357604 658976 357610
rect 658924 357546 658976 357552
rect 651562 351656 651618 351665
rect 651562 351591 651618 351600
rect 651576 350606 651604 351591
rect 651564 350600 651616 350606
rect 651564 350542 651616 350548
rect 651654 338328 651710 338337
rect 651654 338263 651710 338272
rect 651668 338162 651696 338263
rect 651656 338156 651708 338162
rect 651656 338098 651708 338104
rect 651562 325000 651618 325009
rect 651562 324935 651618 324944
rect 651576 324358 651604 324935
rect 651564 324352 651616 324358
rect 651564 324294 651616 324300
rect 659028 312050 659056 444382
rect 660304 430636 660356 430642
rect 660304 430578 660356 430584
rect 659016 312044 659068 312050
rect 659016 311986 659068 311992
rect 651562 311808 651618 311817
rect 651562 311743 651618 311752
rect 651576 310622 651604 311743
rect 651564 310616 651616 310622
rect 651564 310558 651616 310564
rect 652022 298480 652078 298489
rect 652022 298415 652078 298424
rect 651562 285288 651618 285297
rect 651562 285223 651618 285232
rect 651576 284374 651604 285223
rect 651564 284368 651616 284374
rect 651564 284310 651616 284316
rect 651472 213308 651524 213314
rect 651472 213250 651524 213256
rect 651380 213036 651432 213042
rect 651380 212978 651432 212984
rect 652036 210458 652064 298415
rect 656900 278180 656952 278186
rect 656900 278122 656952 278128
rect 654140 231396 654192 231402
rect 654140 231338 654192 231344
rect 652760 231260 652812 231266
rect 652760 231202 652812 231208
rect 652024 210452 652076 210458
rect 652024 210394 652076 210400
rect 651668 210310 651972 210338
rect 651668 210066 651696 210310
rect 650472 210038 650808 210066
rect 650932 210038 651696 210066
rect 651944 210066 651972 210310
rect 652772 210202 652800 231202
rect 653048 210310 653352 210338
rect 653048 210202 653076 210310
rect 652740 210174 653076 210202
rect 653324 210066 653352 210310
rect 654152 210202 654180 231338
rect 655520 231192 655572 231198
rect 655520 231134 655572 231140
rect 654428 210310 654732 210338
rect 654428 210202 654456 210310
rect 654120 210174 654456 210202
rect 654704 210066 654732 210310
rect 655532 210202 655560 231134
rect 655808 210310 656112 210338
rect 655808 210202 655836 210310
rect 655500 210174 655836 210202
rect 656084 210066 656112 210310
rect 656912 210202 656940 278122
rect 658280 278044 658332 278050
rect 658280 277986 658332 277992
rect 657188 210310 657492 210338
rect 657188 210202 657216 210310
rect 656880 210174 657216 210202
rect 657464 210066 657492 210310
rect 658292 210202 658320 277986
rect 660316 267782 660344 430578
rect 660408 403170 660436 536794
rect 661696 534274 661724 629274
rect 661776 550656 661828 550662
rect 661776 550598 661828 550604
rect 661684 534268 661736 534274
rect 661684 534210 661736 534216
rect 661684 510672 661736 510678
rect 661684 510614 661736 510620
rect 660488 484424 660540 484430
rect 660488 484366 660540 484372
rect 660396 403164 660448 403170
rect 660396 403106 660448 403112
rect 660396 364404 660448 364410
rect 660396 364346 660448 364352
rect 660304 267776 660356 267782
rect 660304 267718 660356 267724
rect 660408 222222 660436 364346
rect 660500 357746 660528 484366
rect 661696 357882 661724 510614
rect 661788 403306 661816 550598
rect 663076 535634 663104 656882
rect 664548 625394 664576 763166
rect 664536 625388 664588 625394
rect 664536 625330 664588 625336
rect 664444 590708 664496 590714
rect 664444 590650 664496 590656
rect 663064 535628 663116 535634
rect 663064 535570 663116 535576
rect 663248 523048 663300 523054
rect 663248 522990 663300 522996
rect 663156 456816 663208 456822
rect 663156 456758 663208 456764
rect 663064 416832 663116 416838
rect 663064 416774 663116 416780
rect 661868 404388 661920 404394
rect 661868 404330 661920 404336
rect 661776 403300 661828 403306
rect 661776 403242 661828 403248
rect 661684 357876 661736 357882
rect 661684 357818 661736 357824
rect 660488 357740 660540 357746
rect 660488 357682 660540 357688
rect 661880 267986 661908 404330
rect 662420 278112 662472 278118
rect 662420 278054 662472 278060
rect 661868 267980 661920 267986
rect 661868 267922 661920 267928
rect 661040 231464 661092 231470
rect 661040 231406 661092 231412
rect 661052 229094 661080 231406
rect 661052 229066 661172 229094
rect 660396 222216 660448 222222
rect 660396 222158 660448 222164
rect 659752 218748 659804 218754
rect 659752 218690 659804 218696
rect 658568 210310 658872 210338
rect 658568 210202 658596 210310
rect 658260 210174 658596 210202
rect 658844 210066 658872 210310
rect 659764 210202 659792 218690
rect 660040 210310 660344 210338
rect 660040 210202 660068 210310
rect 659732 210174 660068 210202
rect 660316 210066 660344 210310
rect 661144 210202 661172 229066
rect 662432 210338 662460 278054
rect 663076 268122 663104 416774
rect 663168 313410 663196 456758
rect 663260 403442 663288 522990
rect 664456 491706 664484 590650
rect 664444 491700 664496 491706
rect 664444 491642 664496 491648
rect 664536 470620 664588 470626
rect 664536 470562 664588 470568
rect 663248 403436 663300 403442
rect 663248 403378 663300 403384
rect 664444 390584 664496 390590
rect 664444 390526 664496 390532
rect 663156 313404 663208 313410
rect 663156 313346 663208 313352
rect 663064 268116 663116 268122
rect 663064 268058 663116 268064
rect 662512 264240 662564 264246
rect 662512 264182 662564 264188
rect 662524 214606 662552 264182
rect 663800 231668 663852 231674
rect 663800 231610 663852 231616
rect 662604 231124 662656 231130
rect 662604 231066 662656 231072
rect 662512 214600 662564 214606
rect 662512 214542 662564 214548
rect 661420 210310 661724 210338
rect 662432 210310 662552 210338
rect 661420 210202 661448 210310
rect 661112 210174 661448 210202
rect 661696 210066 661724 210310
rect 662524 210202 662552 210310
rect 662492 210174 662552 210202
rect 662616 210066 662644 231066
rect 663812 214606 663840 231610
rect 663892 231600 663944 231606
rect 663892 231542 663944 231548
rect 663904 229094 663932 231542
rect 663904 229066 664024 229094
rect 663890 218648 663946 218657
rect 663890 218583 663946 218592
rect 663064 214600 663116 214606
rect 663064 214542 663116 214548
rect 663800 214600 663852 214606
rect 663800 214542 663852 214548
rect 663076 210066 663104 214542
rect 663904 210202 663932 218583
rect 663872 210174 663932 210202
rect 663996 210066 664024 229066
rect 664456 222426 664484 390526
rect 664548 313546 664576 470562
rect 664536 313540 664588 313546
rect 664536 313482 664588 313488
rect 664444 222420 664496 222426
rect 664444 222362 664496 222368
rect 664444 214600 664496 214606
rect 664444 214542 664496 214548
rect 664456 210066 664484 214542
rect 665272 214396 665324 214402
rect 665272 214338 665324 214344
rect 665284 210202 665312 214338
rect 665252 210174 665312 210202
rect 651944 210038 652280 210066
rect 653324 210038 653660 210066
rect 654704 210038 655040 210066
rect 656084 210038 656420 210066
rect 657464 210038 657800 210066
rect 658844 210038 659272 210066
rect 660316 210038 660652 210066
rect 661696 210038 662032 210066
rect 662616 210038 662952 210066
rect 663076 210038 663412 210066
rect 663996 210038 664332 210066
rect 664456 210038 664792 210066
rect 665468 209817 665496 984846
rect 665824 815652 665876 815658
rect 665824 815594 665876 815600
rect 665836 670954 665864 815594
rect 665824 670948 665876 670954
rect 665824 670890 665876 670896
rect 665824 378208 665876 378214
rect 665824 378150 665876 378156
rect 665836 222562 665864 378150
rect 665824 222556 665876 222562
rect 665824 222498 665876 222504
rect 665732 214124 665784 214130
rect 665732 214066 665784 214072
rect 665744 210202 665772 214066
rect 666192 214056 666244 214062
rect 666192 213998 666244 214004
rect 666204 210202 666232 213998
rect 665712 210174 665772 210202
rect 666172 210174 666232 210202
rect 665454 209808 665510 209817
rect 665454 209743 665510 209752
rect 666572 194041 666600 991442
rect 666652 984972 666704 984978
rect 666652 984914 666704 984920
rect 666558 194032 666614 194041
rect 666558 193967 666614 193976
rect 666572 190641 666600 193967
rect 666558 190632 666614 190641
rect 666558 190567 666614 190576
rect 666664 190454 666692 984914
rect 666756 199073 666784 992870
rect 669964 990208 670016 990214
rect 669964 990150 670016 990156
rect 666836 990140 666888 990146
rect 666836 990082 666888 990088
rect 666848 204241 666876 990082
rect 669976 938602 670004 990150
rect 671344 975724 671396 975730
rect 671344 975666 671396 975672
rect 671356 938738 671384 975666
rect 675772 966521 675800 966723
rect 675758 966512 675814 966521
rect 675758 966447 675814 966456
rect 675758 966240 675814 966249
rect 675758 966175 675814 966184
rect 675772 966076 675800 966175
rect 675772 965025 675800 965435
rect 675758 965016 675814 965025
rect 675758 964951 675814 964960
rect 675404 963393 675432 963595
rect 675390 963384 675446 963393
rect 675390 963319 675446 963328
rect 675496 962742 675524 963016
rect 674840 962736 674892 962742
rect 674840 962678 674892 962684
rect 675484 962736 675536 962742
rect 675484 962678 675536 962684
rect 674746 959032 674802 959041
rect 674852 959018 674880 962678
rect 675404 962062 675432 962404
rect 675024 962056 675076 962062
rect 675024 961998 675076 962004
rect 675392 962056 675444 962062
rect 675392 961998 675444 962004
rect 674802 958990 674880 959018
rect 674746 958967 674802 958976
rect 673276 958384 673328 958390
rect 673276 958326 673328 958332
rect 672356 956548 672408 956554
rect 672356 956490 672408 956496
rect 671344 938732 671396 938738
rect 671344 938674 671396 938680
rect 669964 938596 670016 938602
rect 669964 938538 670016 938544
rect 669964 927444 670016 927450
rect 669964 927386 670016 927392
rect 668584 749420 668636 749426
rect 668584 749362 668636 749368
rect 668596 625530 668624 749362
rect 668676 723172 668728 723178
rect 668676 723114 668728 723120
rect 668688 688702 668716 723114
rect 668676 688696 668728 688702
rect 668676 688638 668728 688644
rect 668676 643136 668728 643142
rect 668676 643078 668728 643084
rect 668584 625524 668636 625530
rect 668584 625466 668636 625472
rect 668688 535770 668716 643078
rect 668676 535764 668728 535770
rect 668676 535706 668728 535712
rect 668584 475856 668636 475862
rect 668584 475798 668636 475804
rect 668124 214260 668176 214266
rect 668124 214202 668176 214208
rect 667204 210452 667256 210458
rect 667204 210394 667256 210400
rect 666834 204232 666890 204241
rect 666834 204167 666890 204176
rect 666848 200841 666876 204167
rect 666834 200832 666890 200841
rect 666834 200767 666890 200776
rect 666742 199064 666798 199073
rect 666742 198999 666798 199008
rect 666572 190426 666692 190454
rect 666572 189009 666600 190426
rect 666558 189000 666614 189009
rect 666558 188935 666614 188944
rect 666572 185609 666600 188935
rect 666558 185600 666614 185609
rect 666558 185535 666614 185544
rect 666558 153368 666614 153377
rect 666558 153303 666614 153312
rect 666572 151881 666600 153303
rect 666558 151872 666614 151881
rect 666558 151807 666614 151816
rect 666558 151600 666614 151609
rect 666558 151535 666614 151544
rect 666572 149977 666600 151535
rect 666558 149968 666614 149977
rect 666558 149903 666614 149912
rect 666558 142080 666614 142089
rect 666558 142015 666614 142024
rect 666572 139777 666600 142015
rect 666558 139768 666614 139777
rect 666558 139703 666614 139712
rect 667216 132666 667244 210394
rect 667938 209264 667994 209273
rect 667938 209199 667994 209208
rect 667952 205873 667980 209199
rect 667938 205864 667994 205873
rect 667938 205799 667994 205808
rect 667938 199064 667994 199073
rect 667938 198999 667994 199008
rect 667952 195673 667980 198999
rect 667938 195664 667994 195673
rect 667938 195599 667994 195608
rect 667940 183932 667992 183938
rect 667940 183874 667992 183880
rect 667952 183841 667980 183874
rect 667938 183832 667994 183841
rect 667938 183767 667994 183776
rect 667952 180794 667980 183767
rect 667952 180766 668072 180794
rect 668044 180441 668072 180766
rect 668030 180432 668086 180441
rect 668030 180367 668086 180376
rect 667940 178832 667992 178838
rect 667938 178800 667940 178809
rect 667992 178800 667994 178809
rect 667938 178735 667994 178744
rect 667952 175409 667980 178735
rect 667938 175400 667994 175409
rect 667938 175335 667994 175344
rect 667938 173632 667994 173641
rect 667938 173567 667994 173576
rect 667952 171193 667980 173567
rect 667938 171184 667994 171193
rect 667938 171119 667994 171128
rect 667940 163872 667992 163878
rect 667940 163814 667992 163820
rect 667952 163577 667980 163814
rect 667938 163568 667994 163577
rect 667938 163503 667994 163512
rect 667952 161537 667980 163503
rect 667938 161528 667994 161537
rect 667938 161463 667994 161472
rect 667938 158400 667994 158409
rect 667938 158335 667994 158344
rect 667952 155009 667980 158335
rect 667938 155000 667994 155009
rect 667938 154935 667994 154944
rect 667940 143472 667992 143478
rect 667940 143414 667992 143420
rect 667952 143177 667980 143414
rect 667938 143168 667994 143177
rect 667938 143103 667994 143112
rect 667940 138236 667992 138242
rect 667940 138178 667992 138184
rect 667952 138145 667980 138178
rect 667938 138136 667994 138145
rect 667938 138071 667994 138080
rect 667952 134745 667980 138071
rect 667938 134736 667994 134745
rect 667938 134671 667994 134680
rect 667204 132660 667256 132666
rect 667204 132602 667256 132608
rect 666558 132424 666614 132433
rect 666558 132359 666614 132368
rect 666572 129577 666600 132359
rect 666558 129568 666614 129577
rect 666558 129503 666614 129512
rect 667940 127968 667992 127974
rect 667938 127936 667940 127945
rect 667992 127936 667994 127945
rect 667938 127871 667994 127880
rect 667952 124545 667980 127871
rect 667938 124536 667994 124545
rect 667938 124471 667994 124480
rect 667940 124092 667992 124098
rect 667940 124034 667992 124040
rect 667952 122913 667980 124034
rect 667938 122904 667994 122913
rect 667938 122839 667994 122848
rect 666558 122768 666614 122777
rect 666558 122703 666614 122712
rect 666572 119513 666600 122703
rect 666558 119504 666614 119513
rect 666558 119439 666614 119448
rect 667940 117768 667992 117774
rect 667938 117736 667940 117745
rect 667992 117736 667994 117745
rect 667938 117671 667994 117680
rect 667940 109336 667992 109342
rect 667938 109304 667940 109313
rect 667992 109304 667994 109313
rect 667938 109239 667994 109248
rect 668136 107545 668164 214202
rect 668308 173800 668360 173806
rect 668308 173742 668360 173748
rect 668320 173641 668348 173742
rect 668306 173632 668362 173641
rect 668306 173567 668362 173576
rect 668308 168700 668360 168706
rect 668308 168642 668360 168648
rect 668320 168609 668348 168642
rect 668306 168600 668362 168609
rect 668306 168535 668362 168544
rect 668320 165209 668348 168535
rect 668306 165200 668362 165209
rect 668306 165135 668362 165144
rect 668596 153377 668624 475798
rect 668676 474564 668728 474570
rect 668676 474506 668728 474512
rect 668688 158409 668716 474506
rect 668768 338156 668820 338162
rect 668768 338098 668820 338104
rect 668780 178226 668808 338098
rect 668860 214328 668912 214334
rect 668860 214270 668912 214276
rect 668768 178220 668820 178226
rect 668768 178162 668820 178168
rect 668674 158400 668730 158409
rect 668674 158335 668730 158344
rect 668582 153368 668638 153377
rect 668582 153303 668638 153312
rect 668308 148436 668360 148442
rect 668308 148378 668360 148384
rect 668320 148209 668348 148378
rect 668306 148200 668362 148209
rect 668306 148135 668362 148144
rect 668320 144945 668348 148135
rect 668306 144936 668362 144945
rect 668306 144871 668362 144880
rect 668584 133000 668636 133006
rect 668582 132968 668584 132977
rect 668636 132968 668638 132977
rect 668582 132903 668638 132912
rect 668872 132494 668900 214270
rect 668952 214192 669004 214198
rect 668952 214134 669004 214140
rect 668780 132466 668900 132494
rect 668676 131164 668728 131170
rect 668676 131106 668728 131112
rect 668584 129804 668636 129810
rect 668584 129746 668636 129752
rect 668400 117020 668452 117026
rect 668400 116962 668452 116968
rect 668412 116113 668440 116962
rect 668398 116104 668454 116113
rect 668398 116039 668454 116048
rect 668308 111784 668360 111790
rect 668308 111726 668360 111732
rect 668320 110945 668348 111726
rect 668306 110936 668362 110945
rect 668306 110871 668362 110880
rect 668122 107536 668178 107545
rect 668122 107471 668178 107480
rect 668596 100881 668624 129746
rect 668688 104145 668716 131106
rect 668780 128382 668808 132466
rect 668964 129810 668992 214134
rect 669044 213988 669096 213994
rect 669044 213930 669096 213936
rect 669056 131170 669084 213930
rect 669976 183938 670004 927386
rect 671988 879096 672040 879102
rect 671988 879038 672040 879044
rect 671344 869440 671396 869446
rect 671344 869382 671396 869388
rect 670516 775600 670568 775606
rect 670516 775542 670568 775548
rect 670056 749420 670108 749426
rect 670056 749362 670108 749368
rect 669964 183932 670016 183938
rect 669964 183874 670016 183880
rect 670068 178838 670096 749362
rect 670528 711686 670556 775542
rect 670608 743844 670660 743850
rect 670608 743786 670660 743792
rect 670516 711680 670568 711686
rect 670516 711622 670568 711628
rect 670620 665378 670648 743786
rect 671356 716174 671384 869382
rect 671896 780768 671948 780774
rect 671896 780710 671948 780716
rect 671804 730516 671856 730522
rect 671804 730458 671856 730464
rect 671344 716168 671396 716174
rect 671344 716110 671396 716116
rect 671436 709368 671488 709374
rect 671436 709310 671488 709316
rect 670608 665372 670660 665378
rect 670608 665314 670660 665320
rect 670516 640348 670568 640354
rect 670516 640290 670568 640296
rect 670528 575618 670556 640290
rect 671344 614168 671396 614174
rect 671344 614110 671396 614116
rect 670608 608048 670660 608054
rect 670608 607990 670660 607996
rect 670516 575612 670568 575618
rect 670516 575554 670568 575560
rect 670620 530058 670648 607990
rect 670608 530052 670660 530058
rect 670608 529994 670660 530000
rect 670148 392012 670200 392018
rect 670148 391954 670200 391960
rect 670056 178832 670108 178838
rect 670056 178774 670108 178780
rect 669964 168292 670016 168298
rect 669964 168234 670016 168240
rect 669044 131164 669096 131170
rect 669044 131106 669096 131112
rect 668952 129804 669004 129810
rect 668952 129746 669004 129752
rect 668768 128376 668820 128382
rect 668768 128318 668820 128324
rect 668674 104136 668730 104145
rect 668674 104071 668730 104080
rect 668780 102513 668808 128318
rect 668860 122868 668912 122874
rect 668860 122810 668912 122816
rect 668872 112713 668900 122810
rect 669976 117774 670004 168234
rect 670160 143478 670188 391954
rect 670240 324352 670292 324358
rect 670240 324294 670292 324300
rect 670252 176866 670280 324294
rect 670332 211200 670384 211206
rect 670332 211142 670384 211148
rect 670240 176860 670292 176866
rect 670240 176802 670292 176808
rect 670148 143472 670200 143478
rect 670148 143414 670200 143420
rect 670344 124098 670372 211142
rect 671356 163878 671384 614110
rect 671448 579970 671476 709310
rect 671816 665514 671844 730458
rect 671908 710462 671936 780710
rect 672000 755002 672028 879038
rect 671988 754996 672040 755002
rect 671988 754938 672040 754944
rect 672172 712428 672224 712434
rect 672172 712370 672224 712376
rect 671896 710456 671948 710462
rect 671896 710398 671948 710404
rect 671988 698216 672040 698222
rect 671988 698158 672040 698164
rect 671804 665508 671856 665514
rect 671804 665450 671856 665456
rect 671896 652792 671948 652798
rect 671896 652734 671948 652740
rect 671804 651568 671856 651574
rect 671804 651510 671856 651516
rect 671436 579964 671488 579970
rect 671436 579906 671488 579912
rect 671816 575754 671844 651510
rect 671908 575890 671936 652734
rect 672000 621178 672028 698158
rect 672184 666738 672212 712370
rect 672264 697400 672316 697406
rect 672264 697342 672316 697348
rect 672172 666732 672224 666738
rect 672172 666674 672224 666680
rect 671988 621172 672040 621178
rect 671988 621114 672040 621120
rect 672276 618458 672304 697342
rect 672368 669089 672396 956490
rect 672632 937168 672684 937174
rect 672632 937110 672684 937116
rect 672540 779340 672592 779346
rect 672540 779282 672592 779288
rect 672448 773628 672500 773634
rect 672448 773570 672500 773576
rect 672460 710054 672488 773570
rect 672448 710048 672500 710054
rect 672448 709990 672500 709996
rect 672552 708014 672580 779282
rect 672644 759354 672672 937110
rect 673184 937100 673236 937106
rect 673184 937042 673236 937048
rect 673092 873588 673144 873594
rect 673092 873530 673144 873536
rect 673000 869644 673052 869650
rect 673000 869586 673052 869592
rect 672908 869032 672960 869038
rect 672908 868974 672960 868980
rect 672816 862844 672868 862850
rect 672816 862786 672868 862792
rect 672724 855636 672776 855642
rect 672724 855578 672776 855584
rect 672632 759348 672684 759354
rect 672632 759290 672684 759296
rect 672632 733916 672684 733922
rect 672632 733858 672684 733864
rect 672540 708008 672592 708014
rect 672540 707950 672592 707956
rect 672448 669384 672500 669390
rect 672448 669326 672500 669332
rect 672354 669080 672410 669089
rect 672354 669015 672410 669024
rect 672460 624170 672488 669326
rect 672540 667956 672592 667962
rect 672540 667898 672592 667904
rect 672448 624164 672500 624170
rect 672448 624106 672500 624112
rect 672552 623966 672580 667898
rect 672644 661162 672672 733858
rect 672736 716582 672764 855578
rect 672828 755138 672856 862786
rect 672816 755132 672868 755138
rect 672816 755074 672868 755080
rect 672920 752282 672948 868974
rect 673012 752418 673040 869586
rect 673104 753642 673132 873530
rect 673196 759218 673224 937042
rect 673288 930306 673316 958326
rect 674840 957840 674892 957846
rect 674840 957782 674892 957788
rect 674748 957024 674800 957030
rect 674748 956966 674800 956972
rect 674564 955732 674616 955738
rect 674564 955674 674616 955680
rect 674196 948116 674248 948122
rect 674196 948058 674248 948064
rect 674208 939214 674236 948058
rect 674196 939208 674248 939214
rect 674196 939150 674248 939156
rect 673644 936692 673696 936698
rect 673644 936634 673696 936640
rect 673276 930300 673328 930306
rect 673276 930242 673328 930248
rect 673276 780020 673328 780026
rect 673276 779962 673328 779968
rect 673184 759212 673236 759218
rect 673184 759154 673236 759160
rect 673092 753636 673144 753642
rect 673092 753578 673144 753584
rect 673000 752412 673052 752418
rect 673000 752354 673052 752360
rect 672908 752276 672960 752282
rect 672908 752218 672960 752224
rect 673184 742552 673236 742558
rect 673184 742494 673236 742500
rect 673000 739152 673052 739158
rect 673000 739094 673052 739100
rect 672908 735004 672960 735010
rect 672908 734946 672960 734952
rect 672724 716576 672776 716582
rect 672724 716518 672776 716524
rect 672724 703860 672776 703866
rect 672724 703802 672776 703808
rect 672632 661156 672684 661162
rect 672632 661098 672684 661104
rect 672540 623960 672592 623966
rect 672540 623902 672592 623908
rect 672448 623892 672500 623898
rect 672448 623834 672500 623840
rect 672264 618452 672316 618458
rect 672264 618394 672316 618400
rect 672460 580106 672488 623834
rect 672540 623824 672592 623830
rect 672540 623766 672592 623772
rect 672448 580100 672500 580106
rect 672448 580042 672500 580048
rect 672552 578474 672580 623766
rect 672632 593428 672684 593434
rect 672632 593370 672684 593376
rect 672540 578468 672592 578474
rect 672540 578410 672592 578416
rect 672448 578332 672500 578338
rect 672448 578274 672500 578280
rect 671896 575884 671948 575890
rect 671896 575826 671948 575832
rect 671804 575748 671856 575754
rect 671804 575690 671856 575696
rect 671436 568608 671488 568614
rect 671436 568550 671488 568556
rect 671448 474570 671476 568550
rect 671988 561944 672040 561950
rect 671988 561886 672040 561892
rect 672000 485246 672028 561886
rect 672460 534546 672488 578274
rect 672540 578264 672592 578270
rect 672540 578206 672592 578212
rect 672448 534540 672500 534546
rect 672448 534482 672500 534488
rect 672552 534410 672580 578206
rect 672540 534404 672592 534410
rect 672540 534346 672592 534352
rect 672644 528698 672672 593370
rect 672632 528692 672684 528698
rect 672632 528634 672684 528640
rect 671988 485240 672040 485246
rect 671988 485182 672040 485188
rect 672078 474872 672134 474881
rect 672078 474807 672134 474816
rect 671436 474564 671488 474570
rect 671436 474506 671488 474512
rect 671528 350600 671580 350606
rect 671528 350542 671580 350548
rect 671436 346452 671488 346458
rect 671436 346394 671488 346400
rect 671344 163872 671396 163878
rect 671344 163814 671396 163820
rect 671448 138242 671476 346394
rect 671540 178362 671568 350542
rect 671620 256760 671672 256766
rect 671620 256702 671672 256708
rect 671528 178356 671580 178362
rect 671528 178298 671580 178304
rect 671528 167884 671580 167890
rect 671528 167826 671580 167832
rect 671436 138236 671488 138242
rect 671436 138178 671488 138184
rect 670332 124092 670384 124098
rect 670332 124034 670384 124040
rect 671344 121508 671396 121514
rect 671344 121450 671396 121456
rect 670056 120760 670108 120766
rect 670056 120702 670108 120708
rect 669964 117768 670016 117774
rect 669964 117710 670016 117716
rect 669228 114368 669280 114374
rect 669226 114336 669228 114345
rect 669280 114336 669282 114345
rect 669226 114271 669282 114280
rect 668858 112704 668914 112713
rect 668858 112639 668914 112648
rect 670068 109342 670096 120702
rect 671356 111790 671384 121450
rect 671540 117026 671568 167826
rect 671632 127974 671660 256702
rect 671620 127968 671672 127974
rect 671620 127910 671672 127916
rect 671528 117020 671580 117026
rect 671528 116962 671580 116968
rect 671344 111784 671396 111790
rect 671344 111726 671396 111732
rect 670056 109336 670108 109342
rect 670056 109278 670108 109284
rect 669228 106140 669280 106146
rect 669228 106082 669280 106088
rect 669240 105913 669268 106082
rect 669226 105904 669282 105913
rect 669226 105839 669282 105848
rect 668766 102504 668822 102513
rect 668766 102439 668822 102448
rect 668582 100872 668638 100881
rect 668582 100807 668638 100816
rect 605852 100014 606740 100042
rect 605748 77988 605800 77994
rect 605748 77930 605800 77936
rect 600964 57248 601016 57254
rect 600964 57190 601016 57196
rect 580264 55684 580316 55690
rect 580264 55626 580316 55632
rect 579068 53100 579120 53106
rect 579068 53042 579120 53048
rect 576122 47560 576178 47569
rect 576122 47495 576178 47504
rect 605852 44985 605880 100014
rect 607370 99770 607398 100028
rect 607324 99742 607398 99770
rect 607692 100014 608028 100042
rect 607220 95532 607272 95538
rect 607220 95474 607272 95480
rect 605838 44976 605894 44985
rect 605838 44911 605894 44920
rect 607232 43489 607260 95474
rect 607324 45121 607352 99742
rect 607692 95538 607720 100014
rect 608658 99770 608686 100028
rect 608612 99742 608686 99770
rect 608796 100014 609316 100042
rect 609960 100014 610020 100042
rect 607680 95532 607732 95538
rect 607680 95474 607732 95480
rect 607310 45112 607366 45121
rect 607310 45047 607366 45056
rect 608612 44849 608640 99742
rect 608796 53174 608824 100014
rect 608784 53168 608836 53174
rect 608784 53110 608836 53116
rect 608598 44840 608654 44849
rect 608598 44775 608654 44784
rect 607218 43480 607274 43489
rect 607218 43415 607274 43424
rect 518622 42392 518678 42401
rect 518678 42350 518834 42378
rect 518622 42327 518678 42336
rect 514850 42120 514906 42129
rect 520370 42120 520426 42129
rect 514906 42078 515154 42106
rect 514850 42055 514906 42064
rect 521750 42120 521806 42129
rect 520426 42078 520674 42106
rect 520370 42055 520426 42064
rect 529662 42120 529718 42129
rect 521806 42078 521870 42106
rect 529322 42078 529662 42106
rect 521750 42055 521806 42064
rect 529662 42055 529718 42064
rect 525890 41848 525946 41857
rect 525946 41806 526194 41834
rect 525890 41783 525946 41792
rect 478786 41576 478842 41585
rect 478786 41511 478842 41520
rect 609992 41449 610020 100014
rect 610176 100014 610604 100042
rect 610912 100014 611248 100042
rect 611464 100014 611892 100042
rect 612200 100014 612536 100042
rect 612752 100014 613180 100042
rect 613488 100014 613916 100042
rect 614560 100014 614896 100042
rect 615204 100014 615448 100042
rect 615848 100014 616184 100042
rect 616492 100014 616736 100042
rect 617136 100014 617472 100042
rect 617780 100014 618116 100042
rect 618424 100014 618760 100042
rect 619068 100014 619496 100042
rect 619712 100014 620048 100042
rect 620448 100014 620784 100042
rect 621092 100014 621428 100042
rect 621736 100014 622072 100042
rect 622380 100014 622716 100042
rect 623024 100014 623544 100042
rect 623668 100014 623728 100042
rect 624312 100014 624648 100042
rect 624956 100014 625108 100042
rect 625600 100014 625936 100042
rect 626244 100014 626396 100042
rect 610072 96960 610124 96966
rect 610072 96902 610124 96908
rect 610084 45257 610112 96902
rect 610176 46209 610204 100014
rect 610912 96966 610940 100014
rect 610900 96960 610952 96966
rect 610900 96902 610952 96908
rect 611360 96960 611412 96966
rect 611360 96902 611412 96908
rect 611372 46617 611400 96902
rect 611358 46608 611414 46617
rect 611358 46543 611414 46552
rect 611464 46345 611492 100014
rect 612200 96966 612228 100014
rect 612188 96960 612240 96966
rect 612188 96902 612240 96908
rect 612752 46481 612780 100014
rect 613488 84194 613516 100014
rect 614868 97510 614896 100014
rect 614856 97504 614908 97510
rect 614856 97446 614908 97452
rect 612844 84166 613516 84194
rect 612844 47705 612872 84166
rect 615420 75206 615448 100014
rect 616156 96966 616184 100014
rect 616144 96960 616196 96966
rect 616144 96902 616196 96908
rect 616708 89690 616736 100014
rect 617444 96966 617472 100014
rect 616788 96960 616840 96966
rect 616788 96902 616840 96908
rect 617432 96960 617484 96966
rect 617432 96902 617484 96908
rect 616696 89684 616748 89690
rect 616696 89626 616748 89632
rect 616800 88330 616828 96902
rect 616788 88324 616840 88330
rect 616788 88266 616840 88272
rect 618088 84114 618116 100014
rect 618168 96960 618220 96966
rect 618168 96902 618220 96908
rect 618180 84182 618208 96902
rect 618732 96898 618760 100014
rect 618720 96892 618772 96898
rect 618720 96834 618772 96840
rect 619468 86290 619496 100014
rect 620020 96898 620048 100014
rect 620756 97442 620784 100014
rect 620744 97436 620796 97442
rect 620744 97378 620796 97384
rect 621400 97238 621428 100014
rect 621664 97504 621716 97510
rect 621664 97446 621716 97452
rect 621388 97232 621440 97238
rect 621388 97174 621440 97180
rect 619548 96892 619600 96898
rect 619548 96834 619600 96840
rect 620008 96892 620060 96898
rect 620008 96834 620060 96840
rect 620928 96892 620980 96898
rect 620928 96834 620980 96840
rect 619456 86284 619508 86290
rect 619456 86226 619508 86232
rect 619560 85542 619588 96834
rect 620940 88262 620968 96834
rect 620928 88256 620980 88262
rect 620928 88198 620980 88204
rect 619548 85536 619600 85542
rect 619548 85478 619600 85484
rect 618168 84176 618220 84182
rect 618168 84118 618220 84124
rect 618076 84108 618128 84114
rect 618076 84050 618128 84056
rect 617524 75268 617576 75274
rect 617524 75210 617576 75216
rect 615408 75200 615460 75206
rect 615408 75142 615460 75148
rect 617536 62150 617564 75210
rect 617524 62144 617576 62150
rect 617524 62086 617576 62092
rect 614764 62076 614816 62082
rect 614764 62018 614816 62024
rect 614776 52494 614804 62018
rect 621676 57254 621704 97446
rect 622044 97306 622072 100014
rect 622032 97300 622084 97306
rect 622032 97242 622084 97248
rect 622688 96830 622716 100014
rect 622676 96824 622728 96830
rect 622676 96766 622728 96772
rect 623516 93854 623544 100014
rect 623700 96966 623728 100014
rect 624620 97986 624648 100014
rect 624608 97980 624660 97986
rect 624608 97922 624660 97928
rect 623688 96960 623740 96966
rect 623688 96902 623740 96908
rect 624424 96960 624476 96966
rect 624424 96902 624476 96908
rect 623688 96824 623740 96830
rect 623688 96766 623740 96772
rect 623516 93826 623636 93854
rect 623608 79354 623636 93826
rect 623596 79348 623648 79354
rect 623596 79290 623648 79296
rect 623700 76566 623728 96766
rect 624436 80714 624464 96902
rect 625080 90001 625108 100014
rect 625804 97980 625856 97986
rect 625804 97922 625856 97928
rect 625066 89992 625122 90001
rect 625066 89927 625122 89936
rect 625816 89729 625844 97922
rect 625908 96966 625936 100014
rect 625896 96960 625948 96966
rect 625896 96902 625948 96908
rect 626368 92585 626396 100014
rect 626552 100014 626980 100042
rect 627624 100014 627868 100042
rect 628268 100014 628328 100042
rect 626448 96960 626500 96966
rect 626448 96902 626500 96908
rect 626354 92576 626410 92585
rect 626354 92511 626410 92520
rect 626460 91633 626488 96902
rect 626552 93537 626580 100014
rect 627840 94489 627868 100014
rect 628300 95985 628328 100014
rect 628760 100014 628912 100042
rect 629556 100014 629708 100042
rect 630200 100014 630628 100042
rect 630844 100014 631180 100042
rect 631488 100014 631824 100042
rect 632132 100014 632468 100042
rect 632776 100014 633112 100042
rect 633512 100014 633848 100042
rect 634156 100014 634492 100042
rect 634800 100014 635136 100042
rect 635444 100014 635780 100042
rect 636088 100014 636148 100042
rect 636732 100014 637068 100042
rect 637376 100014 637528 100042
rect 638020 100014 638356 100042
rect 638664 100014 638908 100042
rect 639308 100014 639644 100042
rect 639952 100014 640104 100042
rect 640688 100014 641024 100042
rect 641332 100014 641668 100042
rect 628286 95976 628342 95985
rect 628286 95911 628342 95920
rect 628760 95826 628788 100014
rect 628728 95798 628788 95826
rect 629680 95826 629708 100014
rect 630600 96642 630628 100014
rect 631152 97646 631180 100014
rect 631140 97640 631192 97646
rect 631140 97582 631192 97588
rect 631796 97170 631824 100014
rect 632152 97640 632204 97646
rect 632152 97582 632204 97588
rect 631784 97164 631836 97170
rect 631784 97106 631836 97112
rect 630600 96614 630720 96642
rect 630692 95826 630720 96614
rect 629680 95798 629832 95826
rect 630692 95798 631028 95826
rect 632164 95690 632192 97582
rect 632440 96898 632468 100014
rect 633084 97918 633112 100014
rect 633820 97986 633848 100014
rect 633808 97980 633860 97986
rect 633808 97922 633860 97928
rect 633072 97912 633124 97918
rect 633072 97854 633124 97860
rect 634464 97714 634492 100014
rect 635108 97782 635136 100014
rect 635280 97912 635332 97918
rect 635280 97854 635332 97860
rect 635096 97776 635148 97782
rect 635096 97718 635148 97724
rect 634452 97708 634504 97714
rect 634452 97650 634504 97656
rect 632980 97164 633032 97170
rect 632980 97106 633032 97112
rect 632428 96892 632480 96898
rect 632428 96834 632480 96840
rect 632992 95826 633020 97106
rect 634084 96892 634136 96898
rect 634084 96834 634136 96840
rect 634096 95826 634124 96834
rect 635292 95826 635320 97854
rect 635752 97646 635780 100014
rect 635740 97640 635792 97646
rect 635740 97582 635792 97588
rect 636120 96762 636148 100014
rect 636384 97980 636436 97986
rect 636384 97922 636436 97928
rect 636108 96756 636160 96762
rect 636108 96698 636160 96704
rect 636396 95826 636424 97922
rect 637040 97578 637068 100014
rect 637500 97918 637528 100014
rect 637488 97912 637540 97918
rect 637488 97854 637540 97860
rect 638328 97850 638356 100014
rect 638316 97844 638368 97850
rect 638316 97786 638368 97792
rect 637580 97708 637632 97714
rect 637580 97650 637632 97656
rect 637028 97572 637080 97578
rect 637028 97514 637080 97520
rect 637592 95826 637620 97650
rect 632992 95798 633328 95826
rect 634096 95798 634432 95826
rect 635292 95798 635628 95826
rect 636396 95798 636732 95826
rect 637592 95798 637928 95826
rect 632132 95662 632192 95690
rect 638880 95606 638908 100014
rect 639052 97776 639104 97782
rect 639052 97718 639104 97724
rect 639064 95690 639092 97718
rect 639616 96626 639644 100014
rect 639880 97640 639932 97646
rect 639880 97582 639932 97588
rect 639604 96620 639656 96626
rect 639604 96562 639656 96568
rect 639892 95826 639920 97582
rect 640076 95946 640104 100014
rect 640996 96898 641024 100014
rect 640984 96892 641036 96898
rect 640984 96834 641036 96840
rect 640984 96756 641036 96762
rect 640984 96698 641036 96704
rect 640064 95940 640116 95946
rect 640064 95882 640116 95888
rect 640996 95826 641024 96698
rect 639892 95798 640228 95826
rect 640996 95798 641332 95826
rect 639032 95662 639092 95690
rect 641640 95674 641668 100014
rect 641732 100014 641976 100042
rect 642284 100014 642620 100042
rect 643264 100014 643600 100042
rect 643908 100014 644428 100042
rect 644552 100014 644888 100042
rect 645196 100014 645532 100042
rect 645840 100014 646176 100042
rect 646484 100014 646820 100042
rect 647220 100014 647556 100042
rect 647864 100014 648200 100042
rect 648508 100014 648568 100042
rect 649152 100014 649488 100042
rect 649796 100014 649948 100042
rect 650440 100014 650776 100042
rect 651084 100014 651236 100042
rect 651728 100014 652064 100042
rect 652372 100014 652708 100042
rect 653016 100014 653352 100042
rect 653752 100014 653996 100042
rect 654396 100014 654732 100042
rect 655040 100014 655376 100042
rect 655684 100014 656020 100042
rect 656328 100014 656664 100042
rect 656972 100014 657308 100042
rect 641732 95849 641760 100014
rect 642180 97572 642232 97578
rect 642180 97514 642232 97520
rect 641718 95840 641774 95849
rect 642192 95826 642220 97514
rect 642284 96529 642312 100014
rect 643572 97510 643600 100014
rect 643560 97504 643612 97510
rect 643560 97446 643612 97452
rect 643284 96892 643336 96898
rect 643284 96834 643336 96840
rect 643100 96620 643152 96626
rect 643100 96562 643152 96568
rect 642270 96520 642326 96529
rect 642270 96455 642326 96464
rect 642192 95798 642528 95826
rect 641718 95775 641774 95784
rect 641628 95668 641680 95674
rect 641628 95610 641680 95616
rect 638868 95600 638920 95606
rect 638868 95542 638920 95548
rect 627826 94480 627882 94489
rect 627826 94415 627882 94424
rect 626538 93528 626594 93537
rect 626538 93463 626594 93472
rect 626446 91624 626502 91633
rect 626446 91559 626502 91568
rect 625802 89720 625858 89729
rect 625802 89655 625858 89664
rect 626448 89684 626500 89690
rect 626448 89626 626500 89632
rect 626460 88913 626488 89626
rect 626446 88904 626502 88913
rect 626446 88839 626502 88848
rect 626448 88324 626500 88330
rect 626448 88266 626500 88272
rect 626356 88256 626408 88262
rect 626356 88198 626408 88204
rect 626368 87009 626396 88198
rect 626460 87961 626488 88266
rect 626446 87952 626502 87961
rect 626446 87887 626502 87896
rect 643112 87689 643140 96562
rect 643098 87680 643154 87689
rect 643098 87615 643154 87624
rect 626354 87000 626410 87009
rect 626354 86935 626410 86944
rect 626448 86284 626500 86290
rect 626448 86226 626500 86232
rect 626460 86057 626488 86226
rect 626446 86048 626502 86057
rect 626446 85983 626502 85992
rect 626448 85536 626500 85542
rect 626448 85478 626500 85484
rect 626460 85105 626488 85478
rect 626446 85096 626502 85105
rect 626446 85031 626502 85040
rect 626080 84176 626132 84182
rect 625618 84144 625674 84153
rect 626080 84118 626132 84124
rect 625618 84079 625620 84088
rect 625672 84079 625674 84088
rect 625620 84050 625672 84056
rect 626092 83201 626120 84118
rect 626078 83192 626134 83201
rect 626078 83127 626134 83136
rect 643296 82249 643324 96834
rect 644400 92478 644428 100014
rect 644664 97912 644716 97918
rect 644664 97854 644716 97860
rect 644572 95940 644624 95946
rect 644572 95882 644624 95888
rect 644480 95600 644532 95606
rect 644480 95542 644532 95548
rect 644388 92472 644440 92478
rect 644388 92414 644440 92420
rect 644492 89729 644520 95542
rect 644478 89720 644534 89729
rect 644478 89655 644534 89664
rect 644584 84697 644612 95882
rect 644676 94625 644704 97854
rect 644756 97844 644808 97850
rect 644756 97786 644808 97792
rect 644662 94616 644718 94625
rect 644662 94551 644718 94560
rect 644768 92177 644796 97786
rect 644860 96626 644888 100014
rect 645504 96966 645532 100014
rect 646044 97436 646096 97442
rect 646044 97378 646096 97384
rect 645492 96960 645544 96966
rect 645492 96902 645544 96908
rect 644848 96620 644900 96626
rect 644848 96562 644900 96568
rect 645952 95668 646004 95674
rect 645952 95610 646004 95616
rect 644754 92168 644810 92177
rect 644754 92103 644810 92112
rect 644570 84688 644626 84697
rect 644570 84623 644626 84632
rect 626446 82240 626502 82249
rect 626446 82175 626502 82184
rect 643282 82240 643338 82249
rect 643282 82175 643338 82184
rect 624424 80708 624476 80714
rect 624424 80650 624476 80656
rect 626460 78198 626488 82175
rect 631520 80974 631856 81002
rect 638972 80974 639308 81002
rect 629206 80880 629262 80889
rect 629206 80815 629262 80824
rect 626448 78192 626500 78198
rect 626448 78134 626500 78140
rect 629220 78062 629248 80815
rect 631048 78124 631100 78130
rect 631048 78066 631100 78072
rect 629208 78056 629260 78062
rect 629208 77998 629260 78004
rect 628380 77648 628432 77654
rect 628380 77590 628432 77596
rect 628392 77382 628420 77590
rect 628380 77376 628432 77382
rect 628380 77318 628432 77324
rect 623688 76560 623740 76566
rect 623688 76502 623740 76508
rect 628392 75290 628420 77318
rect 631060 77314 631088 78066
rect 631520 77654 631548 80974
rect 638972 78130 639000 80974
rect 642456 78192 642508 78198
rect 642456 78134 642508 78140
rect 638960 78124 639012 78130
rect 638960 78066 639012 78072
rect 636752 77988 636804 77994
rect 636752 77930 636804 77936
rect 633898 77752 633954 77761
rect 633898 77687 633954 77696
rect 631508 77648 631560 77654
rect 631508 77590 631560 77596
rect 631048 77308 631100 77314
rect 631048 77250 631100 77256
rect 631060 75290 631088 77250
rect 633912 75993 633940 77687
rect 631138 75984 631194 75993
rect 631138 75919 631194 75928
rect 633898 75984 633954 75993
rect 633898 75919 633954 75928
rect 628176 75262 628420 75290
rect 631028 75262 631088 75290
rect 631152 75274 631180 75919
rect 633912 75290 633940 75919
rect 636764 75290 636792 77930
rect 639602 77752 639658 77761
rect 639602 77687 639658 77696
rect 639616 75290 639644 77687
rect 642468 75290 642496 78134
rect 645308 78056 645360 78062
rect 645308 77998 645360 78004
rect 645320 75290 645348 77998
rect 631140 75268 631192 75274
rect 633880 75262 633940 75290
rect 636732 75262 636792 75290
rect 639584 75276 639644 75290
rect 639570 75262 639644 75276
rect 642436 75262 642496 75290
rect 645288 75262 645348 75290
rect 631140 75210 631192 75216
rect 639234 75168 639290 75177
rect 639570 75154 639598 75262
rect 639290 75140 639598 75154
rect 639290 75126 639584 75140
rect 639234 75103 639290 75112
rect 645964 64874 645992 95610
rect 646056 66042 646084 97378
rect 646148 95946 646176 100014
rect 646504 96960 646556 96966
rect 646504 96902 646556 96908
rect 646136 95940 646188 95946
rect 646136 95882 646188 95888
rect 646516 87038 646544 96902
rect 646792 96082 646820 100014
rect 647528 97850 647556 100014
rect 647516 97844 647568 97850
rect 647516 97786 647568 97792
rect 648172 97442 648200 100014
rect 648160 97436 648212 97442
rect 648160 97378 648212 97384
rect 647424 97232 647476 97238
rect 647424 97174 647476 97180
rect 646780 96076 646832 96082
rect 646780 96018 646832 96024
rect 646504 87032 646556 87038
rect 646504 86974 646556 86980
rect 647332 79348 647384 79354
rect 647332 79290 647384 79296
rect 646136 76560 646188 76566
rect 646136 76502 646188 76508
rect 646148 70417 646176 76502
rect 646872 75200 646924 75206
rect 646872 75142 646924 75148
rect 646884 74497 646912 75142
rect 646870 74488 646926 74497
rect 646870 74423 646926 74432
rect 647344 71505 647372 79290
rect 647330 71496 647386 71505
rect 647330 71431 647386 71440
rect 646134 70408 646190 70417
rect 646134 70343 646190 70352
rect 647436 67017 647464 97174
rect 648540 86766 648568 100014
rect 649460 97918 649488 100014
rect 649448 97912 649500 97918
rect 649448 97854 649500 97860
rect 648620 97300 648672 97306
rect 648620 97242 648672 97248
rect 648632 93854 648660 97242
rect 648632 93826 648844 93854
rect 648528 86760 648580 86766
rect 648528 86702 648580 86708
rect 648712 80708 648764 80714
rect 648712 80650 648764 80656
rect 648724 73001 648752 80650
rect 648710 72992 648766 73001
rect 648710 72927 648766 72936
rect 648816 68513 648844 93826
rect 649920 86834 649948 100014
rect 650748 96898 650776 100014
rect 650736 96892 650788 96898
rect 650736 96834 650788 96840
rect 651208 86970 651236 100014
rect 652036 97374 652064 100014
rect 652024 97368 652076 97374
rect 652024 97310 652076 97316
rect 651288 96892 651340 96898
rect 651288 96834 651340 96840
rect 651196 86964 651248 86970
rect 651196 86906 651248 86912
rect 651300 86902 651328 96834
rect 651932 96620 651984 96626
rect 651932 96562 651984 96568
rect 651944 90982 651972 96562
rect 651932 90976 651984 90982
rect 651932 90918 651984 90924
rect 651288 86896 651340 86902
rect 651288 86838 651340 86844
rect 649908 86828 649960 86834
rect 649908 86770 649960 86776
rect 652680 86630 652708 100014
rect 653324 96014 653352 100014
rect 653312 96008 653364 96014
rect 653312 95950 653364 95956
rect 653968 86698 653996 100014
rect 654704 97238 654732 100014
rect 654784 97844 654836 97850
rect 654784 97786 654836 97792
rect 654692 97232 654744 97238
rect 654692 97174 654744 97180
rect 654796 92585 654824 97786
rect 655348 93401 655376 100014
rect 655992 97374 656020 100014
rect 655980 97368 656032 97374
rect 655980 97310 656032 97316
rect 655428 96960 655480 96966
rect 655428 96902 655480 96908
rect 655334 93392 655390 93401
rect 655334 93327 655390 93336
rect 654782 92576 654838 92585
rect 654782 92511 654838 92520
rect 654324 92472 654376 92478
rect 654324 92414 654376 92420
rect 654336 91497 654364 92414
rect 654322 91488 654378 91497
rect 654322 91423 654378 91432
rect 654324 90976 654376 90982
rect 654324 90918 654376 90924
rect 654336 90681 654364 90918
rect 654322 90672 654378 90681
rect 654322 90607 654378 90616
rect 655440 89865 655468 96902
rect 656636 96218 656664 100014
rect 656808 96620 656860 96626
rect 656808 96562 656860 96568
rect 656624 96212 656676 96218
rect 656624 96154 656676 96160
rect 655426 89856 655482 89865
rect 655426 89791 655482 89800
rect 656820 88874 656848 96562
rect 657280 95266 657308 100014
rect 657372 100014 657616 100042
rect 658260 100014 658320 100042
rect 658904 100014 659240 100042
rect 657268 95260 657320 95266
rect 657268 95202 657320 95208
rect 657372 94761 657400 100014
rect 657728 97300 657780 97306
rect 657728 97242 657780 97248
rect 657740 95132 657768 97242
rect 658292 96626 658320 100014
rect 658832 97912 658884 97918
rect 658832 97854 658884 97860
rect 658372 97232 658424 97238
rect 658372 97174 658424 97180
rect 658280 96620 658332 96626
rect 658280 96562 658332 96568
rect 658384 95146 658412 97174
rect 658306 95118 658412 95146
rect 658844 95132 658872 97854
rect 659212 96830 659240 100014
rect 659304 100014 659548 100042
rect 660284 100014 660620 100042
rect 659304 96966 659332 100014
rect 660396 97504 660448 97510
rect 660396 97446 660448 97452
rect 660120 97436 660172 97442
rect 660120 97378 660172 97384
rect 659568 97368 659620 97374
rect 659568 97310 659620 97316
rect 659292 96960 659344 96966
rect 659292 96902 659344 96908
rect 659200 96824 659252 96830
rect 659200 96766 659252 96772
rect 659580 95132 659608 97310
rect 660132 95132 660160 97378
rect 660408 95146 660436 97446
rect 660592 97238 660620 100014
rect 660684 100014 660928 100042
rect 661572 100014 661908 100042
rect 662216 100014 662368 100042
rect 662860 100014 663104 100042
rect 660684 97306 660712 100014
rect 660672 97300 660724 97306
rect 660672 97242 660724 97248
rect 660580 97232 660632 97238
rect 660580 97174 660632 97180
rect 661408 97232 661460 97238
rect 661408 97174 661460 97180
rect 660408 95118 660698 95146
rect 661420 95132 661448 97174
rect 661880 96898 661908 100014
rect 662340 97170 662368 100014
rect 663076 97986 663104 100014
rect 663168 100014 663504 100042
rect 663064 97980 663116 97986
rect 663064 97922 663116 97928
rect 661960 97164 662012 97170
rect 661960 97106 662012 97112
rect 662328 97164 662380 97170
rect 662328 97106 662380 97112
rect 661868 96892 661920 96898
rect 661868 96834 661920 96840
rect 661972 95132 662000 97106
rect 663064 96892 663116 96898
rect 663064 96834 663116 96840
rect 662512 96824 662564 96830
rect 662512 96766 662564 96772
rect 662524 95132 662552 96766
rect 663076 95132 663104 96834
rect 657358 94752 657414 94761
rect 657358 94687 657414 94696
rect 658108 88874 658306 88890
rect 656808 88868 656860 88874
rect 656808 88810 656860 88816
rect 658096 88868 658306 88874
rect 658148 88862 658306 88868
rect 661986 88874 662368 88890
rect 661986 88868 662380 88874
rect 661986 88862 662328 88868
rect 658096 88810 658148 88816
rect 662328 88810 662380 88816
rect 659488 88330 659594 88346
rect 663168 88330 663196 100014
rect 665364 97980 665416 97986
rect 665364 97922 665416 97928
rect 663984 97164 664036 97170
rect 663984 97106 664036 97112
rect 663892 96212 663944 96218
rect 663892 96154 663944 96160
rect 663800 96076 663852 96082
rect 663800 96018 663852 96024
rect 663812 92585 663840 96018
rect 663798 92576 663854 92585
rect 663798 92511 663854 92520
rect 663904 90681 663932 96154
rect 663890 90672 663946 90681
rect 663890 90607 663946 90616
rect 663996 88874 664024 97106
rect 665272 96008 665324 96014
rect 665272 95950 665324 95956
rect 665180 95940 665232 95946
rect 665180 95882 665232 95888
rect 664076 95260 664128 95266
rect 664076 95202 664128 95208
rect 664088 89049 664116 95202
rect 665192 91769 665220 95882
rect 665178 91760 665234 91769
rect 665178 91695 665234 91704
rect 665284 89865 665312 95950
rect 665376 93401 665404 97922
rect 665362 93392 665418 93401
rect 665362 93327 665418 93336
rect 665270 89856 665326 89865
rect 665270 89791 665326 89800
rect 664074 89040 664130 89049
rect 664074 88975 664130 88984
rect 663984 88868 664036 88874
rect 663984 88810 664036 88816
rect 659476 88324 659594 88330
rect 659528 88318 659594 88324
rect 663156 88324 663208 88330
rect 659476 88266 659528 88272
rect 663156 88266 663208 88272
rect 657188 86970 657216 88196
rect 657176 86964 657228 86970
rect 657176 86906 657228 86912
rect 657740 86902 657768 88196
rect 657728 86896 657780 86902
rect 657728 86838 657780 86844
rect 658844 86698 658872 88196
rect 660132 87038 660160 88196
rect 660120 87032 660172 87038
rect 660120 86974 660172 86980
rect 660684 86834 660712 88196
rect 660672 86828 660724 86834
rect 660672 86770 660724 86776
rect 661420 86766 661448 88196
rect 661408 86760 661460 86766
rect 661408 86702 661460 86708
rect 653956 86692 654008 86698
rect 653956 86634 654008 86640
rect 658832 86692 658884 86698
rect 658832 86634 658884 86640
rect 662524 86630 662552 88196
rect 652668 86624 652720 86630
rect 652668 86566 652720 86572
rect 662512 86624 662564 86630
rect 662512 86566 662564 86572
rect 648802 68504 648858 68513
rect 648802 68439 648858 68448
rect 647422 67008 647478 67017
rect 647422 66943 647478 66952
rect 646134 66056 646190 66065
rect 646056 66014 646134 66042
rect 646134 65991 646190 66000
rect 645964 64846 646176 64874
rect 646148 64433 646176 64846
rect 646134 64424 646190 64433
rect 646134 64359 646190 64368
rect 621664 57248 621716 57254
rect 621664 57190 621716 57196
rect 662420 57248 662472 57254
rect 662420 57190 662472 57196
rect 614764 52488 614816 52494
rect 614764 52430 614816 52436
rect 612830 47696 612886 47705
rect 612830 47631 612886 47640
rect 661130 47560 661186 47569
rect 661130 47495 661186 47504
rect 661144 46898 661172 47495
rect 662432 47433 662460 57190
rect 672092 49570 672120 474807
rect 672632 220244 672684 220250
rect 672632 220186 672684 220192
rect 672644 175710 672672 220186
rect 672632 175704 672684 175710
rect 672632 175646 672684 175652
rect 672736 173806 672764 703802
rect 672816 689376 672868 689382
rect 672816 689318 672868 689324
rect 672828 616894 672856 689318
rect 672920 661298 672948 734946
rect 673012 663814 673040 739094
rect 673092 738676 673144 738682
rect 673092 738618 673144 738624
rect 673000 663808 673052 663814
rect 673000 663750 673052 663756
rect 673104 662454 673132 738618
rect 673196 664018 673224 742494
rect 673288 706722 673316 779962
rect 673656 758878 673684 936634
rect 674576 932006 674604 955674
rect 674656 935876 674708 935882
rect 674656 935818 674708 935824
rect 674564 932000 674616 932006
rect 674564 931942 674616 931948
rect 674380 869848 674432 869854
rect 674380 869790 674432 869796
rect 674288 787364 674340 787370
rect 674288 787306 674340 787312
rect 674196 784304 674248 784310
rect 674196 784246 674248 784252
rect 674012 782944 674064 782950
rect 674012 782886 674064 782892
rect 673736 778660 673788 778666
rect 673736 778602 673788 778608
rect 673644 758872 673696 758878
rect 673644 758814 673696 758820
rect 673552 758260 673604 758266
rect 673552 758202 673604 758208
rect 673368 756288 673420 756294
rect 673368 756230 673420 756236
rect 673380 712910 673408 756230
rect 673564 713726 673592 758202
rect 673644 738268 673696 738274
rect 673644 738210 673696 738216
rect 673552 713720 673604 713726
rect 673552 713662 673604 713668
rect 673368 712904 673420 712910
rect 673368 712846 673420 712852
rect 673276 706716 673328 706722
rect 673276 706658 673328 706664
rect 673552 693048 673604 693054
rect 673552 692990 673604 692996
rect 673368 690464 673420 690470
rect 673368 690406 673420 690412
rect 673184 664012 673236 664018
rect 673184 663954 673236 663960
rect 673092 662448 673144 662454
rect 673092 662390 673144 662396
rect 672908 661292 672960 661298
rect 672908 661234 672960 661240
rect 673184 647760 673236 647766
rect 673184 647702 673236 647708
rect 673000 645040 673052 645046
rect 673000 644982 673052 644988
rect 672816 616888 672868 616894
rect 672816 616830 672868 616836
rect 672816 600432 672868 600438
rect 672816 600374 672868 600380
rect 672828 530194 672856 600374
rect 672908 597780 672960 597786
rect 672908 597722 672960 597728
rect 672816 530188 672868 530194
rect 672816 530130 672868 530136
rect 672920 527474 672948 597722
rect 673012 571538 673040 644982
rect 673092 643408 673144 643414
rect 673092 643350 673144 643356
rect 673000 571532 673052 571538
rect 673000 571474 673052 571480
rect 673104 569974 673132 643350
rect 673196 571674 673224 647702
rect 673276 639124 673328 639130
rect 673276 639066 673328 639072
rect 673288 574258 673316 639066
rect 673380 619818 673408 690406
rect 673460 623076 673512 623082
rect 673460 623018 673512 623024
rect 673368 619812 673420 619818
rect 673368 619754 673420 619760
rect 673368 607640 673420 607646
rect 673368 607582 673420 607588
rect 673276 574252 673328 574258
rect 673276 574194 673328 574200
rect 673184 571668 673236 571674
rect 673184 571610 673236 571616
rect 673092 569968 673144 569974
rect 673092 569910 673144 569916
rect 673276 559156 673328 559162
rect 673276 559098 673328 559104
rect 673184 557592 673236 557598
rect 673184 557534 673236 557540
rect 673092 554804 673144 554810
rect 673092 554746 673144 554752
rect 672908 527468 672960 527474
rect 672908 527410 672960 527416
rect 673104 482798 673132 554746
rect 673196 483206 673224 557534
rect 673288 484838 673316 559098
rect 673380 528834 673408 607582
rect 673472 578202 673500 623018
rect 673564 617438 673592 692990
rect 673656 662386 673684 738210
rect 673748 706790 673776 778602
rect 673920 777368 673972 777374
rect 673920 777310 673972 777316
rect 673828 759076 673880 759082
rect 673828 759018 673880 759024
rect 673840 714542 673868 759018
rect 673828 714536 673880 714542
rect 673828 714478 673880 714484
rect 673828 714060 673880 714066
rect 673828 714002 673880 714008
rect 673736 706784 673788 706790
rect 673736 706726 673788 706732
rect 673840 669526 673868 714002
rect 673932 708422 673960 777310
rect 673920 708416 673972 708422
rect 673920 708358 673972 708364
rect 674024 707606 674052 782886
rect 674208 709238 674236 784246
rect 674300 709646 674328 787306
rect 674392 755614 674420 869790
rect 674564 868080 674616 868086
rect 674564 868022 674616 868028
rect 674472 866856 674524 866862
rect 674472 866798 674524 866804
rect 674380 755608 674432 755614
rect 674380 755550 674432 755556
rect 674484 753438 674512 866798
rect 674472 753432 674524 753438
rect 674472 753374 674524 753380
rect 674576 751942 674604 868022
rect 674668 759121 674696 935818
rect 674760 930209 674788 956966
rect 674852 955534 674880 957782
rect 675036 957681 675064 961998
rect 675772 961353 675800 961755
rect 675758 961344 675814 961353
rect 675758 961279 675814 961288
rect 675680 959177 675708 959276
rect 675666 959168 675722 959177
rect 675666 959103 675722 959112
rect 675404 958390 675432 958732
rect 675392 958384 675444 958390
rect 675392 958326 675444 958332
rect 675496 957817 675524 958052
rect 675482 957808 675538 957817
rect 675482 957743 675538 957752
rect 675022 957672 675078 957681
rect 675022 957607 675078 957616
rect 675404 957030 675432 957440
rect 675392 957024 675444 957030
rect 675392 956966 675444 956972
rect 675036 956554 675142 956570
rect 675024 956548 675142 956554
rect 675076 956542 675142 956548
rect 675024 956490 675076 956496
rect 675496 955738 675524 956216
rect 675484 955732 675536 955738
rect 675484 955674 675536 955680
rect 674840 955528 674892 955534
rect 674840 955470 674892 955476
rect 675484 955528 675536 955534
rect 675484 955470 675536 955476
rect 675496 955060 675524 955470
rect 675772 954009 675800 954380
rect 675758 954000 675814 954009
rect 675758 953935 675814 953944
rect 675772 952066 675800 952544
rect 675760 952060 675812 952066
rect 675760 952002 675812 952008
rect 675760 951788 675812 951794
rect 675760 951730 675812 951736
rect 675772 949482 675800 951730
rect 677506 951008 677562 951017
rect 677506 950943 677562 950952
rect 677414 950872 677470 950881
rect 677414 950807 677470 950816
rect 675760 949476 675812 949482
rect 675760 949418 675812 949424
rect 676034 939992 676090 940001
rect 676034 939927 676090 939936
rect 676048 939826 676076 939927
rect 676036 939820 676088 939826
rect 676036 939762 676088 939768
rect 676218 939312 676274 939321
rect 676218 939247 676274 939256
rect 676036 939208 676088 939214
rect 676034 939176 676036 939185
rect 676088 939176 676090 939185
rect 676034 939111 676090 939120
rect 676034 938768 676090 938777
rect 676232 938738 676260 939247
rect 676034 938703 676090 938712
rect 676220 938732 676272 938738
rect 676048 938602 676076 938703
rect 676220 938674 676272 938680
rect 676036 938596 676088 938602
rect 676036 938538 676088 938544
rect 676126 938088 676182 938097
rect 676126 938023 676182 938032
rect 676034 937544 676090 937553
rect 676034 937479 676090 937488
rect 676048 937106 676076 937479
rect 676140 937174 676168 938023
rect 676218 937680 676274 937689
rect 676218 937615 676274 937624
rect 676232 937378 676260 937615
rect 676220 937372 676272 937378
rect 676220 937314 676272 937320
rect 676218 937272 676274 937281
rect 676218 937207 676220 937216
rect 676272 937207 676274 937216
rect 676220 937178 676272 937184
rect 676128 937168 676180 937174
rect 676128 937110 676180 937116
rect 676036 937100 676088 937106
rect 676036 937042 676088 937048
rect 676034 936728 676090 936737
rect 676034 936663 676036 936672
rect 676088 936663 676090 936672
rect 676036 936634 676088 936640
rect 676218 936048 676274 936057
rect 676218 935983 676274 935992
rect 676034 935912 676090 935921
rect 676034 935847 676036 935856
rect 676088 935847 676090 935856
rect 676036 935818 676088 935824
rect 676232 935678 676260 935983
rect 676220 935672 676272 935678
rect 676220 935614 676272 935620
rect 677428 934833 677456 950807
rect 677414 934824 677470 934833
rect 677414 934759 677470 934768
rect 677520 933201 677548 950943
rect 681002 949784 681058 949793
rect 681002 949719 681058 949728
rect 679806 949648 679862 949657
rect 679806 949583 679862 949592
rect 679622 949512 679678 949521
rect 678244 949476 678296 949482
rect 679622 949447 679678 949456
rect 678244 949418 678296 949424
rect 678256 933609 678284 949418
rect 678242 933600 678298 933609
rect 678242 933535 678298 933544
rect 677506 933192 677562 933201
rect 677506 933127 677562 933136
rect 676220 932000 676272 932006
rect 676218 931968 676220 931977
rect 676272 931968 676274 931977
rect 676218 931903 676274 931912
rect 679636 931161 679664 949447
rect 679820 931569 679848 949583
rect 681016 934425 681044 949719
rect 681094 948832 681150 948841
rect 681094 948767 681150 948776
rect 681002 934416 681058 934425
rect 681002 934351 681058 934360
rect 681108 934017 681136 948767
rect 682382 948016 682438 948025
rect 682382 947951 682438 947960
rect 682396 935241 682424 947951
rect 703694 940508 703722 940644
rect 704154 940508 704182 940644
rect 704614 940508 704642 940644
rect 705074 940508 705102 940644
rect 705534 940508 705562 940644
rect 705994 940508 706022 940644
rect 706454 940508 706482 940644
rect 706914 940508 706942 940644
rect 707374 940508 707402 940644
rect 707834 940508 707862 940644
rect 708294 940508 708322 940644
rect 708754 940508 708782 940644
rect 709214 940508 709242 940644
rect 682382 935232 682438 935241
rect 682382 935167 682438 935176
rect 681094 934008 681150 934017
rect 681094 933943 681150 933952
rect 679806 931560 679862 931569
rect 679806 931495 679862 931504
rect 679622 931152 679678 931161
rect 679622 931087 679678 931096
rect 676218 930336 676274 930345
rect 676218 930271 676220 930280
rect 676272 930271 676274 930280
rect 676220 930242 676272 930248
rect 674746 930200 674802 930209
rect 674746 930135 674802 930144
rect 683118 929520 683174 929529
rect 683118 929455 683174 929464
rect 683132 928713 683160 929455
rect 683118 928704 683174 928713
rect 683118 928639 683174 928648
rect 683132 927450 683160 928639
rect 683120 927444 683172 927450
rect 683120 927386 683172 927392
rect 675300 879096 675352 879102
rect 675300 879038 675352 879044
rect 675312 877418 675340 879038
rect 675404 877418 675432 877540
rect 675312 877390 675432 877418
rect 675772 876625 675800 876860
rect 675758 876616 675814 876625
rect 675758 876551 675814 876560
rect 675298 876480 675354 876489
rect 675298 876415 675354 876424
rect 675312 876262 675340 876415
rect 675312 876234 675418 876262
rect 675772 874177 675800 874412
rect 675758 874168 675814 874177
rect 675758 874103 675814 874112
rect 675404 873594 675432 873868
rect 675392 873588 675444 873594
rect 675392 873530 675444 873536
rect 675772 872817 675800 873188
rect 675758 872808 675814 872817
rect 675758 872743 675814 872752
rect 675404 872273 675432 872576
rect 675390 872264 675446 872273
rect 675390 872199 675446 872208
rect 675404 869854 675432 870060
rect 675392 869848 675444 869854
rect 675392 869790 675444 869796
rect 675392 869644 675444 869650
rect 675392 869586 675444 869592
rect 675404 869516 675432 869586
rect 675392 869032 675444 869038
rect 675392 868974 675444 868980
rect 675404 868875 675432 868974
rect 674932 868692 674984 868698
rect 674932 868634 674984 868640
rect 674944 866250 674972 868634
rect 675404 868086 675432 868224
rect 675392 868080 675444 868086
rect 675392 868022 675444 868028
rect 675404 866862 675432 867035
rect 675392 866856 675444 866862
rect 675392 866798 675444 866804
rect 674932 866244 674984 866250
rect 674932 866186 674984 866192
rect 675392 866244 675444 866250
rect 675392 866186 675444 866192
rect 675404 865844 675432 866186
rect 675772 864793 675800 865195
rect 675758 864784 675814 864793
rect 675758 864719 675814 864728
rect 675496 862850 675524 863328
rect 675484 862844 675536 862850
rect 675484 862786 675536 862792
rect 675404 788089 675432 788324
rect 675390 788080 675446 788089
rect 675390 788015 675446 788024
rect 675404 787370 675432 787679
rect 675392 787364 675444 787370
rect 675392 787306 675444 787312
rect 675772 786729 675800 787032
rect 675758 786720 675814 786729
rect 675758 786655 675814 786664
rect 675496 784825 675524 785196
rect 675482 784816 675538 784825
rect 675482 784751 675538 784760
rect 675404 784310 675432 784652
rect 675392 784304 675444 784310
rect 675392 784246 675444 784252
rect 675758 784136 675814 784145
rect 675758 784071 675814 784080
rect 675772 783972 675800 784071
rect 675496 782950 675524 783360
rect 675484 782944 675536 782950
rect 675484 782886 675536 782892
rect 675496 780774 675524 780844
rect 675484 780768 675536 780774
rect 675484 780710 675536 780716
rect 675496 780026 675524 780300
rect 675484 780020 675536 780026
rect 675484 779962 675536 779968
rect 675404 779346 675432 779688
rect 675392 779340 675444 779346
rect 675392 779282 675444 779288
rect 674748 779000 674800 779006
rect 674748 778942 674800 778948
rect 674760 777102 674788 778942
rect 675496 778666 675524 779008
rect 675484 778660 675536 778666
rect 675484 778602 675536 778608
rect 675404 777374 675432 777852
rect 675392 777368 675444 777374
rect 675392 777310 675444 777316
rect 674748 777096 674800 777102
rect 674748 777038 674800 777044
rect 675392 777096 675444 777102
rect 675392 777038 675444 777044
rect 675404 776628 675432 777038
rect 675404 775606 675432 776016
rect 675392 775600 675444 775606
rect 675392 775542 675444 775548
rect 675206 773936 675262 773945
rect 675206 773871 675262 773880
rect 675220 766630 675248 773871
rect 675496 773634 675524 774180
rect 675484 773628 675536 773634
rect 675484 773570 675536 773576
rect 675482 773392 675538 773401
rect 675482 773327 675538 773336
rect 675666 773392 675722 773401
rect 675666 773327 675722 773336
rect 675208 766624 675260 766630
rect 675496 766601 675524 773327
rect 675680 770054 675708 773327
rect 677414 773120 677470 773129
rect 677414 773055 677470 773064
rect 675588 770026 675708 770054
rect 675208 766566 675260 766572
rect 675482 766592 675538 766601
rect 675482 766527 675538 766536
rect 675588 765105 675616 770026
rect 675668 766624 675720 766630
rect 675666 766592 675668 766601
rect 675720 766592 675722 766601
rect 675666 766527 675722 766536
rect 675574 765096 675630 765105
rect 675574 765031 675630 765040
rect 676126 761288 676182 761297
rect 676126 761223 676182 761232
rect 676034 760744 676090 760753
rect 676140 760714 676168 761223
rect 676218 760880 676274 760889
rect 676218 760815 676220 760824
rect 676272 760815 676274 760824
rect 676220 760786 676272 760792
rect 676034 760679 676090 760688
rect 676128 760708 676180 760714
rect 676048 760578 676076 760679
rect 676128 760650 676180 760656
rect 676036 760572 676088 760578
rect 676036 760514 676088 760520
rect 676218 760064 676274 760073
rect 676218 759999 676274 760008
rect 674746 759928 674802 759937
rect 674746 759863 674802 759872
rect 674654 759112 674710 759121
rect 674654 759047 674710 759056
rect 674564 751936 674616 751942
rect 674564 751878 674616 751884
rect 674380 735684 674432 735690
rect 674380 735626 674432 735632
rect 674288 709640 674340 709646
rect 674288 709582 674340 709588
rect 674196 709232 674248 709238
rect 674196 709174 674248 709180
rect 674012 707600 674064 707606
rect 674012 707542 674064 707548
rect 674012 690056 674064 690062
rect 674012 689998 674064 690004
rect 673920 684276 673972 684282
rect 673920 684218 673972 684224
rect 673828 669520 673880 669526
rect 673828 669462 673880 669468
rect 673828 667276 673880 667282
rect 673828 667218 673880 667224
rect 673644 662380 673696 662386
rect 673644 662322 673696 662328
rect 673736 645448 673788 645454
rect 673736 645390 673788 645396
rect 673552 617432 673604 617438
rect 673552 617374 673604 617380
rect 673552 603084 673604 603090
rect 673552 603026 673604 603032
rect 673460 578196 673512 578202
rect 673460 578138 673512 578144
rect 673368 528828 673420 528834
rect 673368 528770 673420 528776
rect 673564 527134 673592 603026
rect 673644 576972 673696 576978
rect 673644 576914 673696 576920
rect 673656 532710 673684 576914
rect 673748 575006 673776 645390
rect 673840 622878 673868 667218
rect 673828 622872 673880 622878
rect 673828 622814 673880 622820
rect 673828 622260 673880 622266
rect 673828 622202 673880 622208
rect 673840 577454 673868 622202
rect 673932 619886 673960 684218
rect 673920 619880 673972 619886
rect 673920 619822 673972 619828
rect 674024 617030 674052 689998
rect 674196 688764 674248 688770
rect 674196 688706 674248 688712
rect 674208 683114 674236 688706
rect 674288 688696 674340 688702
rect 674288 688638 674340 688644
rect 674300 687070 674328 688638
rect 674288 687064 674340 687070
rect 674288 687006 674340 687012
rect 674208 683086 674328 683114
rect 674196 659728 674248 659734
rect 674196 659670 674248 659676
rect 674012 617024 674064 617030
rect 674012 616966 674064 616972
rect 674012 598460 674064 598466
rect 674012 598402 674064 598408
rect 673920 577652 673972 577658
rect 673920 577594 673972 577600
rect 673828 577448 673880 577454
rect 673828 577390 673880 577396
rect 673736 575000 673788 575006
rect 673736 574942 673788 574948
rect 673932 533322 673960 577594
rect 673920 533316 673972 533322
rect 673920 533258 673972 533264
rect 673644 532704 673696 532710
rect 673644 532646 673696 532652
rect 673552 527128 673604 527134
rect 673552 527070 673604 527076
rect 674024 526590 674052 598402
rect 674012 526584 674064 526590
rect 674012 526526 674064 526532
rect 673276 484832 673328 484838
rect 673276 484774 673328 484780
rect 673184 483200 673236 483206
rect 673184 483142 673236 483148
rect 673092 482792 673144 482798
rect 673092 482734 673144 482740
rect 673276 401668 673328 401674
rect 673276 401610 673328 401616
rect 673184 393372 673236 393378
rect 673184 393314 673236 393320
rect 673196 376650 673224 393314
rect 673184 376644 673236 376650
rect 673184 376586 673236 376592
rect 673288 357542 673316 401610
rect 673368 400240 673420 400246
rect 673368 400182 673420 400188
rect 673276 357536 673328 357542
rect 673276 357478 673328 357484
rect 673276 357060 673328 357066
rect 673276 357002 673328 357008
rect 673000 356244 673052 356250
rect 673000 356186 673052 356192
rect 673012 310690 673040 356186
rect 673184 350600 673236 350606
rect 673184 350542 673236 350548
rect 673092 348900 673144 348906
rect 673092 348842 673144 348848
rect 673104 331634 673132 348842
rect 673092 331628 673144 331634
rect 673092 331570 673144 331576
rect 673196 328438 673224 350542
rect 673184 328432 673236 328438
rect 673184 328374 673236 328380
rect 673288 312186 673316 357002
rect 673380 356726 673408 400182
rect 673368 356720 673420 356726
rect 673368 356662 673420 356668
rect 673276 312180 673328 312186
rect 673276 312122 673328 312128
rect 673368 311908 673420 311914
rect 673368 311850 673420 311856
rect 673000 310684 673052 310690
rect 673000 310626 673052 310632
rect 673276 310548 673328 310554
rect 673276 310490 673328 310496
rect 673184 303816 673236 303822
rect 673184 303758 673236 303764
rect 673092 303748 673144 303754
rect 673092 303690 673144 303696
rect 673000 303680 673052 303686
rect 673000 303622 673052 303628
rect 673012 291106 673040 303622
rect 673000 291100 673052 291106
rect 673000 291042 673052 291048
rect 673104 287978 673132 303690
rect 673092 287972 673144 287978
rect 673092 287914 673144 287920
rect 673196 286618 673224 303758
rect 673184 286612 673236 286618
rect 673184 286554 673236 286560
rect 672816 284368 672868 284374
rect 672816 284310 672868 284316
rect 672724 173800 672776 173806
rect 672724 173742 672776 173748
rect 672828 132802 672856 284310
rect 673288 266490 673316 310490
rect 673380 266626 673408 311850
rect 674104 310616 674156 310622
rect 674104 310558 674156 310564
rect 673920 267028 673972 267034
rect 673920 266970 673972 266976
rect 673368 266620 673420 266626
rect 673368 266562 673420 266568
rect 673276 266484 673328 266490
rect 673276 266426 673328 266432
rect 673368 264988 673420 264994
rect 673368 264930 673420 264936
rect 673276 263628 673328 263634
rect 673276 263570 673328 263576
rect 673000 260908 673052 260914
rect 673000 260850 673052 260856
rect 673012 247042 673040 260850
rect 673184 258188 673236 258194
rect 673184 258130 673236 258136
rect 673092 258120 673144 258126
rect 673092 258062 673144 258068
rect 673000 247036 673052 247042
rect 673000 246978 673052 246984
rect 673104 241670 673132 258062
rect 673092 241664 673144 241670
rect 673092 241606 673144 241612
rect 673196 241126 673224 258130
rect 673184 241120 673236 241126
rect 673184 241062 673236 241068
rect 673288 219910 673316 263570
rect 673380 220726 673408 264930
rect 673932 222290 673960 266970
rect 674012 266076 674064 266082
rect 674012 266018 674064 266024
rect 673920 222284 673972 222290
rect 673920 222226 673972 222232
rect 674024 221542 674052 266018
rect 674012 221536 674064 221542
rect 674012 221478 674064 221484
rect 673368 220720 673420 220726
rect 673368 220662 673420 220668
rect 673276 219904 673328 219910
rect 673276 219846 673328 219852
rect 673368 219496 673420 219502
rect 673368 219438 673420 219444
rect 673000 216164 673052 216170
rect 673000 216106 673052 216112
rect 673012 201890 673040 216106
rect 673184 214124 673236 214130
rect 673184 214066 673236 214072
rect 673092 213716 673144 213722
rect 673092 213658 673144 213664
rect 673000 201884 673052 201890
rect 673000 201826 673052 201832
rect 673104 196586 673132 213658
rect 673196 197470 673224 214066
rect 673184 197464 673236 197470
rect 673184 197406 673236 197412
rect 673092 196580 673144 196586
rect 673092 196522 673144 196528
rect 672908 176724 672960 176730
rect 672908 176666 672960 176672
rect 672816 132796 672868 132802
rect 672816 132738 672868 132744
rect 672920 131442 672948 176666
rect 673184 176044 673236 176050
rect 673184 175986 673236 175992
rect 673000 169516 673052 169522
rect 673000 169458 673052 169464
rect 673012 155514 673040 169458
rect 673092 168632 673144 168638
rect 673092 168574 673144 168580
rect 673000 155508 673052 155514
rect 673000 155450 673052 155456
rect 673104 151434 673132 168574
rect 673092 151428 673144 151434
rect 673092 151370 673144 151376
rect 672908 131436 672960 131442
rect 672908 131378 672960 131384
rect 673196 131306 673224 175986
rect 673276 175228 673328 175234
rect 673276 175170 673328 175176
rect 673184 131300 673236 131306
rect 673184 131242 673236 131248
rect 673288 130014 673316 175170
rect 673380 174894 673408 219438
rect 673368 174888 673420 174894
rect 673368 174830 673420 174836
rect 674116 133074 674144 310558
rect 674208 168706 674236 659670
rect 674300 616758 674328 683086
rect 674392 665310 674420 735626
rect 674656 734868 674708 734874
rect 674656 734810 674708 734816
rect 674668 732086 674696 734810
rect 674656 732080 674708 732086
rect 674656 732022 674708 732028
rect 674656 728680 674708 728686
rect 674656 728622 674708 728628
rect 674564 713244 674616 713250
rect 674564 713186 674616 713192
rect 674472 694340 674524 694346
rect 674472 694282 674524 694288
rect 674380 665304 674432 665310
rect 674380 665246 674432 665252
rect 674380 649120 674432 649126
rect 674380 649062 674432 649068
rect 674288 616752 674340 616758
rect 674288 616694 674340 616700
rect 674288 599820 674340 599826
rect 674288 599762 674340 599768
rect 674300 526998 674328 599762
rect 674392 573782 674420 649062
rect 674484 619070 674512 694282
rect 674576 668574 674604 713186
rect 674564 668568 674616 668574
rect 674564 668510 674616 668516
rect 674668 665038 674696 728622
rect 674760 715329 674788 759863
rect 676232 759354 676260 759999
rect 676220 759348 676272 759354
rect 676220 759290 676272 759296
rect 676218 759248 676274 759257
rect 676218 759183 676220 759192
rect 676272 759183 676274 759192
rect 676220 759154 676272 759160
rect 676034 759112 676090 759121
rect 676034 759047 676036 759056
rect 676088 759047 676090 759056
rect 676036 759018 676088 759024
rect 676220 758872 676272 758878
rect 676218 758840 676220 758849
rect 676272 758840 676274 758849
rect 676218 758775 676274 758784
rect 676034 758296 676090 758305
rect 676034 758231 676036 758240
rect 676088 758231 676090 758240
rect 676036 758202 676088 758208
rect 677428 757217 677456 773055
rect 677506 772984 677562 772993
rect 677506 772919 677562 772928
rect 676218 757208 676274 757217
rect 676218 757143 676274 757152
rect 677414 757208 677470 757217
rect 677414 757143 677470 757152
rect 676232 756294 676260 757143
rect 676220 756288 676272 756294
rect 676220 756230 676272 756236
rect 676126 755984 676182 755993
rect 676126 755919 676182 755928
rect 676140 755002 676168 755919
rect 676220 755608 676272 755614
rect 676218 755576 676220 755585
rect 676272 755576 676274 755585
rect 676218 755511 676274 755520
rect 676218 755168 676274 755177
rect 676218 755103 676220 755112
rect 676272 755103 676274 755112
rect 676220 755074 676272 755080
rect 676128 754996 676180 755002
rect 676128 754938 676180 754944
rect 677520 754769 677548 772919
rect 681002 772712 681058 772721
rect 681002 772647 681058 772656
rect 681016 755993 681044 772647
rect 703694 762076 703722 762212
rect 704154 762076 704182 762212
rect 704614 762076 704642 762212
rect 705074 762076 705102 762212
rect 705534 762076 705562 762212
rect 705994 762076 706022 762212
rect 706454 762076 706482 762212
rect 706914 762076 706942 762212
rect 707374 762076 707402 762212
rect 707834 762076 707862 762212
rect 708294 762076 708322 762212
rect 708754 762076 708782 762212
rect 709214 762076 709242 762212
rect 681002 755984 681058 755993
rect 681002 755919 681058 755928
rect 677506 754760 677562 754769
rect 677506 754695 677562 754704
rect 676218 753944 676274 753953
rect 676218 753879 676274 753888
rect 676232 753642 676260 753879
rect 676220 753636 676272 753642
rect 676220 753578 676272 753584
rect 676036 753432 676088 753438
rect 676034 753400 676036 753409
rect 676088 753400 676090 753409
rect 676034 753335 676090 753344
rect 676126 752720 676182 752729
rect 676126 752655 676182 752664
rect 676140 752282 676168 752655
rect 676220 752412 676272 752418
rect 676220 752354 676272 752360
rect 676232 752321 676260 752354
rect 676218 752312 676274 752321
rect 676128 752276 676180 752282
rect 676218 752247 676274 752256
rect 676128 752218 676180 752224
rect 676220 751936 676272 751942
rect 676218 751904 676220 751913
rect 676272 751904 676274 751913
rect 676218 751839 676274 751848
rect 683118 751088 683174 751097
rect 683118 751023 683174 751032
rect 683132 750281 683160 751023
rect 683118 750272 683174 750281
rect 683118 750207 683174 750216
rect 683132 749426 683160 750207
rect 683120 749420 683172 749426
rect 683120 749362 683172 749368
rect 675392 743776 675444 743782
rect 675392 743718 675444 743724
rect 675404 743308 675432 743718
rect 675404 742558 675432 742696
rect 675392 742552 675444 742558
rect 675392 742494 675444 742500
rect 675680 741713 675708 742016
rect 675666 741704 675722 741713
rect 675666 741639 675722 741648
rect 675404 739974 675432 740180
rect 674840 739968 674892 739974
rect 674840 739910 674892 739916
rect 675392 739968 675444 739974
rect 675392 739910 675444 739916
rect 674852 736137 674880 739910
rect 675404 739158 675432 739636
rect 675392 739152 675444 739158
rect 675392 739094 675444 739100
rect 675404 738682 675432 739024
rect 675392 738676 675444 738682
rect 675392 738618 675444 738624
rect 675404 738274 675432 738344
rect 675392 738268 675444 738274
rect 675392 738210 675444 738216
rect 674838 736128 674894 736137
rect 674838 736063 674894 736072
rect 675404 735690 675432 735896
rect 675392 735684 675444 735690
rect 675392 735626 675444 735632
rect 675404 735010 675432 735319
rect 675392 735004 675444 735010
rect 675392 734946 675444 734952
rect 675772 734369 675800 734672
rect 675758 734360 675814 734369
rect 675758 734295 675814 734304
rect 675404 733922 675432 734031
rect 675392 733916 675444 733922
rect 675392 733858 675444 733864
rect 675758 733000 675814 733009
rect 675758 732935 675814 732944
rect 675772 732836 675800 732935
rect 675392 732080 675444 732086
rect 675392 732022 675444 732028
rect 675404 731612 675432 732022
rect 675404 730522 675432 731000
rect 675392 730516 675444 730522
rect 675392 730458 675444 730464
rect 675496 728686 675524 729164
rect 675484 728680 675536 728686
rect 675484 728622 675536 728628
rect 675482 728376 675538 728385
rect 675482 728311 675538 728320
rect 675666 728376 675722 728385
rect 675666 728311 675722 728320
rect 675496 721565 675524 728311
rect 675680 721565 675708 728311
rect 678242 727288 678298 727297
rect 678242 727223 678298 727232
rect 675482 721556 675538 721565
rect 675482 721491 675538 721500
rect 675666 721556 675722 721565
rect 675666 721491 675722 721500
rect 676036 716576 676088 716582
rect 676034 716544 676036 716553
rect 676088 716544 676090 716553
rect 676034 716479 676090 716488
rect 676036 716168 676088 716174
rect 676034 716136 676036 716145
rect 676088 716136 676090 716145
rect 676034 716071 676090 716080
rect 676034 715728 676090 715737
rect 676034 715663 676090 715672
rect 674746 715320 674802 715329
rect 674746 715255 674802 715264
rect 676048 715018 676076 715663
rect 676036 715012 676088 715018
rect 676036 714954 676088 714960
rect 674746 714912 674802 714921
rect 674746 714847 674802 714856
rect 674760 670177 674788 714847
rect 676036 714536 676088 714542
rect 676034 714504 676036 714513
rect 676088 714504 676090 714513
rect 676034 714439 676090 714448
rect 676034 714096 676090 714105
rect 676034 714031 676036 714040
rect 676088 714031 676090 714040
rect 676036 714002 676088 714008
rect 676036 713720 676088 713726
rect 676034 713688 676036 713697
rect 676088 713688 676090 713697
rect 676034 713623 676090 713632
rect 676954 713488 677010 713497
rect 676954 713423 677010 713432
rect 676034 713280 676090 713289
rect 676034 713215 676036 713224
rect 676088 713215 676090 713224
rect 676036 713186 676088 713192
rect 676036 712904 676088 712910
rect 676034 712872 676036 712881
rect 676088 712872 676090 712881
rect 676034 712807 676090 712816
rect 676034 712464 676090 712473
rect 676034 712399 676036 712408
rect 676088 712399 676090 712408
rect 676036 712370 676088 712376
rect 676036 711680 676088 711686
rect 676034 711648 676036 711657
rect 676088 711648 676090 711657
rect 676034 711583 676090 711592
rect 676036 710456 676088 710462
rect 676034 710424 676036 710433
rect 676088 710424 676090 710433
rect 676034 710359 676090 710368
rect 676036 710048 676088 710054
rect 676034 710016 676036 710025
rect 676088 710016 676090 710025
rect 676034 709951 676090 709960
rect 676036 709640 676088 709646
rect 676034 709608 676036 709617
rect 676088 709608 676090 709617
rect 676034 709543 676090 709552
rect 676036 709232 676088 709238
rect 676034 709200 676036 709209
rect 676088 709200 676090 709209
rect 676034 709135 676090 709144
rect 676968 709102 676996 713423
rect 678256 712065 678284 727223
rect 681002 726608 681058 726617
rect 681002 726543 681058 726552
rect 679622 724432 679678 724441
rect 679622 724367 679678 724376
rect 678242 712056 678298 712065
rect 678242 711991 678298 712000
rect 679636 711249 679664 724367
rect 679622 711240 679678 711249
rect 679622 711175 679678 711184
rect 681016 710841 681044 726543
rect 703694 717196 703722 717264
rect 704154 717196 704182 717264
rect 704614 717196 704642 717264
rect 705074 717196 705102 717264
rect 705534 717196 705562 717264
rect 705994 717196 706022 717264
rect 706454 717196 706482 717264
rect 706914 717196 706942 717264
rect 707374 717196 707402 717264
rect 707834 717196 707862 717264
rect 708294 717196 708322 717264
rect 708754 717196 708782 717264
rect 709214 717196 709242 717264
rect 681002 710832 681058 710841
rect 681002 710767 681058 710776
rect 676036 709096 676088 709102
rect 676036 709038 676088 709044
rect 676956 709096 677008 709102
rect 676956 709038 677008 709044
rect 676048 708801 676076 709038
rect 676034 708792 676090 708801
rect 676034 708727 676090 708736
rect 676036 708416 676088 708422
rect 676034 708384 676036 708393
rect 676088 708384 676090 708393
rect 676034 708319 676090 708328
rect 676036 708008 676088 708014
rect 676034 707976 676036 707985
rect 676088 707976 676090 707985
rect 676034 707911 676090 707920
rect 676036 707600 676088 707606
rect 676034 707568 676036 707577
rect 676088 707568 676090 707577
rect 676034 707503 676090 707512
rect 676034 707160 676090 707169
rect 676034 707095 676090 707104
rect 675944 706784 675996 706790
rect 675942 706752 675944 706761
rect 675996 706752 675998 706761
rect 676048 706722 676076 707095
rect 675942 706687 675998 706696
rect 676036 706716 676088 706722
rect 676036 706658 676088 706664
rect 676034 706344 676090 706353
rect 676034 706279 676090 706288
rect 676048 705129 676076 706279
rect 676034 705120 676090 705129
rect 676034 705055 676090 705064
rect 676048 703866 676076 705055
rect 676036 703860 676088 703866
rect 676036 703802 676088 703808
rect 675404 698222 675432 698323
rect 675392 698216 675444 698222
rect 675392 698158 675444 698164
rect 675404 697406 675432 697680
rect 675392 697400 675444 697406
rect 675392 697342 675444 697348
rect 675404 696969 675432 697035
rect 675390 696960 675446 696969
rect 675390 696895 675446 696904
rect 675496 694793 675524 695195
rect 675482 694784 675538 694793
rect 675482 694719 675538 694728
rect 675496 694346 675524 694620
rect 675484 694340 675536 694346
rect 675484 694282 675536 694288
rect 675758 694240 675814 694249
rect 675758 694175 675814 694184
rect 675772 694008 675800 694175
rect 675496 693054 675524 693328
rect 675484 693048 675536 693054
rect 675484 692990 675536 692996
rect 675404 690470 675432 690880
rect 675392 690464 675444 690470
rect 675392 690406 675444 690412
rect 675404 690062 675432 690336
rect 675392 690056 675444 690062
rect 675392 689998 675444 690004
rect 675496 689382 675524 689656
rect 675484 689376 675536 689382
rect 675484 689318 675536 689324
rect 675404 688770 675432 689044
rect 675392 688764 675444 688770
rect 675392 688706 675444 688712
rect 675772 687449 675800 687820
rect 675758 687440 675814 687449
rect 675758 687375 675814 687384
rect 675484 687064 675536 687070
rect 675484 687006 675536 687012
rect 675496 686664 675524 687006
rect 675666 686216 675722 686225
rect 675666 686151 675722 686160
rect 675680 685984 675708 686151
rect 675392 684276 675444 684282
rect 675392 684218 675444 684224
rect 675404 684148 675432 684218
rect 675390 683360 675446 683369
rect 675390 683295 675446 683304
rect 675758 683360 675814 683369
rect 675758 683295 675814 683304
rect 675404 676433 675432 683295
rect 675482 683224 675538 683233
rect 675482 683159 675538 683168
rect 675390 676424 675446 676433
rect 675390 676359 675446 676368
rect 674746 670168 674802 670177
rect 674746 670103 674802 670112
rect 674746 668128 674802 668137
rect 674746 668063 674802 668072
rect 674656 665032 674708 665038
rect 674656 664974 674708 664980
rect 674656 652180 674708 652186
rect 674656 652122 674708 652128
rect 674564 643748 674616 643754
rect 674564 643690 674616 643696
rect 674576 641918 674604 643690
rect 674564 641912 674616 641918
rect 674564 641854 674616 641860
rect 674472 619064 674524 619070
rect 674472 619006 674524 619012
rect 674472 604376 674524 604382
rect 674472 604318 674524 604324
rect 674380 573776 674432 573782
rect 674380 573718 674432 573724
rect 674380 553444 674432 553450
rect 674380 553386 674432 553392
rect 674392 548049 674420 553386
rect 674378 548040 674434 548049
rect 674378 547975 674434 547984
rect 674380 547936 674432 547942
rect 674380 547878 674432 547884
rect 674288 526992 674340 526998
rect 674288 526934 674340 526940
rect 674392 486062 674420 547878
rect 674484 529038 674512 604318
rect 674564 603288 674616 603294
rect 674564 603230 674616 603236
rect 674472 529032 674524 529038
rect 674472 528974 674524 528980
rect 674576 528426 674604 603230
rect 674668 574190 674696 652122
rect 674760 623694 674788 668063
rect 675496 653818 675524 683159
rect 675772 676433 675800 683295
rect 676494 683088 676550 683097
rect 676494 683023 676550 683032
rect 676508 676433 676536 683023
rect 679622 681864 679678 681873
rect 679622 681799 679678 681808
rect 675758 676424 675814 676433
rect 675758 676359 675814 676368
rect 676494 676424 676550 676433
rect 676494 676359 676550 676368
rect 676218 671120 676274 671129
rect 676218 671055 676274 671064
rect 676034 670984 676090 670993
rect 676034 670919 676036 670928
rect 676088 670919 676090 670928
rect 676036 670890 676088 670896
rect 676232 670818 676260 671055
rect 676220 670812 676272 670818
rect 676220 670754 676272 670760
rect 676126 670304 676182 670313
rect 676126 670239 676182 670248
rect 676036 669520 676088 669526
rect 676036 669462 676088 669468
rect 676048 669361 676076 669462
rect 676140 669458 676168 670239
rect 676218 669488 676274 669497
rect 676128 669452 676180 669458
rect 676218 669423 676274 669432
rect 676128 669394 676180 669400
rect 676232 669390 676260 669423
rect 676220 669384 676272 669390
rect 676034 669352 676090 669361
rect 676220 669326 676272 669332
rect 676034 669287 676090 669296
rect 676218 668672 676274 668681
rect 676218 668607 676274 668616
rect 676036 668568 676088 668574
rect 676034 668536 676036 668545
rect 676088 668536 676090 668545
rect 676034 668471 676090 668480
rect 676232 667962 676260 668607
rect 676220 667956 676272 667962
rect 676220 667898 676272 667904
rect 676218 667448 676274 667457
rect 676218 667383 676274 667392
rect 676034 667312 676090 667321
rect 676034 667247 676036 667256
rect 676088 667247 676090 667256
rect 676036 667218 676088 667224
rect 676232 666738 676260 667383
rect 679636 667049 679664 681799
rect 679714 678328 679770 678337
rect 679714 678263 679770 678272
rect 679622 667040 679678 667049
rect 679622 666975 679678 666984
rect 676220 666732 676272 666738
rect 676220 666674 676272 666680
rect 676126 666224 676182 666233
rect 676126 666159 676182 666168
rect 676140 665514 676168 666159
rect 679728 665825 679756 678263
rect 703694 671908 703722 672044
rect 704154 671908 704182 672044
rect 704614 671908 704642 672044
rect 705074 671908 705102 672044
rect 705534 671908 705562 672044
rect 705994 671908 706022 672044
rect 706454 671908 706482 672044
rect 706914 671908 706942 672044
rect 707374 671908 707402 672044
rect 707834 671908 707862 672044
rect 708294 671908 708322 672044
rect 708754 671908 708782 672044
rect 709214 671908 709242 672044
rect 676218 665816 676274 665825
rect 676218 665751 676274 665760
rect 679714 665816 679770 665825
rect 679714 665751 679770 665760
rect 676128 665508 676180 665514
rect 676128 665450 676180 665456
rect 676232 665378 676260 665751
rect 676220 665372 676272 665378
rect 676220 665314 676272 665320
rect 676036 665304 676088 665310
rect 676034 665272 676036 665281
rect 676088 665272 676090 665281
rect 676034 665207 676090 665216
rect 676220 665032 676272 665038
rect 676218 665000 676220 665009
rect 676272 665000 676274 665009
rect 676218 664935 676274 664944
rect 676218 664184 676274 664193
rect 676218 664119 676274 664128
rect 676232 664018 676260 664119
rect 676220 664012 676272 664018
rect 676220 663954 676272 663960
rect 676220 663808 676272 663814
rect 676218 663776 676220 663785
rect 676272 663776 676274 663785
rect 676218 663711 676274 663720
rect 676218 663368 676274 663377
rect 676218 663303 676274 663312
rect 676232 662454 676260 663303
rect 676220 662448 676272 662454
rect 676034 662416 676090 662425
rect 676220 662390 676272 662396
rect 676034 662351 676036 662360
rect 676088 662351 676090 662360
rect 676036 662322 676088 662328
rect 676218 661736 676274 661745
rect 676218 661671 676274 661680
rect 676126 661328 676182 661337
rect 676232 661298 676260 661671
rect 676126 661263 676182 661272
rect 676220 661292 676272 661298
rect 676140 661162 676168 661263
rect 676220 661234 676272 661240
rect 676128 661156 676180 661162
rect 676128 661098 676180 661104
rect 683118 660920 683174 660929
rect 683118 660855 683174 660864
rect 683132 660113 683160 660855
rect 683118 660104 683174 660113
rect 683118 660039 683174 660048
rect 683132 659734 683160 660039
rect 683120 659728 683172 659734
rect 683120 659670 683172 659676
rect 675208 653812 675260 653818
rect 675208 653754 675260 653760
rect 675484 653812 675536 653818
rect 675484 653754 675536 653760
rect 675220 645969 675248 653754
rect 675404 652798 675432 653140
rect 675392 652792 675444 652798
rect 675392 652734 675444 652740
rect 675496 652186 675524 652460
rect 675484 652180 675536 652186
rect 675484 652122 675536 652128
rect 675404 651574 675432 651848
rect 675392 651568 675444 651574
rect 675392 651510 675444 651516
rect 675404 649913 675432 650012
rect 675390 649904 675446 649913
rect 675390 649839 675446 649848
rect 675404 649126 675432 649468
rect 675392 649120 675444 649126
rect 675392 649062 675444 649068
rect 675772 648689 675800 648788
rect 675758 648680 675814 648689
rect 675758 648615 675814 648624
rect 675496 647766 675524 648176
rect 675484 647760 675536 647766
rect 675484 647702 675536 647708
rect 675206 645960 675262 645969
rect 675206 645895 675262 645904
rect 675404 645454 675432 645660
rect 675392 645448 675444 645454
rect 675392 645390 675444 645396
rect 675404 645046 675432 645116
rect 675392 645040 675444 645046
rect 675392 644982 675444 644988
rect 675758 644736 675814 644745
rect 675758 644671 675814 644680
rect 675772 644475 675800 644671
rect 675404 643414 675432 643824
rect 675392 643408 675444 643414
rect 675392 643350 675444 643356
rect 675666 643104 675722 643113
rect 675666 643039 675722 643048
rect 675680 642635 675708 643039
rect 675392 641912 675444 641918
rect 675392 641854 675444 641860
rect 675404 641444 675432 641854
rect 675404 640354 675432 640795
rect 675392 640348 675444 640354
rect 675392 640290 675444 640296
rect 675392 639124 675444 639130
rect 675392 639066 675444 639072
rect 675404 638928 675432 639066
rect 675206 638752 675262 638761
rect 675206 638687 675262 638696
rect 675220 631417 675248 638687
rect 675482 638208 675538 638217
rect 675482 638143 675538 638152
rect 675496 633826 675524 638143
rect 676862 637936 676918 637945
rect 676862 637871 676918 637880
rect 677506 637936 677562 637945
rect 677506 637871 677562 637880
rect 675484 633820 675536 633826
rect 675484 633762 675536 633768
rect 676876 631417 676904 637871
rect 675206 631408 675262 631417
rect 675206 631343 675262 631352
rect 676862 631408 676918 631417
rect 676862 631343 676918 631352
rect 676126 626104 676182 626113
rect 676126 626039 676182 626048
rect 676140 625530 676168 626039
rect 676218 625696 676274 625705
rect 676218 625631 676274 625640
rect 676128 625524 676180 625530
rect 676128 625466 676180 625472
rect 676232 625394 676260 625631
rect 676220 625388 676272 625394
rect 676220 625330 676272 625336
rect 676218 625288 676274 625297
rect 676218 625223 676274 625232
rect 676232 625190 676260 625223
rect 676220 625184 676272 625190
rect 676220 625126 676272 625132
rect 676218 624880 676274 624889
rect 676218 624815 676274 624824
rect 676126 624472 676182 624481
rect 676126 624407 676182 624416
rect 676034 623928 676090 623937
rect 676140 623898 676168 624407
rect 676232 624170 676260 624815
rect 676220 624164 676272 624170
rect 676220 624106 676272 624112
rect 676218 624064 676274 624073
rect 676218 623999 676274 624008
rect 676232 623966 676260 623999
rect 676220 623960 676272 623966
rect 676220 623902 676272 623908
rect 676034 623863 676090 623872
rect 676128 623892 676180 623898
rect 676048 623830 676076 623863
rect 676128 623834 676180 623840
rect 676036 623824 676088 623830
rect 676036 623766 676088 623772
rect 674748 623688 674800 623694
rect 676220 623688 676272 623694
rect 674748 623630 674800 623636
rect 676218 623656 676220 623665
rect 676272 623656 676274 623665
rect 676218 623591 676274 623600
rect 676034 623112 676090 623121
rect 676034 623047 676036 623056
rect 676088 623047 676090 623056
rect 676036 623018 676088 623024
rect 676220 622872 676272 622878
rect 676218 622840 676220 622849
rect 676272 622840 676274 622849
rect 676218 622775 676274 622784
rect 676034 622296 676090 622305
rect 676034 622231 676036 622240
rect 676088 622231 676090 622240
rect 676036 622202 676088 622208
rect 676218 621208 676274 621217
rect 676218 621143 676220 621152
rect 676272 621143 676274 621152
rect 676220 621114 676272 621120
rect 676218 619984 676274 619993
rect 676218 619919 676274 619928
rect 676036 619880 676088 619886
rect 676034 619848 676036 619857
rect 676088 619848 676090 619857
rect 676232 619818 676260 619919
rect 676034 619783 676090 619792
rect 676220 619812 676272 619818
rect 676220 619754 676272 619760
rect 676218 619168 676274 619177
rect 676218 619103 676274 619112
rect 676036 619064 676088 619070
rect 676034 619032 676036 619041
rect 676088 619032 676090 619041
rect 676034 618967 676090 618976
rect 676232 618458 676260 619103
rect 677520 618769 677548 637871
rect 681002 637528 681058 637537
rect 681002 637463 681058 637472
rect 679622 637392 679678 637401
rect 679622 637327 679678 637336
rect 679636 622033 679664 637327
rect 679622 622024 679678 622033
rect 679622 621959 679678 621968
rect 681016 620809 681044 637463
rect 681096 633820 681148 633826
rect 681096 633762 681148 633768
rect 681108 621625 681136 633762
rect 703694 626892 703722 627028
rect 704154 626892 704182 627028
rect 704614 626892 704642 627028
rect 705074 626892 705102 627028
rect 705534 626892 705562 627028
rect 705994 626892 706022 627028
rect 706454 626892 706482 627028
rect 706914 626892 706942 627028
rect 707374 626892 707402 627028
rect 707834 626892 707862 627028
rect 708294 626892 708322 627028
rect 708754 626892 708782 627028
rect 709214 626892 709242 627028
rect 681094 621616 681150 621625
rect 681094 621551 681150 621560
rect 681002 620800 681058 620809
rect 681002 620735 681058 620744
rect 677506 618760 677562 618769
rect 677506 618695 677562 618704
rect 676220 618452 676272 618458
rect 676220 618394 676272 618400
rect 676218 617536 676274 617545
rect 676218 617471 676274 617480
rect 676036 617432 676088 617438
rect 676034 617400 676036 617409
rect 676088 617400 676090 617409
rect 676034 617335 676090 617344
rect 676036 617024 676088 617030
rect 676034 616992 676036 617001
rect 676088 616992 676090 617001
rect 676034 616927 676090 616936
rect 676232 616894 676260 617471
rect 676220 616888 676272 616894
rect 676220 616830 676272 616836
rect 676220 616752 676272 616758
rect 676218 616720 676220 616729
rect 676272 616720 676274 616729
rect 676218 616655 676274 616664
rect 683118 615904 683174 615913
rect 683118 615839 683174 615848
rect 683132 615097 683160 615839
rect 683118 615088 683174 615097
rect 683118 615023 683174 615032
rect 683132 614174 683160 615023
rect 683120 614168 683172 614174
rect 683120 614110 683172 614116
rect 675404 608054 675432 608124
rect 675392 608048 675444 608054
rect 675392 607990 675444 607996
rect 675392 607640 675444 607646
rect 675392 607582 675444 607588
rect 675404 607479 675432 607582
rect 675404 606529 675432 606832
rect 675390 606520 675446 606529
rect 675390 606455 675446 606464
rect 675404 604586 675432 604996
rect 675208 604580 675260 604586
rect 675208 604522 675260 604528
rect 675392 604580 675444 604586
rect 675392 604522 675444 604528
rect 675220 600953 675248 604522
rect 675404 604382 675432 604452
rect 675392 604376 675444 604382
rect 675392 604318 675444 604324
rect 675496 603294 675524 603772
rect 675484 603288 675536 603294
rect 675484 603230 675536 603236
rect 675404 603090 675432 603160
rect 675392 603084 675444 603090
rect 675392 603026 675444 603032
rect 675206 600944 675262 600953
rect 675206 600879 675262 600888
rect 675496 600438 675524 600644
rect 675484 600432 675536 600438
rect 675484 600374 675536 600380
rect 675496 599826 675524 600100
rect 675484 599820 675536 599826
rect 675484 599762 675536 599768
rect 674748 599616 674800 599622
rect 674748 599558 674800 599564
rect 674760 596902 674788 599558
rect 675772 599049 675800 599488
rect 675758 599040 675814 599049
rect 675758 598975 675814 598984
rect 675496 598466 675524 598808
rect 675484 598460 675536 598466
rect 675484 598402 675536 598408
rect 675484 597780 675536 597786
rect 675484 597722 675536 597728
rect 675496 597652 675524 597722
rect 674748 596896 674800 596902
rect 674748 596838 674800 596844
rect 675392 596896 675444 596902
rect 675392 596838 675444 596844
rect 675404 596428 675432 596838
rect 675588 595377 675616 595816
rect 675574 595368 675630 595377
rect 675574 595303 675630 595312
rect 675496 593434 675524 593980
rect 675484 593428 675536 593434
rect 675484 593370 675536 593376
rect 675758 593192 675814 593201
rect 675758 593127 675814 593136
rect 675574 593056 675630 593065
rect 675574 592991 675630 593000
rect 675482 592104 675538 592113
rect 675482 592039 675538 592048
rect 675496 584633 675524 592039
rect 675588 586265 675616 592991
rect 675772 586514 675800 593127
rect 677506 592104 677562 592113
rect 677506 592039 677562 592048
rect 675772 586486 675892 586514
rect 675864 586265 675892 586486
rect 675574 586256 675630 586265
rect 675574 586191 675630 586200
rect 675850 586256 675906 586265
rect 675850 586191 675906 586200
rect 675482 584624 675538 584633
rect 675482 584559 675538 584568
rect 676034 581088 676090 581097
rect 676034 581023 676036 581032
rect 676088 581023 676090 581032
rect 676036 580994 676088 581000
rect 676126 580544 676182 580553
rect 676126 580479 676182 580488
rect 676034 580272 676090 580281
rect 676034 580207 676090 580216
rect 676048 579834 676076 580207
rect 676140 579970 676168 580479
rect 676218 580136 676274 580145
rect 676218 580071 676220 580080
rect 676272 580071 676274 580080
rect 676220 580042 676272 580048
rect 676128 579964 676180 579970
rect 676128 579906 676180 579912
rect 676036 579828 676088 579834
rect 676036 579770 676088 579776
rect 676310 579320 676366 579329
rect 676310 579255 676366 579264
rect 676218 578912 676274 578921
rect 676218 578847 676274 578856
rect 676126 578504 676182 578513
rect 676232 578474 676260 578847
rect 676126 578439 676182 578448
rect 676220 578468 676272 578474
rect 676140 578270 676168 578439
rect 676220 578410 676272 578416
rect 676324 578338 676352 579255
rect 676312 578332 676364 578338
rect 676312 578274 676364 578280
rect 676128 578264 676180 578270
rect 676034 578232 676090 578241
rect 676128 578206 676180 578212
rect 676034 578167 676036 578176
rect 676088 578167 676090 578176
rect 676036 578138 676088 578144
rect 676218 577688 676274 577697
rect 676218 577623 676220 577632
rect 676272 577623 676274 577632
rect 676220 577594 676272 577600
rect 676036 577448 676088 577454
rect 676034 577416 676036 577425
rect 676088 577416 676090 577425
rect 676034 577351 676090 577360
rect 676034 577008 676090 577017
rect 676034 576943 676036 576952
rect 676088 576943 676090 576952
rect 676036 576914 676088 576920
rect 676126 576464 676182 576473
rect 676126 576399 676182 576408
rect 676036 575884 676088 575890
rect 676036 575826 676088 575832
rect 676048 575793 676076 575826
rect 676034 575784 676090 575793
rect 676140 575754 676168 576399
rect 676218 576056 676274 576065
rect 676218 575991 676274 576000
rect 676034 575719 676090 575728
rect 676128 575748 676180 575754
rect 676128 575690 676180 575696
rect 676232 575618 676260 575991
rect 676220 575612 676272 575618
rect 676220 575554 676272 575560
rect 676036 575000 676088 575006
rect 676034 574968 676036 574977
rect 676088 574968 676090 574977
rect 676034 574903 676090 574912
rect 676218 574424 676274 574433
rect 676218 574359 676274 574368
rect 676232 574258 676260 574359
rect 676220 574252 676272 574258
rect 676220 574194 676272 574200
rect 674656 574184 674708 574190
rect 676036 574184 676088 574190
rect 674656 574126 674708 574132
rect 676034 574152 676036 574161
rect 676088 574152 676090 574161
rect 676034 574087 676090 574096
rect 676036 573776 676088 573782
rect 676034 573744 676036 573753
rect 676088 573744 676090 573753
rect 676034 573679 676090 573688
rect 677520 573617 677548 592039
rect 682382 591424 682438 591433
rect 682382 591359 682438 591368
rect 682396 575657 682424 591359
rect 703694 581740 703722 581876
rect 704154 581740 704182 581876
rect 704614 581740 704642 581876
rect 705074 581740 705102 581876
rect 705534 581740 705562 581876
rect 705994 581740 706022 581876
rect 706454 581740 706482 581876
rect 706914 581740 706942 581876
rect 707374 581740 707402 581876
rect 707834 581740 707862 581876
rect 708294 581740 708322 581876
rect 708754 581740 708782 581876
rect 709214 581740 709242 581876
rect 682382 575648 682438 575657
rect 682382 575583 682438 575592
rect 677506 573608 677562 573617
rect 677506 573543 677562 573552
rect 676218 571976 676274 571985
rect 676218 571911 676274 571920
rect 676232 571674 676260 571911
rect 676220 571668 676272 571674
rect 676220 571610 676272 571616
rect 676218 571568 676274 571577
rect 676218 571503 676220 571512
rect 676272 571503 676274 571512
rect 676220 571474 676272 571480
rect 676218 571160 676274 571169
rect 676218 571095 676274 571104
rect 676232 569974 676260 571095
rect 683118 570752 683174 570761
rect 683118 570687 683174 570696
rect 676220 569968 676272 569974
rect 683132 569945 683160 570687
rect 676220 569910 676272 569916
rect 683118 569936 683174 569945
rect 683118 569871 683174 569880
rect 683132 568614 683160 569871
rect 683120 568608 683172 568614
rect 683120 568550 683172 568556
rect 675772 562737 675800 562904
rect 675758 562728 675814 562737
rect 675758 562663 675814 562672
rect 675404 561950 675432 562292
rect 675392 561944 675444 561950
rect 675392 561886 675444 561892
rect 675496 561241 675524 561612
rect 675482 561232 675538 561241
rect 675482 561167 675538 561176
rect 675588 559609 675616 559776
rect 675574 559600 675630 559609
rect 675574 559535 675630 559544
rect 675404 559162 675432 559232
rect 675392 559156 675444 559162
rect 675392 559098 675444 559104
rect 675758 558920 675814 558929
rect 675758 558855 675814 558864
rect 675772 558620 675800 558855
rect 675496 557598 675524 557940
rect 675484 557592 675536 557598
rect 675484 557534 675536 557540
rect 675404 555286 675432 555492
rect 674748 555280 674800 555286
rect 674748 555222 674800 555228
rect 675392 555280 675444 555286
rect 675392 555222 675444 555228
rect 674656 549364 674708 549370
rect 674656 549306 674708 549312
rect 674668 548010 674696 549306
rect 674760 548486 674788 555222
rect 675312 554905 675418 554933
rect 674930 554840 674986 554849
rect 675312 554810 675340 554905
rect 674930 554775 674986 554784
rect 675300 554804 675352 554810
rect 674944 549370 674972 554775
rect 675300 554746 675352 554752
rect 675300 554056 675352 554062
rect 675772 554033 675800 554268
rect 675300 553998 675352 554004
rect 675758 554024 675814 554033
rect 675312 551253 675340 553998
rect 675758 553959 675814 553968
rect 675404 553450 675432 553656
rect 675392 553444 675444 553450
rect 675392 553386 675444 553392
rect 675772 551993 675800 552432
rect 675758 551984 675814 551993
rect 675758 551919 675814 551928
rect 675312 551225 675418 551253
rect 675312 550582 675418 550610
rect 675022 550352 675078 550361
rect 675022 550287 675078 550296
rect 674932 549364 674984 549370
rect 674932 549306 674984 549312
rect 674932 549228 674984 549234
rect 674932 549170 674984 549176
rect 674748 548480 674800 548486
rect 674748 548422 674800 548428
rect 674748 548344 674800 548350
rect 674748 548286 674800 548292
rect 674656 548004 674708 548010
rect 674656 547946 674708 547952
rect 674654 547904 674710 547913
rect 674654 547839 674710 547848
rect 674564 528420 674616 528426
rect 674564 528362 674616 528368
rect 674472 524476 674524 524482
rect 674472 524418 674524 524424
rect 674380 486056 674432 486062
rect 674380 485998 674432 486004
rect 674288 480276 674340 480282
rect 674288 480218 674340 480224
rect 674196 168700 674248 168706
rect 674196 168642 674248 168648
rect 674196 167068 674248 167074
rect 674196 167010 674248 167016
rect 674104 133068 674156 133074
rect 674104 133010 674156 133016
rect 673276 130008 673328 130014
rect 673276 129950 673328 129956
rect 672724 129872 672776 129878
rect 672724 129814 672776 129820
rect 672736 106146 672764 129814
rect 674208 114374 674236 167010
rect 674300 148442 674328 480218
rect 674484 475862 674512 524418
rect 674668 482361 674696 547839
rect 674760 485625 674788 548286
rect 674944 498302 674972 549170
rect 675036 500954 675064 550287
rect 675312 549234 675340 550582
rect 675300 549228 675352 549234
rect 675300 549170 675352 549176
rect 675312 548746 675418 548774
rect 675312 548350 675340 548746
rect 675300 548344 675352 548350
rect 675300 548286 675352 548292
rect 675760 548004 675812 548010
rect 675760 547946 675812 547952
rect 675024 500948 675076 500954
rect 675024 500890 675076 500896
rect 674932 498296 674984 498302
rect 674932 498238 674984 498244
rect 675772 498234 675800 547946
rect 678242 546816 678298 546825
rect 678242 546751 678298 546760
rect 677506 546544 677562 546553
rect 677506 546479 677562 546488
rect 676218 535936 676274 535945
rect 676218 535871 676274 535880
rect 676232 535770 676260 535871
rect 676220 535764 676272 535770
rect 676034 535732 676090 535741
rect 676220 535706 676272 535712
rect 676034 535667 676090 535676
rect 676048 535634 676076 535667
rect 676036 535628 676088 535634
rect 676036 535570 676088 535576
rect 676126 535120 676182 535129
rect 676126 535055 676182 535064
rect 675942 534508 675998 534517
rect 675942 534443 675998 534452
rect 675852 528420 675904 528426
rect 675850 528388 675852 528397
rect 675904 528388 675906 528397
rect 675850 528323 675906 528332
rect 675850 527164 675906 527173
rect 675850 527099 675852 527108
rect 675904 527099 675906 527108
rect 675852 527070 675904 527076
rect 675760 498228 675812 498234
rect 675760 498170 675812 498176
rect 675956 495258 675984 534443
rect 676140 534274 676168 535055
rect 676218 534712 676274 534721
rect 676218 534647 676274 534656
rect 676232 534546 676260 534647
rect 676220 534540 676272 534546
rect 676220 534482 676272 534488
rect 676220 534404 676272 534410
rect 676220 534346 676272 534352
rect 676232 534313 676260 534346
rect 676218 534304 676274 534313
rect 676128 534268 676180 534274
rect 676218 534239 676274 534248
rect 676128 534210 676180 534216
rect 676036 533316 676088 533322
rect 676034 533284 676036 533293
rect 676088 533284 676090 533293
rect 676034 533219 676090 533228
rect 676034 532876 676090 532885
rect 676034 532811 676090 532820
rect 675772 495230 675984 495258
rect 675772 490929 675800 495230
rect 675850 492144 675906 492153
rect 675850 492079 675906 492088
rect 675864 491706 675892 492079
rect 675942 491736 675998 491745
rect 675852 491700 675904 491706
rect 675942 491671 675998 491680
rect 675852 491642 675904 491648
rect 675956 491570 675984 491671
rect 675944 491564 675996 491570
rect 675944 491506 675996 491512
rect 675944 491428 675996 491434
rect 675944 491370 675996 491376
rect 675956 491337 675984 491370
rect 675942 491328 675998 491337
rect 675942 491263 675998 491272
rect 675758 490920 675814 490929
rect 675758 490855 675814 490864
rect 675942 490512 675998 490521
rect 675942 490447 675998 490456
rect 675956 490210 675984 490447
rect 675944 490204 675996 490210
rect 675944 490146 675996 490152
rect 675850 489696 675906 489705
rect 675850 489631 675906 489640
rect 675864 485774 675892 489631
rect 676048 489297 676076 532811
rect 676220 532704 676272 532710
rect 676218 532672 676220 532681
rect 676272 532672 676274 532681
rect 676218 532607 676274 532616
rect 677230 531856 677286 531865
rect 677230 531791 677286 531800
rect 676126 530632 676182 530641
rect 676126 530567 676182 530576
rect 676140 530058 676168 530567
rect 676218 530224 676274 530233
rect 676218 530159 676220 530168
rect 676272 530159 676274 530168
rect 676220 530130 676272 530136
rect 676128 530052 676180 530058
rect 676128 529994 676180 530000
rect 676126 529408 676182 529417
rect 676126 529343 676182 529352
rect 676140 528698 676168 529343
rect 676404 529032 676456 529038
rect 676218 529000 676274 529009
rect 676218 528935 676274 528944
rect 676402 529000 676404 529009
rect 676456 529000 676458 529009
rect 676402 528935 676458 528944
rect 676232 528834 676260 528935
rect 676220 528828 676272 528834
rect 676220 528770 676272 528776
rect 676128 528692 676180 528698
rect 676128 528634 676180 528640
rect 676218 527776 676274 527785
rect 676218 527711 676274 527720
rect 676232 527474 676260 527711
rect 676220 527468 676272 527474
rect 676220 527410 676272 527416
rect 676220 526992 676272 526998
rect 676218 526960 676220 526969
rect 676272 526960 676274 526969
rect 676218 526895 676274 526904
rect 676220 526584 676272 526590
rect 676218 526552 676220 526561
rect 676272 526552 676274 526561
rect 676218 526487 676274 526496
rect 676128 490204 676180 490210
rect 676128 490146 676180 490152
rect 676034 489288 676090 489297
rect 676034 489223 676090 489232
rect 676034 488880 676090 488889
rect 676034 488815 676036 488824
rect 676088 488815 676090 488824
rect 676036 488786 676088 488792
rect 676036 488504 676088 488510
rect 676034 488472 676036 488481
rect 676088 488472 676090 488481
rect 676034 488407 676090 488416
rect 676034 488064 676090 488073
rect 676034 487999 676036 488008
rect 676088 487999 676090 488008
rect 676036 487970 676088 487976
rect 676036 486872 676088 486878
rect 676034 486840 676036 486849
rect 676088 486840 676090 486849
rect 676034 486775 676090 486784
rect 676036 486056 676088 486062
rect 676034 486024 676036 486033
rect 676088 486024 676090 486033
rect 676034 485959 676090 485968
rect 675864 485746 676076 485774
rect 674746 485616 674802 485625
rect 674746 485551 674802 485560
rect 675944 485240 675996 485246
rect 675942 485208 675944 485217
rect 675996 485208 675998 485217
rect 675942 485143 675998 485152
rect 675944 484832 675996 484838
rect 675942 484800 675944 484809
rect 675996 484800 675998 484809
rect 675942 484735 675998 484744
rect 675944 483200 675996 483206
rect 675942 483168 675944 483177
rect 675996 483168 675998 483177
rect 675942 483103 675998 483112
rect 675944 482792 675996 482798
rect 675942 482760 675944 482769
rect 675996 482760 675998 482769
rect 675942 482695 675998 482704
rect 674654 482352 674710 482361
rect 674654 482287 674710 482296
rect 674472 475856 674524 475862
rect 674472 475798 674524 475804
rect 676048 401849 676076 485746
rect 676140 402937 676168 490146
rect 677244 488510 677272 531791
rect 677324 520328 677376 520334
rect 677324 520270 677376 520276
rect 677336 489937 677364 520270
rect 677520 518810 677548 546479
rect 678256 531457 678284 546751
rect 679622 546680 679678 546689
rect 679622 546615 679678 546624
rect 678334 543008 678390 543017
rect 678334 542943 678390 542952
rect 678242 531448 678298 531457
rect 678242 531383 678298 531392
rect 678348 530641 678376 542943
rect 679636 531865 679664 546615
rect 683302 543688 683358 543697
rect 683302 543623 683358 543632
rect 679622 531856 679678 531865
rect 679622 531791 679678 531800
rect 678334 530632 678390 530641
rect 678334 530567 678390 530576
rect 683316 527785 683344 543623
rect 703694 536724 703722 536860
rect 704154 536724 704182 536860
rect 704614 536724 704642 536860
rect 705074 536724 705102 536860
rect 705534 536724 705562 536860
rect 705994 536724 706022 536860
rect 706454 536724 706482 536860
rect 706914 536724 706942 536860
rect 707374 536724 707402 536860
rect 707834 536724 707862 536860
rect 708294 536724 708322 536860
rect 708754 536724 708782 536860
rect 709214 536724 709242 536860
rect 683854 533488 683910 533497
rect 683854 533423 683910 533432
rect 683302 527776 683358 527785
rect 683302 527711 683358 527720
rect 683118 525736 683174 525745
rect 683118 525671 683174 525680
rect 683132 524929 683160 525671
rect 683118 524920 683174 524929
rect 683118 524855 683174 524864
rect 683132 524482 683160 524855
rect 683120 524476 683172 524482
rect 683120 524418 683172 524424
rect 683868 520334 683896 533423
rect 683856 520328 683908 520334
rect 683856 520270 683908 520276
rect 677510 518774 677548 518810
rect 677510 513812 677538 518774
rect 677510 513778 677548 513812
rect 677520 508904 677548 513778
rect 677512 508872 677548 508904
rect 677512 503714 677540 508872
rect 677512 503686 677548 503714
rect 677414 492416 677470 492425
rect 677414 492351 677470 492360
rect 677322 489928 677378 489937
rect 677322 489863 677378 489872
rect 677324 488844 677376 488850
rect 677324 488786 677376 488792
rect 677232 488504 677284 488510
rect 677232 488446 677284 488452
rect 677232 488028 677284 488034
rect 677232 487970 677284 487976
rect 676310 403744 676366 403753
rect 676310 403679 676366 403688
rect 676218 403336 676274 403345
rect 676218 403271 676220 403280
rect 676272 403271 676274 403280
rect 676220 403242 676272 403248
rect 676324 403170 676352 403679
rect 676404 403436 676456 403442
rect 676404 403378 676456 403384
rect 676416 403345 676444 403378
rect 676402 403336 676458 403345
rect 676402 403271 676458 403280
rect 676312 403164 676364 403170
rect 676312 403106 676364 403112
rect 676126 402928 676182 402937
rect 676126 402863 676182 402872
rect 676218 402112 676274 402121
rect 676218 402047 676274 402056
rect 676034 401840 676090 401849
rect 676034 401775 676090 401784
rect 676232 401674 676260 402047
rect 676220 401668 676272 401674
rect 676220 401610 676272 401616
rect 676218 401296 676274 401305
rect 676218 401231 676274 401240
rect 674746 400616 674802 400625
rect 674746 400551 674802 400560
rect 674656 399628 674708 399634
rect 674656 399570 674708 399576
rect 674564 394324 674616 394330
rect 674564 394266 674616 394272
rect 674576 378010 674604 394266
rect 674564 378004 674616 378010
rect 674564 377946 674616 377952
rect 674668 355094 674696 399570
rect 674760 355881 674788 400551
rect 676232 400246 676260 401231
rect 677244 400489 677272 487970
rect 677336 401305 677364 488786
rect 677428 484401 677456 492351
rect 677520 486878 677548 503686
rect 681004 500948 681056 500954
rect 681004 500890 681056 500896
rect 679716 498296 679768 498302
rect 679716 498238 679768 498244
rect 679624 498228 679676 498234
rect 679624 498170 679676 498176
rect 677508 486872 677560 486878
rect 677508 486814 677560 486820
rect 679636 486441 679664 498170
rect 679728 487257 679756 498238
rect 681016 487665 681044 500890
rect 703694 492796 703722 492864
rect 704154 492796 704182 492864
rect 704614 492796 704642 492864
rect 705074 492796 705102 492864
rect 705534 492796 705562 492864
rect 705994 492796 706022 492864
rect 706454 492796 706482 492864
rect 706914 492796 706942 492864
rect 707374 492796 707402 492864
rect 707834 492796 707862 492864
rect 708294 492796 708322 492864
rect 708754 492796 708782 492864
rect 709214 492796 709242 492864
rect 681002 487656 681058 487665
rect 681002 487591 681058 487600
rect 679714 487248 679770 487257
rect 679714 487183 679770 487192
rect 679622 486432 679678 486441
rect 679622 486367 679678 486376
rect 677414 484392 677470 484401
rect 677414 484327 677470 484336
rect 678978 480720 679034 480729
rect 678978 480655 679034 480664
rect 678992 480282 679020 480655
rect 678980 480276 679032 480282
rect 678980 480218 679032 480224
rect 703694 404532 703722 404668
rect 704154 404532 704182 404668
rect 704614 404532 704642 404668
rect 705074 404532 705102 404668
rect 705534 404532 705562 404668
rect 705994 404532 706022 404668
rect 706454 404532 706482 404668
rect 706914 404532 706942 404668
rect 707374 404532 707402 404668
rect 707834 404532 707862 404668
rect 708294 404532 708322 404668
rect 708754 404532 708782 404668
rect 709214 404532 709242 404668
rect 677322 401296 677378 401305
rect 677322 401231 677378 401240
rect 677230 400480 677286 400489
rect 677230 400415 677286 400424
rect 676220 400240 676272 400246
rect 676220 400182 676272 400188
rect 676218 399664 676274 399673
rect 676218 399599 676220 399608
rect 676272 399599 676274 399608
rect 676220 399570 676272 399576
rect 676034 398576 676090 398585
rect 676034 398511 676090 398520
rect 676048 398274 676076 398511
rect 675024 398268 675076 398274
rect 675024 398210 675076 398216
rect 676036 398268 676088 398274
rect 676036 398210 676088 398216
rect 674932 397520 674984 397526
rect 674932 397462 674984 397468
rect 674944 383110 674972 397462
rect 675036 386170 675064 398210
rect 676034 398168 676090 398177
rect 676034 398103 676090 398112
rect 676048 397526 676076 398103
rect 676862 397624 676918 397633
rect 676862 397559 676918 397568
rect 676036 397520 676088 397526
rect 676036 397462 676088 397468
rect 676402 395584 676458 395593
rect 676402 395519 676458 395528
rect 676218 394360 676274 394369
rect 676218 394295 676220 394304
rect 676272 394295 676274 394304
rect 676220 394266 676272 394272
rect 676218 393952 676274 393961
rect 676218 393887 676274 393896
rect 676232 393378 676260 393887
rect 676220 393372 676272 393378
rect 676220 393314 676272 393320
rect 675208 389156 675260 389162
rect 675208 389098 675260 389104
rect 675116 387592 675168 387598
rect 675116 387534 675168 387540
rect 675024 386164 675076 386170
rect 675024 386106 675076 386112
rect 675024 386028 675076 386034
rect 675024 385970 675076 385976
rect 675036 383926 675064 385970
rect 675024 383920 675076 383926
rect 675024 383862 675076 383868
rect 674932 383104 674984 383110
rect 674932 383046 674984 383052
rect 675128 381138 675156 387534
rect 675220 385642 675248 389098
rect 676416 387705 676444 395519
rect 676494 394768 676550 394777
rect 676494 394703 676550 394712
rect 676402 387696 676458 387705
rect 676402 387631 676458 387640
rect 676508 387598 676536 394703
rect 676876 388521 676904 397559
rect 676954 396808 677010 396817
rect 676954 396743 677010 396752
rect 676968 389162 676996 396743
rect 678334 396400 678390 396409
rect 678334 396335 678390 396344
rect 678242 395992 678298 396001
rect 678242 395927 678298 395936
rect 676956 389156 677008 389162
rect 676956 389098 677008 389104
rect 676862 388512 676918 388521
rect 676862 388447 676918 388456
rect 676496 387592 676548 387598
rect 676496 387534 676548 387540
rect 678256 387122 678284 395927
rect 678348 387569 678376 396335
rect 683118 393544 683174 393553
rect 683118 393479 683174 393488
rect 683132 392329 683160 393479
rect 683118 392320 683174 392329
rect 683118 392255 683174 392264
rect 683132 392018 683160 392255
rect 683120 392012 683172 392018
rect 683120 391954 683172 391960
rect 678334 387560 678390 387569
rect 678334 387495 678390 387504
rect 675300 387116 675352 387122
rect 675300 387058 675352 387064
rect 678244 387116 678296 387122
rect 678244 387058 678296 387064
rect 675312 386034 675340 387058
rect 675392 386164 675444 386170
rect 675392 386106 675444 386112
rect 675300 386028 675352 386034
rect 675300 385970 675352 385976
rect 675404 385696 675432 386106
rect 675220 385614 675432 385642
rect 675404 385084 675432 385614
rect 675758 384976 675814 384985
rect 675758 384911 675814 384920
rect 675772 384435 675800 384911
rect 675300 383920 675352 383926
rect 675300 383862 675352 383868
rect 675312 381426 675340 383862
rect 675392 383104 675444 383110
rect 675392 383046 675444 383052
rect 675404 382568 675432 383046
rect 675390 382256 675446 382265
rect 675390 382191 675446 382200
rect 675404 382024 675432 382191
rect 675312 381398 675418 381426
rect 675116 381132 675168 381138
rect 675116 381074 675168 381080
rect 675392 381132 675444 381138
rect 675392 381074 675444 381080
rect 675404 380732 675432 381074
rect 675482 378720 675538 378729
rect 675482 378655 675538 378664
rect 675496 378284 675524 378655
rect 675484 378004 675536 378010
rect 675484 377946 675536 377952
rect 675496 377740 675524 377946
rect 675758 377632 675814 377641
rect 675758 377567 675814 377576
rect 675772 377060 675800 377567
rect 675484 376644 675536 376650
rect 675484 376586 675536 376592
rect 675496 376448 675524 376586
rect 675758 375456 675814 375465
rect 675758 375391 675814 375400
rect 675772 375224 675800 375391
rect 675758 373688 675814 373697
rect 675758 373623 675814 373632
rect 675772 373388 675800 373623
rect 675758 372056 675814 372065
rect 675758 371991 675814 372000
rect 675772 371552 675800 371991
rect 703694 359380 703722 359516
rect 704154 359380 704182 359516
rect 704614 359380 704642 359516
rect 705074 359380 705102 359516
rect 705534 359380 705562 359516
rect 705994 359380 706022 359516
rect 706454 359380 706482 359516
rect 706914 359380 706942 359516
rect 707374 359380 707402 359516
rect 707834 359380 707862 359516
rect 708294 359380 708322 359516
rect 708754 359380 708782 359516
rect 709214 359380 709242 359516
rect 675850 358728 675906 358737
rect 675850 358663 675906 358672
rect 675864 357610 675892 358663
rect 675942 358320 675998 358329
rect 675942 358255 675998 358264
rect 675956 357882 675984 358255
rect 676034 357912 676090 357921
rect 675944 357876 675996 357882
rect 676034 357847 676090 357856
rect 675944 357818 675996 357824
rect 676048 357746 676076 357847
rect 676036 357740 676088 357746
rect 676036 357682 676088 357688
rect 675852 357604 675904 357610
rect 675852 357546 675904 357552
rect 676036 357536 676088 357542
rect 676034 357504 676036 357513
rect 676088 357504 676090 357513
rect 676034 357439 676090 357448
rect 676034 357096 676090 357105
rect 676034 357031 676036 357040
rect 676088 357031 676090 357040
rect 676036 357002 676088 357008
rect 676036 356720 676088 356726
rect 676034 356688 676036 356697
rect 676088 356688 676090 356697
rect 676034 356623 676090 356632
rect 676034 356280 676090 356289
rect 676034 356215 676036 356224
rect 676088 356215 676090 356224
rect 676036 356186 676088 356192
rect 674746 355872 674802 355881
rect 674746 355807 674802 355816
rect 674746 355464 674802 355473
rect 674746 355399 674802 355408
rect 674656 355088 674708 355094
rect 674656 355030 674708 355036
rect 674656 354612 674708 354618
rect 674656 354554 674708 354560
rect 674472 350940 674524 350946
rect 674472 350882 674524 350888
rect 674484 336598 674512 350882
rect 674564 349308 674616 349314
rect 674564 349250 674616 349256
rect 674472 336592 674524 336598
rect 674472 336534 674524 336540
rect 674576 332654 674604 349250
rect 674564 332648 674616 332654
rect 674564 332590 674616 332596
rect 674668 310078 674696 354554
rect 674760 310865 674788 355399
rect 676036 355088 676088 355094
rect 676034 355056 676036 355065
rect 676088 355056 676090 355065
rect 676034 354991 676090 355000
rect 676034 354648 676090 354657
rect 676034 354583 676036 354592
rect 676088 354583 676090 354592
rect 676036 354554 676088 354560
rect 678242 352608 678298 352617
rect 678242 352543 678298 352552
rect 676034 351792 676090 351801
rect 676090 351750 676260 351778
rect 676034 351727 676090 351736
rect 676232 351150 676260 351750
rect 676220 351144 676272 351150
rect 676220 351086 676272 351092
rect 676864 351144 676916 351150
rect 676864 351086 676916 351092
rect 676034 350976 676090 350985
rect 676034 350911 676036 350920
rect 676088 350911 676090 350920
rect 676036 350882 676088 350888
rect 676036 350600 676088 350606
rect 676034 350568 676036 350577
rect 676088 350568 676090 350577
rect 676034 350503 676090 350512
rect 675942 350160 675998 350169
rect 675942 350095 675998 350104
rect 675956 346633 675984 350095
rect 676034 349752 676090 349761
rect 676090 349710 676168 349738
rect 676034 349687 676090 349696
rect 676034 349344 676090 349353
rect 676034 349279 676036 349288
rect 676088 349279 676090 349288
rect 676036 349250 676088 349256
rect 676034 348936 676090 348945
rect 676034 348871 676036 348880
rect 676088 348871 676090 348880
rect 676036 348842 676088 348848
rect 676034 348528 676090 348537
rect 676034 348463 676090 348472
rect 676048 347313 676076 348463
rect 676034 347304 676090 347313
rect 676034 347239 676090 347248
rect 675942 346624 675998 346633
rect 675942 346559 675998 346568
rect 676048 346458 676076 347239
rect 676140 346497 676168 349710
rect 676126 346488 676182 346497
rect 676036 346452 676088 346458
rect 676126 346423 676182 346432
rect 676036 346394 676088 346400
rect 676876 342281 676904 351086
rect 678256 343641 678284 352543
rect 678242 343632 678298 343641
rect 678242 343567 678298 343576
rect 675298 342272 675354 342281
rect 675298 342207 675354 342216
rect 676862 342272 676918 342281
rect 676862 342207 676918 342216
rect 675312 339878 675340 342207
rect 675666 340776 675722 340785
rect 675666 340711 675722 340720
rect 675680 340544 675708 340711
rect 675312 339850 675418 339878
rect 675758 339416 675814 339425
rect 675758 339351 675814 339360
rect 675772 339252 675800 339351
rect 675758 337920 675814 337929
rect 675758 337855 675814 337864
rect 675772 337416 675800 337855
rect 675404 336326 675432 336843
rect 675484 336592 675536 336598
rect 675484 336534 675536 336540
rect 674840 336320 674892 336326
rect 674840 336262 674892 336268
rect 675392 336320 675444 336326
rect 675392 336262 675444 336268
rect 674852 335345 674880 336262
rect 675496 336192 675524 336534
rect 675758 335880 675814 335889
rect 675758 335815 675814 335824
rect 675772 335580 675800 335815
rect 674838 335336 674894 335345
rect 674838 335271 674894 335280
rect 675482 333568 675538 333577
rect 675482 333503 675538 333512
rect 675496 333064 675524 333503
rect 675392 332648 675444 332654
rect 675392 332590 675444 332596
rect 675404 332520 675432 332590
rect 675758 332208 675814 332217
rect 675758 332143 675814 332152
rect 675772 331875 675800 332143
rect 675392 331628 675444 331634
rect 675392 331570 675444 331576
rect 675404 331228 675432 331570
rect 675404 329526 675432 330035
rect 674840 329520 674892 329526
rect 674840 329462 674892 329468
rect 675392 329520 675444 329526
rect 675392 329462 675444 329468
rect 674852 328438 674880 329462
rect 674840 328432 674892 328438
rect 674840 328374 674892 328380
rect 675496 327690 675524 328168
rect 675116 327684 675168 327690
rect 675116 327626 675168 327632
rect 675484 327684 675536 327690
rect 675484 327626 675536 327632
rect 675128 325689 675156 327626
rect 675772 325854 675800 326332
rect 675760 325848 675812 325854
rect 675760 325790 675812 325796
rect 675114 325680 675170 325689
rect 675114 325615 675170 325624
rect 675760 325644 675812 325650
rect 675760 325586 675812 325592
rect 675772 325553 675800 325586
rect 675758 325544 675814 325553
rect 675758 325479 675814 325488
rect 703694 314364 703722 314500
rect 704154 314364 704182 314500
rect 704614 314364 704642 314500
rect 705074 314364 705102 314500
rect 705534 314364 705562 314500
rect 705994 314364 706022 314500
rect 706454 314364 706482 314500
rect 706914 314364 706942 314500
rect 707374 314364 707402 314500
rect 707834 314364 707862 314500
rect 708294 314364 708322 314500
rect 708754 314364 708782 314500
rect 709214 314364 709242 314500
rect 676034 313712 676090 313721
rect 676034 313647 676090 313656
rect 676048 313410 676076 313647
rect 676218 313576 676274 313585
rect 676218 313511 676220 313520
rect 676272 313511 676274 313520
rect 676220 313482 676272 313488
rect 676036 313404 676088 313410
rect 676036 313346 676088 313352
rect 676126 312760 676182 312769
rect 676126 312695 676182 312704
rect 676140 312050 676168 312695
rect 676218 312352 676274 312361
rect 676218 312287 676274 312296
rect 676232 312186 676260 312287
rect 676220 312180 676272 312186
rect 676220 312122 676272 312128
rect 676128 312044 676180 312050
rect 676128 311986 676180 311992
rect 676218 311944 676274 311953
rect 676218 311879 676220 311888
rect 676272 311879 676274 311888
rect 676220 311850 676272 311856
rect 676218 311536 676274 311545
rect 676218 311471 676274 311480
rect 676126 311128 676182 311137
rect 676126 311063 676182 311072
rect 674746 310856 674802 310865
rect 674746 310791 674802 310800
rect 676140 310554 676168 311063
rect 676232 310690 676260 311471
rect 676220 310684 676272 310690
rect 676220 310626 676272 310632
rect 676128 310548 676180 310554
rect 676128 310490 676180 310496
rect 676218 310312 676274 310321
rect 674748 310276 674800 310282
rect 676218 310247 676220 310256
rect 674748 310218 674800 310224
rect 676272 310247 676274 310256
rect 676220 310218 676272 310224
rect 674656 310072 674708 310078
rect 674656 310014 674708 310020
rect 674760 309618 674788 310218
rect 676036 310072 676088 310078
rect 676034 310040 676036 310049
rect 676088 310040 676090 310049
rect 676034 309975 676090 309984
rect 674668 309590 674788 309618
rect 674380 302252 674432 302258
rect 674380 302194 674432 302200
rect 674288 148436 674340 148442
rect 674288 148378 674340 148384
rect 674392 133006 674420 302194
rect 674668 265878 674696 309590
rect 676218 309496 676274 309505
rect 674748 309460 674800 309466
rect 676218 309431 676220 309440
rect 674748 309402 674800 309408
rect 676272 309431 676274 309440
rect 676220 309402 676272 309408
rect 674656 265872 674708 265878
rect 674656 265814 674708 265820
rect 674760 265033 674788 309402
rect 679622 309088 679678 309097
rect 679622 309023 679678 309032
rect 678242 308272 678298 308281
rect 678242 308207 678298 308216
rect 676862 306640 676918 306649
rect 676862 306575 676918 306584
rect 676402 306232 676458 306241
rect 676402 306167 676458 306176
rect 676310 304600 676366 304609
rect 676310 304535 676366 304544
rect 676126 304192 676182 304201
rect 676126 304127 676182 304136
rect 676140 303754 676168 304127
rect 676220 303816 676272 303822
rect 676218 303784 676220 303793
rect 676272 303784 676274 303793
rect 676128 303748 676180 303754
rect 676218 303719 676274 303728
rect 676128 303690 676180 303696
rect 676324 303686 676352 304535
rect 676312 303680 676364 303686
rect 676312 303622 676364 303628
rect 675208 298104 675260 298110
rect 675208 298046 675260 298052
rect 675116 297424 675168 297430
rect 675116 297366 675168 297372
rect 675128 294098 675156 297366
rect 675220 295458 675248 298046
rect 675760 298036 675812 298042
rect 675760 297978 675812 297984
rect 675772 296206 675800 297978
rect 676416 297401 676444 306167
rect 676494 305824 676550 305833
rect 676494 305759 676550 305768
rect 676508 297430 676536 305759
rect 676876 298110 676904 306575
rect 676864 298104 676916 298110
rect 676864 298046 676916 298052
rect 678256 298042 678284 308207
rect 679636 299441 679664 309023
rect 679714 307456 679770 307465
rect 679714 307391 679770 307400
rect 679622 299432 679678 299441
rect 679622 299367 679678 299376
rect 678244 298036 678296 298042
rect 678244 297978 678296 297984
rect 679728 297945 679756 307391
rect 683118 303376 683174 303385
rect 683118 303311 683174 303320
rect 683132 302569 683160 303311
rect 683118 302560 683174 302569
rect 683118 302495 683174 302504
rect 683132 302258 683160 302495
rect 683120 302252 683172 302258
rect 683120 302194 683172 302200
rect 679714 297936 679770 297945
rect 679714 297871 679770 297880
rect 676496 297424 676548 297430
rect 676402 297392 676458 297401
rect 676496 297366 676548 297372
rect 676402 297327 676458 297336
rect 675760 296200 675812 296206
rect 675760 296142 675812 296148
rect 675760 295996 675812 296002
rect 675760 295938 675812 295944
rect 675772 295528 675800 295938
rect 675208 295452 675260 295458
rect 675208 295394 675260 295400
rect 675392 295452 675444 295458
rect 675392 295394 675444 295400
rect 675404 294879 675432 295394
rect 675758 294808 675814 294817
rect 675758 294743 675814 294752
rect 675772 294236 675800 294743
rect 675116 294092 675168 294098
rect 675116 294034 675168 294040
rect 675024 294024 675076 294030
rect 675024 293966 675076 293972
rect 675036 291786 675064 293966
rect 675482 292632 675538 292641
rect 675482 292567 675538 292576
rect 675496 292400 675524 292567
rect 675390 292088 675446 292097
rect 675390 292023 675446 292032
rect 675404 291856 675432 292023
rect 675024 291780 675076 291786
rect 675024 291722 675076 291728
rect 675392 291780 675444 291786
rect 675392 291722 675444 291728
rect 675404 291176 675432 291722
rect 675392 291100 675444 291106
rect 675392 291042 675444 291048
rect 675404 290564 675432 291042
rect 675666 288416 675722 288425
rect 675666 288351 675722 288360
rect 675680 288048 675708 288351
rect 675392 287972 675444 287978
rect 675392 287914 675444 287920
rect 675404 287504 675432 287914
rect 675758 287328 675814 287337
rect 675758 287263 675814 287272
rect 675772 286892 675800 287263
rect 675392 286612 675444 286618
rect 675392 286554 675444 286560
rect 675404 286212 675432 286554
rect 675758 285560 675814 285569
rect 675758 285495 675814 285504
rect 675772 285056 675800 285495
rect 675758 283656 675814 283665
rect 675758 283591 675814 283600
rect 675772 283220 675800 283591
rect 675758 281480 675814 281489
rect 675758 281415 675814 281424
rect 675772 281355 675800 281415
rect 703694 269348 703722 269484
rect 704154 269348 704182 269484
rect 704614 269348 704642 269484
rect 705074 269348 705102 269484
rect 705534 269348 705562 269484
rect 705994 269348 706022 269484
rect 706454 269348 706482 269484
rect 706914 269348 706942 269484
rect 707374 269348 707402 269484
rect 707834 269348 707862 269484
rect 708294 269348 708322 269484
rect 708754 269348 708782 269484
rect 709214 269348 709242 269484
rect 676218 268560 676274 268569
rect 676218 268495 676274 268504
rect 676126 268152 676182 268161
rect 676232 268122 676260 268495
rect 676126 268087 676182 268096
rect 676220 268116 676272 268122
rect 676140 267782 676168 268087
rect 676220 268058 676272 268064
rect 676220 267980 676272 267986
rect 676220 267922 676272 267928
rect 676128 267776 676180 267782
rect 676232 267753 676260 267922
rect 676128 267718 676180 267724
rect 676218 267744 676274 267753
rect 676218 267679 676274 267688
rect 676218 267336 676274 267345
rect 676218 267271 676274 267280
rect 676034 267064 676090 267073
rect 676034 266999 676036 267008
rect 676088 266999 676090 267008
rect 676036 266970 676088 266976
rect 676232 266626 676260 267271
rect 676220 266620 676272 266626
rect 676220 266562 676272 266568
rect 676218 266520 676274 266529
rect 676218 266455 676220 266464
rect 676272 266455 676274 266464
rect 676220 266426 676272 266432
rect 676218 266112 676274 266121
rect 676218 266047 676220 266056
rect 676272 266047 676274 266056
rect 676220 266018 676272 266024
rect 676036 265872 676088 265878
rect 676034 265840 676036 265849
rect 676088 265840 676090 265849
rect 676034 265775 676090 265784
rect 676218 265296 676274 265305
rect 676218 265231 676274 265240
rect 674746 265024 674802 265033
rect 676232 264994 676260 265231
rect 674746 264959 674802 264968
rect 676220 264988 676272 264994
rect 676220 264930 676272 264936
rect 676218 264480 676274 264489
rect 676218 264415 676274 264424
rect 676232 263634 676260 264415
rect 676310 264072 676366 264081
rect 676310 264007 676366 264016
rect 676220 263628 676272 263634
rect 676220 263570 676272 263576
rect 675390 263392 675446 263401
rect 675390 263327 675446 263336
rect 675024 262676 675076 262682
rect 675024 262618 675076 262624
rect 674472 261996 674524 262002
rect 674472 261938 674524 261944
rect 674484 245721 674512 261938
rect 674748 261588 674800 261594
rect 674748 261530 674800 261536
rect 674564 259956 674616 259962
rect 674564 259898 674616 259904
rect 674470 245712 674526 245721
rect 674470 245647 674526 245656
rect 674576 242214 674604 259898
rect 674656 251728 674708 251734
rect 674656 251670 674708 251676
rect 674668 249626 674696 251670
rect 674760 250238 674788 261530
rect 675036 251734 675064 262618
rect 675208 262268 675260 262274
rect 675208 262210 675260 262216
rect 675024 251728 675076 251734
rect 675024 251670 675076 251676
rect 675024 251592 675076 251598
rect 675024 251534 675076 251540
rect 674748 250232 674800 250238
rect 674748 250174 674800 250180
rect 675036 249762 675064 251534
rect 675024 249756 675076 249762
rect 675024 249698 675076 249704
rect 674656 249620 674708 249626
rect 674656 249562 674708 249568
rect 675024 249620 675076 249626
rect 675024 249562 675076 249568
rect 675036 247926 675064 249562
rect 675220 248538 675248 262210
rect 675404 251258 675432 263327
rect 676034 262984 676090 262993
rect 676034 262919 676090 262928
rect 676048 262682 676076 262919
rect 676036 262676 676088 262682
rect 676036 262618 676088 262624
rect 676034 262576 676090 262585
rect 676034 262511 676090 262520
rect 676048 262274 676076 262511
rect 676036 262268 676088 262274
rect 676036 262210 676088 262216
rect 676218 262032 676274 262041
rect 676218 261967 676220 261976
rect 676272 261967 676274 261976
rect 676220 261938 676272 261944
rect 676218 261624 676274 261633
rect 676218 261559 676220 261568
rect 676272 261559 676274 261568
rect 676220 261530 676272 261536
rect 676218 261216 676274 261225
rect 676218 261151 676274 261160
rect 676232 260914 676260 261151
rect 676220 260908 676272 260914
rect 676220 260850 676272 260856
rect 676218 259992 676274 260001
rect 676218 259927 676220 259936
rect 676272 259927 676274 259936
rect 676220 259898 676272 259904
rect 676324 259418 676352 264007
rect 676862 263664 676918 263673
rect 676862 263599 676918 263608
rect 675484 259412 675536 259418
rect 675484 259354 675536 259360
rect 676312 259412 676364 259418
rect 676312 259354 676364 259360
rect 675496 251598 675524 259354
rect 676126 259176 676182 259185
rect 676126 259111 676182 259120
rect 676140 258126 676168 259111
rect 676218 258768 676274 258777
rect 676218 258703 676274 258712
rect 676232 258194 676260 258703
rect 676220 258188 676272 258194
rect 676220 258130 676272 258136
rect 676128 258120 676180 258126
rect 676128 258062 676180 258068
rect 675484 251592 675536 251598
rect 676876 251569 676904 263599
rect 683118 258360 683174 258369
rect 683118 258295 683174 258304
rect 683132 257553 683160 258295
rect 683118 257544 683174 257553
rect 683118 257479 683174 257488
rect 683132 256766 683160 257479
rect 683120 256760 683172 256766
rect 683120 256702 683172 256708
rect 675484 251534 675536 251540
rect 676862 251560 676918 251569
rect 676862 251495 676918 251504
rect 675392 251252 675444 251258
rect 675392 251194 675444 251200
rect 675392 250980 675444 250986
rect 675392 250922 675444 250928
rect 675404 250512 675432 250922
rect 675484 250232 675536 250238
rect 675484 250174 675536 250180
rect 675496 249900 675524 250174
rect 675392 249756 675444 249762
rect 675392 249698 675444 249704
rect 675404 249220 675432 249698
rect 675208 248532 675260 248538
rect 675208 248474 675260 248480
rect 675208 248328 675260 248334
rect 675114 248296 675170 248305
rect 675208 248270 675260 248276
rect 675114 248231 675170 248240
rect 675024 247920 675076 247926
rect 675024 247862 675076 247868
rect 675128 243914 675156 248231
rect 675220 243914 675248 248270
rect 675484 247920 675536 247926
rect 675484 247862 675536 247868
rect 675496 247384 675524 247862
rect 675392 247036 675444 247042
rect 675392 246978 675444 246984
rect 675404 246840 675432 246978
rect 675758 246664 675814 246673
rect 675758 246599 675814 246608
rect 675772 246199 675800 246599
rect 675772 245449 675800 245548
rect 675758 245440 675814 245449
rect 675758 245375 675814 245384
rect 674748 243908 674800 243914
rect 674748 243850 674800 243856
rect 675116 243908 675168 243914
rect 675116 243850 675168 243856
rect 675208 243908 675260 243914
rect 675208 243850 675260 243856
rect 674564 242208 674616 242214
rect 674564 242150 674616 242156
rect 674760 238814 674788 243850
rect 675300 243636 675352 243642
rect 675300 243578 675352 243584
rect 675312 243085 675340 243578
rect 675312 243057 675418 243085
rect 675312 242505 675418 242533
rect 675312 241670 675340 242505
rect 675392 242208 675444 242214
rect 675392 242150 675444 242156
rect 675404 241876 675432 242150
rect 675300 241664 675352 241670
rect 675300 241606 675352 241612
rect 675312 241217 675418 241245
rect 675312 241126 675340 241217
rect 675300 241120 675352 241126
rect 675300 241062 675352 241068
rect 675312 240026 675418 240054
rect 674748 238808 674800 238814
rect 674748 238750 674800 238756
rect 675312 238649 675340 240026
rect 675392 238740 675444 238746
rect 675392 238682 675444 238688
rect 675298 238640 675354 238649
rect 675298 238575 675354 238584
rect 675404 238204 675432 238682
rect 675758 236872 675814 236881
rect 675758 236807 675814 236816
rect 675772 236368 675800 236807
rect 703694 224196 703722 224264
rect 704154 224196 704182 224264
rect 704614 224196 704642 224264
rect 705074 224196 705102 224264
rect 705534 224196 705562 224264
rect 705994 224196 706022 224264
rect 706454 224196 706482 224264
rect 706914 224196 706942 224264
rect 707374 224196 707402 224264
rect 707834 224196 707862 224264
rect 708294 224196 708322 224264
rect 708754 224196 708782 224264
rect 709214 224196 709242 224264
rect 675942 223544 675998 223553
rect 675942 223479 675998 223488
rect 675850 222728 675906 222737
rect 675850 222663 675906 222672
rect 675864 222222 675892 222663
rect 675956 222562 675984 223479
rect 676034 223136 676090 223145
rect 676034 223071 676090 223080
rect 675944 222556 675996 222562
rect 675944 222498 675996 222504
rect 676048 222426 676076 223071
rect 676036 222420 676088 222426
rect 676036 222362 676088 222368
rect 676034 222320 676090 222329
rect 676034 222255 676036 222264
rect 676088 222255 676090 222264
rect 676036 222226 676088 222232
rect 675852 222216 675904 222222
rect 675852 222158 675904 222164
rect 676034 221912 676090 221921
rect 674656 221876 674708 221882
rect 676034 221847 676036 221856
rect 674656 221818 674708 221824
rect 676088 221847 676090 221856
rect 676036 221818 676088 221824
rect 674564 215756 674616 215762
rect 674564 215698 674616 215704
rect 674576 201482 674604 215698
rect 674564 201476 674616 201482
rect 674564 201418 674616 201424
rect 674668 177342 674696 221818
rect 676036 221536 676088 221542
rect 676034 221504 676036 221513
rect 676088 221504 676090 221513
rect 676034 221439 676090 221448
rect 674746 221096 674802 221105
rect 674746 221031 674802 221040
rect 674656 177336 674708 177342
rect 674656 177278 674708 177284
rect 674760 176497 674788 221031
rect 676036 220720 676088 220726
rect 676034 220688 676036 220697
rect 676088 220688 676090 220697
rect 676034 220623 676090 220632
rect 676034 220280 676090 220289
rect 676034 220215 676036 220224
rect 676088 220215 676090 220224
rect 676036 220186 676088 220192
rect 676036 219904 676088 219910
rect 676034 219872 676036 219881
rect 676088 219872 676090 219881
rect 676034 219807 676090 219816
rect 676036 219496 676088 219502
rect 676034 219464 676036 219473
rect 676088 219464 676090 219473
rect 676034 219399 676090 219408
rect 676034 219056 676090 219065
rect 676090 219014 676352 219042
rect 676034 218991 676090 219000
rect 675850 217016 675906 217025
rect 675850 216951 675906 216960
rect 675864 211313 675892 216951
rect 676034 216608 676090 216617
rect 676090 216566 676260 216594
rect 676034 216543 676090 216552
rect 676034 216200 676090 216209
rect 676034 216135 676036 216144
rect 676088 216135 676090 216144
rect 676036 216106 676088 216112
rect 676034 215792 676090 215801
rect 676034 215727 676036 215736
rect 676088 215727 676090 215736
rect 676036 215698 676088 215704
rect 676232 215558 676260 216566
rect 676220 215552 676272 215558
rect 676220 215494 676272 215500
rect 675942 214976 675998 214985
rect 675942 214911 675998 214920
rect 675956 211449 675984 214911
rect 676034 214160 676090 214169
rect 676034 214095 676036 214104
rect 676088 214095 676090 214104
rect 676036 214066 676088 214072
rect 676034 214024 676090 214033
rect 676324 214010 676352 219014
rect 679622 217424 679678 217433
rect 679622 217359 679678 217368
rect 676864 215552 676916 215558
rect 676864 215494 676916 215500
rect 676090 213982 676352 214010
rect 676034 213959 676090 213968
rect 676034 213752 676090 213761
rect 676034 213687 676036 213696
rect 676088 213687 676090 213696
rect 676036 213658 676088 213664
rect 676034 213344 676090 213353
rect 676034 213279 676090 213288
rect 676048 212129 676076 213279
rect 676034 212120 676090 212129
rect 676034 212055 676090 212064
rect 675942 211440 675998 211449
rect 675942 211375 675998 211384
rect 675850 211304 675906 211313
rect 675850 211239 675906 211248
rect 676048 211206 676076 212055
rect 676036 211200 676088 211206
rect 676036 211142 676088 211148
rect 676876 208321 676904 215494
rect 676862 208312 676918 208321
rect 676862 208247 676918 208256
rect 679636 207233 679664 217359
rect 679622 207224 679678 207233
rect 679622 207159 679678 207168
rect 675758 205592 675814 205601
rect 675758 205527 675814 205536
rect 675772 205323 675800 205527
rect 675758 205048 675814 205057
rect 675758 204983 675814 204992
rect 675772 204680 675800 204983
rect 675758 204232 675814 204241
rect 675758 204167 675814 204176
rect 675772 204035 675800 204167
rect 675114 202872 675170 202881
rect 675114 202807 675170 202816
rect 674838 201376 674894 201385
rect 674838 201311 674894 201320
rect 674852 197062 674880 201311
rect 675128 200734 675156 202807
rect 675482 202736 675538 202745
rect 675482 202671 675538 202680
rect 675496 202195 675524 202671
rect 675392 201884 675444 201890
rect 675392 201826 675444 201832
rect 675404 201620 675432 201826
rect 675392 201476 675444 201482
rect 675392 201418 675444 201424
rect 675404 201008 675432 201418
rect 675116 200728 675168 200734
rect 675116 200670 675168 200676
rect 675392 200728 675444 200734
rect 675392 200670 675444 200676
rect 675404 200328 675432 200670
rect 675758 198384 675814 198393
rect 675758 198319 675814 198328
rect 675772 197880 675800 198319
rect 675484 197464 675536 197470
rect 675484 197406 675536 197412
rect 675496 197336 675524 197406
rect 674840 197056 674892 197062
rect 674840 196998 674892 197004
rect 675392 197056 675444 197062
rect 675392 196998 675444 197004
rect 675404 196656 675432 196998
rect 675392 196580 675444 196586
rect 675392 196522 675444 196528
rect 675404 196044 675432 196522
rect 675758 195392 675814 195401
rect 675758 195327 675814 195336
rect 675772 194820 675800 195327
rect 675404 192506 675432 192984
rect 674840 192500 674892 192506
rect 674840 192442 674892 192448
rect 675392 192500 675444 192506
rect 675392 192442 675444 192448
rect 674852 190233 674880 192442
rect 675772 190670 675800 191148
rect 675760 190664 675812 190670
rect 675760 190606 675812 190612
rect 675760 190392 675812 190398
rect 675758 190360 675760 190369
rect 675812 190360 675814 190369
rect 675758 190295 675814 190304
rect 674838 190224 674894 190233
rect 674838 190159 674894 190168
rect 703694 179180 703722 179316
rect 704154 179180 704182 179316
rect 704614 179180 704642 179316
rect 705074 179180 705102 179316
rect 705534 179180 705562 179316
rect 705994 179180 706022 179316
rect 706454 179180 706482 179316
rect 706914 179180 706942 179316
rect 707374 179180 707402 179316
rect 707834 179180 707862 179316
rect 708294 179180 708322 179316
rect 708754 179180 708782 179316
rect 709214 179180 709242 179316
rect 675942 178528 675998 178537
rect 675942 178463 675998 178472
rect 675956 178226 675984 178463
rect 676036 178356 676088 178362
rect 676036 178298 676088 178304
rect 675944 178220 675996 178226
rect 675944 178162 675996 178168
rect 676048 178129 676076 178298
rect 676034 178120 676090 178129
rect 676034 178055 676090 178064
rect 675942 177712 675998 177721
rect 675942 177647 675998 177656
rect 675956 176866 675984 177647
rect 676036 177336 676088 177342
rect 676034 177304 676036 177313
rect 676088 177304 676090 177313
rect 676034 177239 676090 177248
rect 676034 176896 676090 176905
rect 675944 176860 675996 176866
rect 676034 176831 676090 176840
rect 675944 176802 675996 176808
rect 676048 176730 676076 176831
rect 676036 176724 676088 176730
rect 676036 176666 676088 176672
rect 674746 176488 674802 176497
rect 674746 176423 674802 176432
rect 676034 176080 676090 176089
rect 676034 176015 676036 176024
rect 676088 176015 676090 176024
rect 676036 175986 676088 175992
rect 676036 175704 676088 175710
rect 676034 175672 676036 175681
rect 676088 175672 676090 175681
rect 676034 175607 676090 175616
rect 676034 175264 676090 175273
rect 676034 175199 676036 175208
rect 676088 175199 676090 175208
rect 676036 175170 676088 175176
rect 676036 174888 676088 174894
rect 676034 174856 676036 174865
rect 676088 174856 676090 174865
rect 676034 174791 676090 174800
rect 674746 174448 674802 174457
rect 674746 174383 674802 174392
rect 674656 170332 674708 170338
rect 674656 170274 674708 170280
rect 674564 169108 674616 169114
rect 674564 169050 674616 169056
rect 674576 152590 674604 169050
rect 674564 152584 674616 152590
rect 674564 152526 674616 152532
rect 674668 150414 674696 170274
rect 674656 150408 674708 150414
rect 674656 150350 674708 150356
rect 674380 133000 674432 133006
rect 674380 132942 674432 132948
rect 674760 129713 674788 174383
rect 678242 173224 678298 173233
rect 678242 173159 678298 173168
rect 676034 172816 676090 172825
rect 676090 172774 676352 172802
rect 676034 172751 676090 172760
rect 676034 172408 676090 172417
rect 676090 172366 676260 172394
rect 676034 172343 676090 172352
rect 676232 171290 676260 172366
rect 676220 171284 676272 171290
rect 676220 171226 676272 171232
rect 676034 171184 676090 171193
rect 676090 171154 676260 171170
rect 676090 171148 676272 171154
rect 676090 171142 676220 171148
rect 676034 171119 676090 171128
rect 676220 171090 676272 171096
rect 676034 170368 676090 170377
rect 676034 170303 676036 170312
rect 676088 170303 676090 170312
rect 676036 170274 676088 170280
rect 676034 169688 676090 169697
rect 676324 169674 676352 172774
rect 676770 171592 676826 171601
rect 676770 171527 676826 171536
rect 676586 169960 676642 169969
rect 676586 169895 676642 169904
rect 676090 169646 676352 169674
rect 676034 169623 676090 169632
rect 676034 169552 676090 169561
rect 676034 169487 676036 169496
rect 676088 169487 676090 169496
rect 676036 169458 676088 169464
rect 676034 169144 676090 169153
rect 676034 169079 676036 169088
rect 676088 169079 676090 169088
rect 676036 169050 676088 169056
rect 676034 168736 676090 168745
rect 676034 168671 676090 168680
rect 676048 168638 676076 168671
rect 676036 168632 676088 168638
rect 676036 168574 676088 168580
rect 676034 168328 676090 168337
rect 676034 168263 676036 168272
rect 676088 168263 676090 168272
rect 676036 168234 676088 168240
rect 676034 167920 676090 167929
rect 676034 167855 676036 167864
rect 676088 167855 676090 167864
rect 676036 167826 676088 167832
rect 676034 167104 676090 167113
rect 676034 167039 676036 167048
rect 676088 167039 676090 167048
rect 676036 167010 676088 167016
rect 676600 166433 676628 169895
rect 676784 166433 676812 171527
rect 677048 171284 677100 171290
rect 677048 171226 677100 171232
rect 676864 171148 676916 171154
rect 676864 171090 676916 171096
rect 676586 166424 676642 166433
rect 676586 166359 676642 166368
rect 676770 166424 676826 166433
rect 676770 166359 676826 166368
rect 675760 162852 675812 162858
rect 675760 162794 675812 162800
rect 675772 161022 675800 162794
rect 676876 162625 676904 171090
rect 677060 162761 677088 171226
rect 678256 162858 678284 173159
rect 678244 162852 678296 162858
rect 678244 162794 678296 162800
rect 677046 162752 677102 162761
rect 677046 162687 677102 162696
rect 676862 162616 676918 162625
rect 676862 162551 676918 162560
rect 675760 161016 675812 161022
rect 675760 160958 675812 160964
rect 675760 160812 675812 160818
rect 675760 160754 675812 160760
rect 675772 160344 675800 160754
rect 675758 160032 675814 160041
rect 675758 159967 675814 159976
rect 675772 159664 675800 159967
rect 675482 159488 675538 159497
rect 675482 159423 675538 159432
rect 675496 159052 675524 159423
rect 675666 157448 675722 157457
rect 675666 157383 675722 157392
rect 675680 157216 675708 157383
rect 675482 157040 675538 157049
rect 675482 156975 675538 156984
rect 675496 156643 675524 156975
rect 675758 156360 675814 156369
rect 675758 156295 675814 156304
rect 675772 155992 675800 156295
rect 675484 155508 675536 155514
rect 675484 155450 675536 155456
rect 675496 155380 675524 155450
rect 675758 153096 675814 153105
rect 675758 153031 675814 153040
rect 675772 152864 675800 153031
rect 675392 152584 675444 152590
rect 675392 152526 675444 152532
rect 675404 152320 675432 152526
rect 675772 151609 675800 151675
rect 675758 151600 675814 151609
rect 675758 151535 675814 151544
rect 675392 151428 675444 151434
rect 675392 151370 675444 151376
rect 675404 151028 675432 151370
rect 675392 150408 675444 150414
rect 675392 150350 675444 150356
rect 675404 149835 675432 150350
rect 675758 148472 675814 148481
rect 675758 148407 675814 148416
rect 675772 147968 675800 148407
rect 675758 146296 675814 146305
rect 675758 146231 675814 146240
rect 675772 146132 675800 146231
rect 703694 133892 703722 134028
rect 704154 133892 704182 134028
rect 704614 133892 704642 134028
rect 705074 133892 705102 134028
rect 705534 133892 705562 134028
rect 705994 133892 706022 134028
rect 706454 133892 706482 134028
rect 706914 133892 706942 134028
rect 707374 133892 707402 134028
rect 707834 133892 707862 134028
rect 708294 133892 708322 134028
rect 708754 133892 708782 134028
rect 709214 133892 709242 134028
rect 676126 133104 676182 133113
rect 676036 133068 676088 133074
rect 676126 133039 676182 133048
rect 676036 133010 676088 133016
rect 676048 132977 676076 133010
rect 676034 132968 676090 132977
rect 676034 132903 676090 132912
rect 676140 132666 676168 133039
rect 676220 132796 676272 132802
rect 676220 132738 676272 132744
rect 676232 132705 676260 132738
rect 676218 132696 676274 132705
rect 676128 132660 676180 132666
rect 676218 132631 676274 132640
rect 676128 132602 676180 132608
rect 676218 131880 676274 131889
rect 676218 131815 676274 131824
rect 676126 131472 676182 131481
rect 676232 131442 676260 131815
rect 676126 131407 676182 131416
rect 676220 131436 676272 131442
rect 676034 131336 676090 131345
rect 676034 131271 676036 131280
rect 676088 131271 676090 131280
rect 676036 131242 676088 131248
rect 676140 131170 676168 131407
rect 676220 131378 676272 131384
rect 676128 131164 676180 131170
rect 676128 131106 676180 131112
rect 676126 130656 676182 130665
rect 676126 130591 676182 130600
rect 676140 129878 676168 130591
rect 676218 130248 676274 130257
rect 676218 130183 676274 130192
rect 676232 130014 676260 130183
rect 676220 130008 676272 130014
rect 676220 129950 676272 129956
rect 676128 129872 676180 129878
rect 676128 129814 676180 129820
rect 676218 129840 676274 129849
rect 676218 129775 676220 129784
rect 676272 129775 676274 129784
rect 676220 129746 676272 129752
rect 674746 129704 674802 129713
rect 674746 129639 674802 129648
rect 676218 129024 676274 129033
rect 676218 128959 676274 128968
rect 676232 128382 676260 128959
rect 676220 128376 676272 128382
rect 676220 128318 676272 128324
rect 683670 128208 683726 128217
rect 683670 128143 683726 128152
rect 676034 128072 676090 128081
rect 676034 128007 676090 128016
rect 676048 127022 676076 128007
rect 683118 127392 683174 127401
rect 683118 127327 683174 127336
rect 675116 127016 675168 127022
rect 675116 126958 675168 126964
rect 676036 127016 676088 127022
rect 676036 126958 676088 126964
rect 676862 126984 676918 126993
rect 674656 123956 674708 123962
rect 674656 123898 674708 123904
rect 674196 114368 674248 114374
rect 674196 114310 674248 114316
rect 674668 107574 674696 123898
rect 674746 123584 674802 123593
rect 674746 123519 674802 123528
rect 674656 107568 674708 107574
rect 674656 107510 674708 107516
rect 674760 106282 674788 123519
rect 675128 115598 675156 126958
rect 676862 126919 676918 126928
rect 676402 125352 676458 125361
rect 676402 125287 676458 125296
rect 676034 123992 676090 124001
rect 676034 123927 676036 123936
rect 676088 123927 676090 123936
rect 676036 123898 676088 123904
rect 676218 122904 676274 122913
rect 676218 122839 676220 122848
rect 676272 122839 676274 122848
rect 676220 122810 676272 122816
rect 676126 122496 676182 122505
rect 676126 122431 676182 122440
rect 676140 121514 676168 122431
rect 676218 121680 676274 121689
rect 676218 121615 676274 121624
rect 676128 121508 676180 121514
rect 676128 121450 676180 121456
rect 676232 120766 676260 121615
rect 676220 120760 676272 120766
rect 676220 120702 676272 120708
rect 676416 117337 676444 125287
rect 676876 118017 676904 126919
rect 679622 125760 679678 125769
rect 679622 125695 679678 125704
rect 678242 125352 678298 125361
rect 678242 125287 678298 125296
rect 677598 124128 677654 124137
rect 677598 124063 677654 124072
rect 676862 118008 676918 118017
rect 676862 117943 676918 117952
rect 676402 117328 676458 117337
rect 676402 117263 676458 117272
rect 677612 116754 677640 124063
rect 675484 116748 675536 116754
rect 675484 116690 675536 116696
rect 677600 116748 677652 116754
rect 677600 116690 677652 116696
rect 675208 116612 675260 116618
rect 675208 116554 675260 116560
rect 675116 115592 675168 115598
rect 675116 115534 675168 115540
rect 675116 115456 675168 115462
rect 675116 115398 675168 115404
rect 675128 114730 675156 115398
rect 675220 114850 675248 116554
rect 675496 115802 675524 116690
rect 678256 116210 678284 125287
rect 679636 117201 679664 125695
rect 683132 124953 683160 127327
rect 683302 126168 683358 126177
rect 683302 126103 683358 126112
rect 683118 124944 683174 124953
rect 683118 124879 683174 124888
rect 679622 117192 679678 117201
rect 679622 117127 679678 117136
rect 683316 116618 683344 126103
rect 683684 121689 683712 128143
rect 683670 121680 683726 121689
rect 683670 121615 683726 121624
rect 683304 116612 683356 116618
rect 683304 116554 683356 116560
rect 678244 116204 678296 116210
rect 678244 116146 678296 116152
rect 675484 115796 675536 115802
rect 675484 115738 675536 115744
rect 675392 115592 675444 115598
rect 675392 115534 675444 115540
rect 675404 115124 675432 115534
rect 675208 114844 675260 114850
rect 675208 114786 675260 114792
rect 675392 114844 675444 114850
rect 675392 114786 675444 114792
rect 675128 114702 675248 114730
rect 675116 114640 675168 114646
rect 675116 114582 675168 114588
rect 675128 110702 675156 114582
rect 675220 111178 675248 114702
rect 675404 114479 675432 114786
rect 675390 114200 675446 114209
rect 675390 114135 675446 114144
rect 675404 113832 675432 114135
rect 675666 112568 675722 112577
rect 675666 112503 675722 112512
rect 675680 111996 675708 112503
rect 675482 111752 675538 111761
rect 675482 111687 675538 111696
rect 675496 111452 675524 111687
rect 675208 111172 675260 111178
rect 675208 111114 675260 111120
rect 675392 111172 675444 111178
rect 675392 111114 675444 111120
rect 675404 110772 675432 111114
rect 675116 110696 675168 110702
rect 675116 110638 675168 110644
rect 675392 110696 675444 110702
rect 675392 110638 675444 110644
rect 675404 110160 675432 110638
rect 675114 109032 675170 109041
rect 675114 108967 675170 108976
rect 675128 106758 675156 108967
rect 675758 108216 675814 108225
rect 675758 108151 675814 108160
rect 675772 107644 675800 108151
rect 675392 107568 675444 107574
rect 675392 107510 675444 107516
rect 675404 107100 675432 107510
rect 675116 106752 675168 106758
rect 675116 106694 675168 106700
rect 675392 106752 675444 106758
rect 675392 106694 675444 106700
rect 675404 106488 675432 106694
rect 674748 106276 674800 106282
rect 674748 106218 674800 106224
rect 675392 106276 675444 106282
rect 675392 106218 675444 106224
rect 672724 106140 672776 106146
rect 672724 106082 672776 106088
rect 675404 105808 675432 106218
rect 675758 104816 675814 104825
rect 675758 104751 675814 104760
rect 675772 104652 675800 104751
rect 675758 103184 675814 103193
rect 675758 103119 675814 103128
rect 675772 102816 675800 103119
rect 675758 101416 675814 101425
rect 675758 101351 675814 101360
rect 675772 100980 675800 101351
rect 664260 49564 664312 49570
rect 664260 49506 664312 49512
rect 672080 49564 672132 49570
rect 672080 49506 672132 49512
rect 664272 48521 664300 49506
rect 664258 48512 664314 48521
rect 664258 48447 664314 48456
rect 662418 47424 662474 47433
rect 662418 47359 662474 47368
rect 661144 46870 661512 46898
rect 612738 46472 612794 46481
rect 612738 46407 612794 46416
rect 611450 46336 611506 46345
rect 611450 46271 611506 46280
rect 661484 46238 661512 46870
rect 661472 46232 661524 46238
rect 610162 46200 610218 46209
rect 661472 46174 661524 46180
rect 610162 46135 610218 46144
rect 610070 45248 610126 45257
rect 610070 45183 610126 45192
rect 609978 41440 610034 41449
rect 609978 41375 610034 41384
rect 141698 40352 141754 40361
rect 141698 40287 141754 40296
rect 141712 39984 141740 40287
<< via2 >>
rect 203890 1007140 203946 1007176
rect 203890 1007120 203892 1007140
rect 203892 1007120 203944 1007140
rect 203944 1007120 203946 1007140
rect 99930 1006596 99986 1006632
rect 99930 1006576 99932 1006596
rect 99932 1006576 99984 1006596
rect 99984 1006576 99986 1006596
rect 86498 995696 86554 995752
rect 89626 995696 89682 995752
rect 92518 996512 92574 996568
rect 82358 995560 82414 995616
rect 85946 995560 86002 995616
rect 84658 995424 84714 995480
rect 80150 995016 80206 995072
rect 92610 995424 92666 995480
rect 93214 996376 93270 996432
rect 93122 995560 93178 995616
rect 104346 1006460 104402 1006496
rect 104346 1006440 104348 1006460
rect 104348 1006440 104400 1006460
rect 104400 1006440 104402 1006460
rect 104806 1006476 104808 1006496
rect 104808 1006476 104860 1006496
rect 104860 1006476 104862 1006496
rect 104806 1006440 104862 1006476
rect 100666 1006324 100722 1006360
rect 149702 1006340 149704 1006360
rect 149704 1006340 149756 1006360
rect 149756 1006340 149758 1006360
rect 100666 1006304 100668 1006324
rect 100668 1006304 100720 1006324
rect 100720 1006304 100722 1006324
rect 103610 1006188 103666 1006224
rect 103610 1006168 103612 1006188
rect 103612 1006168 103664 1006188
rect 103664 1006168 103666 1006188
rect 98274 1006068 98276 1006088
rect 98276 1006068 98328 1006088
rect 98328 1006068 98330 1006088
rect 98274 1006032 98330 1006068
rect 99102 1006068 99104 1006088
rect 99104 1006068 99156 1006088
rect 99156 1006068 99158 1006088
rect 99102 1006032 99158 1006068
rect 99470 1003332 99526 1003368
rect 99470 1003312 99472 1003332
rect 99472 1003312 99524 1003332
rect 99524 1003312 99526 1003332
rect 101494 1002244 101550 1002280
rect 101494 1002224 101496 1002244
rect 101496 1002224 101548 1002244
rect 101548 1002224 101550 1002244
rect 97262 996240 97318 996296
rect 100298 1002108 100354 1002144
rect 100298 1002088 100300 1002108
rect 100300 1002088 100352 1002108
rect 100352 1002088 100354 1002108
rect 102322 1002124 102324 1002144
rect 102324 1002124 102376 1002144
rect 102376 1002124 102378 1002144
rect 102322 1002088 102378 1002124
rect 101126 1001988 101128 1002008
rect 101128 1001988 101180 1002008
rect 101180 1001988 101182 1002008
rect 101126 1001952 101182 1001988
rect 101954 1001972 102010 1002008
rect 101954 1001952 101956 1001972
rect 101956 1001952 102008 1001972
rect 102008 1001952 102010 1001972
rect 92702 995016 92758 995072
rect 41786 968768 41842 968824
rect 41786 967272 41842 967328
rect 42062 965096 42118 965152
rect 41786 963328 41842 963384
rect 41786 962104 41842 962160
rect 41786 958296 41842 958352
rect 42062 957752 42118 957808
rect 32402 951632 32458 951688
rect 31022 938168 31078 938224
rect 34518 943744 34574 943800
rect 35806 943064 35862 943120
rect 35714 942656 35770 942712
rect 32402 937352 32458 937408
rect 37922 952176 37978 952232
rect 36542 936536 36598 936592
rect 41786 951632 41842 951688
rect 41970 951768 42026 951824
rect 41878 941840 41934 941896
rect 41786 941024 41842 941080
rect 37922 936128 37978 936184
rect 39946 933272 40002 933328
rect 41234 817944 41290 818000
rect 41326 817264 41382 817320
rect 40682 816856 40738 816912
rect 41694 940072 41750 940128
rect 41694 939256 41750 939312
rect 41970 937760 42026 937816
rect 42154 938984 42210 939040
rect 42062 935312 42118 935368
rect 42982 935720 43038 935776
rect 44822 941432 44878 941488
rect 47582 940616 47638 940672
rect 48962 942248 49018 942304
rect 103150 1006052 103206 1006088
rect 103150 1006032 103152 1006052
rect 103152 1006032 103204 1006052
rect 103204 1006032 103206 1006052
rect 108854 1006068 108856 1006088
rect 108856 1006068 108908 1006088
rect 108908 1006068 108910 1006088
rect 108854 1006032 108910 1006068
rect 103150 1004692 103206 1004728
rect 103150 1004672 103152 1004692
rect 103152 1004672 103204 1004692
rect 103204 1004672 103206 1004692
rect 106830 1002380 106886 1002416
rect 106830 1002360 106832 1002380
rect 106832 1002360 106884 1002380
rect 106884 1002360 106886 1002380
rect 106002 1002244 106058 1002280
rect 108486 1002260 108488 1002280
rect 108488 1002260 108540 1002280
rect 108540 1002260 108542 1002280
rect 106002 1002224 106004 1002244
rect 106004 1002224 106056 1002244
rect 106056 1002224 106058 1002244
rect 105634 1002124 105636 1002144
rect 105636 1002124 105688 1002144
rect 105688 1002124 105690 1002144
rect 105634 1002088 105690 1002124
rect 104346 1001988 104348 1002008
rect 104348 1001988 104400 1002008
rect 104400 1001988 104402 1002008
rect 104346 1001952 104402 1001988
rect 108486 1002224 108542 1002260
rect 107658 1002108 107714 1002144
rect 108026 1002124 108028 1002144
rect 108028 1002124 108080 1002144
rect 108080 1002124 108082 1002144
rect 107658 1002088 107660 1002108
rect 107660 1002088 107712 1002108
rect 107712 1002088 107714 1002108
rect 106462 1001972 106518 1002008
rect 107198 1001988 107200 1002008
rect 107200 1001988 107252 1002008
rect 107252 1001988 107254 1002008
rect 106462 1001952 106464 1001972
rect 106464 1001952 106516 1001972
rect 106516 1001952 106518 1001972
rect 107198 1001952 107254 1001988
rect 108026 1002088 108082 1002124
rect 108486 1001972 108542 1002008
rect 108486 1001952 108488 1001972
rect 108488 1001952 108540 1001972
rect 108540 1001952 108542 1001972
rect 109682 1001988 109684 1002008
rect 109684 1001988 109736 1002008
rect 109736 1001988 109738 1002008
rect 109682 1001952 109738 1001988
rect 117226 997056 117282 997112
rect 116306 996920 116362 996976
rect 149702 1006304 149758 1006340
rect 150898 1006340 150900 1006360
rect 150900 1006340 150952 1006360
rect 150952 1006340 150954 1006360
rect 150898 1006304 150954 1006340
rect 154118 1006324 154174 1006360
rect 154118 1006304 154120 1006324
rect 154120 1006304 154172 1006324
rect 154172 1006304 154174 1006324
rect 131762 995696 131818 995752
rect 133050 995696 133106 995752
rect 137926 995696 137982 995752
rect 142894 995696 142950 995752
rect 144826 997056 144882 997112
rect 144734 996920 144790 996976
rect 144182 995560 144238 995616
rect 137374 995424 137430 995480
rect 143998 995424 144054 995480
rect 136454 995288 136510 995344
rect 151726 1006204 151728 1006224
rect 151728 1006204 151780 1006224
rect 151780 1006204 151782 1006224
rect 151726 1006168 151782 1006204
rect 152094 1006188 152150 1006224
rect 152094 1006168 152096 1006188
rect 152096 1006168 152148 1006188
rect 152148 1006168 152150 1006188
rect 150898 1006052 150954 1006088
rect 150898 1006032 150900 1006052
rect 150900 1006032 150952 1006052
rect 150952 1006032 150954 1006052
rect 146942 995696 146998 995752
rect 148874 996240 148930 996296
rect 151266 998028 151322 998064
rect 151266 998008 151268 998028
rect 151268 998008 151320 998028
rect 151320 998008 151322 998028
rect 148322 995288 148378 995344
rect 132130 995152 132186 995208
rect 152554 997892 152610 997928
rect 152554 997872 152556 997892
rect 152556 997872 152608 997892
rect 152608 997872 152610 997892
rect 152922 998044 152924 998064
rect 152924 998044 152976 998064
rect 152976 998044 152978 998064
rect 152922 998008 152978 998044
rect 153750 997908 153752 997928
rect 153752 997908 153804 997928
rect 153804 997908 153806 997928
rect 153750 997872 153806 997908
rect 153382 997772 153384 997792
rect 153384 997772 153436 997792
rect 153436 997772 153438 997792
rect 153382 997736 153438 997772
rect 152738 995832 152794 995888
rect 151266 995152 151322 995208
rect 128450 995016 128506 995072
rect 159086 1006052 159142 1006088
rect 159086 1006032 159088 1006052
rect 159088 1006032 159140 1006052
rect 159140 1006032 159142 1006052
rect 160650 1006068 160652 1006088
rect 160652 1006068 160704 1006088
rect 160704 1006068 160706 1006088
rect 160650 1006032 160706 1006068
rect 159454 1004828 159510 1004864
rect 159454 1004808 159456 1004828
rect 159456 1004808 159508 1004828
rect 159508 1004808 159510 1004828
rect 159822 1004844 159824 1004864
rect 159824 1004844 159876 1004864
rect 159876 1004844 159878 1004864
rect 159822 1004808 159878 1004844
rect 160282 1004708 160284 1004728
rect 160284 1004708 160336 1004728
rect 160336 1004708 160338 1004728
rect 160282 1004672 160338 1004708
rect 160650 1004692 160706 1004728
rect 160650 1004672 160652 1004692
rect 160652 1004672 160704 1004692
rect 160704 1004672 160706 1004692
rect 154578 1002532 154580 1002552
rect 154580 1002532 154632 1002552
rect 154632 1002532 154634 1002552
rect 154578 1002496 154634 1002532
rect 158258 1002244 158314 1002280
rect 158258 1002224 158260 1002244
rect 158260 1002224 158312 1002244
rect 158312 1002224 158314 1002244
rect 157430 1002108 157486 1002144
rect 157430 1002088 157432 1002108
rect 157432 1002088 157484 1002108
rect 157484 1002088 157486 1002108
rect 157798 1002124 157800 1002144
rect 157800 1002124 157852 1002144
rect 157852 1002124 157854 1002144
rect 157798 1002088 157854 1002124
rect 156970 1001972 157026 1002008
rect 156970 1001952 156972 1001972
rect 156972 1001952 157024 1001972
rect 157024 1001952 157026 1001972
rect 158626 1001988 158628 1002008
rect 158628 1001988 158680 1002008
rect 158680 1001988 158682 1002008
rect 158626 1001952 158682 1001988
rect 154946 1000592 155002 1000648
rect 155774 999796 155830 999832
rect 155774 999776 155776 999796
rect 155776 999776 155828 999796
rect 155828 999776 155830 999796
rect 156142 997736 156198 997792
rect 167642 997192 167698 997248
rect 167550 996920 167606 996976
rect 184938 995696 184994 995752
rect 188802 995696 188858 995752
rect 189446 995696 189502 995752
rect 195242 996920 195298 996976
rect 195242 995832 195298 995888
rect 258170 1006476 258172 1006496
rect 258172 1006476 258224 1006496
rect 258224 1006476 258226 1006496
rect 195426 995968 195482 996024
rect 195058 995696 195114 995752
rect 179832 995288 179888 995344
rect 183834 995424 183890 995480
rect 182960 995152 183016 995208
rect 188158 995560 188214 995616
rect 194322 995560 194378 995616
rect 195978 995424 196034 995480
rect 202694 1006324 202750 1006360
rect 202694 1006304 202696 1006324
rect 202696 1006304 202748 1006324
rect 202748 1006304 202750 1006324
rect 210054 1006324 210110 1006360
rect 210054 1006304 210056 1006324
rect 210056 1006304 210108 1006324
rect 210108 1006304 210110 1006324
rect 204350 1006204 204352 1006224
rect 204352 1006204 204404 1006224
rect 204404 1006204 204406 1006224
rect 204350 1006168 204406 1006204
rect 201038 1006068 201040 1006088
rect 201040 1006068 201092 1006088
rect 201092 1006068 201094 1006088
rect 201038 1006032 201094 1006068
rect 201866 1006068 201868 1006088
rect 201868 1006068 201920 1006088
rect 201920 1006068 201922 1006088
rect 201866 1006032 201922 1006068
rect 202234 1004692 202290 1004728
rect 202234 1004672 202236 1004692
rect 202236 1004672 202288 1004692
rect 202288 1004672 202290 1004692
rect 200210 997228 200212 997248
rect 200212 997228 200264 997248
rect 200264 997228 200266 997248
rect 200210 997192 200266 997228
rect 200210 996240 200266 996296
rect 202050 995288 202106 995344
rect 191746 995016 191802 995072
rect 203522 1002124 203524 1002144
rect 203524 1002124 203576 1002144
rect 203576 1002124 203578 1002144
rect 203522 1002088 203578 1002124
rect 203062 1001988 203064 1002008
rect 203064 1001988 203116 1002008
rect 203116 1001988 203118 1002008
rect 203062 1001952 203118 1001988
rect 204718 1001972 204774 1002008
rect 204718 1001952 204720 1001972
rect 204720 1001952 204772 1001972
rect 204772 1001952 204774 1001972
rect 207202 1006068 207204 1006088
rect 207204 1006068 207256 1006088
rect 207256 1006068 207258 1006088
rect 207202 1006032 207258 1006068
rect 207570 1006052 207626 1006088
rect 207570 1006032 207572 1006052
rect 207572 1006032 207624 1006052
rect 207624 1006032 207626 1006052
rect 205178 1002244 205234 1002280
rect 205178 1002224 205180 1002244
rect 205180 1002224 205232 1002244
rect 205232 1002224 205234 1002244
rect 205914 1002108 205970 1002144
rect 205914 1002088 205916 1002108
rect 205916 1002088 205968 1002108
rect 205968 1002088 205970 1002108
rect 205546 1001988 205548 1002008
rect 205548 1001988 205600 1002008
rect 205600 1001988 205602 1002008
rect 205546 1001952 205602 1001988
rect 206742 1001972 206798 1002008
rect 206742 1001952 206744 1001972
rect 206744 1001952 206796 1001972
rect 206796 1001952 206798 1001972
rect 210422 1006188 210478 1006224
rect 210422 1006168 210424 1006188
rect 210424 1006168 210476 1006188
rect 210476 1006168 210478 1006188
rect 209594 1006068 209596 1006088
rect 209596 1006068 209648 1006088
rect 209648 1006068 209650 1006088
rect 209594 1006032 209650 1006068
rect 208766 1004828 208822 1004864
rect 208766 1004808 208768 1004828
rect 208768 1004808 208820 1004828
rect 208820 1004808 208822 1004828
rect 208398 1004692 208454 1004728
rect 208398 1004672 208400 1004692
rect 208400 1004672 208452 1004692
rect 208452 1004672 208454 1004692
rect 209226 1004708 209228 1004728
rect 209228 1004708 209280 1004728
rect 209280 1004708 209282 1004728
rect 209226 1004672 209282 1004708
rect 210422 1002124 210424 1002144
rect 210424 1002124 210476 1002144
rect 210476 1002124 210478 1002144
rect 210422 1002088 210478 1002124
rect 211618 1002244 211674 1002280
rect 211618 1002224 211620 1002244
rect 211620 1002224 211672 1002244
rect 211672 1002224 211674 1002244
rect 211250 1002108 211306 1002144
rect 211250 1002088 211252 1002108
rect 211252 1002088 211304 1002108
rect 211304 1002088 211306 1002108
rect 212078 1001972 212134 1002008
rect 212078 1001952 212080 1001972
rect 212080 1001952 212132 1001972
rect 212132 1001952 212134 1001972
rect 212538 1001988 212540 1002008
rect 212540 1001988 212592 1002008
rect 212592 1001988 212594 1002008
rect 212538 1001952 212594 1001988
rect 203522 995560 203578 995616
rect 215298 995016 215354 995072
rect 218886 996920 218942 996976
rect 246578 996920 246634 996976
rect 238574 995696 238630 995752
rect 240230 995696 240286 995752
rect 243818 995696 243874 995752
rect 247038 996240 247094 996296
rect 248326 997328 248382 997384
rect 236550 995560 236606 995616
rect 234388 995152 234444 995208
rect 232870 995016 232926 995072
rect 258170 1006440 258226 1006476
rect 254858 1006340 254860 1006360
rect 254860 1006340 254912 1006360
rect 254912 1006340 254914 1006360
rect 254858 1006304 254914 1006340
rect 255318 1006188 255374 1006224
rect 255318 1006168 255320 1006188
rect 255320 1006168 255372 1006188
rect 255372 1006168 255374 1006188
rect 257342 1006204 257344 1006224
rect 257344 1006204 257396 1006224
rect 257396 1006204 257398 1006224
rect 257342 1006168 257398 1006204
rect 252466 1006052 252522 1006088
rect 252466 1006032 252468 1006052
rect 252468 1006032 252520 1006052
rect 252520 1006032 252522 1006052
rect 253294 1006052 253350 1006088
rect 253294 1006032 253296 1006052
rect 253296 1006032 253348 1006052
rect 253348 1006032 253350 1006052
rect 254490 1002244 254546 1002280
rect 254490 1002224 254492 1002244
rect 254492 1002224 254544 1002244
rect 254544 1002224 254546 1002244
rect 249154 997192 249210 997248
rect 249706 996376 249762 996432
rect 254122 1001972 254178 1002008
rect 254122 1001952 254124 1001972
rect 254124 1001952 254176 1001972
rect 254176 1001952 254178 1001972
rect 253662 997772 253664 997792
rect 253664 997772 253716 997792
rect 253716 997772 253718 997792
rect 253662 997736 253718 997772
rect 256974 1006052 257030 1006088
rect 258538 1006068 258540 1006088
rect 258540 1006068 258592 1006088
rect 258592 1006068 258594 1006088
rect 256974 1006032 256976 1006052
rect 256976 1006032 257028 1006052
rect 257028 1006032 257030 1006052
rect 258538 1006032 258594 1006068
rect 258998 1006052 259054 1006088
rect 258998 1006032 259000 1006052
rect 259000 1006032 259052 1006052
rect 259052 1006032 259054 1006052
rect 261022 1006052 261078 1006088
rect 261022 1006032 261024 1006052
rect 261024 1006032 261076 1006052
rect 261076 1006032 261078 1006052
rect 255686 1002108 255742 1002144
rect 255686 1002088 255688 1002108
rect 255688 1002088 255740 1002108
rect 255740 1002088 255742 1002108
rect 256146 1002124 256148 1002144
rect 256148 1002124 256200 1002144
rect 256200 1002124 256202 1002144
rect 256146 1002088 256202 1002124
rect 256514 1001972 256570 1002008
rect 256514 1001952 256516 1001972
rect 256516 1001952 256568 1001972
rect 256568 1001952 256570 1001972
rect 261482 1002244 261538 1002280
rect 261482 1002224 261484 1002244
rect 261484 1002224 261536 1002244
rect 261536 1002224 261538 1002244
rect 261850 1002260 261852 1002280
rect 261852 1002260 261904 1002280
rect 261904 1002260 261906 1002280
rect 261850 1002224 261906 1002260
rect 259826 1002108 259882 1002144
rect 261850 1002124 261852 1002144
rect 261852 1002124 261904 1002144
rect 261904 1002124 261906 1002144
rect 259826 1002088 259828 1002108
rect 259828 1002088 259880 1002108
rect 259880 1002088 259882 1002108
rect 260194 1001988 260196 1002008
rect 260196 1001988 260248 1002008
rect 260248 1001988 260250 1002008
rect 260194 1001952 260250 1001988
rect 260654 1001972 260710 1002008
rect 260654 1001952 260656 1001972
rect 260656 1001952 260708 1001972
rect 260708 1001952 260710 1001972
rect 261850 1002088 261906 1002124
rect 262678 1002124 262680 1002144
rect 262680 1002124 262732 1002144
rect 262732 1002124 262734 1002144
rect 262678 1002088 262734 1002124
rect 263506 1002108 263562 1002144
rect 263506 1002088 263508 1002108
rect 263508 1002088 263560 1002108
rect 263560 1002088 263562 1002108
rect 263046 1001988 263048 1002008
rect 263048 1001988 263100 1002008
rect 263100 1001988 263102 1002008
rect 263046 1001952 263102 1001988
rect 263874 1001972 263930 1002008
rect 263874 1001952 263876 1001972
rect 263876 1001952 263928 1001972
rect 263928 1001952 263930 1001972
rect 257342 995016 257398 995072
rect 270406 996920 270462 996976
rect 298190 997736 298246 997792
rect 293498 995696 293554 995752
rect 298466 998144 298522 998200
rect 291750 995560 291806 995616
rect 298558 995560 298614 995616
rect 298742 996920 298798 996976
rect 300214 998144 300270 998200
rect 307298 1006460 307354 1006496
rect 307298 1006440 307300 1006460
rect 307300 1006440 307352 1006460
rect 307352 1006440 307354 1006460
rect 308126 1006476 308128 1006496
rect 308128 1006476 308180 1006496
rect 308180 1006476 308182 1006496
rect 308126 1006440 308182 1006476
rect 358174 1006460 358230 1006496
rect 358174 1006440 358176 1006460
rect 358176 1006440 358228 1006460
rect 358228 1006440 358230 1006460
rect 427542 1006460 427598 1006496
rect 427542 1006440 427544 1006460
rect 427544 1006440 427596 1006460
rect 427596 1006440 427598 1006460
rect 428370 1006476 428372 1006496
rect 428372 1006476 428424 1006496
rect 428424 1006476 428426 1006496
rect 428370 1006440 428426 1006476
rect 310610 1006324 310666 1006360
rect 310610 1006304 310612 1006324
rect 310612 1006304 310664 1006324
rect 310664 1006304 310666 1006324
rect 356058 1006340 356060 1006360
rect 356060 1006340 356112 1006360
rect 356112 1006340 356114 1006360
rect 356058 1006304 356114 1006340
rect 357714 1006324 357770 1006360
rect 357714 1006304 357716 1006324
rect 357716 1006304 357768 1006324
rect 357768 1006304 357770 1006324
rect 306470 1006204 306472 1006224
rect 306472 1006204 306524 1006224
rect 306524 1006204 306526 1006224
rect 306470 1006168 306526 1006204
rect 358910 1006204 358912 1006224
rect 358912 1006204 358964 1006224
rect 358964 1006204 358966 1006224
rect 358910 1006168 358966 1006204
rect 504546 1006340 504548 1006360
rect 504548 1006340 504600 1006360
rect 504600 1006340 504602 1006360
rect 304078 1006068 304080 1006088
rect 304080 1006068 304132 1006088
rect 304132 1006068 304134 1006088
rect 303250 997772 303252 997792
rect 303252 997772 303304 997792
rect 303304 997772 303306 997792
rect 303250 997736 303306 997772
rect 303250 996412 303252 996432
rect 303252 996412 303304 996432
rect 303304 996412 303306 996432
rect 303250 996376 303306 996412
rect 285954 995016 286010 995072
rect 304078 1006032 304134 1006068
rect 304906 1006068 304908 1006088
rect 304908 1006068 304960 1006088
rect 304960 1006068 304962 1006088
rect 304906 1006032 304962 1006068
rect 305274 1006052 305330 1006088
rect 305274 1006032 305276 1006052
rect 305276 1006032 305328 1006052
rect 305328 1006032 305330 1006052
rect 315118 1006052 315174 1006088
rect 315118 1006032 315120 1006052
rect 315120 1006032 315172 1006052
rect 315172 1006032 315174 1006052
rect 354494 1006052 354550 1006088
rect 354494 1006032 354496 1006052
rect 354496 1006032 354548 1006052
rect 354548 1006032 354550 1006052
rect 355230 1006032 355286 1006088
rect 356886 1006068 356888 1006088
rect 356888 1006068 356940 1006088
rect 356940 1006068 356942 1006088
rect 356886 1006032 356942 1006068
rect 358542 1006052 358598 1006088
rect 361394 1006068 361396 1006088
rect 361396 1006068 361448 1006088
rect 361448 1006068 361450 1006088
rect 358542 1006032 358544 1006052
rect 358544 1006032 358596 1006052
rect 358596 1006032 358598 1006052
rect 306930 1004828 306986 1004864
rect 306930 1004808 306932 1004828
rect 306932 1004808 306984 1004828
rect 306984 1004808 306986 1004828
rect 313830 1004828 313886 1004864
rect 313830 1004808 313832 1004828
rect 313832 1004808 313884 1004828
rect 313884 1004808 313886 1004828
rect 305734 1001972 305790 1002008
rect 305734 1001952 305736 1001972
rect 305736 1001952 305788 1001972
rect 305788 1001952 305790 1001972
rect 307758 1004692 307814 1004728
rect 307758 1004672 307760 1004692
rect 307760 1004672 307812 1004692
rect 307812 1004672 307814 1004692
rect 308586 1004708 308588 1004728
rect 308588 1004708 308640 1004728
rect 308640 1004708 308642 1004728
rect 308586 1004672 308642 1004708
rect 314658 1004708 314660 1004728
rect 314660 1004708 314712 1004728
rect 314712 1004708 314714 1004728
rect 314658 1004672 314714 1004708
rect 315486 1004692 315542 1004728
rect 315486 1004672 315488 1004692
rect 315488 1004672 315540 1004692
rect 315540 1004672 315542 1004692
rect 308954 1004572 308956 1004592
rect 308956 1004572 309008 1004592
rect 309008 1004572 309010 1004592
rect 308954 1004536 309010 1004572
rect 310150 1002108 310206 1002144
rect 310150 1002088 310152 1002108
rect 310152 1002088 310204 1002108
rect 310204 1002088 310206 1002108
rect 306102 1001988 306104 1002008
rect 306104 1001988 306156 1002008
rect 306156 1001988 306158 1002008
rect 306102 1001952 306158 1001988
rect 309322 1001988 309324 1002008
rect 309324 1001988 309376 1002008
rect 309376 1001988 309378 1002008
rect 309322 1001952 309378 1001988
rect 310150 1001952 310206 1002008
rect 311438 1001972 311494 1002008
rect 311438 1001952 311440 1001972
rect 311440 1001952 311492 1001972
rect 311492 1001952 311494 1001972
rect 312266 1001988 312268 1002008
rect 312268 1001988 312320 1002008
rect 312320 1001988 312322 1002008
rect 312266 1001952 312322 1001988
rect 313002 1001952 313058 1002008
rect 307022 995016 307078 995072
rect 360566 1005372 360622 1005408
rect 360566 1005352 360568 1005372
rect 360568 1005352 360620 1005372
rect 360620 1005352 360622 1005372
rect 360198 1005252 360200 1005272
rect 360200 1005252 360252 1005272
rect 360252 1005252 360254 1005272
rect 360198 1005216 360254 1005252
rect 356058 1004692 356114 1004728
rect 356058 1004672 356060 1004692
rect 356060 1004672 356112 1004692
rect 356112 1004672 356114 1004692
rect 356886 1004708 356888 1004728
rect 356888 1004708 356940 1004728
rect 356940 1004708 356942 1004728
rect 356886 1004672 356942 1004708
rect 358910 1001972 358966 1002008
rect 358910 1001952 358912 1001972
rect 358912 1001952 358964 1001972
rect 358964 1001952 358966 1001972
rect 359370 1001988 359372 1002008
rect 359372 1001988 359424 1002008
rect 359424 1001988 359426 1002008
rect 359370 1001952 359426 1001988
rect 361394 1006032 361450 1006068
rect 361026 1005388 361028 1005408
rect 361028 1005388 361080 1005408
rect 361080 1005388 361082 1005408
rect 361026 1005352 361082 1005388
rect 361854 1004708 361856 1004728
rect 361856 1004708 361908 1004728
rect 361908 1004708 361910 1004728
rect 361854 1004672 361910 1004708
rect 363418 1004844 363420 1004864
rect 363420 1004844 363472 1004864
rect 363472 1004844 363474 1004864
rect 363418 1004808 363474 1004844
rect 364246 1004828 364302 1004864
rect 364246 1004808 364248 1004828
rect 364248 1004808 364300 1004828
rect 364300 1004808 364302 1004828
rect 362590 1004692 362646 1004728
rect 362590 1004672 362592 1004692
rect 362592 1004672 362644 1004692
rect 362644 1004672 362646 1004692
rect 365074 1002108 365130 1002144
rect 365074 1002088 365076 1002108
rect 365076 1002088 365128 1002108
rect 365128 1002088 365130 1002108
rect 365442 1001972 365498 1002008
rect 365442 1001952 365444 1001972
rect 365444 1001952 365496 1001972
rect 365496 1001952 365498 1001972
rect 365902 1001988 365904 1002008
rect 365904 1001988 365956 1002008
rect 365956 1001988 365958 1002008
rect 365902 1001952 365958 1001988
rect 372434 997056 372490 997112
rect 372526 996920 372582 996976
rect 372342 996376 372398 996432
rect 374642 995560 374698 995616
rect 376022 995288 376078 995344
rect 504546 1006304 504602 1006340
rect 425150 1006188 425206 1006224
rect 425150 1006168 425152 1006188
rect 425152 1006168 425204 1006188
rect 425204 1006168 425206 1006188
rect 422666 1006068 422668 1006088
rect 422668 1006068 422720 1006088
rect 422720 1006068 422722 1006088
rect 380898 995424 380954 995480
rect 380162 995152 380218 995208
rect 422666 1006032 422722 1006068
rect 423494 1006052 423550 1006088
rect 428002 1006068 428004 1006088
rect 428004 1006068 428056 1006088
rect 428056 1006068 428058 1006088
rect 423494 1006032 423496 1006052
rect 423496 1006032 423548 1006052
rect 423548 1006032 423550 1006052
rect 428002 1006032 428058 1006068
rect 430026 1006052 430082 1006088
rect 430026 1006032 430028 1006052
rect 430028 1006032 430080 1006052
rect 430080 1006032 430082 1006052
rect 423862 1004572 423864 1004592
rect 423864 1004572 423916 1004592
rect 423916 1004572 423918 1004592
rect 421470 1001972 421526 1002008
rect 421470 1001952 421472 1001972
rect 421472 1001952 421524 1001972
rect 421524 1001952 421526 1001972
rect 383566 997464 383622 997520
rect 383658 997328 383714 997384
rect 381542 995696 381598 995752
rect 399942 997056 399998 997112
rect 400034 996920 400090 996976
rect 387890 995696 387946 995752
rect 388166 995696 388222 995752
rect 396630 995696 396686 995752
rect 394882 995560 394938 995616
rect 389362 995424 389418 995480
rect 385314 995288 385370 995344
rect 393962 995152 394018 995208
rect 423862 1004536 423918 1004572
rect 424690 1004028 424692 1004048
rect 424692 1004028 424744 1004048
rect 424744 1004028 424746 1004048
rect 424690 1003992 424746 1004028
rect 423494 1003892 423496 1003912
rect 423496 1003892 423548 1003912
rect 423548 1003892 423550 1003912
rect 423494 1003856 423550 1003892
rect 425978 1002532 425980 1002552
rect 425980 1002532 426032 1002552
rect 426032 1002532 426034 1002552
rect 425978 1002496 426034 1002532
rect 425978 1002108 426034 1002144
rect 425978 1002088 425980 1002108
rect 425980 1002088 426032 1002108
rect 426032 1002088 426034 1002108
rect 425150 1001972 425206 1002008
rect 426346 1001988 426348 1002008
rect 426348 1001988 426400 1002008
rect 426400 1001988 426402 1002008
rect 425150 1001952 425152 1001972
rect 425152 1001952 425204 1001972
rect 425204 1001952 425206 1001972
rect 426346 1001952 426402 1001988
rect 426806 1001972 426862 1002008
rect 426806 1001952 426808 1001972
rect 426808 1001952 426860 1001972
rect 426860 1001952 426862 1001972
rect 428830 999796 428886 999832
rect 428830 999776 428832 999796
rect 428832 999776 428884 999796
rect 428884 999776 428886 999796
rect 430854 998164 430910 998200
rect 430854 998144 430856 998164
rect 430856 998144 430908 998164
rect 430908 998144 430910 998164
rect 429658 998028 429714 998064
rect 429658 998008 429660 998028
rect 429660 998008 429712 998028
rect 429712 998008 429714 998028
rect 431682 998044 431684 998064
rect 431684 998044 431736 998064
rect 431736 998044 431738 998064
rect 431682 998008 431738 998044
rect 430394 997892 430450 997928
rect 430394 997872 430396 997892
rect 430396 997872 430448 997892
rect 430448 997872 430450 997892
rect 430854 997908 430856 997928
rect 430856 997908 430908 997928
rect 430908 997908 430910 997928
rect 430854 997872 430910 997908
rect 429198 997772 429200 997792
rect 429200 997772 429252 997792
rect 429252 997772 429254 997792
rect 429198 997736 429254 997772
rect 432418 997892 432474 997928
rect 432418 997872 432420 997892
rect 432420 997872 432472 997892
rect 432472 997872 432474 997892
rect 432878 997908 432880 997928
rect 432880 997908 432932 997928
rect 432932 997908 432934 997928
rect 432878 997872 432934 997908
rect 432050 997772 432052 997792
rect 432052 997772 432104 997792
rect 432104 997772 432106 997792
rect 432050 997736 432106 997772
rect 435362 997736 435418 997792
rect 432050 995832 432106 995888
rect 439686 996920 439742 996976
rect 439778 995732 439780 995752
rect 439780 995732 439832 995752
rect 439832 995732 439834 995752
rect 439778 995696 439834 995732
rect 505006 1006188 505062 1006224
rect 505006 1006168 505008 1006188
rect 505008 1006168 505060 1006188
rect 505060 1006168 505062 1006188
rect 505374 1006204 505376 1006224
rect 505376 1006204 505428 1006224
rect 505428 1006204 505430 1006224
rect 505374 1006168 505430 1006204
rect 459558 998280 459614 998336
rect 456062 995424 456118 995480
rect 499670 1006052 499726 1006088
rect 499670 1006032 499672 1006052
rect 499672 1006032 499724 1006052
rect 499724 1006032 499726 1006052
rect 500498 1006052 500554 1006088
rect 500498 1006032 500500 1006052
rect 500500 1006032 500552 1006052
rect 500552 1006032 500554 1006052
rect 502522 1006068 502524 1006088
rect 502524 1006068 502576 1006088
rect 502576 1006068 502578 1006088
rect 502522 1006032 502578 1006068
rect 462962 996240 463018 996296
rect 503350 1005252 503352 1005272
rect 503352 1005252 503404 1005272
rect 503404 1005252 503406 1005272
rect 503350 1005216 503406 1005252
rect 501326 1004828 501382 1004864
rect 501326 1004808 501328 1004828
rect 501328 1004808 501380 1004828
rect 501380 1004808 501382 1004828
rect 469402 998416 469458 998472
rect 472438 998416 472494 998472
rect 472714 998280 472770 998336
rect 472622 997192 472678 997248
rect 488906 996920 488962 996976
rect 472714 996376 472770 996432
rect 480810 995696 480866 995752
rect 482006 995696 482062 995752
rect 485594 995696 485650 995752
rect 482650 995560 482706 995616
rect 476394 995424 476450 995480
rect 459650 995288 459706 995344
rect 484122 995288 484178 995344
rect 454314 995152 454370 995208
rect 481638 995152 481694 995208
rect 449806 995016 449862 995072
rect 485962 995016 486018 995072
rect 446494 991480 446550 991536
rect 498474 1001952 498530 1002008
rect 500498 1004692 500554 1004728
rect 500498 1004672 500500 1004692
rect 500500 1004672 500552 1004692
rect 500552 1004672 500554 1004692
rect 500866 1004708 500868 1004728
rect 500868 1004708 500920 1004728
rect 500920 1004708 500922 1004728
rect 500866 1004672 500922 1004708
rect 503718 1003892 503720 1003912
rect 503720 1003892 503772 1003912
rect 503772 1003892 503774 1003912
rect 503718 1003856 503774 1003892
rect 501694 1001952 501750 1002008
rect 502522 1002224 502578 1002280
rect 503718 1002108 503774 1002144
rect 503718 1002088 503720 1002108
rect 503720 1002088 503772 1002108
rect 503772 1002088 503774 1002108
rect 508686 1005100 508742 1005136
rect 508686 1005080 508688 1005100
rect 508688 1005080 508740 1005100
rect 508740 1005080 508742 1005100
rect 507030 1004980 507032 1005000
rect 507032 1004980 507084 1005000
rect 507084 1004980 507086 1005000
rect 507030 1004944 507086 1004980
rect 508226 1004964 508282 1005000
rect 508226 1004944 508228 1004964
rect 508228 1004944 508280 1004964
rect 508280 1004944 508282 1004964
rect 507858 1004828 507914 1004864
rect 507858 1004808 507860 1004828
rect 507860 1004808 507912 1004828
rect 507912 1004808 507914 1004828
rect 507398 1004692 507454 1004728
rect 507398 1004672 507400 1004692
rect 507400 1004672 507452 1004692
rect 507452 1004672 507454 1004692
rect 509054 1004708 509056 1004728
rect 509056 1004708 509108 1004728
rect 509108 1004708 509110 1004728
rect 509054 1004672 509110 1004708
rect 505834 1001988 505836 1002008
rect 505836 1001988 505888 1002008
rect 505888 1001988 505890 1002008
rect 505834 1001952 505890 1001988
rect 506202 1001972 506258 1002008
rect 506202 1001952 506204 1001972
rect 506204 1001952 506256 1001972
rect 506256 1001952 506258 1001972
rect 506570 1001952 506626 1002008
rect 509514 1002108 509570 1002144
rect 509514 1002088 509516 1002108
rect 509516 1002088 509568 1002108
rect 509568 1002088 509570 1002108
rect 509882 1001988 509884 1002008
rect 509884 1001988 509936 1002008
rect 509936 1001988 509938 1002008
rect 509882 1001952 509938 1001988
rect 510342 1001972 510398 1002008
rect 510342 1001952 510344 1001972
rect 510344 1001952 510396 1001972
rect 510396 1001952 510398 1001972
rect 511078 992296 511134 992352
rect 555974 1006324 556030 1006360
rect 555974 1006304 555976 1006324
rect 555976 1006304 556028 1006324
rect 556028 1006304 556030 1006324
rect 557170 1006188 557226 1006224
rect 557170 1006168 557172 1006188
rect 557172 1006168 557224 1006188
rect 557224 1006168 557226 1006188
rect 550270 1006052 550326 1006088
rect 550270 1006032 550272 1006052
rect 550272 1006032 550324 1006052
rect 550324 1006032 550326 1006052
rect 551098 1006052 551154 1006088
rect 551098 1006032 551100 1006052
rect 551100 1006032 551152 1006052
rect 551152 1006032 551154 1006052
rect 552294 1006052 552350 1006088
rect 552294 1006032 552296 1006052
rect 552296 1006032 552348 1006052
rect 552348 1006032 552350 1006052
rect 556802 1006052 556858 1006088
rect 556802 1006032 556804 1006052
rect 556804 1006032 556856 1006052
rect 556856 1006032 556858 1006052
rect 516782 996920 516838 996976
rect 516690 996376 516746 996432
rect 516874 995560 516930 995616
rect 519266 995424 519322 995480
rect 516966 995152 517022 995208
rect 520186 996512 520242 996568
rect 524050 997192 524106 997248
rect 540886 996920 540942 996976
rect 526166 995696 526222 995752
rect 528006 995696 528062 995752
rect 532146 995696 532202 995752
rect 536562 995696 536618 995752
rect 529846 995560 529902 995616
rect 522394 995288 522450 995344
rect 534354 995288 534410 995344
rect 533066 995152 533122 995208
rect 538954 995424 539010 995480
rect 556342 1004708 556344 1004728
rect 556344 1004708 556396 1004728
rect 556396 1004708 556398 1004728
rect 556342 1004672 556398 1004708
rect 554778 1003312 554834 1003368
rect 552294 1002108 552350 1002144
rect 552294 1002088 552296 1002108
rect 552296 1002088 552348 1002108
rect 552348 1002088 552350 1002108
rect 553122 1002124 553124 1002144
rect 553124 1002124 553176 1002144
rect 553176 1002124 553178 1002144
rect 553122 1002088 553178 1002124
rect 551466 1001972 551522 1002008
rect 552662 1001988 552664 1002008
rect 552664 1001988 552716 1002008
rect 552716 1001988 552718 1002008
rect 551466 1001952 551468 1001972
rect 551468 1001952 551520 1001972
rect 551520 1001952 551522 1001972
rect 552662 1001952 552718 1001988
rect 553950 1002652 554006 1002688
rect 553950 1002632 553952 1002652
rect 553952 1002632 554004 1002652
rect 554004 1002632 554006 1002652
rect 554318 1002532 554320 1002552
rect 554320 1002532 554372 1002552
rect 554372 1002532 554374 1002552
rect 554318 1002496 554374 1002532
rect 553490 1001972 553546 1002008
rect 553490 1001952 553492 1001972
rect 553492 1001952 553544 1001972
rect 553544 1001952 553546 1001972
rect 555146 1001988 555148 1002008
rect 555148 1001988 555200 1002008
rect 555200 1001988 555202 1002008
rect 555146 1001952 555202 1001988
rect 557630 1004692 557686 1004728
rect 557630 1004672 557632 1004692
rect 557632 1004672 557684 1004692
rect 557684 1004672 557686 1004692
rect 559194 1002396 559196 1002416
rect 559196 1002396 559248 1002416
rect 559248 1002396 559250 1002416
rect 559194 1002360 559250 1002396
rect 558458 1002260 558460 1002280
rect 558460 1002260 558512 1002280
rect 558512 1002260 558514 1002280
rect 558458 1002224 558514 1002260
rect 557998 1001988 558000 1002008
rect 558000 1001988 558052 1002008
rect 558052 1001988 558054 1002008
rect 557998 1001952 558054 1001988
rect 558826 1001972 558882 1002008
rect 558826 1001952 558828 1001972
rect 558828 1001952 558880 1001972
rect 558880 1001952 558882 1001972
rect 557538 995852 557594 995888
rect 557538 995832 557540 995852
rect 557540 995832 557592 995852
rect 557592 995832 557594 995852
rect 559654 1002244 559710 1002280
rect 559654 1002224 559656 1002244
rect 559656 1002224 559708 1002244
rect 559708 1002224 559710 1002244
rect 560850 1002380 560906 1002416
rect 560850 1002360 560852 1002380
rect 560852 1002360 560904 1002380
rect 560904 1002360 560906 1002380
rect 560022 1002108 560078 1002144
rect 560022 1002088 560024 1002108
rect 560024 1002088 560076 1002108
rect 560076 1002088 560078 1002108
rect 560482 1002124 560484 1002144
rect 560484 1002124 560536 1002144
rect 560536 1002124 560538 1002144
rect 560482 1002088 560538 1002124
rect 561310 1001972 561366 1002008
rect 561310 1001952 561312 1001972
rect 561312 1001952 561364 1001972
rect 561364 1001952 561366 1001972
rect 561678 1001988 561680 1002008
rect 561680 1001988 561732 1002008
rect 561732 1001988 561734 1002008
rect 561678 1001952 561734 1001988
rect 568210 995696 568266 995752
rect 590566 996648 590622 996704
rect 590566 996512 590622 996568
rect 590566 996376 590622 996432
rect 618166 995152 618222 995208
rect 622398 996104 622454 996160
rect 627918 995696 627974 995752
rect 630310 995696 630366 995752
rect 631598 995696 631654 995752
rect 635186 995560 635242 995616
rect 626860 995152 626916 995208
rect 620282 995016 620338 995072
rect 629666 995016 629722 995072
rect 576306 990936 576362 990992
rect 62118 975976 62174 976032
rect 62118 962920 62174 962976
rect 62118 949864 62174 949920
rect 50342 939800 50398 939856
rect 62118 936980 62120 937000
rect 62120 936980 62172 937000
rect 62172 936980 62174 937000
rect 62118 936944 62174 936980
rect 44178 934496 44234 934552
rect 42890 934088 42946 934144
rect 42798 933680 42854 933736
rect 41878 932084 41880 932104
rect 41880 932084 41932 932104
rect 41932 932084 41934 932104
rect 41878 932048 41934 932084
rect 43442 932048 43498 932104
rect 41970 816448 42026 816504
rect 41786 815632 41842 815688
rect 41786 814852 41788 814872
rect 41788 814852 41840 814872
rect 41840 814852 41842 814872
rect 41786 814816 41842 814852
rect 41878 814000 41934 814056
rect 42154 812776 42210 812832
rect 33782 812368 33838 812424
rect 33046 810328 33102 810384
rect 32402 809104 32458 809160
rect 33046 802440 33102 802496
rect 35162 811960 35218 812016
rect 34426 810736 34482 810792
rect 40682 811552 40738 811608
rect 35254 808696 35310 808752
rect 35162 802712 35218 802768
rect 34426 802576 34482 802632
rect 35806 807272 35862 807328
rect 33782 800944 33838 801000
rect 42062 809512 42118 809568
rect 41786 807880 41842 807936
rect 41878 806248 41934 806304
rect 41786 804752 41842 804808
rect 42338 811144 42394 811200
rect 42430 796728 42486 796784
rect 42338 791968 42394 792024
rect 42154 788704 42210 788760
rect 42706 788160 42762 788216
rect 42430 788024 42486 788080
rect 41878 786936 41934 786992
rect 35806 774288 35862 774344
rect 42798 771976 42854 772032
rect 33782 769392 33838 769448
rect 32402 768576 32458 768632
rect 31022 767760 31078 767816
rect 30378 764088 30434 764144
rect 30378 763272 30434 763328
rect 32494 766536 32550 766592
rect 40682 768984 40738 769040
rect 33874 767352 33930 767408
rect 33874 758240 33930 758296
rect 41510 762864 41566 762920
rect 40682 757696 40738 757752
rect 41786 757016 41842 757072
rect 42430 757016 42486 757072
rect 41878 754840 41934 754896
rect 42614 754160 42670 754216
rect 41786 753072 41842 753128
rect 41786 750352 41842 750408
rect 42706 749264 42762 749320
rect 42614 746544 42670 746600
rect 41786 742328 41842 742384
rect 31482 731040 31538 731096
rect 31666 731040 31722 731096
rect 31574 730632 31630 730688
rect 31390 730224 31446 730280
rect 42890 769936 42946 769992
rect 42982 768304 43038 768360
rect 43258 765856 43314 765912
rect 42798 729272 42854 729328
rect 31022 726552 31078 726608
rect 40682 726144 40738 726200
rect 39302 725736 39358 725792
rect 35806 723696 35862 723752
rect 35714 723288 35770 723344
rect 39302 716080 39358 716136
rect 31022 715400 31078 715456
rect 42062 725192 42118 725248
rect 40774 724512 40830 724568
rect 40866 723288 40922 723344
rect 41510 720840 41566 720896
rect 41510 719652 41512 719672
rect 41512 719652 41564 719672
rect 41564 719652 41566 719672
rect 41510 719616 41566 719652
rect 42982 722744 43038 722800
rect 42062 713768 42118 713824
rect 42430 713224 42486 713280
rect 42522 710776 42578 710832
rect 42522 708464 42578 708520
rect 42062 706696 42118 706752
rect 42246 705064 42302 705120
rect 42522 705064 42578 705120
rect 42430 703704 42486 703760
rect 41786 702344 41842 702400
rect 41786 699352 41842 699408
rect 35622 688336 35678 688392
rect 35806 687656 35862 687712
rect 30286 687248 30342 687304
rect 39302 683576 39358 683632
rect 32402 682760 32458 682816
rect 31022 681536 31078 681592
rect 30470 676864 30526 676866
rect 30470 676812 30472 676864
rect 30472 676812 30524 676864
rect 30524 676812 30526 676864
rect 30470 676810 30526 676812
rect 35162 680312 35218 680368
rect 32402 671336 32458 671392
rect 41694 683052 41750 683088
rect 41694 683032 41696 683052
rect 41696 683032 41748 683052
rect 41748 683032 41750 683052
rect 39302 670928 39358 670984
rect 41694 681828 41750 681864
rect 41694 681808 41696 681828
rect 41696 681808 41748 681828
rect 41748 681808 41750 681828
rect 42798 681128 42854 681184
rect 41970 680720 42026 680776
rect 41786 670656 41842 670712
rect 42062 670656 42118 670712
rect 42430 670112 42486 670168
rect 41878 668480 41934 668536
rect 42890 679088 42946 679144
rect 41786 665352 41842 665408
rect 41786 664536 41842 664592
rect 42062 663312 42118 663368
rect 42706 661272 42762 661328
rect 42154 660456 42210 660512
rect 42522 660320 42578 660376
rect 42338 658280 42394 658336
rect 35622 644680 35678 644736
rect 35806 644680 35862 644736
rect 35162 640192 35218 640248
rect 32402 638152 32458 638208
rect 33782 637744 33838 637800
rect 33782 629856 33838 629912
rect 39302 639784 39358 639840
rect 40682 638968 40738 639024
rect 42890 638560 42946 638616
rect 40866 637336 40922 637392
rect 42798 635704 42854 635760
rect 40866 629176 40922 629232
rect 40682 629040 40738 629096
rect 35162 628496 35218 628552
rect 42522 625096 42578 625152
rect 42522 623736 42578 623792
rect 41786 621424 41842 621480
rect 42246 618976 42302 619032
rect 42154 616664 42210 616720
rect 42522 616800 42578 616856
rect 42522 614080 42578 614136
rect 41786 613400 41842 613456
rect 35806 601840 35862 601896
rect 35806 601432 35862 601488
rect 35714 601024 35770 601080
rect 35622 600616 35678 600672
rect 42798 599256 42854 599312
rect 39302 596944 39358 597000
rect 31666 594904 31722 594960
rect 33782 594904 33838 594960
rect 32402 593272 32458 593328
rect 31666 587152 31722 587208
rect 40866 596536 40922 596592
rect 40682 596128 40738 596184
rect 39302 585112 39358 585168
rect 42062 595992 42118 596048
rect 41510 591232 41566 591288
rect 41510 590008 41566 590064
rect 40866 585384 40922 585440
rect 40682 584588 40738 584644
rect 41602 584452 41658 584508
rect 42154 593952 42210 594008
rect 42154 584160 42210 584216
rect 41786 581712 41842 581768
rect 41786 580216 41842 580272
rect 41786 578992 41842 579048
rect 41786 577496 41842 577552
rect 42338 573960 42394 574016
rect 42154 573824 42210 573880
rect 42706 571512 42762 571568
rect 42154 570424 42210 570480
rect 35622 558320 35678 558376
rect 35806 558320 35862 558376
rect 35714 557912 35770 557968
rect 42890 594360 42946 594416
rect 42798 556416 42854 556472
rect 42798 556008 42854 556064
rect 40866 553832 40922 553888
rect 40682 553424 40738 553480
rect 32402 552608 32458 552664
rect 31022 551792 31078 551848
rect 31666 548120 31722 548176
rect 35806 546896 35862 546952
rect 32402 542816 32458 542872
rect 40774 552200 40830 552256
rect 40958 553016 41014 553072
rect 40866 545128 40922 545184
rect 40958 542952 41014 543008
rect 40774 542272 40830 542328
rect 42614 535880 42670 535936
rect 41786 534520 41842 534576
rect 42614 533840 42670 533896
rect 42338 532616 42394 532672
rect 41786 531392 41842 531448
rect 42338 529488 42394 529544
rect 42614 529352 42670 529408
rect 41786 430480 41842 430536
rect 42890 551520 42946 551576
rect 43074 549888 43130 549944
rect 43166 430888 43222 430944
rect 42798 428848 42854 428904
rect 42798 428440 42854 428496
rect 32402 425992 32458 426048
rect 31022 422320 31078 422376
rect 35162 425176 35218 425232
rect 32494 424360 32550 424416
rect 41786 419484 41842 419520
rect 41786 419464 41788 419484
rect 41788 419464 41840 419484
rect 41840 419464 41842 419484
rect 35162 414704 35218 414760
rect 32402 414568 32458 414624
rect 41878 411168 41934 411224
rect 41786 409400 41842 409456
rect 41786 406272 41842 406328
rect 42062 402464 42118 402520
rect 41786 401784 41842 401840
rect 41786 400016 41842 400072
rect 41786 399608 41842 399664
rect 41786 398792 41842 398848
rect 35622 387096 35678 387152
rect 35806 387504 35862 387560
rect 35806 387096 35862 387152
rect 35714 386688 35770 386744
rect 42890 423136 42946 423192
rect 42982 421504 43038 421560
rect 42798 385600 42854 385656
rect 42798 383560 42854 383616
rect 40866 382608 40922 382664
rect 37922 381384 37978 381440
rect 31022 380976 31078 381032
rect 33782 378120 33838 378176
rect 35806 377304 35862 377360
rect 33782 371864 33838 371920
rect 40682 379344 40738 379400
rect 37922 371320 37978 371376
rect 41510 376100 41566 376136
rect 41510 376080 41512 376100
rect 41512 376080 41564 376100
rect 41564 376080 41566 376100
rect 41786 370232 41842 370288
rect 41878 366288 41934 366344
rect 41970 363704 42026 363760
rect 41786 362888 41842 362944
rect 41786 360032 41842 360088
rect 41786 358672 41842 358728
rect 41786 356904 41842 356960
rect 41786 355680 41842 355736
rect 27618 344664 27674 344720
rect 35806 344256 35862 344312
rect 35714 343848 35770 343904
rect 43166 380704 43222 380760
rect 42982 380296 43038 380352
rect 43074 378664 43130 378720
rect 42890 341264 42946 341320
rect 42798 340856 42854 340912
rect 42798 340448 42854 340504
rect 31022 339360 31078 339416
rect 30378 334056 30434 334112
rect 30378 333260 30434 333296
rect 30378 333240 30380 333260
rect 30380 333240 30432 333260
rect 30432 333240 30434 333260
rect 32402 338136 32458 338192
rect 32402 327800 32458 327856
rect 31022 327664 31078 327720
rect 41786 324808 41842 324864
rect 41786 321136 41842 321192
rect 41786 319912 41842 319968
rect 41786 317328 41842 317384
rect 41786 315832 41842 315888
rect 41970 315424 42026 315480
rect 41878 313792 41934 313848
rect 41786 313112 41842 313168
rect 41786 312296 41842 312352
rect 35806 301552 35862 301608
rect 35806 300908 35808 300928
rect 35808 300908 35860 300928
rect 35860 300908 35862 300928
rect 35806 300872 35862 300908
rect 42982 336776 43038 336832
rect 43074 335144 43130 335200
rect 42890 298424 42946 298480
rect 42798 297608 42854 297664
rect 42798 297200 42854 297256
rect 35162 296384 35218 296440
rect 32402 294752 32458 294808
rect 35162 284824 35218 284880
rect 41786 281424 41842 281480
rect 41786 279792 41842 279848
rect 41786 278024 41842 278080
rect 41786 272992 41842 273048
rect 41786 272176 41842 272232
rect 41970 270408 42026 270464
rect 41786 269728 41842 269784
rect 41786 269048 41842 269104
rect 28354 258304 28410 258360
rect 31482 257488 31538 257544
rect 31666 257488 31722 257544
rect 31574 257080 31630 257136
rect 42890 295160 42946 295216
rect 42982 292304 43038 292360
rect 43166 291896 43222 291952
rect 62118 923752 62174 923808
rect 43534 806248 43590 806304
rect 42890 256400 42946 256456
rect 42798 254360 42854 254416
rect 31022 253408 31078 253464
rect 32402 253000 32458 253056
rect 31114 252184 31170 252240
rect 35806 246472 35862 246528
rect 41970 240624 42026 240680
rect 42706 238720 42762 238776
rect 41970 238448 42026 238504
rect 42706 237360 42762 237416
rect 41786 236680 41842 236736
rect 42430 232872 42486 232928
rect 42154 228928 42210 228984
rect 41970 227296 42026 227352
rect 28722 215056 28778 215112
rect 35806 214648 35862 214704
rect 35806 214240 35862 214296
rect 31022 210160 31078 210216
rect 43350 255584 43406 255640
rect 42982 252728 43038 252784
rect 43166 251912 43222 251968
rect 43074 250688 43130 250744
rect 43258 249056 43314 249112
rect 42890 213696 42946 213752
rect 41510 213424 41566 213480
rect 44178 815224 44234 815280
rect 43626 773608 43682 773664
rect 44270 813592 44326 813648
rect 44178 772384 44234 772440
rect 44362 809920 44418 809976
rect 44454 808288 44510 808344
rect 44546 772792 44602 772848
rect 44270 770752 44326 770808
rect 44362 767080 44418 767136
rect 44454 765448 44510 765504
rect 44730 770344 44786 770400
rect 44270 728864 44326 728920
rect 44178 721928 44234 721984
rect 44730 727640 44786 727696
rect 44546 727232 44602 727288
rect 44362 724376 44418 724432
rect 44454 722336 44510 722392
rect 44270 686024 44326 686080
rect 44270 685616 44326 685672
rect 44178 679904 44234 679960
rect 44178 643184 44234 643240
rect 44638 686432 44694 686488
rect 44546 684392 44602 684448
rect 44362 683984 44418 684040
rect 44270 643048 44326 643104
rect 44454 678680 44510 678736
rect 62118 910696 62174 910752
rect 62118 897776 62174 897832
rect 62118 884720 62174 884776
rect 62118 871664 62174 871720
rect 50434 773880 50490 773936
rect 44638 643728 44694 643784
rect 44638 642232 44694 642288
rect 44362 641416 44418 641472
rect 44454 636928 44510 636984
rect 44546 635296 44602 635352
rect 44178 600072 44234 600128
rect 44730 640600 44786 640656
rect 44638 599664 44694 599720
rect 44730 598032 44786 598088
rect 44270 597624 44326 597680
rect 44178 557232 44234 557288
rect 44362 595584 44418 595640
rect 44638 593136 44694 593192
rect 44454 592728 44510 592784
rect 44638 556824 44694 556880
rect 44362 555192 44418 555248
rect 44270 554784 44326 554840
rect 44270 554376 44326 554432
rect 44178 550296 44234 550352
rect 43626 430072 43682 430128
rect 44178 429256 44234 429312
rect 44454 551112 44510 551168
rect 44546 548664 44602 548720
rect 44638 429664 44694 429720
rect 44362 428032 44418 428088
rect 44362 427624 44418 427680
rect 44270 427216 44326 427272
rect 44178 385192 44234 385248
rect 44546 426808 44602 426864
rect 44454 421912 44510 421968
rect 44362 384784 44418 384840
rect 44638 421096 44694 421152
rect 44638 386008 44694 386064
rect 44546 383968 44602 384024
rect 44454 379072 44510 379128
rect 44546 377848 44602 377904
rect 44730 384376 44786 384432
rect 44638 343304 44694 343360
rect 44270 342896 44326 342952
rect 44178 342488 44234 342544
rect 44178 338000 44234 338056
rect 44546 342080 44602 342136
rect 44362 336368 44418 336424
rect 44454 334736 44510 334792
rect 44270 300056 44326 300112
rect 44362 299648 44418 299704
rect 44270 298832 44326 298888
rect 43534 231104 43590 231160
rect 44178 298016 44234 298072
rect 43902 290672 43958 290728
rect 44730 341672 44786 341728
rect 44546 299240 44602 299296
rect 44454 293528 44510 293584
rect 44546 291488 44602 291544
rect 44270 255992 44326 256048
rect 44178 255176 44234 255232
rect 44270 254768 44326 254824
rect 44178 251504 44234 251560
rect 43350 212880 43406 212936
rect 44730 253952 44786 254008
rect 44362 251096 44418 251152
rect 44546 249464 44602 249520
rect 44638 248240 44694 248296
rect 44270 212064 44326 212120
rect 41326 211792 41382 211848
rect 45006 300464 45062 300520
rect 45006 291080 45062 291136
rect 44914 248648 44970 248704
rect 54482 633392 54538 633448
rect 51814 289856 51870 289912
rect 62118 858608 62174 858664
rect 62118 845552 62174 845608
rect 62118 832496 62174 832552
rect 62118 819440 62174 819496
rect 62118 806520 62174 806576
rect 62118 793600 62174 793656
rect 62118 780408 62174 780464
rect 62118 767372 62174 767408
rect 62118 767352 62120 767372
rect 62120 767352 62172 767372
rect 62172 767352 62174 767372
rect 62118 754296 62174 754352
rect 62118 741240 62174 741296
rect 62118 728184 62174 728240
rect 62118 715264 62174 715320
rect 62762 702208 62818 702264
rect 62118 689152 62174 689208
rect 62118 676096 62174 676152
rect 62118 663040 62174 663096
rect 62118 649984 62174 650040
rect 62762 643456 62818 643512
rect 62118 637064 62174 637120
rect 62118 624008 62174 624064
rect 62118 610952 62174 611008
rect 62118 597896 62174 597952
rect 62118 584840 62174 584896
rect 62118 571784 62174 571840
rect 62118 558728 62174 558784
rect 62118 545808 62174 545864
rect 62118 532772 62174 532808
rect 62118 532752 62120 532772
rect 62120 532752 62172 532772
rect 62172 532752 62174 532772
rect 62118 519696 62174 519752
rect 62118 506640 62174 506696
rect 62118 493584 62174 493640
rect 62118 480528 62174 480584
rect 62118 467472 62174 467528
rect 62118 454552 62174 454608
rect 62118 441496 62174 441552
rect 62118 428440 62174 428496
rect 62118 415420 62120 415440
rect 62120 415420 62172 415440
rect 62172 415420 62174 415440
rect 62118 415384 62174 415420
rect 62118 402328 62174 402384
rect 62118 389272 62174 389328
rect 62118 376216 62174 376272
rect 62118 363296 62174 363352
rect 62118 350240 62174 350296
rect 62118 337184 62174 337240
rect 62118 324128 62174 324184
rect 62118 311072 62174 311128
rect 62118 298172 62174 298208
rect 62118 298152 62120 298172
rect 62120 298152 62172 298172
rect 62172 298152 62174 298172
rect 62118 285096 62174 285152
rect 371238 275304 371294 275360
rect 376482 270000 376538 270056
rect 379334 271224 379390 271280
rect 382186 274080 382242 274136
rect 383382 272720 383438 272776
rect 386050 269864 386106 269920
rect 388258 265784 388314 265840
rect 389178 267008 389234 267064
rect 391938 275440 391994 275496
rect 395710 271088 395766 271144
rect 394974 269728 395030 269784
rect 398470 268640 398526 268696
rect 401046 273944 401102 274000
rect 402518 268368 402574 268424
rect 402058 266464 402114 266520
rect 404174 272584 404230 272640
rect 404358 267008 404414 267064
rect 404726 266328 404782 266384
rect 405186 265648 405242 265704
rect 406106 271360 406162 271416
rect 405738 268504 405794 268560
rect 405738 266464 405794 266520
rect 406934 272448 406990 272504
rect 409694 275168 409750 275224
rect 407394 267280 407450 267336
rect 407854 265512 407910 265568
rect 411902 273808 411958 273864
rect 410982 267144 411038 267200
rect 412270 267008 412326 267064
rect 411902 266328 411958 266384
rect 448978 271360 449034 271416
rect 457994 267280 458050 267336
rect 537574 275304 537630 275360
rect 544658 275440 544714 275496
rect 554778 270000 554834 270056
rect 562414 271224 562470 271280
rect 569498 274080 569554 274136
rect 572994 272720 573050 272776
rect 579618 269864 579674 269920
rect 585138 265784 585194 265840
rect 604918 271088 604974 271144
rect 603078 269728 603134 269784
rect 396998 264152 397054 264208
rect 401230 264172 401286 264208
rect 612738 268640 612794 268696
rect 401230 264152 401232 264172
rect 401232 264152 401284 264172
rect 401284 264152 401286 264172
rect 619086 273944 619142 274000
rect 622398 268504 622454 268560
rect 629758 273808 629814 273864
rect 628562 272584 628618 272640
rect 623778 268368 623834 268424
rect 635646 272448 635702 272504
rect 630678 265648 630734 265704
rect 640430 275168 640486 275224
rect 645858 267144 645914 267200
rect 637578 265512 637634 265568
rect 415306 262268 415362 262304
rect 415306 262248 415308 262268
rect 415308 262248 415360 262268
rect 415360 262248 415362 262268
rect 414202 259120 414258 259176
rect 189078 258576 189134 258632
rect 415306 255856 415362 255912
rect 185214 253136 185270 253192
rect 414386 252728 414442 252784
rect 414202 249464 414258 249520
rect 190366 247968 190422 248024
rect 189722 247152 189778 247208
rect 64142 229880 64198 229936
rect 57886 229744 57942 229800
rect 47214 212472 47270 212528
rect 44730 211248 44786 211304
rect 50066 210568 50122 210624
rect 42798 209208 42854 209264
rect 39302 208528 39358 208584
rect 31298 204856 31354 204912
rect 31114 204448 31170 204504
rect 35806 203224 35862 203280
rect 31022 199280 31078 199336
rect 39302 197648 39358 197704
rect 41878 197104 41934 197160
rect 41786 195200 41842 195256
rect 41786 190168 41842 190224
rect 42154 187312 42210 187368
rect 44178 207984 44234 208040
rect 42890 207576 42946 207632
rect 43350 206760 43406 206816
rect 43166 206352 43222 206408
rect 42982 205944 43038 206000
rect 43258 205128 43314 205184
rect 43442 205536 43498 205592
rect 41878 184184 41934 184240
rect 41786 182960 41842 183016
rect 55126 222808 55182 222864
rect 56874 221448 56930 221504
rect 59266 226888 59322 226944
rect 58622 222944 58678 223000
rect 62762 227024 62818 227080
rect 61934 224168 61990 224224
rect 72974 227160 73030 227216
rect 72054 224440 72110 224496
rect 69478 224304 69534 224360
rect 66994 221584 67050 221640
rect 67546 220088 67602 220144
rect 70214 221720 70270 221776
rect 73710 221856 73766 221912
rect 90546 228384 90602 228440
rect 86866 228248 86922 228304
rect 74446 220224 74502 220280
rect 78494 224576 78550 224632
rect 89534 225528 89590 225584
rect 93030 225664 93086 225720
rect 92294 223080 92350 223136
rect 99010 223216 99066 223272
rect 175002 241596 175058 241632
rect 175002 241576 175004 241596
rect 175004 241576 175056 241596
rect 175056 241576 175058 241596
rect 189078 237396 189080 237416
rect 189080 237396 189132 237416
rect 189132 237396 189134 237416
rect 189078 237360 189134 237396
rect 117962 218592 118018 218648
rect 191102 247288 191158 247344
rect 415306 246336 415362 246392
rect 414386 243072 414442 243128
rect 414938 239944 414994 240000
rect 414202 236680 414258 236736
rect 415306 233552 415362 233608
rect 192390 222808 192446 222864
rect 194046 222944 194102 223000
rect 193402 221448 193458 221504
rect 194782 229744 194838 229800
rect 196162 229880 196218 229936
rect 195794 226888 195850 226944
rect 195426 224168 195482 224224
rect 196622 230288 196678 230344
rect 197266 227024 197322 227080
rect 197726 221584 197782 221640
rect 196622 220088 196678 220144
rect 199014 230288 199070 230344
rect 199750 224440 199806 224496
rect 200118 224304 200174 224360
rect 199106 221720 199162 221776
rect 201498 227160 201554 227216
rect 200578 221856 200634 221912
rect 202602 224576 202658 224632
rect 201590 220224 201646 220280
rect 206558 228248 206614 228304
rect 207938 228384 207994 228440
rect 208030 223080 208086 223136
rect 208674 225528 208730 225584
rect 210054 225664 210110 225720
rect 211158 223216 211214 223272
rect 375838 230016 375894 230072
rect 376942 230288 376998 230344
rect 378690 229880 378746 229936
rect 377678 224712 377734 224768
rect 376206 223216 376262 223272
rect 379058 223080 379114 223136
rect 380162 229744 380218 229800
rect 380530 227296 380586 227352
rect 380346 220360 380402 220416
rect 381542 230152 381598 230208
rect 381910 224576 381966 224632
rect 383014 227160 383070 227216
rect 382186 220224 382242 220280
rect 384026 224440 384082 224496
rect 384854 220088 384910 220144
rect 386234 225936 386290 225992
rect 387246 228656 387302 228712
rect 388350 227024 388406 227080
rect 389178 220496 389234 220552
rect 389362 222944 389418 223000
rect 390466 222808 390522 222864
rect 394054 225800 394110 225856
rect 392858 221720 392914 221776
rect 396446 225664 396502 225720
rect 397182 221584 397238 221640
rect 399390 228520 399446 228576
rect 400494 225528 400550 225584
rect 402610 228384 402666 228440
rect 401138 224304 401194 224360
rect 400678 221856 400734 221912
rect 405002 221448 405058 221504
rect 406106 224168 406162 224224
rect 407946 226888 408002 226944
rect 428646 230288 428702 230344
rect 411074 228248 411130 228304
rect 478142 230152 478198 230208
rect 486422 230016 486478 230072
rect 493322 229880 493378 229936
rect 496082 229744 496138 229800
rect 490194 224712 490250 224768
rect 487802 223216 487858 223272
rect 489458 220360 489514 220416
rect 494150 223080 494206 223136
rect 495622 220496 495678 220552
rect 496910 227296 496966 227352
rect 499578 224576 499634 224632
rect 498658 220224 498714 220280
rect 502522 227160 502578 227216
rect 505374 224440 505430 224496
rect 507214 220088 507270 220144
rect 507214 219408 507270 219464
rect 513378 228656 513434 228712
rect 510710 225936 510766 225992
rect 515494 227024 515550 227080
rect 517978 222944 518034 223000
rect 520462 222808 520518 222864
rect 492586 216824 492642 216880
rect 489090 216688 489146 216744
rect 525890 221720 525946 221776
rect 528926 225800 528982 225856
rect 528098 221856 528154 221912
rect 534078 225664 534134 225720
rect 532974 216960 533030 217016
rect 536010 221584 536066 221640
rect 541530 228520 541586 228576
rect 544014 225528 544070 225584
rect 545762 224304 545818 224360
rect 549258 228384 549314 228440
rect 546682 221448 546738 221504
rect 561678 226888 561734 226944
rect 556710 224168 556766 224224
rect 564438 228248 564494 228304
rect 648618 267008 648674 267064
rect 578882 216144 578938 216200
rect 578422 211656 578478 211712
rect 578514 210160 578570 210216
rect 579250 214648 579306 214704
rect 578974 213152 579030 213208
rect 579526 208664 579582 208720
rect 578790 207168 578846 207224
rect 579434 205672 579490 205728
rect 578882 204176 578938 204232
rect 579250 202680 579306 202736
rect 578238 201184 578294 201240
rect 578422 199688 578478 199744
rect 579066 198192 579122 198248
rect 579526 196696 579582 196752
rect 579526 195236 579528 195256
rect 579528 195236 579580 195256
rect 579580 195236 579582 195256
rect 579526 195200 579582 195236
rect 579526 193568 579582 193624
rect 579526 192072 579582 192128
rect 579250 190576 579306 190632
rect 578238 189080 578294 189136
rect 579250 187584 579306 187640
rect 578882 184592 578938 184648
rect 578238 177112 578294 177168
rect 578330 175616 578386 175672
rect 578882 180104 578938 180160
rect 578422 174120 578478 174176
rect 579526 186088 579582 186144
rect 579434 183096 579490 183152
rect 579526 181600 579582 181656
rect 579342 178608 579398 178664
rect 578790 172624 578846 172680
rect 578698 171128 578754 171184
rect 578606 166504 578662 166560
rect 578238 164328 578294 164384
rect 578882 157528 578938 157584
rect 579158 162016 579214 162072
rect 579434 169496 579490 169552
rect 579342 168000 579398 168056
rect 579526 163512 579582 163568
rect 579250 160520 579306 160576
rect 579066 159024 579122 159080
rect 578974 156032 579030 156088
rect 578330 154536 578386 154592
rect 578514 148588 578516 148608
rect 578516 148588 578568 148608
rect 578568 148588 578570 148608
rect 578514 148552 578570 148588
rect 578698 145424 578754 145480
rect 578698 142432 578754 142488
rect 578882 131960 578938 132016
rect 578330 130500 578332 130520
rect 578332 130500 578384 130520
rect 578384 130500 578386 130520
rect 578330 130464 578386 130500
rect 579158 139440 579214 139496
rect 579526 153040 579582 153096
rect 579434 151580 579436 151600
rect 579436 151580 579488 151600
rect 579488 151580 579490 151600
rect 579434 151544 579490 151580
rect 579434 150048 579490 150104
rect 579526 146956 579528 146976
rect 579528 146956 579580 146976
rect 579580 146956 579582 146976
rect 579526 146920 579582 146956
rect 579526 143928 579582 143984
rect 579342 140936 579398 140992
rect 579526 137964 579582 138000
rect 579526 137944 579528 137964
rect 579528 137944 579580 137964
rect 579580 137944 579582 137964
rect 579526 136484 579528 136504
rect 579528 136484 579580 136504
rect 579580 136484 579582 136504
rect 579526 136448 579582 136484
rect 579250 134952 579306 135008
rect 579066 133456 579122 133512
rect 578974 128968 579030 129024
rect 579526 127472 579582 127528
rect 578698 126012 578700 126032
rect 578700 126012 578752 126032
rect 578752 126012 578754 126032
rect 578698 125976 578754 126012
rect 578422 124480 578478 124536
rect 579250 122848 579306 122904
rect 579250 119856 579306 119912
rect 578514 118360 578570 118416
rect 578698 110880 578754 110936
rect 578790 107888 578846 107944
rect 578238 104896 578294 104952
rect 578330 101904 578386 101960
rect 578698 100308 578700 100328
rect 578700 100308 578752 100328
rect 578752 100308 578754 100328
rect 578698 100272 578754 100308
rect 578698 97280 578754 97336
rect 578514 95784 578570 95840
rect 578606 94288 578662 94344
rect 52182 52400 52238 52456
rect 150300 52400 150356 52456
rect 281446 50496 281502 50552
rect 216126 50360 216182 50416
rect 85118 50224 85174 50280
rect 142342 44240 142398 44296
rect 187514 42064 187570 42120
rect 307298 43424 307354 43480
rect 310104 42336 310160 42392
rect 361946 42064 362002 42120
rect 365074 42064 365130 42120
rect 543002 50224 543058 50280
rect 473174 47640 473230 47696
rect 412454 46688 412510 46744
rect 470138 46416 470194 46472
rect 415122 46144 415178 46200
rect 419722 45192 419778 45248
rect 460570 42064 460626 42120
rect 416686 41792 416742 41848
rect 471610 42064 471666 42120
rect 579526 121388 579528 121408
rect 579528 121388 579580 121408
rect 579580 121388 579582 121408
rect 579526 121352 579582 121388
rect 603078 209480 603134 209536
rect 603170 208528 603226 208584
rect 603078 207440 603134 207496
rect 603078 206488 603134 206544
rect 603078 205400 603134 205456
rect 603170 204448 603226 204504
rect 603078 203360 603134 203416
rect 603078 202408 603134 202464
rect 603078 201320 603134 201376
rect 603170 200368 603226 200424
rect 603078 199280 603134 199336
rect 603078 198328 603134 198384
rect 603078 197240 603134 197296
rect 603170 196288 603226 196344
rect 603078 195236 603080 195256
rect 603080 195236 603132 195256
rect 603132 195236 603134 195256
rect 603078 195200 603134 195236
rect 603078 194248 603134 194304
rect 603078 193160 603134 193216
rect 603078 192208 603134 192264
rect 603078 191120 603134 191176
rect 603170 190168 603226 190224
rect 603078 189116 603080 189136
rect 603080 189116 603132 189136
rect 603132 189116 603134 189136
rect 603078 189080 603134 189116
rect 603078 188128 603134 188184
rect 603078 187040 603134 187096
rect 603170 186088 603226 186144
rect 603078 185000 603134 185056
rect 603078 184048 603134 184104
rect 603078 182960 603134 183016
rect 603170 182008 603226 182064
rect 603078 180920 603134 180976
rect 603078 179968 603134 180024
rect 603078 178880 603134 178936
rect 603170 177928 603226 177984
rect 603078 176840 603134 176896
rect 603078 175888 603134 175944
rect 603078 174800 603134 174856
rect 603722 173848 603778 173904
rect 603078 172760 603134 172816
rect 603078 171808 603134 171864
rect 603170 170720 603226 170776
rect 603078 169788 603134 169824
rect 603078 169768 603080 169788
rect 603080 169768 603132 169788
rect 603132 169768 603134 169788
rect 603078 168680 603134 168736
rect 603078 167728 603134 167784
rect 603078 165688 603134 165744
rect 603078 164600 603134 164656
rect 603814 166640 603870 166696
rect 603078 163648 603134 163704
rect 603078 162560 603134 162616
rect 603722 161608 603778 161664
rect 579526 116864 579582 116920
rect 579434 115368 579490 115424
rect 579250 113872 579306 113928
rect 579526 112376 579582 112432
rect 579526 109384 579582 109440
rect 579434 106392 579490 106448
rect 579342 103436 579344 103456
rect 579344 103436 579396 103456
rect 579396 103436 579398 103456
rect 579342 103400 579398 103436
rect 579526 98776 579582 98832
rect 579526 92792 579582 92848
rect 579526 91296 579582 91352
rect 579526 89800 579582 89856
rect 579526 88304 579582 88360
rect 579526 86808 579582 86864
rect 579526 85312 579582 85368
rect 579526 83816 579582 83872
rect 579158 82320 579214 82376
rect 579526 80860 579528 80880
rect 579528 80860 579580 80880
rect 579580 80860 579582 80880
rect 579526 80824 579582 80860
rect 579066 79328 579122 79384
rect 579526 77832 579582 77888
rect 578974 76200 579030 76256
rect 578882 73208 578938 73264
rect 578698 68720 578754 68776
rect 578698 64232 578754 64288
rect 578698 61240 578754 61296
rect 578882 59744 578938 59800
rect 578882 58248 578938 58304
rect 578238 55256 578294 55312
rect 578882 56752 578938 56808
rect 578330 53760 578386 53816
rect 579526 74704 579582 74760
rect 579526 71732 579582 71768
rect 579526 71712 579528 71732
rect 579528 71712 579580 71732
rect 579580 71712 579582 71732
rect 579250 70252 579252 70272
rect 579252 70252 579304 70272
rect 579304 70252 579306 70272
rect 579250 70216 579306 70252
rect 579526 67224 579582 67280
rect 579526 65728 579582 65784
rect 579526 62736 579582 62792
rect 603078 160520 603134 160576
rect 603078 159568 603134 159624
rect 603170 158480 603226 158536
rect 603078 157528 603134 157584
rect 603078 156440 603134 156496
rect 603078 155488 603134 155544
rect 603170 154400 603226 154456
rect 603078 153448 603134 153504
rect 603078 152360 603134 152416
rect 603078 151408 603134 151464
rect 603078 150320 603134 150376
rect 603078 148280 603134 148336
rect 603078 147328 603134 147384
rect 603906 149368 603962 149424
rect 603170 146240 603226 146296
rect 603722 145288 603778 145344
rect 603078 144200 603134 144256
rect 603078 142180 603134 142216
rect 603078 142160 603080 142180
rect 603080 142160 603132 142180
rect 603132 142160 603134 142180
rect 603078 141208 603134 141264
rect 603078 140120 603134 140176
rect 603170 139168 603226 139224
rect 603078 138100 603134 138136
rect 603078 138080 603080 138100
rect 603080 138080 603132 138100
rect 603132 138080 603134 138100
rect 603078 137128 603134 137184
rect 603078 136040 603134 136096
rect 603170 135088 603226 135144
rect 603078 134000 603134 134056
rect 603814 143248 603870 143304
rect 603078 133048 603134 133104
rect 603078 131960 603134 132016
rect 603170 131008 603226 131064
rect 603078 129920 603134 129976
rect 603078 128968 603134 129024
rect 603078 127880 603134 127936
rect 603170 126928 603226 126984
rect 603078 125840 603134 125896
rect 603078 124888 603134 124944
rect 603078 123800 603134 123856
rect 603170 122884 603172 122904
rect 603172 122884 603224 122904
rect 603224 122884 603226 122904
rect 603170 122848 603226 122884
rect 603078 121760 603134 121816
rect 603078 120808 603134 120864
rect 603078 119720 603134 119776
rect 603722 118768 603778 118824
rect 603078 117680 603134 117736
rect 602342 116728 602398 116784
rect 603078 115640 603134 115696
rect 603170 114688 603226 114744
rect 603078 113600 603134 113656
rect 603078 112648 603134 112704
rect 603078 110608 603134 110664
rect 603078 109520 603134 109576
rect 603078 108568 603134 108624
rect 603170 107480 603226 107536
rect 603078 106528 603134 106584
rect 603078 105440 603134 105496
rect 603078 104488 603134 104544
rect 603170 103400 603226 103456
rect 603078 102448 603134 102504
rect 603078 101360 603134 101416
rect 603446 100408 603502 100464
rect 603814 111560 603870 111616
rect 620926 216688 620982 216744
rect 622030 216824 622086 216880
rect 623962 219408 624018 219464
rect 628930 216960 628986 217016
rect 646134 229608 646190 229664
rect 647146 213016 647202 213072
rect 648526 213016 648582 213072
rect 651654 975840 651710 975896
rect 652022 962512 652078 962568
rect 651562 949320 651618 949376
rect 651562 936128 651618 936184
rect 651562 922664 651618 922720
rect 651562 909492 651618 909528
rect 651562 909472 651564 909492
rect 651564 909472 651616 909492
rect 651616 909472 651618 909492
rect 651562 896144 651618 896200
rect 652022 882816 652078 882872
rect 651562 869624 651618 869680
rect 652574 856296 652630 856352
rect 651562 842968 651618 843024
rect 651562 829776 651618 829832
rect 651562 816448 651618 816504
rect 651562 803256 651618 803312
rect 651654 789928 651710 789984
rect 651562 776600 651618 776656
rect 651562 763272 651618 763328
rect 651562 750080 651618 750136
rect 651562 736752 651618 736808
rect 652022 723424 652078 723480
rect 651562 710232 651618 710288
rect 652022 696904 652078 696960
rect 651838 683576 651894 683632
rect 651562 670384 651618 670440
rect 651562 657056 651618 657112
rect 651562 643728 651618 643784
rect 651562 630536 651618 630592
rect 651562 603880 651618 603936
rect 651562 590708 651618 590744
rect 651562 590688 651564 590708
rect 651564 590688 651616 590708
rect 651616 590688 651618 590708
rect 652390 617208 652446 617264
rect 651562 577360 651618 577416
rect 652114 564032 652170 564088
rect 651562 550840 651618 550896
rect 651562 537512 651618 537568
rect 651562 524184 651618 524240
rect 651562 510992 651618 511048
rect 651562 497664 651618 497720
rect 651562 484472 651618 484528
rect 651654 471144 651710 471200
rect 651562 457816 651618 457872
rect 651562 444488 651618 444544
rect 651562 431296 651618 431352
rect 651562 417968 651618 418024
rect 652022 404640 652078 404696
rect 651562 391448 651618 391504
rect 651562 378156 651564 378176
rect 651564 378156 651616 378176
rect 651616 378156 651618 378176
rect 651562 378120 651618 378156
rect 652022 364792 652078 364848
rect 651562 351600 651618 351656
rect 651654 338272 651710 338328
rect 651562 324944 651618 325000
rect 651562 311752 651618 311808
rect 652022 298424 652078 298480
rect 651562 285232 651618 285288
rect 663890 218592 663946 218648
rect 665454 209752 665510 209808
rect 666558 193976 666614 194032
rect 666558 190576 666614 190632
rect 675758 966456 675814 966512
rect 675758 966184 675814 966240
rect 675758 964960 675814 965016
rect 675390 963328 675446 963384
rect 674746 958976 674802 959032
rect 666834 204176 666890 204232
rect 666834 200776 666890 200832
rect 666742 199008 666798 199064
rect 666558 188944 666614 189000
rect 666558 185544 666614 185600
rect 666558 153312 666614 153368
rect 666558 151816 666614 151872
rect 666558 151544 666614 151600
rect 666558 149912 666614 149968
rect 666558 142024 666614 142080
rect 666558 139712 666614 139768
rect 667938 209208 667994 209264
rect 667938 205808 667994 205864
rect 667938 199008 667994 199064
rect 667938 195608 667994 195664
rect 667938 183776 667994 183832
rect 668030 180376 668086 180432
rect 667938 178780 667940 178800
rect 667940 178780 667992 178800
rect 667992 178780 667994 178800
rect 667938 178744 667994 178780
rect 667938 175344 667994 175400
rect 667938 173576 667994 173632
rect 667938 171128 667994 171184
rect 667938 163512 667994 163568
rect 667938 161472 667994 161528
rect 667938 158344 667994 158400
rect 667938 154944 667994 155000
rect 667938 143112 667994 143168
rect 667938 138080 667994 138136
rect 667938 134680 667994 134736
rect 666558 132368 666614 132424
rect 666558 129512 666614 129568
rect 667938 127916 667940 127936
rect 667940 127916 667992 127936
rect 667992 127916 667994 127936
rect 667938 127880 667994 127916
rect 667938 124480 667994 124536
rect 667938 122848 667994 122904
rect 666558 122712 666614 122768
rect 666558 119448 666614 119504
rect 667938 117716 667940 117736
rect 667940 117716 667992 117736
rect 667992 117716 667994 117736
rect 667938 117680 667994 117716
rect 667938 109284 667940 109304
rect 667940 109284 667992 109304
rect 667992 109284 667994 109304
rect 667938 109248 667994 109284
rect 668306 173576 668362 173632
rect 668306 168544 668362 168600
rect 668306 165144 668362 165200
rect 668674 158344 668730 158400
rect 668582 153312 668638 153368
rect 668306 148144 668362 148200
rect 668306 144880 668362 144936
rect 668582 132948 668584 132968
rect 668584 132948 668636 132968
rect 668636 132948 668638 132968
rect 668582 132912 668638 132948
rect 668398 116048 668454 116104
rect 668306 110880 668362 110936
rect 668122 107480 668178 107536
rect 668674 104080 668730 104136
rect 672354 669024 672410 669080
rect 672078 474816 672134 474872
rect 669226 114316 669228 114336
rect 669228 114316 669280 114336
rect 669280 114316 669282 114336
rect 669226 114280 669282 114316
rect 668858 112648 668914 112704
rect 669226 105848 669282 105904
rect 668766 102448 668822 102504
rect 668582 100816 668638 100872
rect 576122 47504 576178 47560
rect 605838 44920 605894 44976
rect 607310 45056 607366 45112
rect 608598 44784 608654 44840
rect 607218 43424 607274 43480
rect 518622 42336 518678 42392
rect 514850 42064 514906 42120
rect 520370 42064 520426 42120
rect 521750 42064 521806 42120
rect 529662 42064 529718 42120
rect 525890 41792 525946 41848
rect 478786 41520 478842 41576
rect 611358 46552 611414 46608
rect 625066 89936 625122 89992
rect 626354 92520 626410 92576
rect 628286 95920 628342 95976
rect 641718 95784 641774 95840
rect 642270 96464 642326 96520
rect 627826 94424 627882 94480
rect 626538 93472 626594 93528
rect 626446 91568 626502 91624
rect 625802 89664 625858 89720
rect 626446 88848 626502 88904
rect 626446 87896 626502 87952
rect 643098 87624 643154 87680
rect 626354 86944 626410 87000
rect 626446 85992 626502 86048
rect 626446 85040 626502 85096
rect 625618 84108 625674 84144
rect 625618 84088 625620 84108
rect 625620 84088 625672 84108
rect 625672 84088 625674 84108
rect 626078 83136 626134 83192
rect 644478 89664 644534 89720
rect 644662 94560 644718 94616
rect 644754 92112 644810 92168
rect 644570 84632 644626 84688
rect 626446 82184 626502 82240
rect 643282 82184 643338 82240
rect 629206 80824 629262 80880
rect 633898 77696 633954 77752
rect 631138 75928 631194 75984
rect 633898 75928 633954 75984
rect 639602 77696 639658 77752
rect 639234 75112 639290 75168
rect 646870 74432 646926 74488
rect 647330 71440 647386 71496
rect 646134 70352 646190 70408
rect 648710 72936 648766 72992
rect 655334 93336 655390 93392
rect 654782 92520 654838 92576
rect 654322 91432 654378 91488
rect 654322 90616 654378 90672
rect 655426 89800 655482 89856
rect 657358 94696 657414 94752
rect 663798 92520 663854 92576
rect 663890 90616 663946 90672
rect 665178 91704 665234 91760
rect 665362 93336 665418 93392
rect 665270 89800 665326 89856
rect 664074 88984 664130 89040
rect 648802 68448 648858 68504
rect 647422 66952 647478 67008
rect 646134 66000 646190 66056
rect 646134 64368 646190 64424
rect 612830 47640 612886 47696
rect 661130 47504 661186 47560
rect 675758 961288 675814 961344
rect 675666 959112 675722 959168
rect 675482 957752 675538 957808
rect 675022 957616 675078 957672
rect 675758 953944 675814 954000
rect 677506 950952 677562 951008
rect 677414 950816 677470 950872
rect 676034 939936 676090 939992
rect 676218 939256 676274 939312
rect 676034 939156 676036 939176
rect 676036 939156 676088 939176
rect 676088 939156 676090 939176
rect 676034 939120 676090 939156
rect 676034 938712 676090 938768
rect 676126 938032 676182 938088
rect 676034 937488 676090 937544
rect 676218 937624 676274 937680
rect 676218 937236 676274 937272
rect 676218 937216 676220 937236
rect 676220 937216 676272 937236
rect 676272 937216 676274 937236
rect 676034 936692 676090 936728
rect 676034 936672 676036 936692
rect 676036 936672 676088 936692
rect 676088 936672 676090 936692
rect 676218 935992 676274 936048
rect 676034 935876 676090 935912
rect 676034 935856 676036 935876
rect 676036 935856 676088 935876
rect 676088 935856 676090 935876
rect 677414 934768 677470 934824
rect 681002 949728 681058 949784
rect 679806 949592 679862 949648
rect 679622 949456 679678 949512
rect 678242 933544 678298 933600
rect 677506 933136 677562 933192
rect 676218 931948 676220 931968
rect 676220 931948 676272 931968
rect 676272 931948 676274 931968
rect 676218 931912 676274 931948
rect 681094 948776 681150 948832
rect 681002 934360 681058 934416
rect 682382 947960 682438 948016
rect 682382 935176 682438 935232
rect 681094 933952 681150 934008
rect 679806 931504 679862 931560
rect 679622 931096 679678 931152
rect 676218 930300 676274 930336
rect 676218 930280 676220 930300
rect 676220 930280 676272 930300
rect 676272 930280 676274 930300
rect 674746 930144 674802 930200
rect 683118 929464 683174 929520
rect 683118 928648 683174 928704
rect 675758 876560 675814 876616
rect 675298 876424 675354 876480
rect 675758 874112 675814 874168
rect 675758 872752 675814 872808
rect 675390 872208 675446 872264
rect 675758 864728 675814 864784
rect 675390 788024 675446 788080
rect 675758 786664 675814 786720
rect 675482 784760 675538 784816
rect 675758 784080 675814 784136
rect 675206 773880 675262 773936
rect 675482 773336 675538 773392
rect 675666 773336 675722 773392
rect 677414 773064 677470 773120
rect 675482 766536 675538 766592
rect 675666 766572 675668 766592
rect 675668 766572 675720 766592
rect 675720 766572 675722 766592
rect 675666 766536 675722 766572
rect 675574 765040 675630 765096
rect 676126 761232 676182 761288
rect 676034 760688 676090 760744
rect 676218 760844 676274 760880
rect 676218 760824 676220 760844
rect 676220 760824 676272 760844
rect 676272 760824 676274 760844
rect 676218 760008 676274 760064
rect 674746 759872 674802 759928
rect 674654 759056 674710 759112
rect 676218 759212 676274 759248
rect 676218 759192 676220 759212
rect 676220 759192 676272 759212
rect 676272 759192 676274 759212
rect 676034 759076 676090 759112
rect 676034 759056 676036 759076
rect 676036 759056 676088 759076
rect 676088 759056 676090 759076
rect 676218 758820 676220 758840
rect 676220 758820 676272 758840
rect 676272 758820 676274 758840
rect 676218 758784 676274 758820
rect 676034 758260 676090 758296
rect 676034 758240 676036 758260
rect 676036 758240 676088 758260
rect 676088 758240 676090 758260
rect 677506 772928 677562 772984
rect 676218 757152 676274 757208
rect 677414 757152 677470 757208
rect 676126 755928 676182 755984
rect 676218 755556 676220 755576
rect 676220 755556 676272 755576
rect 676272 755556 676274 755576
rect 676218 755520 676274 755556
rect 676218 755132 676274 755168
rect 676218 755112 676220 755132
rect 676220 755112 676272 755132
rect 676272 755112 676274 755132
rect 681002 772656 681058 772712
rect 681002 755928 681058 755984
rect 677506 754704 677562 754760
rect 676218 753888 676274 753944
rect 676034 753380 676036 753400
rect 676036 753380 676088 753400
rect 676088 753380 676090 753400
rect 676034 753344 676090 753380
rect 676126 752664 676182 752720
rect 676218 752256 676274 752312
rect 676218 751884 676220 751904
rect 676220 751884 676272 751904
rect 676272 751884 676274 751904
rect 676218 751848 676274 751884
rect 683118 751032 683174 751088
rect 683118 750216 683174 750272
rect 675666 741648 675722 741704
rect 674838 736072 674894 736128
rect 675758 734304 675814 734360
rect 675758 732944 675814 733000
rect 675482 728320 675538 728376
rect 675666 728320 675722 728376
rect 678242 727232 678298 727288
rect 675482 721500 675538 721556
rect 675666 721500 675722 721556
rect 676034 716524 676036 716544
rect 676036 716524 676088 716544
rect 676088 716524 676090 716544
rect 676034 716488 676090 716524
rect 676034 716116 676036 716136
rect 676036 716116 676088 716136
rect 676088 716116 676090 716136
rect 676034 716080 676090 716116
rect 676034 715672 676090 715728
rect 674746 715264 674802 715320
rect 674746 714856 674802 714912
rect 676034 714484 676036 714504
rect 676036 714484 676088 714504
rect 676088 714484 676090 714504
rect 676034 714448 676090 714484
rect 676034 714060 676090 714096
rect 676034 714040 676036 714060
rect 676036 714040 676088 714060
rect 676088 714040 676090 714060
rect 676034 713668 676036 713688
rect 676036 713668 676088 713688
rect 676088 713668 676090 713688
rect 676034 713632 676090 713668
rect 676954 713432 677010 713488
rect 676034 713244 676090 713280
rect 676034 713224 676036 713244
rect 676036 713224 676088 713244
rect 676088 713224 676090 713244
rect 676034 712852 676036 712872
rect 676036 712852 676088 712872
rect 676088 712852 676090 712872
rect 676034 712816 676090 712852
rect 676034 712428 676090 712464
rect 676034 712408 676036 712428
rect 676036 712408 676088 712428
rect 676088 712408 676090 712428
rect 676034 711628 676036 711648
rect 676036 711628 676088 711648
rect 676088 711628 676090 711648
rect 676034 711592 676090 711628
rect 676034 710404 676036 710424
rect 676036 710404 676088 710424
rect 676088 710404 676090 710424
rect 676034 710368 676090 710404
rect 676034 709996 676036 710016
rect 676036 709996 676088 710016
rect 676088 709996 676090 710016
rect 676034 709960 676090 709996
rect 676034 709588 676036 709608
rect 676036 709588 676088 709608
rect 676088 709588 676090 709608
rect 676034 709552 676090 709588
rect 676034 709180 676036 709200
rect 676036 709180 676088 709200
rect 676088 709180 676090 709200
rect 676034 709144 676090 709180
rect 681002 726552 681058 726608
rect 679622 724376 679678 724432
rect 678242 712000 678298 712056
rect 679622 711184 679678 711240
rect 681002 710776 681058 710832
rect 676034 708736 676090 708792
rect 676034 708364 676036 708384
rect 676036 708364 676088 708384
rect 676088 708364 676090 708384
rect 676034 708328 676090 708364
rect 676034 707956 676036 707976
rect 676036 707956 676088 707976
rect 676088 707956 676090 707976
rect 676034 707920 676090 707956
rect 676034 707548 676036 707568
rect 676036 707548 676088 707568
rect 676088 707548 676090 707568
rect 676034 707512 676090 707548
rect 676034 707104 676090 707160
rect 675942 706732 675944 706752
rect 675944 706732 675996 706752
rect 675996 706732 675998 706752
rect 675942 706696 675998 706732
rect 676034 706288 676090 706344
rect 676034 705064 676090 705120
rect 675390 696904 675446 696960
rect 675482 694728 675538 694784
rect 675758 694184 675814 694240
rect 675758 687384 675814 687440
rect 675666 686160 675722 686216
rect 675390 683304 675446 683360
rect 675758 683304 675814 683360
rect 675482 683168 675538 683224
rect 675390 676368 675446 676424
rect 674746 670112 674802 670168
rect 674746 668072 674802 668128
rect 674378 547984 674434 548040
rect 676494 683032 676550 683088
rect 679622 681808 679678 681864
rect 675758 676368 675814 676424
rect 676494 676368 676550 676424
rect 676218 671064 676274 671120
rect 676034 670948 676090 670984
rect 676034 670928 676036 670948
rect 676036 670928 676088 670948
rect 676088 670928 676090 670948
rect 676126 670248 676182 670304
rect 676218 669432 676274 669488
rect 676034 669296 676090 669352
rect 676218 668616 676274 668672
rect 676034 668516 676036 668536
rect 676036 668516 676088 668536
rect 676088 668516 676090 668536
rect 676034 668480 676090 668516
rect 676218 667392 676274 667448
rect 676034 667276 676090 667312
rect 676034 667256 676036 667276
rect 676036 667256 676088 667276
rect 676088 667256 676090 667276
rect 679714 678272 679770 678328
rect 679622 666984 679678 667040
rect 676126 666168 676182 666224
rect 676218 665760 676274 665816
rect 679714 665760 679770 665816
rect 676034 665252 676036 665272
rect 676036 665252 676088 665272
rect 676088 665252 676090 665272
rect 676034 665216 676090 665252
rect 676218 664980 676220 665000
rect 676220 664980 676272 665000
rect 676272 664980 676274 665000
rect 676218 664944 676274 664980
rect 676218 664128 676274 664184
rect 676218 663756 676220 663776
rect 676220 663756 676272 663776
rect 676272 663756 676274 663776
rect 676218 663720 676274 663756
rect 676218 663312 676274 663368
rect 676034 662380 676090 662416
rect 676034 662360 676036 662380
rect 676036 662360 676088 662380
rect 676088 662360 676090 662380
rect 676218 661680 676274 661736
rect 676126 661272 676182 661328
rect 683118 660864 683174 660920
rect 683118 660048 683174 660104
rect 675390 649848 675446 649904
rect 675758 648624 675814 648680
rect 675206 645904 675262 645960
rect 675758 644680 675814 644736
rect 675666 643048 675722 643104
rect 675206 638696 675262 638752
rect 675482 638152 675538 638208
rect 676862 637880 676918 637936
rect 677506 637880 677562 637936
rect 675206 631352 675262 631408
rect 676862 631352 676918 631408
rect 676126 626048 676182 626104
rect 676218 625640 676274 625696
rect 676218 625232 676274 625288
rect 676218 624824 676274 624880
rect 676126 624416 676182 624472
rect 676034 623872 676090 623928
rect 676218 624008 676274 624064
rect 676218 623636 676220 623656
rect 676220 623636 676272 623656
rect 676272 623636 676274 623656
rect 676218 623600 676274 623636
rect 676034 623076 676090 623112
rect 676034 623056 676036 623076
rect 676036 623056 676088 623076
rect 676088 623056 676090 623076
rect 676218 622820 676220 622840
rect 676220 622820 676272 622840
rect 676272 622820 676274 622840
rect 676218 622784 676274 622820
rect 676034 622260 676090 622296
rect 676034 622240 676036 622260
rect 676036 622240 676088 622260
rect 676088 622240 676090 622260
rect 676218 621172 676274 621208
rect 676218 621152 676220 621172
rect 676220 621152 676272 621172
rect 676272 621152 676274 621172
rect 676218 619928 676274 619984
rect 676034 619828 676036 619848
rect 676036 619828 676088 619848
rect 676088 619828 676090 619848
rect 676034 619792 676090 619828
rect 676218 619112 676274 619168
rect 676034 619012 676036 619032
rect 676036 619012 676088 619032
rect 676088 619012 676090 619032
rect 676034 618976 676090 619012
rect 681002 637472 681058 637528
rect 679622 637336 679678 637392
rect 679622 621968 679678 622024
rect 681094 621560 681150 621616
rect 681002 620744 681058 620800
rect 677506 618704 677562 618760
rect 676218 617480 676274 617536
rect 676034 617380 676036 617400
rect 676036 617380 676088 617400
rect 676088 617380 676090 617400
rect 676034 617344 676090 617380
rect 676034 616972 676036 616992
rect 676036 616972 676088 616992
rect 676088 616972 676090 616992
rect 676034 616936 676090 616972
rect 676218 616700 676220 616720
rect 676220 616700 676272 616720
rect 676272 616700 676274 616720
rect 676218 616664 676274 616700
rect 683118 615848 683174 615904
rect 683118 615032 683174 615088
rect 675390 606464 675446 606520
rect 675206 600888 675262 600944
rect 675758 598984 675814 599040
rect 675574 595312 675630 595368
rect 675758 593136 675814 593192
rect 675574 593000 675630 593056
rect 675482 592048 675538 592104
rect 677506 592048 677562 592104
rect 675574 586200 675630 586256
rect 675850 586200 675906 586256
rect 675482 584568 675538 584624
rect 676034 581052 676090 581088
rect 676034 581032 676036 581052
rect 676036 581032 676088 581052
rect 676088 581032 676090 581052
rect 676126 580488 676182 580544
rect 676034 580216 676090 580272
rect 676218 580100 676274 580136
rect 676218 580080 676220 580100
rect 676220 580080 676272 580100
rect 676272 580080 676274 580100
rect 676310 579264 676366 579320
rect 676218 578856 676274 578912
rect 676126 578448 676182 578504
rect 676034 578196 676090 578232
rect 676034 578176 676036 578196
rect 676036 578176 676088 578196
rect 676088 578176 676090 578196
rect 676218 577652 676274 577688
rect 676218 577632 676220 577652
rect 676220 577632 676272 577652
rect 676272 577632 676274 577652
rect 676034 577396 676036 577416
rect 676036 577396 676088 577416
rect 676088 577396 676090 577416
rect 676034 577360 676090 577396
rect 676034 576972 676090 577008
rect 676034 576952 676036 576972
rect 676036 576952 676088 576972
rect 676088 576952 676090 576972
rect 676126 576408 676182 576464
rect 676034 575728 676090 575784
rect 676218 576000 676274 576056
rect 676034 574948 676036 574968
rect 676036 574948 676088 574968
rect 676088 574948 676090 574968
rect 676034 574912 676090 574948
rect 676218 574368 676274 574424
rect 676034 574132 676036 574152
rect 676036 574132 676088 574152
rect 676088 574132 676090 574152
rect 676034 574096 676090 574132
rect 676034 573724 676036 573744
rect 676036 573724 676088 573744
rect 676088 573724 676090 573744
rect 676034 573688 676090 573724
rect 682382 591368 682438 591424
rect 682382 575592 682438 575648
rect 677506 573552 677562 573608
rect 676218 571920 676274 571976
rect 676218 571532 676274 571568
rect 676218 571512 676220 571532
rect 676220 571512 676272 571532
rect 676272 571512 676274 571532
rect 676218 571104 676274 571160
rect 683118 570696 683174 570752
rect 683118 569880 683174 569936
rect 675758 562672 675814 562728
rect 675482 561176 675538 561232
rect 675574 559544 675630 559600
rect 675758 558864 675814 558920
rect 674930 554784 674986 554840
rect 675758 553968 675814 554024
rect 675758 551928 675814 551984
rect 675022 550296 675078 550352
rect 674654 547848 674710 547904
rect 678242 546760 678298 546816
rect 677506 546488 677562 546544
rect 676218 535880 676274 535936
rect 676034 535676 676090 535732
rect 676126 535064 676182 535120
rect 675942 534452 675998 534508
rect 675850 528368 675852 528388
rect 675852 528368 675904 528388
rect 675904 528368 675906 528388
rect 675850 528332 675906 528368
rect 675850 527128 675906 527164
rect 675850 527108 675852 527128
rect 675852 527108 675904 527128
rect 675904 527108 675906 527128
rect 676218 534656 676274 534712
rect 676218 534248 676274 534304
rect 676034 533264 676036 533284
rect 676036 533264 676088 533284
rect 676088 533264 676090 533284
rect 676034 533228 676090 533264
rect 676034 532820 676090 532876
rect 675850 492088 675906 492144
rect 675942 491680 675998 491736
rect 675942 491272 675998 491328
rect 675758 490864 675814 490920
rect 675942 490456 675998 490512
rect 675850 489640 675906 489696
rect 676218 532652 676220 532672
rect 676220 532652 676272 532672
rect 676272 532652 676274 532672
rect 676218 532616 676274 532652
rect 677230 531800 677286 531856
rect 676126 530576 676182 530632
rect 676218 530188 676274 530224
rect 676218 530168 676220 530188
rect 676220 530168 676272 530188
rect 676272 530168 676274 530188
rect 676126 529352 676182 529408
rect 676218 528944 676274 529000
rect 676402 528980 676404 529000
rect 676404 528980 676456 529000
rect 676456 528980 676458 529000
rect 676402 528944 676458 528980
rect 676218 527720 676274 527776
rect 676218 526940 676220 526960
rect 676220 526940 676272 526960
rect 676272 526940 676274 526960
rect 676218 526904 676274 526940
rect 676218 526532 676220 526552
rect 676220 526532 676272 526552
rect 676272 526532 676274 526552
rect 676218 526496 676274 526532
rect 676034 489232 676090 489288
rect 676034 488844 676090 488880
rect 676034 488824 676036 488844
rect 676036 488824 676088 488844
rect 676088 488824 676090 488844
rect 676034 488452 676036 488472
rect 676036 488452 676088 488472
rect 676088 488452 676090 488472
rect 676034 488416 676090 488452
rect 676034 488028 676090 488064
rect 676034 488008 676036 488028
rect 676036 488008 676088 488028
rect 676088 488008 676090 488028
rect 676034 486820 676036 486840
rect 676036 486820 676088 486840
rect 676088 486820 676090 486840
rect 676034 486784 676090 486820
rect 676034 486004 676036 486024
rect 676036 486004 676088 486024
rect 676088 486004 676090 486024
rect 676034 485968 676090 486004
rect 674746 485560 674802 485616
rect 675942 485188 675944 485208
rect 675944 485188 675996 485208
rect 675996 485188 675998 485208
rect 675942 485152 675998 485188
rect 675942 484780 675944 484800
rect 675944 484780 675996 484800
rect 675996 484780 675998 484800
rect 675942 484744 675998 484780
rect 675942 483148 675944 483168
rect 675944 483148 675996 483168
rect 675996 483148 675998 483168
rect 675942 483112 675998 483148
rect 675942 482740 675944 482760
rect 675944 482740 675996 482760
rect 675996 482740 675998 482760
rect 675942 482704 675998 482740
rect 674654 482296 674710 482352
rect 679622 546624 679678 546680
rect 678334 542952 678390 543008
rect 678242 531392 678298 531448
rect 683302 543632 683358 543688
rect 679622 531800 679678 531856
rect 678334 530576 678390 530632
rect 683854 533432 683910 533488
rect 683302 527720 683358 527776
rect 683118 525680 683174 525736
rect 683118 524864 683174 524920
rect 677414 492360 677470 492416
rect 677322 489872 677378 489928
rect 676310 403688 676366 403744
rect 676218 403300 676274 403336
rect 676218 403280 676220 403300
rect 676220 403280 676272 403300
rect 676272 403280 676274 403300
rect 676402 403280 676458 403336
rect 676126 402872 676182 402928
rect 676218 402056 676274 402112
rect 676034 401784 676090 401840
rect 676218 401240 676274 401296
rect 674746 400560 674802 400616
rect 681002 487600 681058 487656
rect 679714 487192 679770 487248
rect 679622 486376 679678 486432
rect 677414 484336 677470 484392
rect 678978 480664 679034 480720
rect 677322 401240 677378 401296
rect 677230 400424 677286 400480
rect 676218 399628 676274 399664
rect 676218 399608 676220 399628
rect 676220 399608 676272 399628
rect 676272 399608 676274 399628
rect 676034 398520 676090 398576
rect 676034 398112 676090 398168
rect 676862 397568 676918 397624
rect 676402 395528 676458 395584
rect 676218 394324 676274 394360
rect 676218 394304 676220 394324
rect 676220 394304 676272 394324
rect 676272 394304 676274 394324
rect 676218 393896 676274 393952
rect 676494 394712 676550 394768
rect 676402 387640 676458 387696
rect 676954 396752 677010 396808
rect 678334 396344 678390 396400
rect 678242 395936 678298 395992
rect 676862 388456 676918 388512
rect 683118 393488 683174 393544
rect 683118 392264 683174 392320
rect 678334 387504 678390 387560
rect 675758 384920 675814 384976
rect 675390 382200 675446 382256
rect 675482 378664 675538 378720
rect 675758 377576 675814 377632
rect 675758 375400 675814 375456
rect 675758 373632 675814 373688
rect 675758 372000 675814 372056
rect 675850 358672 675906 358728
rect 675942 358264 675998 358320
rect 676034 357856 676090 357912
rect 676034 357484 676036 357504
rect 676036 357484 676088 357504
rect 676088 357484 676090 357504
rect 676034 357448 676090 357484
rect 676034 357060 676090 357096
rect 676034 357040 676036 357060
rect 676036 357040 676088 357060
rect 676088 357040 676090 357060
rect 676034 356668 676036 356688
rect 676036 356668 676088 356688
rect 676088 356668 676090 356688
rect 676034 356632 676090 356668
rect 676034 356244 676090 356280
rect 676034 356224 676036 356244
rect 676036 356224 676088 356244
rect 676088 356224 676090 356244
rect 674746 355816 674802 355872
rect 674746 355408 674802 355464
rect 676034 355036 676036 355056
rect 676036 355036 676088 355056
rect 676088 355036 676090 355056
rect 676034 355000 676090 355036
rect 676034 354612 676090 354648
rect 676034 354592 676036 354612
rect 676036 354592 676088 354612
rect 676088 354592 676090 354612
rect 678242 352552 678298 352608
rect 676034 351736 676090 351792
rect 676034 350940 676090 350976
rect 676034 350920 676036 350940
rect 676036 350920 676088 350940
rect 676088 350920 676090 350940
rect 676034 350548 676036 350568
rect 676036 350548 676088 350568
rect 676088 350548 676090 350568
rect 676034 350512 676090 350548
rect 675942 350104 675998 350160
rect 676034 349696 676090 349752
rect 676034 349308 676090 349344
rect 676034 349288 676036 349308
rect 676036 349288 676088 349308
rect 676088 349288 676090 349308
rect 676034 348900 676090 348936
rect 676034 348880 676036 348900
rect 676036 348880 676088 348900
rect 676088 348880 676090 348900
rect 676034 348472 676090 348528
rect 676034 347248 676090 347304
rect 675942 346568 675998 346624
rect 676126 346432 676182 346488
rect 678242 343576 678298 343632
rect 675298 342216 675354 342272
rect 676862 342216 676918 342272
rect 675666 340720 675722 340776
rect 675758 339360 675814 339416
rect 675758 337864 675814 337920
rect 675758 335824 675814 335880
rect 674838 335280 674894 335336
rect 675482 333512 675538 333568
rect 675758 332152 675814 332208
rect 675114 325624 675170 325680
rect 675758 325488 675814 325544
rect 676034 313656 676090 313712
rect 676218 313540 676274 313576
rect 676218 313520 676220 313540
rect 676220 313520 676272 313540
rect 676272 313520 676274 313540
rect 676126 312704 676182 312760
rect 676218 312296 676274 312352
rect 676218 311908 676274 311944
rect 676218 311888 676220 311908
rect 676220 311888 676272 311908
rect 676272 311888 676274 311908
rect 676218 311480 676274 311536
rect 676126 311072 676182 311128
rect 674746 310800 674802 310856
rect 676218 310276 676274 310312
rect 676218 310256 676220 310276
rect 676220 310256 676272 310276
rect 676272 310256 676274 310276
rect 676034 310020 676036 310040
rect 676036 310020 676088 310040
rect 676088 310020 676090 310040
rect 676034 309984 676090 310020
rect 676218 309460 676274 309496
rect 676218 309440 676220 309460
rect 676220 309440 676272 309460
rect 676272 309440 676274 309460
rect 679622 309032 679678 309088
rect 678242 308216 678298 308272
rect 676862 306584 676918 306640
rect 676402 306176 676458 306232
rect 676310 304544 676366 304600
rect 676126 304136 676182 304192
rect 676218 303764 676220 303784
rect 676220 303764 676272 303784
rect 676272 303764 676274 303784
rect 676218 303728 676274 303764
rect 676494 305768 676550 305824
rect 679714 307400 679770 307456
rect 679622 299376 679678 299432
rect 683118 303320 683174 303376
rect 683118 302504 683174 302560
rect 679714 297880 679770 297936
rect 676402 297336 676458 297392
rect 675758 294752 675814 294808
rect 675482 292576 675538 292632
rect 675390 292032 675446 292088
rect 675666 288360 675722 288416
rect 675758 287272 675814 287328
rect 675758 285504 675814 285560
rect 675758 283600 675814 283656
rect 675758 281424 675814 281480
rect 676218 268504 676274 268560
rect 676126 268096 676182 268152
rect 676218 267688 676274 267744
rect 676218 267280 676274 267336
rect 676034 267028 676090 267064
rect 676034 267008 676036 267028
rect 676036 267008 676088 267028
rect 676088 267008 676090 267028
rect 676218 266484 676274 266520
rect 676218 266464 676220 266484
rect 676220 266464 676272 266484
rect 676272 266464 676274 266484
rect 676218 266076 676274 266112
rect 676218 266056 676220 266076
rect 676220 266056 676272 266076
rect 676272 266056 676274 266076
rect 676034 265820 676036 265840
rect 676036 265820 676088 265840
rect 676088 265820 676090 265840
rect 676034 265784 676090 265820
rect 676218 265240 676274 265296
rect 674746 264968 674802 265024
rect 676218 264424 676274 264480
rect 676310 264016 676366 264072
rect 675390 263336 675446 263392
rect 674470 245656 674526 245712
rect 676034 262928 676090 262984
rect 676034 262520 676090 262576
rect 676218 261996 676274 262032
rect 676218 261976 676220 261996
rect 676220 261976 676272 261996
rect 676272 261976 676274 261996
rect 676218 261588 676274 261624
rect 676218 261568 676220 261588
rect 676220 261568 676272 261588
rect 676272 261568 676274 261588
rect 676218 261160 676274 261216
rect 676218 259956 676274 259992
rect 676218 259936 676220 259956
rect 676220 259936 676272 259956
rect 676272 259936 676274 259956
rect 676862 263608 676918 263664
rect 676126 259120 676182 259176
rect 676218 258712 676274 258768
rect 683118 258304 683174 258360
rect 683118 257488 683174 257544
rect 676862 251504 676918 251560
rect 675114 248240 675170 248296
rect 675758 246608 675814 246664
rect 675758 245384 675814 245440
rect 675298 238584 675354 238640
rect 675758 236816 675814 236872
rect 675942 223488 675998 223544
rect 675850 222672 675906 222728
rect 676034 223080 676090 223136
rect 676034 222284 676090 222320
rect 676034 222264 676036 222284
rect 676036 222264 676088 222284
rect 676088 222264 676090 222284
rect 676034 221876 676090 221912
rect 676034 221856 676036 221876
rect 676036 221856 676088 221876
rect 676088 221856 676090 221876
rect 676034 221484 676036 221504
rect 676036 221484 676088 221504
rect 676088 221484 676090 221504
rect 676034 221448 676090 221484
rect 674746 221040 674802 221096
rect 676034 220668 676036 220688
rect 676036 220668 676088 220688
rect 676088 220668 676090 220688
rect 676034 220632 676090 220668
rect 676034 220244 676090 220280
rect 676034 220224 676036 220244
rect 676036 220224 676088 220244
rect 676088 220224 676090 220244
rect 676034 219852 676036 219872
rect 676036 219852 676088 219872
rect 676088 219852 676090 219872
rect 676034 219816 676090 219852
rect 676034 219444 676036 219464
rect 676036 219444 676088 219464
rect 676088 219444 676090 219464
rect 676034 219408 676090 219444
rect 676034 219000 676090 219056
rect 675850 216960 675906 217016
rect 676034 216552 676090 216608
rect 676034 216164 676090 216200
rect 676034 216144 676036 216164
rect 676036 216144 676088 216164
rect 676088 216144 676090 216164
rect 676034 215756 676090 215792
rect 676034 215736 676036 215756
rect 676036 215736 676088 215756
rect 676088 215736 676090 215756
rect 675942 214920 675998 214976
rect 676034 214124 676090 214160
rect 676034 214104 676036 214124
rect 676036 214104 676088 214124
rect 676088 214104 676090 214124
rect 676034 213968 676090 214024
rect 679622 217368 679678 217424
rect 676034 213716 676090 213752
rect 676034 213696 676036 213716
rect 676036 213696 676088 213716
rect 676088 213696 676090 213716
rect 676034 213288 676090 213344
rect 676034 212064 676090 212120
rect 675942 211384 675998 211440
rect 675850 211248 675906 211304
rect 676862 208256 676918 208312
rect 679622 207168 679678 207224
rect 675758 205536 675814 205592
rect 675758 204992 675814 205048
rect 675758 204176 675814 204232
rect 675114 202816 675170 202872
rect 674838 201320 674894 201376
rect 675482 202680 675538 202736
rect 675758 198328 675814 198384
rect 675758 195336 675814 195392
rect 675758 190340 675760 190360
rect 675760 190340 675812 190360
rect 675812 190340 675814 190360
rect 675758 190304 675814 190340
rect 674838 190168 674894 190224
rect 675942 178472 675998 178528
rect 676034 178064 676090 178120
rect 675942 177656 675998 177712
rect 676034 177284 676036 177304
rect 676036 177284 676088 177304
rect 676088 177284 676090 177304
rect 676034 177248 676090 177284
rect 676034 176840 676090 176896
rect 674746 176432 674802 176488
rect 676034 176044 676090 176080
rect 676034 176024 676036 176044
rect 676036 176024 676088 176044
rect 676088 176024 676090 176044
rect 676034 175652 676036 175672
rect 676036 175652 676088 175672
rect 676088 175652 676090 175672
rect 676034 175616 676090 175652
rect 676034 175228 676090 175264
rect 676034 175208 676036 175228
rect 676036 175208 676088 175228
rect 676088 175208 676090 175228
rect 676034 174836 676036 174856
rect 676036 174836 676088 174856
rect 676088 174836 676090 174856
rect 676034 174800 676090 174836
rect 674746 174392 674802 174448
rect 678242 173168 678298 173224
rect 676034 172760 676090 172816
rect 676034 172352 676090 172408
rect 676034 171128 676090 171184
rect 676034 170332 676090 170368
rect 676034 170312 676036 170332
rect 676036 170312 676088 170332
rect 676088 170312 676090 170332
rect 676034 169632 676090 169688
rect 676770 171536 676826 171592
rect 676586 169904 676642 169960
rect 676034 169516 676090 169552
rect 676034 169496 676036 169516
rect 676036 169496 676088 169516
rect 676088 169496 676090 169516
rect 676034 169108 676090 169144
rect 676034 169088 676036 169108
rect 676036 169088 676088 169108
rect 676088 169088 676090 169108
rect 676034 168680 676090 168736
rect 676034 168292 676090 168328
rect 676034 168272 676036 168292
rect 676036 168272 676088 168292
rect 676088 168272 676090 168292
rect 676034 167884 676090 167920
rect 676034 167864 676036 167884
rect 676036 167864 676088 167884
rect 676088 167864 676090 167884
rect 676034 167068 676090 167104
rect 676034 167048 676036 167068
rect 676036 167048 676088 167068
rect 676088 167048 676090 167068
rect 676586 166368 676642 166424
rect 676770 166368 676826 166424
rect 677046 162696 677102 162752
rect 676862 162560 676918 162616
rect 675758 159976 675814 160032
rect 675482 159432 675538 159488
rect 675666 157392 675722 157448
rect 675482 156984 675538 157040
rect 675758 156304 675814 156360
rect 675758 153040 675814 153096
rect 675758 151544 675814 151600
rect 675758 148416 675814 148472
rect 675758 146240 675814 146296
rect 676126 133048 676182 133104
rect 676034 132912 676090 132968
rect 676218 132640 676274 132696
rect 676218 131824 676274 131880
rect 676126 131416 676182 131472
rect 676034 131300 676090 131336
rect 676034 131280 676036 131300
rect 676036 131280 676088 131300
rect 676088 131280 676090 131300
rect 676126 130600 676182 130656
rect 676218 130192 676274 130248
rect 676218 129804 676274 129840
rect 676218 129784 676220 129804
rect 676220 129784 676272 129804
rect 676272 129784 676274 129804
rect 674746 129648 674802 129704
rect 676218 128968 676274 129024
rect 683670 128152 683726 128208
rect 676034 128016 676090 128072
rect 683118 127336 683174 127392
rect 674746 123528 674802 123584
rect 676862 126928 676918 126984
rect 676402 125296 676458 125352
rect 676034 123956 676090 123992
rect 676034 123936 676036 123956
rect 676036 123936 676088 123956
rect 676088 123936 676090 123956
rect 676218 122868 676274 122904
rect 676218 122848 676220 122868
rect 676220 122848 676272 122868
rect 676272 122848 676274 122868
rect 676126 122440 676182 122496
rect 676218 121624 676274 121680
rect 679622 125704 679678 125760
rect 678242 125296 678298 125352
rect 677598 124072 677654 124128
rect 676862 117952 676918 118008
rect 676402 117272 676458 117328
rect 683302 126112 683358 126168
rect 683118 124888 683174 124944
rect 679622 117136 679678 117192
rect 683670 121624 683726 121680
rect 675390 114144 675446 114200
rect 675666 112512 675722 112568
rect 675482 111696 675538 111752
rect 675114 108976 675170 109032
rect 675758 108160 675814 108216
rect 675758 104760 675814 104816
rect 675758 103128 675814 103184
rect 675758 101360 675814 101416
rect 664258 48456 664314 48512
rect 662418 47368 662474 47424
rect 612738 46416 612794 46472
rect 611450 46280 611506 46336
rect 610162 46144 610218 46200
rect 610070 45192 610126 45248
rect 609978 41384 610034 41440
rect 141698 40296 141754 40352
<< metal3 >>
rect 203885 1007178 203951 1007181
rect 203885 1007176 204148 1007178
rect 203885 1007120 203890 1007176
rect 203946 1007120 204148 1007176
rect 203885 1007118 204148 1007120
rect 203885 1007115 203951 1007118
rect 99925 1006634 99991 1006637
rect 99925 1006632 100096 1006634
rect 99925 1006576 99930 1006632
rect 99986 1006576 100096 1006632
rect 99925 1006574 100096 1006576
rect 99925 1006571 99991 1006574
rect 104341 1006498 104407 1006501
rect 104801 1006498 104867 1006501
rect 258165 1006498 258231 1006501
rect 307293 1006498 307359 1006501
rect 308121 1006498 308187 1006501
rect 358169 1006498 358235 1006501
rect 427537 1006498 427603 1006501
rect 428365 1006498 428431 1006501
rect 104341 1006496 104604 1006498
rect 104341 1006440 104346 1006496
rect 104402 1006440 104604 1006496
rect 104341 1006438 104604 1006440
rect 104801 1006496 104972 1006498
rect 104801 1006440 104806 1006496
rect 104862 1006440 104972 1006496
rect 104801 1006438 104972 1006440
rect 258165 1006496 258428 1006498
rect 258165 1006440 258170 1006496
rect 258226 1006440 258428 1006496
rect 258165 1006438 258428 1006440
rect 307293 1006496 307556 1006498
rect 307293 1006440 307298 1006496
rect 307354 1006440 307556 1006496
rect 307293 1006438 307556 1006440
rect 308121 1006496 308384 1006498
rect 308121 1006440 308126 1006496
rect 308182 1006440 308384 1006496
rect 308121 1006438 308384 1006440
rect 357972 1006496 358235 1006498
rect 357972 1006440 358174 1006496
rect 358230 1006440 358235 1006496
rect 357972 1006438 358235 1006440
rect 427340 1006496 427603 1006498
rect 427340 1006440 427542 1006496
rect 427598 1006440 427603 1006496
rect 427340 1006438 427603 1006440
rect 428260 1006496 428431 1006498
rect 428260 1006440 428370 1006496
rect 428426 1006440 428431 1006496
rect 428260 1006438 428431 1006440
rect 104341 1006435 104407 1006438
rect 104801 1006435 104867 1006438
rect 258165 1006435 258231 1006438
rect 307293 1006435 307359 1006438
rect 308121 1006435 308187 1006438
rect 358169 1006435 358235 1006438
rect 427537 1006435 427603 1006438
rect 428365 1006435 428431 1006438
rect 100661 1006362 100727 1006365
rect 149697 1006362 149763 1006365
rect 150893 1006362 150959 1006365
rect 100661 1006360 100924 1006362
rect 100661 1006304 100666 1006360
rect 100722 1006304 100924 1006360
rect 100661 1006302 100924 1006304
rect 149500 1006360 149763 1006362
rect 149500 1006304 149702 1006360
rect 149758 1006304 149763 1006360
rect 149500 1006302 149763 1006304
rect 150696 1006360 150959 1006362
rect 150696 1006304 150898 1006360
rect 150954 1006304 150959 1006360
rect 150696 1006302 150959 1006304
rect 100661 1006299 100727 1006302
rect 149697 1006299 149763 1006302
rect 150893 1006299 150959 1006302
rect 154113 1006362 154179 1006365
rect 202689 1006362 202755 1006365
rect 210049 1006362 210115 1006365
rect 154113 1006360 154376 1006362
rect 154113 1006304 154118 1006360
rect 154174 1006304 154376 1006360
rect 154113 1006302 154376 1006304
rect 202689 1006360 202952 1006362
rect 202689 1006304 202694 1006360
rect 202750 1006304 202952 1006360
rect 202689 1006302 202952 1006304
rect 209852 1006360 210115 1006362
rect 209852 1006304 210054 1006360
rect 210110 1006304 210115 1006360
rect 209852 1006302 210115 1006304
rect 154113 1006299 154179 1006302
rect 202689 1006299 202755 1006302
rect 210049 1006299 210115 1006302
rect 254853 1006362 254919 1006365
rect 310605 1006362 310671 1006365
rect 356053 1006362 356119 1006365
rect 357709 1006362 357775 1006365
rect 504541 1006362 504607 1006365
rect 555969 1006362 556035 1006365
rect 254853 1006360 255116 1006362
rect 254853 1006304 254858 1006360
rect 254914 1006304 255116 1006360
rect 254853 1006302 255116 1006304
rect 310605 1006360 310868 1006362
rect 310605 1006304 310610 1006360
rect 310666 1006304 310868 1006360
rect 310605 1006302 310868 1006304
rect 355948 1006360 356119 1006362
rect 355948 1006304 356058 1006360
rect 356114 1006304 356119 1006360
rect 355948 1006302 356119 1006304
rect 357604 1006360 357775 1006362
rect 357604 1006304 357714 1006360
rect 357770 1006304 357775 1006360
rect 357604 1006302 357775 1006304
rect 504436 1006360 504607 1006362
rect 504436 1006304 504546 1006360
rect 504602 1006304 504607 1006360
rect 504436 1006302 504607 1006304
rect 555772 1006360 556035 1006362
rect 555772 1006304 555974 1006360
rect 556030 1006304 556035 1006360
rect 555772 1006302 556035 1006304
rect 254853 1006299 254919 1006302
rect 310605 1006299 310671 1006302
rect 356053 1006299 356119 1006302
rect 357709 1006299 357775 1006302
rect 504541 1006299 504607 1006302
rect 555969 1006299 556035 1006302
rect 103605 1006226 103671 1006229
rect 151721 1006226 151787 1006229
rect 152089 1006226 152155 1006229
rect 204345 1006226 204411 1006229
rect 210417 1006226 210483 1006229
rect 255313 1006226 255379 1006229
rect 257337 1006226 257403 1006229
rect 306465 1006226 306531 1006229
rect 358905 1006226 358971 1006229
rect 425145 1006226 425211 1006229
rect 505001 1006226 505067 1006229
rect 505369 1006226 505435 1006229
rect 557165 1006226 557231 1006229
rect 103605 1006224 103776 1006226
rect 103605 1006168 103610 1006224
rect 103666 1006168 103776 1006224
rect 103605 1006166 103776 1006168
rect 151721 1006224 151892 1006226
rect 151721 1006168 151726 1006224
rect 151782 1006168 151892 1006224
rect 151721 1006166 151892 1006168
rect 152089 1006224 152352 1006226
rect 152089 1006168 152094 1006224
rect 152150 1006168 152352 1006224
rect 152089 1006166 152352 1006168
rect 204345 1006224 204516 1006226
rect 204345 1006168 204350 1006224
rect 204406 1006168 204516 1006224
rect 204345 1006166 204516 1006168
rect 210417 1006224 210680 1006226
rect 210417 1006168 210422 1006224
rect 210478 1006168 210680 1006224
rect 210417 1006166 210680 1006168
rect 255313 1006224 255576 1006226
rect 255313 1006168 255318 1006224
rect 255374 1006168 255576 1006224
rect 255313 1006166 255576 1006168
rect 257337 1006224 257600 1006226
rect 257337 1006168 257342 1006224
rect 257398 1006168 257600 1006224
rect 257337 1006166 257600 1006168
rect 306465 1006224 306728 1006226
rect 306465 1006168 306470 1006224
rect 306526 1006168 306728 1006224
rect 306465 1006166 306728 1006168
rect 358800 1006224 358971 1006226
rect 358800 1006168 358910 1006224
rect 358966 1006168 358971 1006224
rect 358800 1006166 358971 1006168
rect 424948 1006224 425211 1006226
rect 424948 1006168 425150 1006224
rect 425206 1006168 425211 1006224
rect 424948 1006166 425211 1006168
rect 504804 1006224 505067 1006226
rect 504804 1006168 505006 1006224
rect 505062 1006168 505067 1006224
rect 504804 1006166 505067 1006168
rect 505172 1006224 505435 1006226
rect 505172 1006168 505374 1006224
rect 505430 1006168 505435 1006224
rect 505172 1006166 505435 1006168
rect 557060 1006224 557231 1006226
rect 557060 1006168 557170 1006224
rect 557226 1006168 557231 1006224
rect 557060 1006166 557231 1006168
rect 103605 1006163 103671 1006166
rect 151721 1006163 151787 1006166
rect 152089 1006163 152155 1006166
rect 204345 1006163 204411 1006166
rect 210417 1006163 210483 1006166
rect 255313 1006163 255379 1006166
rect 257337 1006163 257403 1006166
rect 306465 1006163 306531 1006166
rect 358905 1006163 358971 1006166
rect 425145 1006163 425211 1006166
rect 505001 1006163 505067 1006166
rect 505369 1006163 505435 1006166
rect 557165 1006163 557231 1006166
rect 98269 1006090 98335 1006093
rect 99097 1006090 99163 1006093
rect 103145 1006090 103211 1006093
rect 108849 1006090 108915 1006093
rect 150893 1006090 150959 1006093
rect 159081 1006090 159147 1006093
rect 98072 1006088 98335 1006090
rect 98072 1006032 98274 1006088
rect 98330 1006032 98335 1006088
rect 98072 1006030 98335 1006032
rect 98532 1006030 98900 1006090
rect 99097 1006088 99268 1006090
rect 99097 1006032 99102 1006088
rect 99158 1006032 99268 1006088
rect 99097 1006030 99268 1006032
rect 103145 1006088 103408 1006090
rect 103145 1006032 103150 1006088
rect 103206 1006032 103408 1006088
rect 103145 1006030 103408 1006032
rect 108849 1006088 109112 1006090
rect 108849 1006032 108854 1006088
rect 108910 1006032 109112 1006088
rect 108849 1006030 109112 1006032
rect 149868 1006030 150328 1006090
rect 150893 1006088 151156 1006090
rect 150893 1006032 150898 1006088
rect 150954 1006032 151156 1006088
rect 150893 1006030 151156 1006032
rect 158884 1006088 159147 1006090
rect 158884 1006032 159086 1006088
rect 159142 1006032 159147 1006088
rect 158884 1006030 159147 1006032
rect 98269 1006027 98335 1006030
rect 99097 1006027 99163 1006030
rect 103145 1006027 103211 1006030
rect 108849 1006027 108915 1006030
rect 150893 1006027 150959 1006030
rect 159081 1006027 159147 1006030
rect 160645 1006090 160711 1006093
rect 201033 1006090 201099 1006093
rect 201861 1006090 201927 1006093
rect 207197 1006090 207263 1006093
rect 207565 1006090 207631 1006093
rect 209589 1006090 209655 1006093
rect 252461 1006090 252527 1006093
rect 253289 1006090 253355 1006093
rect 256969 1006090 257035 1006093
rect 258533 1006090 258599 1006093
rect 258993 1006090 259059 1006093
rect 261017 1006090 261083 1006093
rect 304073 1006090 304139 1006093
rect 304901 1006090 304967 1006093
rect 305269 1006090 305335 1006093
rect 315113 1006090 315179 1006093
rect 354489 1006090 354555 1006093
rect 355225 1006090 355291 1006093
rect 356881 1006090 356947 1006093
rect 358537 1006090 358603 1006093
rect 361389 1006090 361455 1006093
rect 422661 1006090 422727 1006093
rect 423489 1006090 423555 1006093
rect 427997 1006090 428063 1006093
rect 430021 1006090 430087 1006093
rect 499665 1006090 499731 1006093
rect 500493 1006090 500559 1006093
rect 502517 1006090 502583 1006093
rect 550265 1006090 550331 1006093
rect 551093 1006090 551159 1006093
rect 552289 1006090 552355 1006093
rect 556797 1006090 556863 1006093
rect 160645 1006088 160908 1006090
rect 160645 1006032 160650 1006088
rect 160706 1006032 160908 1006088
rect 160645 1006030 160908 1006032
rect 200836 1006088 201099 1006090
rect 200836 1006032 201038 1006088
rect 201094 1006032 201099 1006088
rect 200836 1006030 201099 1006032
rect 201296 1006030 201756 1006090
rect 201861 1006088 202124 1006090
rect 201861 1006032 201866 1006088
rect 201922 1006032 202124 1006088
rect 201861 1006030 202124 1006032
rect 207197 1006088 207460 1006090
rect 207197 1006032 207202 1006088
rect 207258 1006032 207460 1006088
rect 207197 1006030 207460 1006032
rect 207565 1006088 207828 1006090
rect 207565 1006032 207570 1006088
rect 207626 1006032 207828 1006088
rect 207565 1006030 207828 1006032
rect 209484 1006088 209655 1006090
rect 209484 1006032 209594 1006088
rect 209650 1006032 209655 1006088
rect 209484 1006030 209655 1006032
rect 252264 1006088 252527 1006090
rect 252264 1006032 252466 1006088
rect 252522 1006032 252527 1006088
rect 252264 1006030 252527 1006032
rect 252724 1006030 253092 1006090
rect 253289 1006088 253460 1006090
rect 253289 1006032 253294 1006088
rect 253350 1006032 253460 1006088
rect 253289 1006030 253460 1006032
rect 256969 1006088 257140 1006090
rect 256969 1006032 256974 1006088
rect 257030 1006032 257140 1006088
rect 256969 1006030 257140 1006032
rect 258533 1006088 258796 1006090
rect 258533 1006032 258538 1006088
rect 258594 1006032 258796 1006088
rect 258533 1006030 258796 1006032
rect 258993 1006088 259164 1006090
rect 258993 1006032 258998 1006088
rect 259054 1006032 259164 1006088
rect 258993 1006030 259164 1006032
rect 260820 1006088 261083 1006090
rect 260820 1006032 261022 1006088
rect 261078 1006032 261083 1006088
rect 260820 1006030 261083 1006032
rect 303876 1006088 304139 1006090
rect 303876 1006032 304078 1006088
rect 304134 1006032 304139 1006088
rect 303876 1006030 304139 1006032
rect 304244 1006030 304704 1006090
rect 304901 1006088 305164 1006090
rect 304901 1006032 304906 1006088
rect 304962 1006032 305164 1006088
rect 304901 1006030 305164 1006032
rect 305269 1006088 305532 1006090
rect 305269 1006032 305274 1006088
rect 305330 1006032 305532 1006088
rect 305269 1006030 305532 1006032
rect 314916 1006088 315179 1006090
rect 314916 1006032 315118 1006088
rect 315174 1006032 315179 1006088
rect 314916 1006030 315179 1006032
rect 354292 1006088 354555 1006090
rect 354292 1006032 354494 1006088
rect 354550 1006032 354555 1006088
rect 354292 1006030 354555 1006032
rect 354660 1006030 355120 1006090
rect 355225 1006088 355488 1006090
rect 355225 1006032 355230 1006088
rect 355286 1006032 355488 1006088
rect 355225 1006030 355488 1006032
rect 356684 1006088 356947 1006090
rect 356684 1006032 356886 1006088
rect 356942 1006032 356947 1006088
rect 356684 1006030 356947 1006032
rect 358340 1006088 358603 1006090
rect 358340 1006032 358542 1006088
rect 358598 1006032 358603 1006088
rect 358340 1006030 358603 1006032
rect 361192 1006088 361455 1006090
rect 361192 1006032 361394 1006088
rect 361450 1006032 361455 1006088
rect 361192 1006030 361455 1006032
rect 422096 1006030 422556 1006090
rect 422661 1006088 422924 1006090
rect 422661 1006032 422666 1006088
rect 422722 1006032 422924 1006088
rect 422661 1006030 422924 1006032
rect 423292 1006088 423555 1006090
rect 423292 1006032 423494 1006088
rect 423550 1006032 423555 1006088
rect 423292 1006030 423555 1006032
rect 427800 1006088 428063 1006090
rect 427800 1006032 428002 1006088
rect 428058 1006032 428063 1006088
rect 427800 1006030 428063 1006032
rect 429824 1006088 430087 1006090
rect 429824 1006032 430026 1006088
rect 430082 1006032 430087 1006088
rect 429824 1006030 430087 1006032
rect 499100 1006030 499468 1006090
rect 499665 1006088 499928 1006090
rect 499665 1006032 499670 1006088
rect 499726 1006032 499928 1006088
rect 499665 1006030 499928 1006032
rect 500296 1006088 500559 1006090
rect 500296 1006032 500498 1006088
rect 500554 1006032 500559 1006088
rect 500296 1006030 500559 1006032
rect 502412 1006088 502583 1006090
rect 502412 1006032 502522 1006088
rect 502578 1006032 502583 1006088
rect 502412 1006030 502583 1006032
rect 550068 1006088 550331 1006090
rect 550068 1006032 550270 1006088
rect 550326 1006032 550331 1006088
rect 550068 1006030 550331 1006032
rect 550436 1006030 550896 1006090
rect 551093 1006088 551356 1006090
rect 551093 1006032 551098 1006088
rect 551154 1006032 551356 1006088
rect 551093 1006030 551356 1006032
rect 552092 1006088 552355 1006090
rect 552092 1006032 552294 1006088
rect 552350 1006032 552355 1006088
rect 552092 1006030 552355 1006032
rect 556600 1006088 556863 1006090
rect 556600 1006032 556802 1006088
rect 556858 1006032 556863 1006088
rect 556600 1006030 556863 1006032
rect 160645 1006027 160711 1006030
rect 201033 1006027 201099 1006030
rect 201861 1006027 201927 1006030
rect 207197 1006027 207263 1006030
rect 207565 1006027 207631 1006030
rect 209589 1006027 209655 1006030
rect 252461 1006027 252527 1006030
rect 253289 1006027 253355 1006030
rect 256969 1006027 257035 1006030
rect 258533 1006027 258599 1006030
rect 258993 1006027 259059 1006030
rect 261017 1006027 261083 1006030
rect 304073 1006027 304139 1006030
rect 304901 1006027 304967 1006030
rect 305269 1006027 305335 1006030
rect 315113 1006027 315179 1006030
rect 354489 1006027 354555 1006030
rect 355225 1006027 355291 1006030
rect 356881 1006027 356947 1006030
rect 358537 1006027 358603 1006030
rect 361389 1006027 361455 1006030
rect 422661 1006027 422727 1006030
rect 423489 1006027 423555 1006030
rect 427997 1006027 428063 1006030
rect 430021 1006027 430087 1006030
rect 499665 1006027 499731 1006030
rect 500493 1006027 500559 1006030
rect 502517 1006027 502583 1006030
rect 550265 1006027 550331 1006030
rect 551093 1006027 551159 1006030
rect 552289 1006027 552355 1006030
rect 556797 1006027 556863 1006030
rect 360561 1005410 360627 1005413
rect 361021 1005410 361087 1005413
rect 360364 1005408 360627 1005410
rect 360364 1005352 360566 1005408
rect 360622 1005352 360627 1005408
rect 360364 1005350 360627 1005352
rect 360824 1005408 361087 1005410
rect 360824 1005352 361026 1005408
rect 361082 1005352 361087 1005408
rect 360824 1005350 361087 1005352
rect 360561 1005347 360627 1005350
rect 361021 1005347 361087 1005350
rect 360193 1005274 360259 1005277
rect 503345 1005274 503411 1005277
rect 359996 1005272 360259 1005274
rect 359996 1005216 360198 1005272
rect 360254 1005216 360259 1005272
rect 359996 1005214 360259 1005216
rect 503148 1005272 503411 1005274
rect 503148 1005216 503350 1005272
rect 503406 1005216 503411 1005272
rect 503148 1005214 503411 1005216
rect 360193 1005211 360259 1005214
rect 503345 1005211 503411 1005214
rect 508681 1005138 508747 1005141
rect 508484 1005136 508747 1005138
rect 508484 1005080 508686 1005136
rect 508742 1005080 508747 1005136
rect 508484 1005078 508747 1005080
rect 508681 1005075 508747 1005078
rect 507025 1005002 507091 1005005
rect 508221 1005002 508287 1005005
rect 506828 1005000 507091 1005002
rect 506828 1004944 507030 1005000
rect 507086 1004944 507091 1005000
rect 506828 1004942 507091 1004944
rect 508116 1005000 508287 1005002
rect 508116 1004944 508226 1005000
rect 508282 1004944 508287 1005000
rect 508116 1004942 508287 1004944
rect 507025 1004939 507091 1004942
rect 508221 1004939 508287 1004942
rect 159449 1004866 159515 1004869
rect 159817 1004866 159883 1004869
rect 208761 1004866 208827 1004869
rect 159252 1004864 159515 1004866
rect 159252 1004808 159454 1004864
rect 159510 1004808 159515 1004864
rect 159252 1004806 159515 1004808
rect 159712 1004864 159883 1004866
rect 159712 1004808 159822 1004864
rect 159878 1004808 159883 1004864
rect 159712 1004806 159883 1004808
rect 208656 1004864 208827 1004866
rect 208656 1004808 208766 1004864
rect 208822 1004808 208827 1004864
rect 208656 1004806 208827 1004808
rect 159449 1004803 159515 1004806
rect 159817 1004803 159883 1004806
rect 208761 1004803 208827 1004806
rect 306925 1004866 306991 1004869
rect 313825 1004866 313891 1004869
rect 363413 1004866 363479 1004869
rect 364241 1004866 364307 1004869
rect 306925 1004864 307188 1004866
rect 306925 1004808 306930 1004864
rect 306986 1004808 307188 1004864
rect 306925 1004806 307188 1004808
rect 313628 1004864 313891 1004866
rect 313628 1004808 313830 1004864
rect 313886 1004808 313891 1004864
rect 313628 1004806 313891 1004808
rect 363308 1004864 363479 1004866
rect 363308 1004808 363418 1004864
rect 363474 1004808 363479 1004864
rect 363308 1004806 363479 1004808
rect 364044 1004864 364307 1004866
rect 364044 1004808 364246 1004864
rect 364302 1004808 364307 1004864
rect 364044 1004806 364307 1004808
rect 306925 1004803 306991 1004806
rect 313825 1004803 313891 1004806
rect 363413 1004803 363479 1004806
rect 364241 1004803 364307 1004806
rect 501321 1004866 501387 1004869
rect 507853 1004866 507919 1004869
rect 501321 1004864 501492 1004866
rect 501321 1004808 501326 1004864
rect 501382 1004808 501492 1004864
rect 501321 1004806 501492 1004808
rect 507656 1004864 507919 1004866
rect 507656 1004808 507858 1004864
rect 507914 1004808 507919 1004864
rect 507656 1004806 507919 1004808
rect 501321 1004803 501387 1004806
rect 507853 1004803 507919 1004806
rect 103145 1004730 103211 1004733
rect 160277 1004730 160343 1004733
rect 160645 1004730 160711 1004733
rect 102948 1004728 103211 1004730
rect 102948 1004672 103150 1004728
rect 103206 1004672 103211 1004728
rect 102948 1004670 103211 1004672
rect 160080 1004728 160343 1004730
rect 160080 1004672 160282 1004728
rect 160338 1004672 160343 1004728
rect 160080 1004670 160343 1004672
rect 160540 1004728 160711 1004730
rect 160540 1004672 160650 1004728
rect 160706 1004672 160711 1004728
rect 160540 1004670 160711 1004672
rect 103145 1004667 103211 1004670
rect 160277 1004667 160343 1004670
rect 160645 1004667 160711 1004670
rect 202229 1004730 202295 1004733
rect 208393 1004730 208459 1004733
rect 209221 1004730 209287 1004733
rect 202229 1004728 202492 1004730
rect 202229 1004672 202234 1004728
rect 202290 1004672 202492 1004728
rect 202229 1004670 202492 1004672
rect 208196 1004728 208459 1004730
rect 208196 1004672 208398 1004728
rect 208454 1004672 208459 1004728
rect 208196 1004670 208459 1004672
rect 209024 1004728 209287 1004730
rect 209024 1004672 209226 1004728
rect 209282 1004672 209287 1004728
rect 209024 1004670 209287 1004672
rect 202229 1004667 202295 1004670
rect 208393 1004667 208459 1004670
rect 209221 1004667 209287 1004670
rect 307753 1004730 307819 1004733
rect 308581 1004730 308647 1004733
rect 314653 1004730 314719 1004733
rect 315481 1004730 315547 1004733
rect 307753 1004728 307924 1004730
rect 307753 1004672 307758 1004728
rect 307814 1004672 307924 1004728
rect 307753 1004670 307924 1004672
rect 308581 1004728 308752 1004730
rect 308581 1004672 308586 1004728
rect 308642 1004672 308752 1004728
rect 308581 1004670 308752 1004672
rect 314548 1004728 314719 1004730
rect 314548 1004672 314658 1004728
rect 314714 1004672 314719 1004728
rect 314548 1004670 314719 1004672
rect 315284 1004728 315547 1004730
rect 315284 1004672 315486 1004728
rect 315542 1004672 315547 1004728
rect 315284 1004670 315547 1004672
rect 307753 1004667 307819 1004670
rect 308581 1004667 308647 1004670
rect 314653 1004667 314719 1004670
rect 315481 1004667 315547 1004670
rect 356053 1004730 356119 1004733
rect 356881 1004730 356947 1004733
rect 361849 1004730 361915 1004733
rect 362585 1004730 362651 1004733
rect 356053 1004728 356316 1004730
rect 356053 1004672 356058 1004728
rect 356114 1004672 356316 1004728
rect 356053 1004670 356316 1004672
rect 356881 1004728 357144 1004730
rect 356881 1004672 356886 1004728
rect 356942 1004672 357144 1004728
rect 356881 1004670 357144 1004672
rect 361652 1004728 361915 1004730
rect 361652 1004672 361854 1004728
rect 361910 1004672 361915 1004728
rect 361652 1004670 361915 1004672
rect 362388 1004728 362651 1004730
rect 362388 1004672 362590 1004728
rect 362646 1004672 362651 1004728
rect 362388 1004670 362651 1004672
rect 356053 1004667 356119 1004670
rect 356881 1004667 356947 1004670
rect 361849 1004667 361915 1004670
rect 362585 1004667 362651 1004670
rect 500493 1004730 500559 1004733
rect 500861 1004730 500927 1004733
rect 507393 1004730 507459 1004733
rect 509049 1004730 509115 1004733
rect 556337 1004730 556403 1004733
rect 557625 1004730 557691 1004733
rect 500493 1004728 500756 1004730
rect 500493 1004672 500498 1004728
rect 500554 1004672 500756 1004728
rect 500493 1004670 500756 1004672
rect 500861 1004728 501124 1004730
rect 500861 1004672 500866 1004728
rect 500922 1004672 501124 1004728
rect 500861 1004670 501124 1004672
rect 507196 1004728 507459 1004730
rect 507196 1004672 507398 1004728
rect 507454 1004672 507459 1004728
rect 507196 1004670 507459 1004672
rect 508852 1004728 509115 1004730
rect 508852 1004672 509054 1004728
rect 509110 1004672 509115 1004728
rect 508852 1004670 509115 1004672
rect 556232 1004728 556403 1004730
rect 556232 1004672 556342 1004728
rect 556398 1004672 556403 1004728
rect 556232 1004670 556403 1004672
rect 557428 1004728 557691 1004730
rect 557428 1004672 557630 1004728
rect 557686 1004672 557691 1004728
rect 557428 1004670 557691 1004672
rect 500493 1004667 500559 1004670
rect 500861 1004667 500927 1004670
rect 507393 1004667 507459 1004670
rect 509049 1004667 509115 1004670
rect 556337 1004667 556403 1004670
rect 557625 1004667 557691 1004670
rect 308949 1004594 309015 1004597
rect 423857 1004594 423923 1004597
rect 308949 1004592 309212 1004594
rect 308949 1004536 308954 1004592
rect 309010 1004536 309212 1004592
rect 308949 1004534 309212 1004536
rect 423857 1004592 424120 1004594
rect 423857 1004536 423862 1004592
rect 423918 1004536 424120 1004592
rect 423857 1004534 424120 1004536
rect 308949 1004531 309015 1004534
rect 423857 1004531 423923 1004534
rect 424685 1004050 424751 1004053
rect 424580 1004048 424751 1004050
rect 424580 1003992 424690 1004048
rect 424746 1003992 424751 1004048
rect 424580 1003990 424751 1003992
rect 424685 1003987 424751 1003990
rect 423489 1003914 423555 1003917
rect 503713 1003914 503779 1003917
rect 423489 1003912 423752 1003914
rect 423489 1003856 423494 1003912
rect 423550 1003856 423752 1003912
rect 423489 1003854 423752 1003856
rect 503608 1003912 503779 1003914
rect 503608 1003856 503718 1003912
rect 503774 1003856 503779 1003912
rect 503608 1003854 503779 1003856
rect 423489 1003851 423555 1003854
rect 503713 1003851 503779 1003854
rect 99465 1003370 99531 1003373
rect 554773 1003370 554839 1003373
rect 99465 1003368 99728 1003370
rect 99465 1003312 99470 1003368
rect 99526 1003312 99728 1003368
rect 99465 1003310 99728 1003312
rect 554773 1003368 555036 1003370
rect 554773 1003312 554778 1003368
rect 554834 1003312 555036 1003368
rect 554773 1003310 555036 1003312
rect 99465 1003307 99531 1003310
rect 554773 1003307 554839 1003310
rect 553945 1002690 554011 1002693
rect 553945 1002688 554116 1002690
rect 553945 1002632 553950 1002688
rect 554006 1002632 554116 1002688
rect 553945 1002630 554116 1002632
rect 553945 1002627 554011 1002630
rect 154573 1002554 154639 1002557
rect 425973 1002554 426039 1002557
rect 154573 1002552 154836 1002554
rect 154573 1002496 154578 1002552
rect 154634 1002496 154836 1002552
rect 154573 1002494 154836 1002496
rect 425776 1002552 426039 1002554
rect 425776 1002496 425978 1002552
rect 426034 1002496 426039 1002552
rect 425776 1002494 426039 1002496
rect 154573 1002491 154639 1002494
rect 425973 1002491 426039 1002494
rect 554313 1002554 554379 1002557
rect 554313 1002552 554576 1002554
rect 554313 1002496 554318 1002552
rect 554374 1002496 554576 1002552
rect 554313 1002494 554576 1002496
rect 554313 1002491 554379 1002494
rect 106825 1002418 106891 1002421
rect 559189 1002418 559255 1002421
rect 560845 1002418 560911 1002421
rect 106628 1002416 106891 1002418
rect 106628 1002360 106830 1002416
rect 106886 1002360 106891 1002416
rect 106628 1002358 106891 1002360
rect 559084 1002416 559255 1002418
rect 559084 1002360 559194 1002416
rect 559250 1002360 559255 1002416
rect 559084 1002358 559255 1002360
rect 560740 1002416 560911 1002418
rect 560740 1002360 560850 1002416
rect 560906 1002360 560911 1002416
rect 560740 1002358 560911 1002360
rect 106825 1002355 106891 1002358
rect 559189 1002355 559255 1002358
rect 560845 1002355 560911 1002358
rect 101489 1002282 101555 1002285
rect 105997 1002282 106063 1002285
rect 101489 1002280 101752 1002282
rect 101489 1002224 101494 1002280
rect 101550 1002224 101752 1002280
rect 101489 1002222 101752 1002224
rect 105892 1002280 106063 1002282
rect 105892 1002224 106002 1002280
rect 106058 1002224 106063 1002280
rect 105892 1002222 106063 1002224
rect 101489 1002219 101555 1002222
rect 105997 1002219 106063 1002222
rect 108481 1002282 108547 1002285
rect 158253 1002282 158319 1002285
rect 108481 1002280 108652 1002282
rect 108481 1002224 108486 1002280
rect 108542 1002224 108652 1002280
rect 108481 1002222 108652 1002224
rect 158056 1002280 158319 1002282
rect 158056 1002224 158258 1002280
rect 158314 1002224 158319 1002280
rect 158056 1002222 158319 1002224
rect 108481 1002219 108547 1002222
rect 158253 1002219 158319 1002222
rect 205173 1002282 205239 1002285
rect 211613 1002282 211679 1002285
rect 205173 1002280 205344 1002282
rect 205173 1002224 205178 1002280
rect 205234 1002224 205344 1002280
rect 205173 1002222 205344 1002224
rect 211508 1002280 211679 1002282
rect 211508 1002224 211618 1002280
rect 211674 1002224 211679 1002280
rect 211508 1002222 211679 1002224
rect 205173 1002219 205239 1002222
rect 211613 1002219 211679 1002222
rect 254485 1002282 254551 1002285
rect 261477 1002282 261543 1002285
rect 261845 1002282 261911 1002285
rect 254485 1002280 254748 1002282
rect 254485 1002224 254490 1002280
rect 254546 1002224 254748 1002280
rect 254485 1002222 254748 1002224
rect 261280 1002280 261543 1002282
rect 261280 1002224 261482 1002280
rect 261538 1002224 261543 1002280
rect 261280 1002222 261543 1002224
rect 261648 1002280 261911 1002282
rect 261648 1002224 261850 1002280
rect 261906 1002224 261911 1002280
rect 261648 1002222 261911 1002224
rect 254485 1002219 254551 1002222
rect 261477 1002219 261543 1002222
rect 261845 1002219 261911 1002222
rect 502517 1002282 502583 1002285
rect 558453 1002282 558519 1002285
rect 559649 1002282 559715 1002285
rect 502517 1002280 502780 1002282
rect 502517 1002224 502522 1002280
rect 502578 1002224 502780 1002280
rect 502517 1002222 502780 1002224
rect 558256 1002280 558519 1002282
rect 558256 1002224 558458 1002280
rect 558514 1002224 558519 1002280
rect 558256 1002222 558519 1002224
rect 559452 1002280 559715 1002282
rect 559452 1002224 559654 1002280
rect 559710 1002224 559715 1002280
rect 559452 1002222 559715 1002224
rect 502517 1002219 502583 1002222
rect 558453 1002219 558519 1002222
rect 559649 1002219 559715 1002222
rect 100293 1002146 100359 1002149
rect 102317 1002146 102383 1002149
rect 105629 1002146 105695 1002149
rect 107653 1002146 107719 1002149
rect 108021 1002146 108087 1002149
rect 157425 1002146 157491 1002149
rect 157793 1002146 157859 1002149
rect 100293 1002144 100556 1002146
rect 100293 1002088 100298 1002144
rect 100354 1002088 100556 1002144
rect 100293 1002086 100556 1002088
rect 102317 1002144 102580 1002146
rect 102317 1002088 102322 1002144
rect 102378 1002088 102580 1002144
rect 102317 1002086 102580 1002088
rect 105432 1002144 105695 1002146
rect 105432 1002088 105634 1002144
rect 105690 1002088 105695 1002144
rect 105432 1002086 105695 1002088
rect 107456 1002144 107719 1002146
rect 107456 1002088 107658 1002144
rect 107714 1002088 107719 1002144
rect 107456 1002086 107719 1002088
rect 107916 1002144 108087 1002146
rect 107916 1002088 108026 1002144
rect 108082 1002088 108087 1002144
rect 107916 1002086 108087 1002088
rect 157228 1002144 157491 1002146
rect 157228 1002088 157430 1002144
rect 157486 1002088 157491 1002144
rect 157228 1002086 157491 1002088
rect 157596 1002144 157859 1002146
rect 157596 1002088 157798 1002144
rect 157854 1002088 157859 1002144
rect 157596 1002086 157859 1002088
rect 100293 1002083 100359 1002086
rect 102317 1002083 102383 1002086
rect 105629 1002083 105695 1002086
rect 107653 1002083 107719 1002086
rect 108021 1002083 108087 1002086
rect 157425 1002083 157491 1002086
rect 157793 1002083 157859 1002086
rect 203517 1002146 203583 1002149
rect 205909 1002146 205975 1002149
rect 210417 1002146 210483 1002149
rect 211245 1002146 211311 1002149
rect 203517 1002144 203780 1002146
rect 203517 1002088 203522 1002144
rect 203578 1002088 203780 1002144
rect 203517 1002086 203780 1002088
rect 205909 1002144 206172 1002146
rect 205909 1002088 205914 1002144
rect 205970 1002088 206172 1002144
rect 205909 1002086 206172 1002088
rect 210220 1002144 210483 1002146
rect 210220 1002088 210422 1002144
rect 210478 1002088 210483 1002144
rect 210220 1002086 210483 1002088
rect 211140 1002144 211311 1002146
rect 211140 1002088 211250 1002144
rect 211306 1002088 211311 1002144
rect 211140 1002086 211311 1002088
rect 203517 1002083 203583 1002086
rect 205909 1002083 205975 1002086
rect 210417 1002083 210483 1002086
rect 211245 1002083 211311 1002086
rect 255681 1002146 255747 1002149
rect 256141 1002146 256207 1002149
rect 259821 1002146 259887 1002149
rect 255681 1002144 255944 1002146
rect 255681 1002088 255686 1002144
rect 255742 1002088 255944 1002144
rect 255681 1002086 255944 1002088
rect 256141 1002144 256404 1002146
rect 256141 1002088 256146 1002144
rect 256202 1002088 256404 1002144
rect 256141 1002086 256404 1002088
rect 259624 1002144 259887 1002146
rect 259624 1002088 259826 1002144
rect 259882 1002088 259887 1002144
rect 259624 1002086 259887 1002088
rect 255681 1002083 255747 1002086
rect 256141 1002083 256207 1002086
rect 259821 1002083 259887 1002086
rect 261845 1002146 261911 1002149
rect 262673 1002146 262739 1002149
rect 263501 1002146 263567 1002149
rect 310145 1002146 310211 1002149
rect 365069 1002146 365135 1002149
rect 261845 1002144 262108 1002146
rect 261845 1002088 261850 1002144
rect 261906 1002088 262108 1002144
rect 261845 1002086 262108 1002088
rect 262476 1002144 262739 1002146
rect 262476 1002088 262678 1002144
rect 262734 1002088 262739 1002144
rect 262476 1002086 262739 1002088
rect 263304 1002144 263567 1002146
rect 263304 1002088 263506 1002144
rect 263562 1002088 263567 1002144
rect 263304 1002086 263567 1002088
rect 309948 1002144 310211 1002146
rect 309948 1002088 310150 1002144
rect 310206 1002088 310211 1002144
rect 309948 1002086 310211 1002088
rect 364872 1002144 365135 1002146
rect 364872 1002088 365074 1002144
rect 365130 1002088 365135 1002144
rect 364872 1002086 365135 1002088
rect 261845 1002083 261911 1002086
rect 262673 1002083 262739 1002086
rect 263501 1002083 263567 1002086
rect 310145 1002083 310211 1002086
rect 365069 1002083 365135 1002086
rect 425973 1002146 426039 1002149
rect 503713 1002146 503779 1002149
rect 509509 1002146 509575 1002149
rect 425973 1002144 426144 1002146
rect 425973 1002088 425978 1002144
rect 426034 1002088 426144 1002144
rect 425973 1002086 426144 1002088
rect 503713 1002144 503976 1002146
rect 503713 1002088 503718 1002144
rect 503774 1002088 503976 1002144
rect 503713 1002086 503976 1002088
rect 509312 1002144 509575 1002146
rect 509312 1002088 509514 1002144
rect 509570 1002088 509575 1002144
rect 509312 1002086 509575 1002088
rect 425973 1002083 426039 1002086
rect 503713 1002083 503779 1002086
rect 509509 1002083 509575 1002086
rect 552289 1002146 552355 1002149
rect 553117 1002146 553183 1002149
rect 560017 1002146 560083 1002149
rect 560477 1002146 560543 1002149
rect 552289 1002144 552552 1002146
rect 552289 1002088 552294 1002144
rect 552350 1002088 552552 1002144
rect 552289 1002086 552552 1002088
rect 553117 1002144 553380 1002146
rect 553117 1002088 553122 1002144
rect 553178 1002088 553380 1002144
rect 553117 1002086 553380 1002088
rect 559820 1002144 560083 1002146
rect 559820 1002088 560022 1002144
rect 560078 1002088 560083 1002144
rect 559820 1002086 560083 1002088
rect 560280 1002144 560543 1002146
rect 560280 1002088 560482 1002144
rect 560538 1002088 560543 1002144
rect 560280 1002086 560543 1002088
rect 552289 1002083 552355 1002086
rect 553117 1002083 553183 1002086
rect 560017 1002083 560083 1002086
rect 560477 1002083 560543 1002086
rect 101121 1002010 101187 1002013
rect 101949 1002010 102015 1002013
rect 104341 1002010 104407 1002013
rect 106457 1002010 106523 1002013
rect 107193 1002010 107259 1002013
rect 108481 1002010 108547 1002013
rect 109677 1002010 109743 1002013
rect 156965 1002010 157031 1002013
rect 158621 1002010 158687 1002013
rect 101121 1002008 101292 1002010
rect 101121 1001952 101126 1002008
rect 101182 1001952 101292 1002008
rect 101121 1001950 101292 1001952
rect 101949 1002008 102212 1002010
rect 101949 1001952 101954 1002008
rect 102010 1001952 102212 1002008
rect 101949 1001950 102212 1001952
rect 104236 1002008 104407 1002010
rect 104236 1001952 104346 1002008
rect 104402 1001952 104407 1002008
rect 104236 1001950 104407 1001952
rect 106260 1002008 106523 1002010
rect 106260 1001952 106462 1002008
rect 106518 1001952 106523 1002008
rect 106260 1001950 106523 1001952
rect 107088 1002008 107259 1002010
rect 107088 1001952 107198 1002008
rect 107254 1001952 107259 1002008
rect 107088 1001950 107259 1001952
rect 108284 1002008 108547 1002010
rect 108284 1001952 108486 1002008
rect 108542 1001952 108547 1002008
rect 108284 1001950 108547 1001952
rect 109480 1002008 109743 1002010
rect 109480 1001952 109682 1002008
rect 109738 1001952 109743 1002008
rect 109480 1001950 109743 1001952
rect 156860 1002008 157031 1002010
rect 156860 1001952 156970 1002008
rect 157026 1001952 157031 1002008
rect 156860 1001950 157031 1001952
rect 158516 1002008 158687 1002010
rect 158516 1001952 158626 1002008
rect 158682 1001952 158687 1002008
rect 158516 1001950 158687 1001952
rect 101121 1001947 101187 1001950
rect 101949 1001947 102015 1001950
rect 104341 1001947 104407 1001950
rect 106457 1001947 106523 1001950
rect 107193 1001947 107259 1001950
rect 108481 1001947 108547 1001950
rect 109677 1001947 109743 1001950
rect 156965 1001947 157031 1001950
rect 158621 1001947 158687 1001950
rect 203057 1002010 203123 1002013
rect 204713 1002010 204779 1002013
rect 205541 1002010 205607 1002013
rect 206737 1002010 206803 1002013
rect 212073 1002010 212139 1002013
rect 212533 1002010 212599 1002013
rect 203057 1002008 203320 1002010
rect 203057 1001952 203062 1002008
rect 203118 1001952 203320 1002008
rect 203057 1001950 203320 1001952
rect 204713 1002008 204976 1002010
rect 204713 1001952 204718 1002008
rect 204774 1001952 204976 1002008
rect 204713 1001950 204976 1001952
rect 205541 1002008 205804 1002010
rect 205541 1001952 205546 1002008
rect 205602 1001952 205804 1002008
rect 205541 1001950 205804 1001952
rect 206737 1002008 207000 1002010
rect 206737 1001952 206742 1002008
rect 206798 1001952 207000 1002008
rect 206737 1001950 207000 1001952
rect 211876 1002008 212139 1002010
rect 211876 1001952 212078 1002008
rect 212134 1001952 212139 1002008
rect 211876 1001950 212139 1001952
rect 212336 1002008 212599 1002010
rect 212336 1001952 212538 1002008
rect 212594 1001952 212599 1002008
rect 212336 1001950 212599 1001952
rect 203057 1001947 203123 1001950
rect 204713 1001947 204779 1001950
rect 205541 1001947 205607 1001950
rect 206737 1001947 206803 1001950
rect 212073 1001947 212139 1001950
rect 212533 1001947 212599 1001950
rect 254117 1002010 254183 1002013
rect 256509 1002010 256575 1002013
rect 260189 1002010 260255 1002013
rect 260649 1002010 260715 1002013
rect 263041 1002010 263107 1002013
rect 263869 1002010 263935 1002013
rect 254117 1002008 254380 1002010
rect 254117 1001952 254122 1002008
rect 254178 1001952 254380 1002008
rect 254117 1001950 254380 1001952
rect 256509 1002008 256772 1002010
rect 256509 1001952 256514 1002008
rect 256570 1001952 256772 1002008
rect 256509 1001950 256772 1001952
rect 260084 1002008 260255 1002010
rect 260084 1001952 260194 1002008
rect 260250 1001952 260255 1002008
rect 260084 1001950 260255 1001952
rect 260452 1002008 260715 1002010
rect 260452 1001952 260654 1002008
rect 260710 1001952 260715 1002008
rect 260452 1001950 260715 1001952
rect 262844 1002008 263107 1002010
rect 262844 1001952 263046 1002008
rect 263102 1001952 263107 1002008
rect 262844 1001950 263107 1001952
rect 263764 1002008 263935 1002010
rect 263764 1001952 263874 1002008
rect 263930 1001952 263935 1002008
rect 263764 1001950 263935 1001952
rect 254117 1001947 254183 1001950
rect 256509 1001947 256575 1001950
rect 260189 1001947 260255 1001950
rect 260649 1001947 260715 1001950
rect 263041 1001947 263107 1001950
rect 263869 1001947 263935 1001950
rect 305729 1002010 305795 1002013
rect 306097 1002010 306163 1002013
rect 309317 1002010 309383 1002013
rect 310145 1002010 310211 1002013
rect 311433 1002010 311499 1002013
rect 312261 1002010 312327 1002013
rect 312997 1002010 313063 1002013
rect 305729 1002008 305900 1002010
rect 305729 1001952 305734 1002008
rect 305790 1001952 305900 1002008
rect 305729 1001950 305900 1001952
rect 306097 1002008 306360 1002010
rect 306097 1001952 306102 1002008
rect 306158 1001952 306360 1002008
rect 306097 1001950 306360 1001952
rect 309317 1002008 309580 1002010
rect 309317 1001952 309322 1002008
rect 309378 1001952 309580 1002008
rect 309317 1001950 309580 1001952
rect 310145 1002008 310408 1002010
rect 310145 1001952 310150 1002008
rect 310206 1001952 310408 1002008
rect 310145 1001950 310408 1001952
rect 311236 1002008 311499 1002010
rect 311236 1001952 311438 1002008
rect 311494 1001952 311499 1002008
rect 311236 1001950 311499 1001952
rect 312064 1002008 312327 1002010
rect 312064 1001952 312266 1002008
rect 312322 1001952 312327 1002008
rect 312064 1001950 312327 1001952
rect 312892 1002008 313063 1002010
rect 312892 1001952 313002 1002008
rect 313058 1001952 313063 1002008
rect 312892 1001950 313063 1001952
rect 305729 1001947 305795 1001950
rect 306097 1001947 306163 1001950
rect 309317 1001947 309383 1001950
rect 310145 1001947 310211 1001950
rect 311433 1001947 311499 1001950
rect 312261 1001947 312327 1001950
rect 312997 1001947 313063 1001950
rect 358905 1002010 358971 1002013
rect 359365 1002010 359431 1002013
rect 365437 1002010 365503 1002013
rect 365897 1002010 365963 1002013
rect 358905 1002008 359168 1002010
rect 358905 1001952 358910 1002008
rect 358966 1001952 359168 1002008
rect 358905 1001950 359168 1001952
rect 359365 1002008 359628 1002010
rect 359365 1001952 359370 1002008
rect 359426 1001952 359628 1002008
rect 359365 1001950 359628 1001952
rect 365332 1002008 365503 1002010
rect 365332 1001952 365442 1002008
rect 365498 1001952 365503 1002008
rect 365332 1001950 365503 1001952
rect 365700 1002008 365963 1002010
rect 365700 1001952 365902 1002008
rect 365958 1001952 365963 1002008
rect 365700 1001950 365963 1001952
rect 358905 1001947 358971 1001950
rect 359365 1001947 359431 1001950
rect 365437 1001947 365503 1001950
rect 365897 1001947 365963 1001950
rect 421465 1002010 421531 1002013
rect 425145 1002010 425211 1002013
rect 426341 1002010 426407 1002013
rect 426801 1002010 426867 1002013
rect 498469 1002010 498535 1002013
rect 501689 1002010 501755 1002013
rect 505829 1002010 505895 1002013
rect 506197 1002010 506263 1002013
rect 506565 1002010 506631 1002013
rect 509877 1002010 509943 1002013
rect 510337 1002010 510403 1002013
rect 421465 1002008 421636 1002010
rect 421465 1001952 421470 1002008
rect 421526 1001952 421636 1002008
rect 421465 1001950 421636 1001952
rect 425145 1002008 425316 1002010
rect 425145 1001952 425150 1002008
rect 425206 1001952 425316 1002008
rect 425145 1001950 425316 1001952
rect 426341 1002008 426604 1002010
rect 426341 1001952 426346 1002008
rect 426402 1001952 426604 1002008
rect 426341 1001950 426604 1001952
rect 426801 1002008 426972 1002010
rect 426801 1001952 426806 1002008
rect 426862 1001952 426972 1002008
rect 426801 1001950 426972 1001952
rect 498469 1002008 498732 1002010
rect 498469 1001952 498474 1002008
rect 498530 1001952 498732 1002008
rect 498469 1001950 498732 1001952
rect 501689 1002008 501952 1002010
rect 501689 1001952 501694 1002008
rect 501750 1001952 501952 1002008
rect 501689 1001950 501952 1001952
rect 505632 1002008 505895 1002010
rect 505632 1001952 505834 1002008
rect 505890 1001952 505895 1002008
rect 505632 1001950 505895 1001952
rect 506000 1002008 506263 1002010
rect 506000 1001952 506202 1002008
rect 506258 1001952 506263 1002008
rect 506000 1001950 506263 1001952
rect 506460 1002008 506631 1002010
rect 506460 1001952 506570 1002008
rect 506626 1001952 506631 1002008
rect 506460 1001950 506631 1001952
rect 509680 1002008 509943 1002010
rect 509680 1001952 509882 1002008
rect 509938 1001952 509943 1002008
rect 509680 1001950 509943 1001952
rect 510140 1002008 510403 1002010
rect 510140 1001952 510342 1002008
rect 510398 1001952 510403 1002008
rect 510140 1001950 510403 1001952
rect 421465 1001947 421531 1001950
rect 425145 1001947 425211 1001950
rect 426341 1001947 426407 1001950
rect 426801 1001947 426867 1001950
rect 498469 1001947 498535 1001950
rect 501689 1001947 501755 1001950
rect 505829 1001947 505895 1001950
rect 506197 1001947 506263 1001950
rect 506565 1001947 506631 1001950
rect 509877 1001947 509943 1001950
rect 510337 1001947 510403 1001950
rect 551461 1002010 551527 1002013
rect 552657 1002010 552723 1002013
rect 553485 1002010 553551 1002013
rect 555141 1002010 555207 1002013
rect 557993 1002010 558059 1002013
rect 558821 1002010 558887 1002013
rect 561305 1002010 561371 1002013
rect 561673 1002010 561739 1002013
rect 551461 1002008 551724 1002010
rect 551461 1001952 551466 1002008
rect 551522 1001952 551724 1002008
rect 551461 1001950 551724 1001952
rect 552657 1002008 552920 1002010
rect 552657 1001952 552662 1002008
rect 552718 1001952 552920 1002008
rect 552657 1001950 552920 1001952
rect 553485 1002008 553748 1002010
rect 553485 1001952 553490 1002008
rect 553546 1001952 553748 1002008
rect 553485 1001950 553748 1001952
rect 555141 1002008 555404 1002010
rect 555141 1001952 555146 1002008
rect 555202 1001952 555404 1002008
rect 555141 1001950 555404 1001952
rect 557796 1002008 558059 1002010
rect 557796 1001952 557998 1002008
rect 558054 1001952 558059 1002008
rect 557796 1001950 558059 1001952
rect 558624 1002008 558887 1002010
rect 558624 1001952 558826 1002008
rect 558882 1001952 558887 1002008
rect 558624 1001950 558887 1001952
rect 561108 1002008 561371 1002010
rect 561108 1001952 561310 1002008
rect 561366 1001952 561371 1002008
rect 561108 1001950 561371 1001952
rect 561476 1002008 561739 1002010
rect 561476 1001952 561678 1002008
rect 561734 1001952 561739 1002008
rect 561476 1001950 561739 1001952
rect 551461 1001947 551527 1001950
rect 552657 1001947 552723 1001950
rect 553485 1001947 553551 1001950
rect 555141 1001947 555207 1001950
rect 557993 1001947 558059 1001950
rect 558821 1001947 558887 1001950
rect 561305 1001947 561371 1001950
rect 561673 1001947 561739 1001950
rect 154941 1000650 155007 1000653
rect 154941 1000648 155204 1000650
rect 154941 1000592 154946 1000648
rect 155002 1000592 155204 1000648
rect 154941 1000590 155204 1000592
rect 154941 1000587 155007 1000590
rect 155769 999834 155835 999837
rect 428825 999834 428891 999837
rect 155769 999832 156032 999834
rect 155769 999776 155774 999832
rect 155830 999776 156032 999832
rect 155769 999774 156032 999776
rect 428628 999832 428891 999834
rect 428628 999776 428830 999832
rect 428886 999776 428891 999832
rect 428628 999774 428891 999776
rect 155769 999771 155835 999774
rect 428825 999771 428891 999774
rect 469397 998474 469463 998477
rect 472433 998474 472499 998477
rect 469397 998472 472499 998474
rect 469397 998416 469402 998472
rect 469458 998416 472438 998472
rect 472494 998416 472499 998472
rect 469397 998414 472499 998416
rect 469397 998411 469463 998414
rect 472433 998411 472499 998414
rect 459553 998338 459619 998341
rect 472709 998338 472775 998341
rect 459553 998336 472775 998338
rect 459553 998280 459558 998336
rect 459614 998280 472714 998336
rect 472770 998280 472775 998336
rect 459553 998278 472775 998280
rect 459553 998275 459619 998278
rect 472709 998275 472775 998278
rect 298461 998202 298527 998205
rect 300209 998202 300275 998205
rect 430849 998202 430915 998205
rect 298461 998200 300275 998202
rect 298461 998144 298466 998200
rect 298522 998144 300214 998200
rect 300270 998144 300275 998200
rect 298461 998142 300275 998144
rect 430652 998200 430915 998202
rect 430652 998144 430854 998200
rect 430910 998144 430915 998200
rect 430652 998142 430915 998144
rect 298461 998139 298527 998142
rect 300209 998139 300275 998142
rect 430849 998139 430915 998142
rect 151261 998066 151327 998069
rect 152917 998066 152983 998069
rect 429653 998066 429719 998069
rect 431677 998066 431743 998069
rect 151261 998064 151524 998066
rect 151261 998008 151266 998064
rect 151322 998008 151524 998064
rect 151261 998006 151524 998008
rect 152917 998064 153180 998066
rect 152917 998008 152922 998064
rect 152978 998008 153180 998064
rect 152917 998006 153180 998008
rect 429456 998064 429719 998066
rect 429456 998008 429658 998064
rect 429714 998008 429719 998064
rect 429456 998006 429719 998008
rect 431480 998064 431743 998066
rect 431480 998008 431682 998064
rect 431738 998008 431743 998064
rect 431480 998006 431743 998008
rect 151261 998003 151327 998006
rect 152917 998003 152983 998006
rect 429653 998003 429719 998006
rect 431677 998003 431743 998006
rect 152549 997930 152615 997933
rect 153745 997930 153811 997933
rect 430389 997930 430455 997933
rect 152549 997928 152720 997930
rect 152549 997872 152554 997928
rect 152610 997872 152720 997928
rect 152549 997870 152720 997872
rect 153745 997928 153916 997930
rect 153745 997872 153750 997928
rect 153806 997872 153916 997928
rect 153745 997870 153916 997872
rect 430284 997928 430455 997930
rect 430284 997872 430394 997928
rect 430450 997872 430455 997928
rect 430284 997870 430455 997872
rect 152549 997867 152615 997870
rect 153745 997867 153811 997870
rect 430389 997867 430455 997870
rect 430849 997930 430915 997933
rect 432413 997930 432479 997933
rect 432873 997930 432939 997933
rect 430849 997928 431020 997930
rect 430849 997872 430854 997928
rect 430910 997872 431020 997928
rect 430849 997870 431020 997872
rect 432308 997928 432479 997930
rect 432308 997872 432418 997928
rect 432474 997872 432479 997928
rect 432308 997870 432479 997872
rect 432676 997928 432939 997930
rect 432676 997872 432878 997928
rect 432934 997872 432939 997928
rect 432676 997870 432939 997872
rect 430849 997867 430915 997870
rect 432413 997867 432479 997870
rect 432873 997867 432939 997870
rect 153377 997794 153443 997797
rect 156137 997794 156203 997797
rect 253657 997794 253723 997797
rect 298185 997794 298251 997797
rect 303245 997794 303311 997797
rect 429193 997794 429259 997797
rect 432045 997794 432111 997797
rect 435357 997794 435423 997797
rect 153377 997792 153548 997794
rect 153377 997736 153382 997792
rect 153438 997736 153548 997792
rect 153377 997734 153548 997736
rect 156137 997792 156400 997794
rect 156137 997736 156142 997792
rect 156198 997736 156400 997792
rect 156137 997734 156400 997736
rect 253657 997792 253920 997794
rect 253657 997736 253662 997792
rect 253718 997736 253920 997792
rect 253657 997734 253920 997736
rect 298185 997792 303311 997794
rect 298185 997736 298190 997792
rect 298246 997736 303250 997792
rect 303306 997736 303311 997792
rect 298185 997734 303311 997736
rect 428996 997792 429259 997794
rect 428996 997736 429198 997792
rect 429254 997736 429259 997792
rect 428996 997734 429259 997736
rect 431940 997792 432111 997794
rect 431940 997736 432050 997792
rect 432106 997736 432111 997792
rect 431940 997734 432111 997736
rect 433136 997792 435423 997794
rect 433136 997736 435362 997792
rect 435418 997736 435423 997792
rect 433136 997734 435423 997736
rect 153377 997731 153443 997734
rect 156137 997731 156203 997734
rect 253657 997731 253723 997734
rect 298185 997731 298251 997734
rect 303245 997731 303311 997734
rect 429193 997731 429259 997734
rect 432045 997731 432111 997734
rect 435357 997731 435423 997734
rect 383561 997522 383627 997525
rect 383561 997520 383670 997522
rect 383561 997464 383566 997520
rect 383622 997464 383670 997520
rect 383561 997459 383670 997464
rect 383610 997389 383670 997459
rect 246430 997324 246436 997388
rect 246500 997386 246506 997388
rect 248321 997386 248387 997389
rect 246500 997384 248387 997386
rect 246500 997328 248326 997384
rect 248382 997328 248387 997384
rect 246500 997326 248387 997328
rect 383610 997384 383719 997389
rect 383610 997328 383658 997384
rect 383714 997328 383719 997384
rect 383610 997326 383719 997328
rect 246500 997324 246506 997326
rect 248321 997323 248387 997326
rect 383653 997323 383719 997326
rect 167637 997250 167703 997253
rect 200205 997250 200271 997253
rect 167637 997248 200271 997250
rect 167637 997192 167642 997248
rect 167698 997192 200210 997248
rect 200266 997192 200271 997248
rect 167637 997190 200271 997192
rect 167637 997187 167703 997190
rect 200205 997187 200271 997190
rect 238518 997188 238524 997252
rect 238588 997250 238594 997252
rect 249149 997250 249215 997253
rect 238588 997248 249215 997250
rect 238588 997192 249154 997248
rect 249210 997192 249215 997248
rect 238588 997190 249215 997192
rect 238588 997188 238594 997190
rect 249149 997187 249215 997190
rect 472617 997250 472683 997253
rect 480662 997250 480668 997252
rect 472617 997248 480668 997250
rect 472617 997192 472622 997248
rect 472678 997192 480668 997248
rect 472617 997190 480668 997192
rect 472617 997187 472683 997190
rect 480662 997188 480668 997190
rect 480732 997188 480738 997252
rect 524045 997250 524111 997253
rect 531998 997250 532004 997252
rect 524045 997248 532004 997250
rect 524045 997192 524050 997248
rect 524106 997192 532004 997248
rect 524045 997190 532004 997192
rect 524045 997187 524111 997190
rect 531998 997188 532004 997190
rect 532068 997188 532074 997252
rect 117221 997114 117287 997117
rect 144821 997114 144887 997117
rect 117221 997112 144887 997114
rect 117221 997056 117226 997112
rect 117282 997056 144826 997112
rect 144882 997056 144887 997112
rect 117221 997054 144887 997056
rect 117221 997051 117287 997054
rect 144821 997051 144887 997054
rect 372429 997114 372495 997117
rect 399937 997114 400003 997117
rect 372429 997112 400003 997114
rect 372429 997056 372434 997112
rect 372490 997056 399942 997112
rect 399998 997056 400003 997112
rect 372429 997054 400003 997056
rect 372429 997051 372495 997054
rect 399937 997051 400003 997054
rect 116301 996978 116367 996981
rect 144729 996978 144795 996981
rect 116301 996976 144795 996978
rect 116301 996920 116306 996976
rect 116362 996920 144734 996976
rect 144790 996920 144795 996976
rect 116301 996918 144795 996920
rect 116301 996915 116367 996918
rect 144729 996915 144795 996918
rect 167545 996978 167611 996981
rect 195237 996978 195303 996981
rect 167545 996976 195303 996978
rect 167545 996920 167550 996976
rect 167606 996920 195242 996976
rect 195298 996920 195303 996976
rect 167545 996918 195303 996920
rect 167545 996915 167611 996918
rect 195237 996915 195303 996918
rect 218881 996978 218947 996981
rect 246573 996978 246639 996981
rect 218881 996976 246639 996978
rect 218881 996920 218886 996976
rect 218942 996920 246578 996976
rect 246634 996920 246639 996976
rect 218881 996918 246639 996920
rect 218881 996915 218947 996918
rect 246573 996915 246639 996918
rect 270401 996978 270467 996981
rect 298737 996978 298803 996981
rect 270401 996976 298803 996978
rect 270401 996920 270406 996976
rect 270462 996920 298742 996976
rect 298798 996920 298803 996976
rect 270401 996918 298803 996920
rect 270401 996915 270467 996918
rect 298737 996915 298803 996918
rect 372521 996978 372587 996981
rect 400029 996978 400095 996981
rect 372521 996976 400095 996978
rect 372521 996920 372526 996976
rect 372582 996920 400034 996976
rect 400090 996920 400095 996976
rect 372521 996918 400095 996920
rect 372521 996915 372587 996918
rect 400029 996915 400095 996918
rect 439681 996978 439747 996981
rect 488901 996978 488967 996981
rect 439681 996976 488967 996978
rect 439681 996920 439686 996976
rect 439742 996920 488906 996976
rect 488962 996920 488967 996976
rect 439681 996918 488967 996920
rect 439681 996915 439747 996918
rect 488901 996915 488967 996918
rect 516777 996978 516843 996981
rect 540881 996978 540947 996981
rect 516777 996976 540947 996978
rect 516777 996920 516782 996976
rect 516838 996920 540886 996976
rect 540942 996920 540947 996976
rect 516777 996918 540947 996920
rect 516777 996915 516843 996918
rect 540881 996915 540947 996918
rect 590561 996706 590627 996709
rect 627862 996706 627868 996708
rect 590561 996704 627868 996706
rect 590561 996648 590566 996704
rect 590622 996648 627868 996704
rect 590561 996646 627868 996648
rect 590561 996643 590627 996646
rect 627862 996644 627868 996646
rect 627932 996644 627938 996708
rect 86534 996508 86540 996572
rect 86604 996570 86610 996572
rect 92513 996570 92579 996573
rect 86604 996568 92579 996570
rect 86604 996512 92518 996568
rect 92574 996512 92579 996568
rect 86604 996510 92579 996512
rect 86604 996508 86610 996510
rect 92513 996507 92579 996510
rect 520181 996570 520247 996573
rect 590561 996570 590627 996573
rect 630254 996570 630260 996572
rect 520181 996568 528018 996570
rect 520181 996512 520186 996568
rect 520242 996512 528018 996568
rect 520181 996510 528018 996512
rect 520181 996507 520247 996510
rect 89662 996372 89668 996436
rect 89732 996434 89738 996436
rect 93209 996434 93275 996437
rect 249701 996434 249767 996437
rect 303245 996434 303311 996437
rect 89732 996432 93275 996434
rect 89732 996376 93214 996432
rect 93270 996376 93275 996432
rect 89732 996374 93275 996376
rect 89732 996372 89738 996374
rect 93209 996371 93275 996374
rect 243862 996432 249767 996434
rect 243862 996376 249706 996432
rect 249762 996376 249767 996432
rect 243862 996374 249767 996376
rect 97257 996298 97323 996301
rect 84150 996296 97323 996298
rect 84150 996240 97262 996296
rect 97318 996240 97323 996296
rect 84150 996238 97323 996240
rect 82353 995618 82419 995621
rect 84150 995618 84210 996238
rect 97257 996235 97323 996238
rect 135294 996236 135300 996300
rect 135364 996298 135370 996300
rect 148869 996298 148935 996301
rect 200205 996298 200271 996301
rect 135364 996296 148935 996298
rect 135364 996240 148874 996296
rect 148930 996240 148935 996296
rect 135364 996238 148935 996240
rect 135364 996236 135370 996238
rect 148869 996235 148935 996238
rect 190410 996296 200271 996298
rect 190410 996240 200210 996296
rect 200266 996240 200271 996296
rect 190410 996238 200271 996240
rect 190410 996162 190470 996238
rect 200205 996235 200271 996238
rect 152733 995890 152799 995893
rect 132450 995888 152799 995890
rect 132450 995832 152738 995888
rect 152794 995832 152799 995888
rect 132450 995830 152799 995832
rect 86493 995756 86559 995757
rect 89621 995756 89687 995757
rect 86493 995754 86540 995756
rect 86448 995752 86540 995754
rect 86448 995696 86498 995752
rect 86448 995694 86540 995696
rect 86493 995692 86540 995694
rect 86604 995692 86610 995756
rect 89621 995754 89668 995756
rect 89576 995752 89668 995754
rect 89576 995696 89626 995752
rect 89576 995694 89668 995696
rect 89621 995692 89668 995694
rect 89732 995692 89738 995756
rect 131757 995754 131823 995757
rect 132450 995754 132510 995830
rect 152733 995827 152799 995830
rect 131757 995752 132510 995754
rect 131757 995696 131762 995752
rect 131818 995696 132510 995752
rect 131757 995694 132510 995696
rect 133045 995754 133111 995757
rect 135294 995754 135300 995756
rect 133045 995752 135300 995754
rect 133045 995696 133050 995752
rect 133106 995696 135300 995752
rect 133045 995694 135300 995696
rect 86493 995691 86559 995692
rect 89621 995691 89687 995692
rect 131757 995691 131823 995694
rect 133045 995691 133111 995694
rect 135294 995692 135300 995694
rect 135364 995692 135370 995756
rect 137921 995754 137987 995757
rect 142889 995754 142955 995757
rect 146937 995754 147003 995757
rect 137921 995752 142170 995754
rect 137921 995696 137926 995752
rect 137982 995696 142170 995752
rect 137921 995694 142170 995696
rect 137921 995691 137987 995694
rect 82353 995616 84210 995618
rect 82353 995560 82358 995616
rect 82414 995560 84210 995616
rect 82353 995558 84210 995560
rect 85941 995618 86007 995621
rect 93117 995618 93183 995621
rect 85941 995616 93183 995618
rect 85941 995560 85946 995616
rect 86002 995560 93122 995616
rect 93178 995560 93183 995616
rect 85941 995558 93183 995560
rect 142110 995618 142170 995694
rect 142889 995752 147003 995754
rect 142889 995696 142894 995752
rect 142950 995696 146942 995752
rect 146998 995696 147003 995752
rect 142889 995694 147003 995696
rect 142889 995691 142955 995694
rect 146937 995691 147003 995694
rect 144177 995618 144243 995621
rect 142110 995616 144243 995618
rect 142110 995560 144182 995616
rect 144238 995560 144243 995616
rect 142110 995558 144243 995560
rect 82353 995555 82419 995558
rect 85941 995555 86007 995558
rect 93117 995555 93183 995558
rect 144177 995555 144243 995558
rect 84653 995482 84719 995485
rect 92605 995482 92671 995485
rect 84653 995480 92671 995482
rect 84653 995424 84658 995480
rect 84714 995424 92610 995480
rect 92666 995424 92671 995480
rect 84653 995422 92671 995424
rect 84653 995419 84719 995422
rect 92605 995419 92671 995422
rect 137369 995482 137435 995485
rect 143993 995482 144059 995485
rect 137369 995480 144059 995482
rect 137369 995424 137374 995480
rect 137430 995424 143998 995480
rect 144054 995424 144059 995480
rect 137369 995422 144059 995424
rect 137369 995419 137435 995422
rect 143993 995419 144059 995422
rect 136449 995346 136515 995349
rect 148317 995346 148383 995349
rect 136449 995344 148383 995346
rect 136449 995288 136454 995344
rect 136510 995288 148322 995344
rect 148378 995288 148383 995344
rect 136449 995286 148383 995288
rect 136449 995283 136515 995286
rect 148317 995283 148383 995286
rect 132125 995210 132191 995213
rect 151261 995210 151327 995213
rect 132125 995208 151327 995210
rect 132125 995152 132130 995208
rect 132186 995152 151266 995208
rect 151322 995152 151327 995208
rect 132125 995150 151327 995152
rect 132125 995147 132191 995150
rect 151261 995147 151327 995150
rect 80145 995074 80211 995077
rect 92697 995074 92763 995077
rect 80145 995072 92763 995074
rect 80145 995016 80150 995072
rect 80206 995016 92702 995072
rect 92758 995016 92763 995072
rect 80145 995014 92763 995016
rect 80145 995011 80211 995014
rect 92697 995011 92763 995014
rect 128445 995074 128511 995077
rect 155542 995074 155602 996132
rect 187558 996102 190470 996162
rect 184933 995754 184999 995757
rect 187558 995754 187618 996102
rect 195421 996026 195487 996029
rect 189582 996024 195487 996026
rect 189582 995968 195426 996024
rect 195482 995968 195487 996024
rect 189582 995966 195487 995968
rect 189582 995890 189642 995966
rect 195421 995963 195487 995966
rect 195237 995890 195303 995893
rect 189214 995830 189642 995890
rect 189766 995888 195303 995890
rect 189766 995832 195242 995888
rect 195298 995832 195303 995888
rect 189766 995830 195303 995832
rect 184933 995752 187618 995754
rect 184933 995696 184938 995752
rect 184994 995696 187618 995752
rect 184933 995694 187618 995696
rect 188797 995754 188863 995757
rect 189214 995754 189274 995830
rect 188797 995752 189274 995754
rect 188797 995696 188802 995752
rect 188858 995696 189274 995752
rect 188797 995694 189274 995696
rect 189441 995754 189507 995757
rect 189766 995754 189826 995830
rect 195237 995827 195303 995830
rect 195053 995754 195119 995757
rect 189441 995752 189826 995754
rect 189441 995696 189446 995752
rect 189502 995696 189826 995752
rect 189441 995694 189826 995696
rect 190410 995752 195119 995754
rect 190410 995696 195058 995752
rect 195114 995696 195119 995752
rect 190410 995694 195119 995696
rect 184933 995691 184999 995694
rect 188797 995691 188863 995694
rect 189441 995691 189507 995694
rect 188153 995618 188219 995621
rect 190410 995618 190470 995694
rect 195053 995691 195119 995694
rect 188153 995616 190470 995618
rect 188153 995560 188158 995616
rect 188214 995560 190470 995616
rect 188153 995558 190470 995560
rect 194317 995618 194383 995621
rect 203517 995618 203583 995621
rect 194317 995616 203583 995618
rect 194317 995560 194322 995616
rect 194378 995560 203522 995616
rect 203578 995560 203583 995616
rect 194317 995558 203583 995560
rect 188153 995555 188219 995558
rect 194317 995555 194383 995558
rect 203517 995555 203583 995558
rect 183829 995482 183895 995485
rect 195973 995482 196039 995485
rect 183829 995480 196039 995482
rect 183829 995424 183834 995480
rect 183890 995424 195978 995480
rect 196034 995424 196039 995480
rect 183829 995422 196039 995424
rect 183829 995419 183895 995422
rect 195973 995419 196039 995422
rect 179827 995346 179893 995349
rect 202045 995346 202111 995349
rect 179827 995344 202111 995346
rect 179827 995288 179832 995344
rect 179888 995288 202050 995344
rect 202106 995288 202111 995344
rect 179827 995286 202111 995288
rect 179827 995283 179893 995286
rect 202045 995283 202111 995286
rect 182955 995210 183021 995213
rect 206510 995210 206570 996132
rect 243862 995757 243922 996374
rect 249701 996371 249767 996374
rect 293542 996432 303311 996434
rect 293542 996376 303250 996432
rect 303306 996376 303311 996432
rect 293542 996374 303311 996376
rect 247033 996298 247099 996301
rect 238569 995756 238635 995757
rect 238518 995692 238524 995756
rect 238588 995754 238635 995756
rect 240225 995754 240291 995757
rect 240358 995754 240364 995756
rect 238588 995752 238680 995754
rect 238630 995696 238680 995752
rect 238588 995694 238680 995696
rect 240225 995752 240364 995754
rect 240225 995696 240230 995752
rect 240286 995696 240364 995752
rect 240225 995694 240364 995696
rect 238588 995692 238635 995694
rect 238569 995691 238635 995692
rect 240225 995691 240291 995694
rect 240358 995692 240364 995694
rect 240428 995692 240434 995756
rect 243813 995752 243922 995757
rect 243813 995696 243818 995752
rect 243874 995696 243922 995752
rect 243813 995694 243922 995696
rect 244230 996296 247099 996298
rect 244230 996240 247038 996296
rect 247094 996240 247099 996296
rect 244230 996238 247099 996240
rect 243813 995691 243879 995694
rect 236545 995618 236611 995621
rect 244230 995618 244290 996238
rect 247033 996235 247099 996238
rect 236545 995616 244290 995618
rect 236545 995560 236550 995616
rect 236606 995560 244290 995616
rect 236545 995558 244290 995560
rect 236545 995555 236611 995558
rect 182955 995208 206570 995210
rect 182955 995152 182960 995208
rect 183016 995152 206570 995208
rect 182955 995150 206570 995152
rect 234383 995210 234449 995213
rect 257938 995210 257998 996132
rect 293542 995757 293602 996374
rect 303245 996371 303311 996374
rect 372337 996434 372403 996437
rect 472709 996434 472775 996437
rect 516685 996434 516751 996437
rect 372337 996432 388178 996434
rect 372337 996376 372342 996432
rect 372398 996376 388178 996432
rect 372337 996374 388178 996376
rect 372337 996371 372403 996374
rect 388118 995757 388178 996374
rect 472709 996432 482018 996434
rect 472709 996376 472714 996432
rect 472770 996376 482018 996432
rect 472709 996374 482018 996376
rect 472709 996371 472775 996374
rect 462957 996298 463023 996301
rect 462957 996296 470610 996298
rect 462957 996240 462962 996296
rect 463018 996240 470610 996296
rect 462957 996238 470610 996240
rect 462957 996235 463023 996238
rect 432045 995890 432111 995893
rect 402930 995888 432111 995890
rect 402930 995832 432050 995888
rect 432106 995832 432111 995888
rect 402930 995830 432111 995832
rect 293493 995752 293602 995757
rect 293493 995696 293498 995752
rect 293554 995696 293602 995752
rect 293493 995694 293602 995696
rect 381537 995754 381603 995757
rect 387885 995754 387951 995757
rect 381537 995752 387951 995754
rect 381537 995696 381542 995752
rect 381598 995696 387890 995752
rect 387946 995696 387951 995752
rect 381537 995694 387951 995696
rect 388118 995752 388227 995757
rect 388118 995696 388166 995752
rect 388222 995696 388227 995752
rect 388118 995694 388227 995696
rect 293493 995691 293559 995694
rect 381537 995691 381603 995694
rect 387885 995691 387951 995694
rect 388161 995691 388227 995694
rect 396625 995754 396691 995757
rect 402930 995754 402990 995830
rect 432045 995827 432111 995830
rect 439773 995756 439839 995757
rect 439773 995754 439820 995756
rect 396625 995752 402990 995754
rect 396625 995696 396630 995752
rect 396686 995696 402990 995752
rect 396625 995694 402990 995696
rect 439728 995752 439820 995754
rect 439728 995696 439778 995752
rect 439728 995694 439820 995696
rect 396625 995691 396691 995694
rect 439773 995692 439820 995694
rect 439884 995692 439890 995756
rect 439773 995691 439839 995692
rect 291745 995618 291811 995621
rect 298553 995618 298619 995621
rect 291745 995616 298619 995618
rect 291745 995560 291750 995616
rect 291806 995560 298558 995616
rect 298614 995560 298619 995616
rect 291745 995558 298619 995560
rect 291745 995555 291811 995558
rect 298553 995555 298619 995558
rect 374637 995618 374703 995621
rect 394877 995618 394943 995621
rect 374637 995616 394943 995618
rect 374637 995560 374642 995616
rect 374698 995560 394882 995616
rect 394938 995560 394943 995616
rect 374637 995558 394943 995560
rect 470550 995618 470610 996238
rect 481958 995757 482018 996374
rect 516685 996432 526178 996434
rect 516685 996376 516690 996432
rect 516746 996376 526178 996432
rect 516685 996374 526178 996376
rect 516685 996371 516751 996374
rect 526118 995757 526178 996374
rect 527958 995757 528018 996510
rect 590561 996568 630260 996570
rect 590561 996512 590566 996568
rect 590622 996512 630260 996568
rect 590561 996510 630260 996512
rect 590561 996507 590627 996510
rect 630254 996508 630260 996510
rect 630324 996508 630330 996572
rect 590561 996434 590627 996437
rect 590561 996432 627746 996434
rect 590561 996376 590566 996432
rect 590622 996376 627746 996432
rect 590561 996374 627746 996376
rect 590561 996371 590627 996374
rect 627686 996298 627746 996374
rect 628054 996374 630138 996434
rect 628054 996298 628114 996374
rect 627686 996238 628114 996298
rect 630078 996298 630138 996374
rect 630446 996374 631610 996434
rect 630446 996298 630506 996374
rect 630078 996238 630506 996298
rect 622393 996162 622459 996165
rect 622393 996160 625170 996162
rect 622393 996104 622398 996160
rect 622454 996104 625170 996160
rect 622393 996102 625170 996104
rect 622393 996099 622459 996102
rect 554630 995828 554636 995892
rect 554700 995890 554706 995892
rect 557533 995890 557599 995893
rect 554700 995888 557599 995890
rect 554700 995832 557538 995888
rect 557594 995832 557599 995888
rect 554700 995830 557599 995832
rect 554700 995828 554706 995830
rect 557533 995827 557599 995830
rect 480662 995692 480668 995756
rect 480732 995754 480738 995756
rect 480805 995754 480871 995757
rect 480732 995752 480871 995754
rect 480732 995696 480810 995752
rect 480866 995696 480871 995752
rect 480732 995694 480871 995696
rect 481958 995752 482067 995757
rect 485589 995756 485655 995757
rect 485589 995754 485636 995756
rect 481958 995696 482006 995752
rect 482062 995696 482067 995752
rect 481958 995694 482067 995696
rect 485544 995752 485636 995754
rect 485544 995696 485594 995752
rect 485544 995694 485636 995696
rect 480732 995692 480738 995694
rect 480805 995691 480871 995694
rect 482001 995691 482067 995694
rect 485589 995692 485636 995694
rect 485700 995692 485706 995756
rect 526118 995752 526227 995757
rect 526118 995696 526166 995752
rect 526222 995696 526227 995752
rect 526118 995694 526227 995696
rect 527958 995752 528067 995757
rect 527958 995696 528006 995752
rect 528062 995696 528067 995752
rect 527958 995694 528067 995696
rect 485589 995691 485655 995692
rect 526161 995691 526227 995694
rect 528001 995691 528067 995694
rect 531998 995692 532004 995756
rect 532068 995754 532074 995756
rect 532141 995754 532207 995757
rect 536557 995756 536623 995757
rect 536557 995754 536604 995756
rect 532068 995752 532207 995754
rect 532068 995696 532146 995752
rect 532202 995696 532207 995752
rect 532068 995694 532207 995696
rect 536512 995752 536604 995754
rect 536512 995696 536562 995752
rect 536512 995694 536604 995696
rect 532068 995692 532074 995694
rect 532141 995691 532207 995694
rect 536557 995692 536604 995694
rect 536668 995692 536674 995756
rect 568205 995754 568271 995757
rect 573214 995754 573220 995756
rect 568205 995752 573220 995754
rect 568205 995696 568210 995752
rect 568266 995696 573220 995752
rect 568205 995694 573220 995696
rect 536557 995691 536623 995692
rect 568205 995691 568271 995694
rect 573214 995692 573220 995694
rect 573284 995692 573290 995756
rect 482645 995618 482711 995621
rect 470550 995616 482711 995618
rect 470550 995560 482650 995616
rect 482706 995560 482711 995616
rect 470550 995558 482711 995560
rect 374637 995555 374703 995558
rect 394877 995555 394943 995558
rect 482645 995555 482711 995558
rect 516869 995618 516935 995621
rect 529841 995618 529907 995621
rect 516869 995616 529907 995618
rect 516869 995560 516874 995616
rect 516930 995560 529846 995616
rect 529902 995560 529907 995616
rect 516869 995558 529907 995560
rect 625110 995618 625170 996102
rect 631550 995757 631610 996374
rect 627913 995756 627979 995757
rect 630305 995756 630371 995757
rect 627862 995692 627868 995756
rect 627932 995754 627979 995756
rect 627932 995752 628024 995754
rect 627974 995696 628024 995752
rect 627932 995694 628024 995696
rect 627932 995692 627979 995694
rect 630254 995692 630260 995756
rect 630324 995754 630371 995756
rect 630324 995752 630416 995754
rect 630366 995696 630416 995752
rect 630324 995694 630416 995696
rect 631550 995752 631659 995757
rect 631550 995696 631598 995752
rect 631654 995696 631659 995752
rect 631550 995694 631659 995696
rect 630324 995692 630371 995694
rect 627913 995691 627979 995692
rect 630305 995691 630371 995692
rect 631593 995691 631659 995694
rect 635181 995618 635247 995621
rect 625110 995616 635247 995618
rect 625110 995560 635186 995616
rect 635242 995560 635247 995616
rect 625110 995558 635247 995560
rect 516869 995555 516935 995558
rect 529841 995555 529907 995558
rect 635181 995555 635247 995558
rect 380893 995482 380959 995485
rect 389357 995482 389423 995485
rect 380893 995480 389423 995482
rect 380893 995424 380898 995480
rect 380954 995424 389362 995480
rect 389418 995424 389423 995480
rect 380893 995422 389423 995424
rect 380893 995419 380959 995422
rect 389357 995419 389423 995422
rect 456057 995482 456123 995485
rect 476389 995482 476455 995485
rect 456057 995480 476455 995482
rect 456057 995424 456062 995480
rect 456118 995424 476394 995480
rect 476450 995424 476455 995480
rect 456057 995422 476455 995424
rect 456057 995419 456123 995422
rect 476389 995419 476455 995422
rect 519261 995482 519327 995485
rect 538949 995482 539015 995485
rect 519261 995480 539015 995482
rect 519261 995424 519266 995480
rect 519322 995424 538954 995480
rect 539010 995424 539015 995480
rect 519261 995422 539015 995424
rect 519261 995419 519327 995422
rect 538949 995419 539015 995422
rect 376017 995346 376083 995349
rect 385309 995346 385375 995349
rect 376017 995344 385375 995346
rect 376017 995288 376022 995344
rect 376078 995288 385314 995344
rect 385370 995288 385375 995344
rect 376017 995286 385375 995288
rect 376017 995283 376083 995286
rect 385309 995283 385375 995286
rect 459645 995346 459711 995349
rect 484117 995346 484183 995349
rect 459645 995344 484183 995346
rect 459645 995288 459650 995344
rect 459706 995288 484122 995344
rect 484178 995288 484183 995344
rect 459645 995286 484183 995288
rect 459645 995283 459711 995286
rect 484117 995283 484183 995286
rect 522389 995346 522455 995349
rect 534349 995346 534415 995349
rect 522389 995344 534415 995346
rect 522389 995288 522394 995344
rect 522450 995288 534354 995344
rect 534410 995288 534415 995344
rect 522389 995286 534415 995288
rect 522389 995283 522455 995286
rect 534349 995283 534415 995286
rect 234383 995208 257998 995210
rect 234383 995152 234388 995208
rect 234444 995152 257998 995208
rect 234383 995150 257998 995152
rect 380157 995210 380223 995213
rect 393957 995210 394023 995213
rect 380157 995208 394023 995210
rect 380157 995152 380162 995208
rect 380218 995152 393962 995208
rect 394018 995152 394023 995208
rect 380157 995150 394023 995152
rect 182955 995147 183021 995150
rect 234383 995147 234449 995150
rect 380157 995147 380223 995150
rect 393957 995147 394023 995150
rect 454309 995210 454375 995213
rect 481633 995210 481699 995213
rect 454309 995208 481699 995210
rect 454309 995152 454314 995208
rect 454370 995152 481638 995208
rect 481694 995152 481699 995208
rect 454309 995150 481699 995152
rect 454309 995147 454375 995150
rect 481633 995147 481699 995150
rect 516961 995210 517027 995213
rect 533061 995210 533127 995213
rect 516961 995208 533127 995210
rect 516961 995152 516966 995208
rect 517022 995152 533066 995208
rect 533122 995152 533127 995208
rect 516961 995150 533127 995152
rect 516961 995147 517027 995150
rect 533061 995147 533127 995150
rect 618161 995210 618227 995213
rect 626855 995210 626921 995213
rect 618161 995208 626921 995210
rect 618161 995152 618166 995208
rect 618222 995152 626860 995208
rect 626916 995152 626921 995208
rect 618161 995150 626921 995152
rect 618161 995147 618227 995150
rect 626855 995147 626921 995150
rect 128445 995072 155602 995074
rect 128445 995016 128450 995072
rect 128506 995016 155602 995072
rect 128445 995014 155602 995016
rect 191741 995074 191807 995077
rect 215293 995074 215359 995077
rect 191741 995072 215359 995074
rect 191741 995016 191746 995072
rect 191802 995016 215298 995072
rect 215354 995016 215359 995072
rect 191741 995014 215359 995016
rect 128445 995011 128511 995014
rect 191741 995011 191807 995014
rect 215293 995011 215359 995014
rect 232865 995074 232931 995077
rect 257337 995074 257403 995077
rect 232865 995072 257403 995074
rect 232865 995016 232870 995072
rect 232926 995016 257342 995072
rect 257398 995016 257403 995072
rect 232865 995014 257403 995016
rect 232865 995011 232931 995014
rect 257337 995011 257403 995014
rect 285949 995074 286015 995077
rect 307017 995074 307083 995077
rect 285949 995072 307083 995074
rect 285949 995016 285954 995072
rect 286010 995016 307022 995072
rect 307078 995016 307083 995072
rect 285949 995014 307083 995016
rect 285949 995011 286015 995014
rect 307017 995011 307083 995014
rect 449801 995074 449867 995077
rect 485957 995074 486023 995077
rect 449801 995072 486023 995074
rect 449801 995016 449806 995072
rect 449862 995016 485962 995072
rect 486018 995016 486023 995072
rect 449801 995014 486023 995016
rect 449801 995011 449867 995014
rect 485957 995011 486023 995014
rect 620277 995074 620343 995077
rect 629661 995074 629727 995077
rect 620277 995072 629727 995074
rect 620277 995016 620282 995072
rect 620338 995016 629666 995072
rect 629722 995016 629727 995072
rect 620277 995014 629727 995016
rect 620277 995011 620343 995014
rect 629661 995011 629727 995014
rect 505134 992292 505140 992356
rect 505204 992354 505210 992356
rect 511073 992354 511139 992357
rect 505204 992352 511139 992354
rect 505204 992296 511078 992352
rect 511134 992296 511139 992352
rect 505204 992294 511139 992296
rect 505204 992292 505210 992294
rect 511073 992291 511139 992294
rect 439814 991476 439820 991540
rect 439884 991538 439890 991540
rect 446489 991538 446555 991541
rect 439884 991536 446555 991538
rect 439884 991480 446494 991536
rect 446550 991480 446555 991536
rect 439884 991478 446555 991480
rect 439884 991476 439890 991478
rect 446489 991475 446555 991478
rect 573214 990932 573220 990996
rect 573284 990994 573290 990996
rect 576301 990994 576367 990997
rect 573284 990992 576367 990994
rect 573284 990936 576306 990992
rect 576362 990936 576367 990992
rect 573284 990934 576367 990936
rect 573284 990932 573290 990934
rect 576301 990931 576367 990934
rect 62113 976034 62179 976037
rect 62113 976032 64492 976034
rect 62113 975976 62118 976032
rect 62174 975976 64492 976032
rect 62113 975974 64492 975976
rect 62113 975971 62179 975974
rect 651649 975898 651715 975901
rect 650164 975896 651715 975898
rect 650164 975840 651654 975896
rect 651710 975840 651715 975896
rect 650164 975838 651715 975840
rect 651649 975835 651715 975838
rect 40534 968764 40540 968828
rect 40604 968826 40610 968828
rect 41781 968826 41847 968829
rect 40604 968824 41847 968826
rect 40604 968768 41786 968824
rect 41842 968768 41847 968824
rect 40604 968766 41847 968768
rect 40604 968764 40610 968766
rect 41781 968763 41847 968766
rect 40718 967268 40724 967332
rect 40788 967330 40794 967332
rect 41781 967330 41847 967333
rect 40788 967328 41847 967330
rect 40788 967272 41786 967328
rect 41842 967272 41847 967328
rect 40788 967270 41847 967272
rect 40788 967268 40794 967270
rect 41781 967267 41847 967270
rect 675753 966514 675819 966517
rect 676806 966514 676812 966516
rect 675753 966512 676812 966514
rect 675753 966456 675758 966512
rect 675814 966456 676812 966512
rect 675753 966454 676812 966456
rect 675753 966451 675819 966454
rect 676806 966452 676812 966454
rect 676876 966452 676882 966516
rect 675753 966242 675819 966245
rect 676438 966242 676444 966244
rect 675753 966240 676444 966242
rect 675753 966184 675758 966240
rect 675814 966184 676444 966240
rect 675753 966182 676444 966184
rect 675753 966179 675819 966182
rect 676438 966180 676444 966182
rect 676508 966180 676514 966244
rect 42057 965156 42123 965157
rect 42006 965154 42012 965156
rect 41966 965094 42012 965154
rect 42076 965152 42123 965156
rect 42118 965096 42123 965152
rect 42006 965092 42012 965094
rect 42076 965092 42123 965096
rect 42057 965091 42123 965092
rect 675753 965018 675819 965021
rect 677174 965018 677180 965020
rect 675753 965016 677180 965018
rect 675753 964960 675758 965016
rect 675814 964960 677180 965016
rect 675753 964958 677180 964960
rect 675753 964955 675819 964958
rect 677174 964956 677180 964958
rect 677244 964956 677250 965020
rect 40350 963324 40356 963388
rect 40420 963386 40426 963388
rect 41781 963386 41847 963389
rect 675385 963388 675451 963389
rect 675334 963386 675340 963388
rect 40420 963384 41847 963386
rect 40420 963328 41786 963384
rect 41842 963328 41847 963384
rect 40420 963326 41847 963328
rect 675294 963326 675340 963386
rect 675404 963384 675451 963388
rect 675446 963328 675451 963384
rect 40420 963324 40426 963326
rect 41781 963323 41847 963326
rect 675334 963324 675340 963326
rect 675404 963324 675451 963328
rect 675385 963323 675451 963324
rect 62113 962978 62179 962981
rect 62113 962976 64492 962978
rect 62113 962920 62118 962976
rect 62174 962920 64492 962976
rect 62113 962918 64492 962920
rect 62113 962915 62179 962918
rect 652017 962570 652083 962573
rect 650164 962568 652083 962570
rect 650164 962512 652022 962568
rect 652078 962512 652083 962568
rect 650164 962510 652083 962512
rect 652017 962507 652083 962510
rect 41454 962100 41460 962164
rect 41524 962162 41530 962164
rect 41781 962162 41847 962165
rect 41524 962160 41847 962162
rect 41524 962104 41786 962160
rect 41842 962104 41847 962160
rect 41524 962102 41847 962104
rect 41524 962100 41530 962102
rect 41781 962099 41847 962102
rect 675753 961346 675819 961349
rect 675886 961346 675892 961348
rect 675753 961344 675892 961346
rect 675753 961288 675758 961344
rect 675814 961288 675892 961344
rect 675753 961286 675892 961288
rect 675753 961283 675819 961286
rect 675886 961284 675892 961286
rect 675956 961284 675962 961348
rect 675661 959172 675727 959173
rect 675661 959168 675708 959172
rect 675772 959170 675778 959172
rect 675661 959112 675666 959168
rect 675661 959108 675708 959112
rect 675772 959110 675818 959170
rect 675772 959108 675778 959110
rect 675661 959107 675727 959108
rect 674741 959034 674807 959037
rect 676990 959034 676996 959036
rect 674741 959032 676996 959034
rect 674741 958976 674746 959032
rect 674802 958976 676996 959032
rect 674741 958974 676996 958976
rect 674741 958971 674807 958974
rect 676990 958972 676996 958974
rect 677060 958972 677066 959036
rect 41638 958292 41644 958356
rect 41708 958354 41714 958356
rect 41781 958354 41847 958357
rect 41708 958352 41847 958354
rect 41708 958296 41786 958352
rect 41842 958296 41847 958352
rect 41708 958294 41847 958296
rect 41708 958292 41714 958294
rect 41781 958291 41847 958294
rect 42057 957810 42123 957813
rect 675477 957812 675543 957813
rect 42190 957810 42196 957812
rect 42057 957808 42196 957810
rect 42057 957752 42062 957808
rect 42118 957752 42196 957808
rect 42057 957750 42196 957752
rect 42057 957747 42123 957750
rect 42190 957748 42196 957750
rect 42260 957748 42266 957812
rect 675477 957808 675524 957812
rect 675588 957810 675594 957812
rect 675477 957752 675482 957808
rect 675477 957748 675524 957752
rect 675588 957750 675634 957810
rect 675588 957748 675594 957750
rect 675477 957747 675543 957748
rect 675017 957674 675083 957677
rect 676622 957674 676628 957676
rect 675017 957672 676628 957674
rect 675017 957616 675022 957672
rect 675078 957616 676628 957672
rect 675017 957614 676628 957616
rect 675017 957611 675083 957614
rect 676622 957612 676628 957614
rect 676692 957612 676698 957676
rect 675753 954002 675819 954005
rect 676070 954002 676076 954004
rect 675753 954000 676076 954002
rect 675753 953944 675758 954000
rect 675814 953944 676076 954000
rect 675753 953942 676076 953944
rect 675753 953939 675819 953942
rect 676070 953940 676076 953942
rect 676140 953940 676146 954004
rect 37917 952234 37983 952237
rect 41638 952234 41644 952236
rect 37917 952232 41644 952234
rect 37917 952176 37922 952232
rect 37978 952176 41644 952232
rect 37917 952174 41644 952176
rect 37917 952171 37983 952174
rect 41638 952172 41644 952174
rect 41708 952172 41714 952236
rect 41965 951826 42031 951829
rect 42190 951826 42196 951828
rect 41965 951824 42196 951826
rect 41965 951768 41970 951824
rect 42026 951768 42196 951824
rect 41965 951766 42196 951768
rect 41965 951763 42031 951766
rect 42190 951764 42196 951766
rect 42260 951764 42266 951828
rect 32397 951690 32463 951693
rect 41454 951690 41460 951692
rect 32397 951688 41460 951690
rect 32397 951632 32402 951688
rect 32458 951632 41460 951688
rect 32397 951630 41460 951632
rect 32397 951627 32463 951630
rect 41454 951628 41460 951630
rect 41524 951628 41530 951692
rect 41781 951690 41847 951693
rect 42006 951690 42012 951692
rect 41781 951688 42012 951690
rect 41781 951632 41786 951688
rect 41842 951632 42012 951688
rect 41781 951630 42012 951632
rect 41781 951627 41847 951630
rect 42006 951628 42012 951630
rect 42076 951628 42082 951692
rect 676438 950948 676444 951012
rect 676508 951010 676514 951012
rect 677501 951010 677567 951013
rect 676508 951008 677567 951010
rect 676508 950952 677506 951008
rect 677562 950952 677567 951008
rect 676508 950950 677567 950952
rect 676508 950948 676514 950950
rect 677501 950947 677567 950950
rect 676806 950812 676812 950876
rect 676876 950874 676882 950876
rect 677409 950874 677475 950877
rect 676876 950872 677475 950874
rect 676876 950816 677414 950872
rect 677470 950816 677475 950872
rect 676876 950814 677475 950816
rect 676876 950812 676882 950814
rect 677409 950811 677475 950814
rect 62113 949922 62179 949925
rect 62113 949920 64492 949922
rect 62113 949864 62118 949920
rect 62174 949864 64492 949920
rect 62113 949862 64492 949864
rect 62113 949859 62179 949862
rect 675334 949724 675340 949788
rect 675404 949786 675410 949788
rect 680997 949786 681063 949789
rect 675404 949784 681063 949786
rect 675404 949728 681002 949784
rect 681058 949728 681063 949784
rect 675404 949726 681063 949728
rect 675404 949724 675410 949726
rect 680997 949723 681063 949726
rect 675518 949588 675524 949652
rect 675588 949650 675594 949652
rect 679801 949650 679867 949653
rect 675588 949648 679867 949650
rect 675588 949592 679806 949648
rect 679862 949592 679867 949648
rect 675588 949590 679867 949592
rect 675588 949588 675594 949590
rect 679801 949587 679867 949590
rect 675886 949452 675892 949516
rect 675956 949514 675962 949516
rect 679617 949514 679683 949517
rect 675956 949512 679683 949514
rect 675956 949456 679622 949512
rect 679678 949456 679683 949512
rect 675956 949454 679683 949456
rect 675956 949452 675962 949454
rect 679617 949451 679683 949454
rect 651557 949378 651623 949381
rect 650164 949376 651623 949378
rect 650164 949320 651562 949376
rect 651618 949320 651623 949376
rect 650164 949318 651623 949320
rect 651557 949315 651623 949318
rect 675702 948772 675708 948836
rect 675772 948834 675778 948836
rect 681089 948834 681155 948837
rect 675772 948832 681155 948834
rect 675772 948776 681094 948832
rect 681150 948776 681155 948832
rect 675772 948774 681155 948776
rect 675772 948772 675778 948774
rect 681089 948771 681155 948774
rect 676070 947956 676076 948020
rect 676140 948018 676146 948020
rect 682377 948018 682443 948021
rect 676140 948016 682443 948018
rect 676140 947960 682382 948016
rect 682438 947960 682443 948016
rect 676140 947958 682443 947960
rect 676140 947956 676146 947958
rect 682377 947955 682443 947958
rect 34513 943802 34579 943805
rect 34470 943800 34579 943802
rect 34470 943744 34518 943800
rect 34574 943744 34579 943800
rect 34470 943739 34579 943744
rect 34470 943500 34530 943739
rect 35801 943122 35867 943125
rect 35788 943120 35867 943122
rect 35788 943064 35806 943120
rect 35862 943064 35867 943120
rect 35788 943062 35867 943064
rect 35801 943059 35867 943062
rect 35709 942714 35775 942717
rect 35709 942712 35788 942714
rect 35709 942656 35714 942712
rect 35770 942656 35788 942712
rect 35709 942654 35788 942656
rect 35709 942651 35775 942654
rect 48957 942306 49023 942309
rect 41492 942304 49023 942306
rect 41492 942248 48962 942304
rect 49018 942248 49023 942304
rect 41492 942246 49023 942248
rect 48957 942243 49023 942246
rect 41873 941898 41939 941901
rect 41492 941896 41939 941898
rect 41492 941840 41878 941896
rect 41934 941840 41939 941896
rect 41492 941838 41939 941840
rect 41873 941835 41939 941838
rect 44817 941490 44883 941493
rect 41492 941488 44883 941490
rect 41492 941432 44822 941488
rect 44878 941432 44883 941488
rect 41492 941430 44883 941432
rect 44817 941427 44883 941430
rect 41781 941082 41847 941085
rect 41492 941080 41847 941082
rect 41492 941024 41786 941080
rect 41842 941024 41847 941080
rect 41492 941022 41847 941024
rect 41781 941019 41847 941022
rect 47577 940674 47643 940677
rect 41492 940672 47643 940674
rect 41492 940616 47582 940672
rect 47638 940616 47643 940672
rect 41492 940614 47643 940616
rect 47577 940611 47643 940614
rect 41492 940206 41752 940266
rect 41692 940133 41752 940206
rect 41689 940128 41755 940133
rect 41689 940072 41694 940128
rect 41750 940072 41755 940128
rect 41689 940067 41755 940072
rect 676029 939994 676095 939997
rect 676029 939992 676292 939994
rect 676029 939936 676034 939992
rect 676090 939936 676292 939992
rect 676029 939934 676292 939936
rect 676029 939931 676095 939934
rect 50337 939858 50403 939861
rect 41492 939856 50403 939858
rect 41492 939800 50342 939856
rect 50398 939800 50403 939856
rect 41492 939798 50403 939800
rect 50337 939795 50403 939798
rect 41492 939390 41752 939450
rect 41692 939317 41752 939390
rect 676262 939317 676322 939556
rect 41689 939312 41755 939317
rect 41689 939256 41694 939312
rect 41750 939256 41755 939312
rect 41689 939251 41755 939256
rect 676213 939312 676322 939317
rect 676213 939256 676218 939312
rect 676274 939256 676322 939312
rect 676213 939254 676322 939256
rect 676213 939251 676279 939254
rect 676029 939178 676095 939181
rect 676029 939176 676292 939178
rect 676029 939120 676034 939176
rect 676090 939120 676292 939176
rect 676029 939118 676292 939120
rect 676029 939115 676095 939118
rect 42149 939042 42215 939045
rect 41492 939040 42215 939042
rect 41492 938984 42154 939040
rect 42210 938984 42215 939040
rect 41492 938982 42215 938984
rect 42149 938979 42215 938982
rect 676029 938770 676095 938773
rect 676029 938768 676292 938770
rect 676029 938712 676034 938768
rect 676090 938712 676292 938768
rect 676029 938710 676292 938712
rect 676029 938707 676095 938710
rect 41822 938634 41828 938636
rect 41492 938574 41828 938634
rect 41822 938572 41828 938574
rect 41892 938572 41898 938636
rect 31017 938226 31083 938229
rect 31004 938224 31083 938226
rect 31004 938168 31022 938224
rect 31078 938168 31083 938224
rect 31004 938166 31083 938168
rect 31017 938163 31083 938166
rect 676121 938090 676187 938093
rect 676262 938090 676322 938332
rect 676121 938088 676322 938090
rect 676121 938032 676126 938088
rect 676182 938032 676322 938088
rect 676121 938030 676322 938032
rect 676121 938027 676187 938030
rect 41965 937818 42031 937821
rect 41492 937816 42031 937818
rect 41492 937760 41970 937816
rect 42026 937760 42031 937816
rect 41492 937758 42031 937760
rect 41965 937755 42031 937758
rect 676262 937685 676322 937924
rect 676213 937680 676322 937685
rect 676213 937624 676218 937680
rect 676274 937624 676322 937680
rect 676213 937622 676322 937624
rect 676213 937619 676279 937622
rect 676029 937546 676095 937549
rect 676029 937544 676292 937546
rect 676029 937488 676034 937544
rect 676090 937488 676292 937544
rect 676029 937486 676292 937488
rect 676029 937483 676095 937486
rect 32397 937410 32463 937413
rect 32397 937408 32476 937410
rect 32397 937352 32402 937408
rect 32458 937352 32476 937408
rect 32397 937350 32476 937352
rect 32397 937347 32463 937350
rect 676213 937274 676279 937277
rect 676213 937272 676322 937274
rect 676213 937216 676218 937272
rect 676274 937216 676322 937272
rect 676213 937211 676322 937216
rect 676262 937108 676322 937211
rect 41822 937002 41828 937004
rect 41492 936942 41828 937002
rect 41822 936940 41828 936942
rect 41892 936940 41898 937004
rect 62113 937002 62179 937005
rect 62113 937000 64492 937002
rect 62113 936944 62118 937000
rect 62174 936944 64492 937000
rect 62113 936942 64492 936944
rect 62113 936939 62179 936942
rect 676029 936730 676095 936733
rect 676029 936728 676292 936730
rect 676029 936672 676034 936728
rect 676090 936672 676292 936728
rect 676029 936670 676292 936672
rect 676029 936667 676095 936670
rect 36537 936594 36603 936597
rect 36524 936592 36603 936594
rect 36524 936536 36542 936592
rect 36598 936536 36603 936592
rect 36524 936534 36603 936536
rect 36537 936531 36603 936534
rect 37917 936186 37983 936189
rect 651557 936186 651623 936189
rect 37917 936184 37996 936186
rect 37917 936128 37922 936184
rect 37978 936128 37996 936184
rect 37917 936126 37996 936128
rect 650164 936184 651623 936186
rect 650164 936128 651562 936184
rect 651618 936128 651623 936184
rect 650164 936126 651623 936128
rect 37917 936123 37983 936126
rect 651557 936123 651623 936126
rect 676262 936053 676322 936292
rect 676213 936048 676322 936053
rect 676213 935992 676218 936048
rect 676274 935992 676322 936048
rect 676213 935990 676322 935992
rect 676213 935987 676279 935990
rect 676029 935914 676095 935917
rect 676029 935912 676292 935914
rect 676029 935856 676034 935912
rect 676090 935856 676292 935912
rect 676029 935854 676292 935856
rect 676029 935851 676095 935854
rect 42977 935778 43043 935781
rect 41492 935776 43043 935778
rect 41492 935720 42982 935776
rect 43038 935720 43043 935776
rect 41492 935718 43043 935720
rect 42977 935715 43043 935718
rect 677174 935580 677180 935644
rect 677244 935580 677250 935644
rect 677182 935476 677242 935580
rect 42057 935370 42123 935373
rect 41492 935368 42123 935370
rect 41492 935312 42062 935368
rect 42118 935312 42123 935368
rect 41492 935310 42123 935312
rect 42057 935307 42123 935310
rect 682377 935234 682443 935237
rect 682334 935232 682443 935234
rect 682334 935176 682382 935232
rect 682438 935176 682443 935232
rect 682334 935171 682443 935176
rect 682334 935068 682394 935171
rect 41822 934962 41828 934964
rect 41492 934902 41828 934962
rect 41822 934900 41828 934902
rect 41892 934900 41898 934964
rect 677409 934826 677475 934829
rect 677366 934824 677475 934826
rect 677366 934768 677414 934824
rect 677470 934768 677475 934824
rect 677366 934763 677475 934768
rect 677366 934660 677426 934763
rect 44173 934554 44239 934557
rect 41492 934552 44239 934554
rect 41492 934496 44178 934552
rect 44234 934496 44239 934552
rect 41492 934494 44239 934496
rect 44173 934491 44239 934494
rect 680997 934418 681063 934421
rect 680997 934416 681106 934418
rect 680997 934360 681002 934416
rect 681058 934360 681106 934416
rect 680997 934355 681106 934360
rect 681046 934252 681106 934355
rect 42885 934146 42951 934149
rect 41492 934144 42951 934146
rect 41492 934088 42890 934144
rect 42946 934088 42951 934144
rect 41492 934086 42951 934088
rect 42885 934083 42951 934086
rect 681089 934010 681155 934013
rect 681046 934008 681155 934010
rect 681046 933952 681094 934008
rect 681150 933952 681155 934008
rect 681046 933947 681155 933952
rect 681046 933844 681106 933947
rect 42793 933738 42859 933741
rect 41492 933736 42859 933738
rect 41492 933680 42798 933736
rect 42854 933680 42859 933736
rect 41492 933678 42859 933680
rect 42793 933675 42859 933678
rect 678237 933602 678303 933605
rect 678237 933600 678346 933602
rect 678237 933544 678242 933600
rect 678298 933544 678346 933600
rect 678237 933539 678346 933544
rect 678286 933436 678346 933539
rect 39941 933330 40007 933333
rect 39941 933328 40020 933330
rect 39941 933272 39946 933328
rect 40002 933272 40020 933328
rect 39941 933270 40020 933272
rect 39941 933267 40007 933270
rect 677501 933194 677567 933197
rect 677501 933192 677610 933194
rect 677501 933136 677506 933192
rect 677562 933136 677610 933192
rect 677501 933131 677610 933136
rect 677550 933028 677610 933131
rect 21774 932484 21834 932910
rect 676990 932724 676996 932788
rect 677060 932724 677066 932788
rect 676998 932620 677058 932724
rect 676622 932316 676628 932380
rect 676692 932316 676698 932380
rect 676630 932212 676690 932316
rect 41873 932106 41939 932109
rect 43437 932106 43503 932109
rect 41492 932104 43503 932106
rect 41492 932048 41878 932104
rect 41934 932048 43442 932104
rect 43498 932048 43503 932104
rect 41492 932046 43503 932048
rect 41873 932043 41939 932046
rect 43437 932043 43503 932046
rect 676213 931970 676279 931973
rect 676213 931968 676322 931970
rect 676213 931912 676218 931968
rect 676274 931912 676322 931968
rect 676213 931907 676322 931912
rect 676262 931804 676322 931907
rect 679801 931562 679867 931565
rect 679758 931560 679867 931562
rect 679758 931504 679806 931560
rect 679862 931504 679867 931560
rect 679758 931499 679867 931504
rect 679758 931396 679818 931499
rect 679617 931154 679683 931157
rect 679574 931152 679683 931154
rect 679574 931096 679622 931152
rect 679678 931096 679683 931152
rect 679574 931091 679683 931096
rect 679574 930988 679634 931091
rect 676262 930341 676322 930580
rect 676213 930336 676322 930341
rect 676213 930280 676218 930336
rect 676274 930280 676322 930336
rect 676213 930278 676322 930280
rect 676213 930275 676279 930278
rect 674741 930202 674807 930205
rect 674741 930200 676292 930202
rect 674741 930144 674746 930200
rect 674802 930144 676292 930200
rect 674741 930142 676292 930144
rect 674741 930139 674807 930142
rect 683070 929525 683130 929764
rect 683070 929520 683179 929525
rect 683070 929464 683118 929520
rect 683174 929464 683179 929520
rect 683070 929462 683179 929464
rect 683113 929459 683179 929462
rect 685830 928948 685890 929356
rect 683113 928706 683179 928709
rect 683070 928704 683179 928706
rect 683070 928648 683118 928704
rect 683174 928648 683179 928704
rect 683070 928643 683179 928648
rect 683070 928540 683130 928643
rect 62113 923810 62179 923813
rect 62113 923808 64492 923810
rect 62113 923752 62118 923808
rect 62174 923752 64492 923808
rect 62113 923750 64492 923752
rect 62113 923747 62179 923750
rect 651557 922722 651623 922725
rect 650164 922720 651623 922722
rect 650164 922664 651562 922720
rect 651618 922664 651623 922720
rect 650164 922662 651623 922664
rect 651557 922659 651623 922662
rect 62113 910754 62179 910757
rect 62113 910752 64492 910754
rect 62113 910696 62118 910752
rect 62174 910696 64492 910752
rect 62113 910694 64492 910696
rect 62113 910691 62179 910694
rect 651557 909530 651623 909533
rect 650164 909528 651623 909530
rect 650164 909472 651562 909528
rect 651618 909472 651623 909528
rect 650164 909470 651623 909472
rect 651557 909467 651623 909470
rect 62113 897834 62179 897837
rect 62113 897832 64492 897834
rect 62113 897776 62118 897832
rect 62174 897776 64492 897832
rect 62113 897774 64492 897776
rect 62113 897771 62179 897774
rect 651557 896202 651623 896205
rect 650164 896200 651623 896202
rect 650164 896144 651562 896200
rect 651618 896144 651623 896200
rect 650164 896142 651623 896144
rect 651557 896139 651623 896142
rect 62113 884778 62179 884781
rect 62113 884776 64492 884778
rect 62113 884720 62118 884776
rect 62174 884720 64492 884776
rect 62113 884718 64492 884720
rect 62113 884715 62179 884718
rect 652017 882874 652083 882877
rect 650164 882872 652083 882874
rect 650164 882816 652022 882872
rect 652078 882816 652083 882872
rect 650164 882814 652083 882816
rect 652017 882811 652083 882814
rect 675753 876618 675819 876621
rect 676622 876618 676628 876620
rect 675753 876616 676628 876618
rect 675753 876560 675758 876616
rect 675814 876560 676628 876616
rect 675753 876558 676628 876560
rect 675753 876555 675819 876558
rect 676622 876556 676628 876558
rect 676692 876556 676698 876620
rect 675293 876482 675359 876485
rect 676806 876482 676812 876484
rect 675293 876480 676812 876482
rect 675293 876424 675298 876480
rect 675354 876424 676812 876480
rect 675293 876422 676812 876424
rect 675293 876419 675359 876422
rect 676806 876420 676812 876422
rect 676876 876420 676882 876484
rect 675753 874170 675819 874173
rect 676070 874170 676076 874172
rect 675753 874168 676076 874170
rect 675753 874112 675758 874168
rect 675814 874112 676076 874168
rect 675753 874110 676076 874112
rect 675753 874107 675819 874110
rect 676070 874108 676076 874110
rect 676140 874108 676146 874172
rect 675753 872810 675819 872813
rect 677174 872810 677180 872812
rect 675753 872808 677180 872810
rect 675753 872752 675758 872808
rect 675814 872752 677180 872808
rect 675753 872750 677180 872752
rect 675753 872747 675819 872750
rect 677174 872748 677180 872750
rect 677244 872748 677250 872812
rect 673862 872204 673868 872268
rect 673932 872266 673938 872268
rect 675385 872266 675451 872269
rect 673932 872264 675451 872266
rect 673932 872208 675390 872264
rect 675446 872208 675451 872264
rect 673932 872206 675451 872208
rect 673932 872204 673938 872206
rect 675385 872203 675451 872206
rect 62113 871722 62179 871725
rect 62113 871720 64492 871722
rect 62113 871664 62118 871720
rect 62174 871664 64492 871720
rect 62113 871662 64492 871664
rect 62113 871659 62179 871662
rect 651557 869682 651623 869685
rect 650164 869680 651623 869682
rect 650164 869624 651562 869680
rect 651618 869624 651623 869680
rect 650164 869622 651623 869624
rect 651557 869619 651623 869622
rect 675753 864786 675819 864789
rect 675886 864786 675892 864788
rect 675753 864784 675892 864786
rect 675753 864728 675758 864784
rect 675814 864728 675892 864784
rect 675753 864726 675892 864728
rect 675753 864723 675819 864726
rect 675886 864724 675892 864726
rect 675956 864724 675962 864788
rect 62113 858666 62179 858669
rect 62113 858664 64492 858666
rect 62113 858608 62118 858664
rect 62174 858608 64492 858664
rect 62113 858606 64492 858608
rect 62113 858603 62179 858606
rect 652569 856354 652635 856357
rect 650164 856352 652635 856354
rect 650164 856296 652574 856352
rect 652630 856296 652635 856352
rect 650164 856294 652635 856296
rect 652569 856291 652635 856294
rect 62113 845610 62179 845613
rect 62113 845608 64492 845610
rect 62113 845552 62118 845608
rect 62174 845552 64492 845608
rect 62113 845550 64492 845552
rect 62113 845547 62179 845550
rect 651557 843026 651623 843029
rect 650164 843024 651623 843026
rect 650164 842968 651562 843024
rect 651618 842968 651623 843024
rect 650164 842966 651623 842968
rect 651557 842963 651623 842966
rect 62113 832554 62179 832557
rect 62113 832552 64492 832554
rect 62113 832496 62118 832552
rect 62174 832496 64492 832552
rect 62113 832494 64492 832496
rect 62113 832491 62179 832494
rect 651557 829834 651623 829837
rect 650164 829832 651623 829834
rect 650164 829776 651562 829832
rect 651618 829776 651623 829832
rect 650164 829774 651623 829776
rect 651557 829771 651623 829774
rect 62113 819498 62179 819501
rect 62113 819496 64492 819498
rect 62113 819440 62118 819496
rect 62174 819440 64492 819496
rect 62113 819438 64492 819440
rect 62113 819435 62179 819438
rect 41229 818002 41295 818005
rect 41229 818000 41338 818002
rect 41229 817944 41234 818000
rect 41290 817944 41338 818000
rect 41229 817939 41338 817944
rect 41278 817700 41338 817939
rect 41321 817322 41387 817325
rect 41308 817320 41387 817322
rect 41308 817264 41326 817320
rect 41382 817264 41387 817320
rect 41308 817262 41387 817264
rect 41321 817259 41387 817262
rect 40677 816914 40743 816917
rect 40677 816912 40756 816914
rect 40677 816856 40682 816912
rect 40738 816856 40756 816912
rect 40677 816854 40756 816856
rect 40677 816851 40743 816854
rect 41965 816506 42031 816509
rect 651557 816506 651623 816509
rect 41492 816504 42031 816506
rect 41492 816448 41970 816504
rect 42026 816448 42031 816504
rect 41492 816446 42031 816448
rect 650164 816504 651623 816506
rect 650164 816448 651562 816504
rect 651618 816448 651623 816504
rect 650164 816446 651623 816448
rect 41965 816443 42031 816446
rect 651557 816443 651623 816446
rect 41822 816098 41828 816100
rect 41492 816038 41828 816098
rect 41822 816036 41828 816038
rect 41892 816036 41898 816100
rect 41781 815690 41847 815693
rect 41492 815688 41847 815690
rect 41492 815632 41786 815688
rect 41842 815632 41847 815688
rect 41492 815630 41847 815632
rect 41781 815627 41847 815630
rect 44173 815282 44239 815285
rect 41492 815280 44239 815282
rect 41492 815224 44178 815280
rect 44234 815224 44239 815280
rect 41492 815222 44239 815224
rect 44173 815219 44239 815222
rect 41781 814874 41847 814877
rect 41492 814872 41847 814874
rect 41492 814816 41786 814872
rect 41842 814816 41847 814872
rect 41492 814814 41847 814816
rect 41781 814811 41847 814814
rect 41492 814406 41752 814466
rect 41692 814332 41752 814406
rect 41684 814268 41690 814332
rect 41754 814268 41760 814332
rect 41873 814058 41939 814061
rect 41492 814056 41939 814058
rect 41492 814000 41878 814056
rect 41934 814000 41939 814056
rect 41492 813998 41939 814000
rect 41873 813995 41939 813998
rect 44265 813650 44331 813653
rect 41492 813648 44331 813650
rect 41492 813592 44270 813648
rect 44326 813592 44331 813648
rect 41492 813590 44331 813592
rect 44265 813587 44331 813590
rect 41822 813242 41828 813244
rect 41492 813182 41828 813242
rect 41822 813180 41828 813182
rect 41892 813180 41898 813244
rect 42149 812834 42215 812837
rect 41492 812832 42215 812834
rect 41492 812776 42154 812832
rect 42210 812776 42215 812832
rect 41492 812774 42215 812776
rect 42149 812771 42215 812774
rect 33777 812426 33843 812429
rect 33764 812424 33843 812426
rect 33764 812368 33782 812424
rect 33838 812368 33843 812424
rect 33764 812366 33843 812368
rect 33777 812363 33843 812366
rect 35157 812018 35223 812021
rect 35157 812016 35236 812018
rect 35157 811960 35162 812016
rect 35218 811960 35236 812016
rect 35157 811958 35236 811960
rect 35157 811955 35223 811958
rect 40677 811610 40743 811613
rect 40677 811608 40756 811610
rect 40677 811552 40682 811608
rect 40738 811552 40756 811608
rect 40677 811550 40756 811552
rect 40677 811547 40743 811550
rect 42333 811202 42399 811205
rect 41492 811200 42399 811202
rect 41492 811144 42338 811200
rect 42394 811144 42399 811200
rect 41492 811142 42399 811144
rect 42333 811139 42399 811142
rect 34421 810794 34487 810797
rect 34421 810792 34500 810794
rect 34421 810736 34426 810792
rect 34482 810736 34500 810792
rect 34421 810734 34500 810736
rect 34421 810731 34487 810734
rect 33041 810386 33107 810389
rect 33028 810384 33107 810386
rect 33028 810328 33046 810384
rect 33102 810328 33107 810384
rect 33028 810326 33107 810328
rect 33041 810323 33107 810326
rect 44357 809978 44423 809981
rect 41492 809976 44423 809978
rect 41492 809920 44362 809976
rect 44418 809920 44423 809976
rect 41492 809918 44423 809920
rect 44357 809915 44423 809918
rect 42057 809570 42123 809573
rect 41492 809568 42123 809570
rect 41492 809512 42062 809568
rect 42118 809512 42123 809568
rect 41492 809510 42123 809512
rect 42057 809507 42123 809510
rect 32397 809162 32463 809165
rect 32397 809160 32476 809162
rect 32397 809104 32402 809160
rect 32458 809104 32476 809160
rect 32397 809102 32476 809104
rect 32397 809099 32463 809102
rect 35249 808754 35315 808757
rect 35236 808752 35315 808754
rect 35236 808696 35254 808752
rect 35310 808696 35315 808752
rect 35236 808694 35315 808696
rect 35249 808691 35315 808694
rect 44449 808346 44515 808349
rect 41492 808344 44515 808346
rect 41492 808288 44454 808344
rect 44510 808288 44515 808344
rect 41492 808286 44515 808288
rect 44449 808283 44515 808286
rect 41781 807938 41847 807941
rect 41492 807936 41847 807938
rect 41492 807880 41786 807936
rect 41842 807880 41847 807936
rect 41492 807878 41847 807880
rect 41781 807875 41847 807878
rect 35758 807333 35818 807500
rect 35758 807328 35867 807333
rect 35758 807272 35806 807328
rect 35862 807272 35867 807328
rect 35758 807270 35867 807272
rect 35801 807267 35867 807270
rect 24902 806684 24962 807092
rect 62113 806578 62179 806581
rect 62113 806576 64492 806578
rect 62113 806520 62118 806576
rect 62174 806520 64492 806576
rect 62113 806518 64492 806520
rect 62113 806515 62179 806518
rect 41873 806306 41939 806309
rect 43529 806306 43595 806309
rect 41492 806304 43595 806306
rect 41492 806248 41878 806304
rect 41934 806248 43534 806304
rect 43590 806248 43595 806304
rect 41492 806246 43595 806248
rect 41873 806243 41939 806246
rect 43529 806243 43595 806246
rect 40534 804748 40540 804812
rect 40604 804810 40610 804812
rect 41781 804810 41847 804813
rect 40604 804808 41847 804810
rect 40604 804752 41786 804808
rect 41842 804752 41847 804808
rect 40604 804750 41847 804752
rect 40604 804748 40610 804750
rect 41781 804747 41847 804750
rect 651557 803314 651623 803317
rect 650164 803312 651623 803314
rect 650164 803256 651562 803312
rect 651618 803256 651623 803312
rect 650164 803254 651623 803256
rect 651557 803251 651623 803254
rect 35157 802770 35223 802773
rect 42190 802770 42196 802772
rect 35157 802768 42196 802770
rect 35157 802712 35162 802768
rect 35218 802712 42196 802768
rect 35157 802710 42196 802712
rect 35157 802707 35223 802710
rect 42190 802708 42196 802710
rect 42260 802708 42266 802772
rect 34421 802634 34487 802637
rect 41638 802634 41644 802636
rect 34421 802632 41644 802634
rect 34421 802576 34426 802632
rect 34482 802576 41644 802632
rect 34421 802574 41644 802576
rect 34421 802571 34487 802574
rect 41638 802572 41644 802574
rect 41708 802572 41714 802636
rect 33041 802498 33107 802501
rect 42006 802498 42012 802500
rect 33041 802496 42012 802498
rect 33041 802440 33046 802496
rect 33102 802440 42012 802496
rect 33041 802438 42012 802440
rect 33041 802435 33107 802438
rect 42006 802436 42012 802438
rect 42076 802436 42082 802500
rect 33777 801002 33843 801005
rect 41822 801002 41828 801004
rect 33777 801000 41828 801002
rect 33777 800944 33782 801000
rect 33838 800944 41828 801000
rect 33777 800942 41828 800944
rect 33777 800939 33843 800942
rect 41822 800940 41828 800942
rect 41892 800940 41898 801004
rect 40534 796724 40540 796788
rect 40604 796786 40610 796788
rect 42425 796786 42491 796789
rect 40604 796784 42491 796786
rect 40604 796728 42430 796784
rect 42486 796728 42491 796784
rect 40604 796726 42491 796728
rect 40604 796724 40610 796726
rect 42425 796723 42491 796726
rect 62113 793658 62179 793661
rect 62113 793656 64492 793658
rect 62113 793600 62118 793656
rect 62174 793600 64492 793656
rect 62113 793598 64492 793600
rect 62113 793595 62179 793598
rect 42006 791964 42012 792028
rect 42076 792026 42082 792028
rect 42333 792026 42399 792029
rect 42076 792024 42399 792026
rect 42076 791968 42338 792024
rect 42394 791968 42399 792024
rect 42076 791966 42399 791968
rect 42076 791964 42082 791966
rect 42333 791963 42399 791966
rect 651649 789986 651715 789989
rect 650164 789984 651715 789986
rect 650164 789928 651654 789984
rect 651710 789928 651715 789984
rect 650164 789926 651715 789928
rect 651649 789923 651715 789926
rect 42149 788764 42215 788765
rect 42149 788762 42196 788764
rect 42104 788760 42196 788762
rect 42104 788704 42154 788760
rect 42104 788702 42196 788704
rect 42149 788700 42196 788702
rect 42260 788700 42266 788764
rect 42149 788699 42215 788700
rect 41822 788156 41828 788220
rect 41892 788218 41898 788220
rect 42701 788218 42767 788221
rect 41892 788216 42767 788218
rect 41892 788160 42706 788216
rect 42762 788160 42767 788216
rect 41892 788158 42767 788160
rect 41892 788156 41898 788158
rect 42701 788155 42767 788158
rect 41638 788020 41644 788084
rect 41708 788082 41714 788084
rect 42425 788082 42491 788085
rect 675385 788084 675451 788085
rect 675334 788082 675340 788084
rect 41708 788080 42491 788082
rect 41708 788024 42430 788080
rect 42486 788024 42491 788080
rect 41708 788022 42491 788024
rect 675294 788022 675340 788082
rect 675404 788080 675451 788084
rect 675446 788024 675451 788080
rect 41708 788020 41714 788022
rect 42425 788019 42491 788022
rect 675334 788020 675340 788022
rect 675404 788020 675451 788024
rect 675385 788019 675451 788020
rect 41454 786932 41460 786996
rect 41524 786994 41530 786996
rect 41873 786994 41939 786997
rect 41524 786992 41939 786994
rect 41524 786936 41878 786992
rect 41934 786936 41939 786992
rect 41524 786934 41939 786936
rect 41524 786932 41530 786934
rect 41873 786931 41939 786934
rect 675753 786724 675819 786725
rect 675702 786722 675708 786724
rect 675662 786662 675708 786722
rect 675772 786720 675819 786724
rect 675814 786664 675819 786720
rect 675702 786660 675708 786662
rect 675772 786660 675819 786664
rect 675753 786659 675819 786660
rect 675477 784820 675543 784821
rect 675477 784816 675524 784820
rect 675588 784818 675594 784820
rect 675477 784760 675482 784816
rect 675477 784756 675524 784760
rect 675588 784758 675634 784818
rect 675588 784756 675594 784758
rect 675477 784755 675543 784756
rect 675753 784138 675819 784141
rect 676990 784138 676996 784140
rect 675753 784136 676996 784138
rect 675753 784080 675758 784136
rect 675814 784080 676996 784136
rect 675753 784078 676996 784080
rect 675753 784075 675819 784078
rect 676990 784076 676996 784078
rect 677060 784076 677066 784140
rect 62113 780466 62179 780469
rect 62113 780464 64492 780466
rect 62113 780408 62118 780464
rect 62174 780408 64492 780464
rect 62113 780406 64492 780408
rect 62113 780403 62179 780406
rect 651557 776658 651623 776661
rect 650164 776656 651623 776658
rect 650164 776600 651562 776656
rect 651618 776600 651623 776656
rect 650164 776598 651623 776600
rect 651557 776595 651623 776598
rect 675886 774828 675892 774892
rect 675956 774890 675962 774892
rect 677174 774890 677180 774892
rect 675956 774830 677180 774890
rect 675956 774828 675962 774830
rect 677174 774828 677180 774830
rect 677244 774828 677250 774892
rect 35758 774349 35818 774452
rect 35758 774344 35867 774349
rect 35758 774288 35806 774344
rect 35862 774288 35867 774344
rect 35758 774286 35867 774288
rect 35801 774283 35867 774286
rect 41462 773938 41522 774044
rect 50429 773938 50495 773941
rect 41462 773936 50495 773938
rect 41462 773880 50434 773936
rect 50490 773880 50495 773936
rect 41462 773878 50495 773880
rect 50429 773875 50495 773878
rect 675201 773938 675267 773941
rect 675334 773938 675340 773940
rect 675201 773936 675340 773938
rect 675201 773880 675206 773936
rect 675262 773880 675340 773936
rect 675201 773878 675340 773880
rect 675201 773875 675267 773878
rect 675334 773876 675340 773878
rect 675404 773876 675410 773940
rect 43621 773666 43687 773669
rect 41492 773664 43687 773666
rect 41492 773608 43626 773664
rect 43682 773608 43687 773664
rect 41492 773606 43687 773608
rect 43621 773603 43687 773606
rect 40166 773468 40172 773532
rect 40236 773468 40242 773532
rect 40174 773228 40234 773468
rect 675477 773396 675543 773397
rect 675661 773396 675727 773397
rect 675477 773394 675524 773396
rect 675432 773392 675524 773394
rect 675432 773336 675482 773392
rect 675432 773334 675524 773336
rect 675477 773332 675524 773334
rect 675588 773332 675594 773396
rect 675661 773392 675708 773396
rect 675772 773394 675778 773396
rect 675661 773336 675666 773392
rect 675661 773332 675708 773336
rect 675772 773334 675818 773394
rect 675772 773332 675778 773334
rect 675477 773331 675543 773332
rect 675661 773331 675727 773332
rect 676806 773060 676812 773124
rect 676876 773122 676882 773124
rect 677409 773122 677475 773125
rect 676876 773120 677475 773122
rect 676876 773064 677414 773120
rect 677470 773064 677475 773120
rect 676876 773062 677475 773064
rect 676876 773060 676882 773062
rect 677409 773059 677475 773062
rect 676622 772924 676628 772988
rect 676692 772986 676698 772988
rect 677501 772986 677567 772989
rect 676692 772984 677567 772986
rect 676692 772928 677506 772984
rect 677562 772928 677567 772984
rect 676692 772926 677567 772928
rect 676692 772924 676698 772926
rect 677501 772923 677567 772926
rect 44541 772850 44607 772853
rect 41492 772848 44607 772850
rect 41492 772792 44546 772848
rect 44602 772792 44607 772848
rect 41492 772790 44607 772792
rect 44541 772787 44607 772790
rect 676070 772652 676076 772716
rect 676140 772714 676146 772716
rect 680997 772714 681063 772717
rect 676140 772712 681063 772714
rect 676140 772656 681002 772712
rect 681058 772656 681063 772712
rect 676140 772654 681063 772656
rect 676140 772652 676146 772654
rect 680997 772651 681063 772654
rect 44173 772442 44239 772445
rect 41492 772440 44239 772442
rect 41492 772384 44178 772440
rect 44234 772384 44239 772440
rect 41492 772382 44239 772384
rect 44173 772379 44239 772382
rect 42793 772034 42859 772037
rect 41492 772032 42859 772034
rect 41492 771976 42798 772032
rect 42854 771976 42859 772032
rect 41492 771974 42859 771976
rect 42793 771971 42859 771974
rect 39982 771836 39988 771900
rect 40052 771836 40058 771900
rect 39990 771596 40050 771836
rect 39990 771084 40050 771188
rect 39982 771020 39988 771084
rect 40052 771020 40058 771084
rect 44265 770810 44331 770813
rect 41492 770808 44331 770810
rect 41492 770752 44270 770808
rect 44326 770752 44331 770808
rect 41492 770750 44331 770752
rect 44265 770747 44331 770750
rect 44725 770402 44791 770405
rect 41492 770400 44791 770402
rect 41492 770344 44730 770400
rect 44786 770344 44791 770400
rect 41492 770342 44791 770344
rect 44725 770339 44791 770342
rect 42885 769994 42951 769997
rect 41492 769992 42951 769994
rect 41492 769936 42890 769992
rect 42946 769936 42951 769992
rect 41492 769934 42951 769936
rect 42885 769931 42951 769934
rect 33734 769453 33794 769556
rect 33734 769448 33843 769453
rect 33734 769392 33782 769448
rect 33838 769392 33843 769448
rect 33734 769390 33843 769392
rect 33777 769387 33843 769390
rect 40726 769045 40786 769148
rect 40677 769040 40786 769045
rect 40677 768984 40682 769040
rect 40738 768984 40786 769040
rect 40677 768982 40786 768984
rect 40677 768979 40743 768982
rect 32446 768637 32506 768740
rect 32397 768632 32506 768637
rect 32397 768576 32402 768632
rect 32458 768576 32506 768632
rect 32397 768574 32506 768576
rect 32397 768571 32463 768574
rect 42977 768362 43043 768365
rect 41492 768360 43043 768362
rect 41492 768304 42982 768360
rect 43038 768304 43043 768360
rect 41492 768302 43043 768304
rect 42977 768299 43043 768302
rect 30974 767821 31034 767924
rect 30974 767816 31083 767821
rect 30974 767760 31022 767816
rect 31078 767760 31083 767816
rect 30974 767758 31083 767760
rect 31017 767755 31083 767758
rect 33918 767413 33978 767516
rect 33869 767408 33978 767413
rect 33869 767352 33874 767408
rect 33930 767352 33978 767408
rect 33869 767350 33978 767352
rect 62113 767410 62179 767413
rect 62113 767408 64492 767410
rect 62113 767352 62118 767408
rect 62174 767352 64492 767408
rect 62113 767350 64492 767352
rect 33869 767347 33935 767350
rect 62113 767347 62179 767350
rect 44357 767138 44423 767141
rect 41492 767136 44423 767138
rect 41492 767080 44362 767136
rect 44418 767080 44423 767136
rect 41492 767078 44423 767080
rect 44357 767075 44423 767078
rect 32446 766597 32506 766700
rect 32446 766592 32555 766597
rect 32446 766536 32494 766592
rect 32550 766536 32555 766592
rect 32446 766534 32555 766536
rect 32489 766531 32555 766534
rect 675150 766532 675156 766596
rect 675220 766594 675226 766596
rect 675477 766594 675543 766597
rect 675220 766592 675543 766594
rect 675220 766536 675482 766592
rect 675538 766536 675543 766592
rect 675220 766534 675543 766536
rect 675220 766532 675226 766534
rect 675477 766531 675543 766534
rect 675661 766594 675727 766597
rect 676070 766594 676076 766596
rect 675661 766592 676076 766594
rect 675661 766536 675666 766592
rect 675722 766536 676076 766592
rect 675661 766534 676076 766536
rect 675661 766531 675727 766534
rect 676070 766532 676076 766534
rect 676140 766532 676146 766596
rect 40910 766188 40970 766292
rect 40902 766124 40908 766188
rect 40972 766124 40978 766188
rect 43253 765914 43319 765917
rect 41492 765912 43319 765914
rect 41492 765856 43258 765912
rect 43314 765856 43319 765912
rect 41492 765854 43319 765856
rect 43253 765851 43319 765854
rect 44449 765506 44515 765509
rect 41492 765504 44515 765506
rect 41492 765448 44454 765504
rect 44510 765448 44515 765504
rect 41492 765446 44515 765448
rect 44449 765443 44515 765446
rect 40542 764964 40602 765068
rect 674966 765036 674972 765100
rect 675036 765098 675042 765100
rect 675569 765098 675635 765101
rect 675036 765096 675635 765098
rect 675036 765040 675574 765096
rect 675630 765040 675635 765096
rect 675036 765038 675635 765040
rect 675036 765036 675042 765038
rect 675569 765035 675635 765038
rect 40534 764900 40540 764964
rect 40604 764900 40610 764964
rect 40726 764556 40786 764660
rect 40718 764492 40724 764556
rect 40788 764492 40794 764556
rect 30422 764149 30482 764252
rect 30373 764144 30482 764149
rect 30373 764088 30378 764144
rect 30434 764088 30482 764144
rect 30373 764086 30482 764088
rect 30373 764083 30439 764086
rect 30422 763436 30482 763844
rect 30373 763330 30439 763333
rect 651557 763330 651623 763333
rect 30373 763328 30482 763330
rect 30373 763272 30378 763328
rect 30434 763272 30482 763328
rect 30373 763267 30482 763272
rect 650164 763328 651623 763330
rect 650164 763272 651562 763328
rect 651618 763272 651623 763328
rect 650164 763270 651623 763272
rect 651557 763267 651623 763270
rect 30422 763028 30482 763267
rect 41462 762925 41522 763028
rect 41462 762920 41571 762925
rect 41462 762864 41510 762920
rect 41566 762864 41571 762920
rect 41462 762862 41571 762864
rect 41505 762859 41571 762862
rect 676121 761290 676187 761293
rect 676262 761290 676322 761532
rect 676121 761288 676322 761290
rect 676121 761232 676126 761288
rect 676182 761232 676322 761288
rect 676121 761230 676322 761232
rect 676121 761227 676187 761230
rect 676262 760885 676322 761124
rect 676213 760880 676322 760885
rect 676213 760824 676218 760880
rect 676274 760824 676322 760880
rect 676213 760822 676322 760824
rect 676213 760819 676279 760822
rect 676029 760746 676095 760749
rect 676029 760744 676292 760746
rect 676029 760688 676034 760744
rect 676090 760688 676292 760744
rect 676029 760686 676292 760688
rect 676029 760683 676095 760686
rect 676262 760069 676322 760308
rect 676213 760064 676322 760069
rect 676213 760008 676218 760064
rect 676274 760008 676322 760064
rect 676213 760006 676322 760008
rect 676213 760003 676279 760006
rect 674741 759930 674807 759933
rect 674741 759928 676292 759930
rect 674741 759872 674746 759928
rect 674802 759872 676292 759928
rect 674741 759870 676292 759872
rect 674741 759867 674807 759870
rect 676262 759253 676322 759492
rect 676213 759248 676322 759253
rect 676213 759192 676218 759248
rect 676274 759192 676322 759248
rect 676213 759190 676322 759192
rect 676213 759187 676279 759190
rect 674649 759114 674715 759117
rect 674782 759114 674788 759116
rect 674649 759112 674788 759114
rect 674649 759056 674654 759112
rect 674710 759056 674788 759112
rect 674649 759054 674788 759056
rect 674649 759051 674715 759054
rect 674782 759052 674788 759054
rect 674852 759052 674858 759116
rect 676029 759114 676095 759117
rect 676029 759112 676292 759114
rect 676029 759056 676034 759112
rect 676090 759056 676292 759112
rect 676029 759054 676292 759056
rect 676029 759051 676095 759054
rect 676213 758842 676279 758845
rect 676213 758840 676322 758842
rect 676213 758784 676218 758840
rect 676274 758784 676322 758840
rect 676213 758779 676322 758784
rect 676262 758676 676322 758779
rect 33869 758298 33935 758301
rect 41638 758298 41644 758300
rect 33869 758296 41644 758298
rect 33869 758240 33874 758296
rect 33930 758240 41644 758296
rect 33869 758238 41644 758240
rect 33869 758235 33935 758238
rect 41638 758236 41644 758238
rect 41708 758236 41714 758300
rect 676029 758298 676095 758301
rect 676029 758296 676292 758298
rect 676029 758240 676034 758296
rect 676090 758240 676292 758296
rect 676029 758238 676292 758240
rect 676029 758235 676095 758238
rect 674782 757828 674788 757892
rect 674852 757890 674858 757892
rect 674852 757830 676292 757890
rect 674852 757828 674858 757830
rect 40677 757754 40743 757757
rect 41454 757754 41460 757756
rect 40677 757752 41460 757754
rect 40677 757696 40682 757752
rect 40738 757696 41460 757752
rect 40677 757694 41460 757696
rect 40677 757691 40743 757694
rect 41454 757692 41460 757694
rect 41524 757692 41530 757756
rect 676262 757213 676322 757452
rect 676213 757208 676322 757213
rect 677409 757210 677475 757213
rect 676213 757152 676218 757208
rect 676274 757152 676322 757208
rect 676213 757150 676322 757152
rect 677366 757208 677475 757210
rect 677366 757152 677414 757208
rect 677470 757152 677475 757208
rect 676213 757147 676279 757150
rect 677366 757147 677475 757152
rect 41781 757076 41847 757077
rect 42425 757076 42491 757077
rect 41781 757074 41828 757076
rect 41736 757072 41828 757074
rect 41736 757016 41786 757072
rect 41736 757014 41828 757016
rect 41781 757012 41828 757014
rect 41892 757012 41898 757076
rect 42374 757012 42380 757076
rect 42444 757074 42491 757076
rect 42444 757072 42536 757074
rect 42486 757016 42536 757072
rect 677366 757044 677426 757147
rect 42444 757014 42536 757016
rect 42444 757012 42491 757014
rect 41781 757011 41847 757012
rect 42425 757011 42491 757012
rect 677174 756740 677180 756804
rect 677244 756740 677250 756804
rect 677182 756636 677242 756740
rect 676121 755986 676187 755989
rect 676262 755986 676322 756228
rect 676121 755984 676322 755986
rect 676121 755928 676126 755984
rect 676182 755928 676322 755984
rect 676121 755926 676322 755928
rect 680997 755986 681063 755989
rect 680997 755984 681106 755986
rect 680997 755928 681002 755984
rect 681058 755928 681106 755984
rect 676121 755923 676187 755926
rect 680997 755923 681106 755928
rect 681046 755820 681106 755923
rect 676213 755578 676279 755581
rect 676213 755576 676322 755578
rect 676213 755520 676218 755576
rect 676274 755520 676322 755576
rect 676213 755515 676322 755520
rect 676262 755412 676322 755515
rect 676213 755170 676279 755173
rect 676213 755168 676322 755170
rect 676213 755112 676218 755168
rect 676274 755112 676322 755168
rect 676213 755107 676322 755112
rect 676262 755004 676322 755107
rect 41873 754900 41939 754901
rect 41822 754898 41828 754900
rect 41782 754838 41828 754898
rect 41892 754896 41939 754900
rect 41934 754840 41939 754896
rect 41822 754836 41828 754838
rect 41892 754836 41939 754840
rect 41873 754835 41939 754836
rect 677501 754762 677567 754765
rect 677501 754760 677610 754762
rect 677501 754704 677506 754760
rect 677562 754704 677610 754760
rect 677501 754699 677610 754704
rect 677550 754596 677610 754699
rect 62113 754354 62179 754357
rect 62113 754352 64492 754354
rect 62113 754296 62118 754352
rect 62174 754296 64492 754352
rect 62113 754294 64492 754296
rect 62113 754291 62179 754294
rect 40718 754156 40724 754220
rect 40788 754218 40794 754220
rect 42609 754218 42675 754221
rect 40788 754216 42675 754218
rect 40788 754160 42614 754216
rect 42670 754160 42675 754216
rect 40788 754158 42675 754160
rect 40788 754156 40794 754158
rect 42609 754155 42675 754158
rect 676262 753949 676322 754188
rect 676213 753944 676322 753949
rect 676213 753888 676218 753944
rect 676274 753888 676322 753944
rect 676213 753886 676322 753888
rect 676213 753883 676279 753886
rect 677358 753884 677364 753948
rect 677428 753884 677434 753948
rect 677366 753780 677426 753884
rect 676029 753402 676095 753405
rect 676029 753400 676292 753402
rect 676029 753344 676034 753400
rect 676090 753344 676292 753400
rect 676029 753342 676292 753344
rect 676029 753339 676095 753342
rect 40902 753068 40908 753132
rect 40972 753130 40978 753132
rect 41781 753130 41847 753133
rect 40972 753128 41847 753130
rect 40972 753072 41786 753128
rect 41842 753072 41847 753128
rect 40972 753070 41847 753072
rect 40972 753068 40978 753070
rect 41781 753067 41847 753070
rect 676121 752722 676187 752725
rect 676262 752722 676322 752964
rect 676121 752720 676322 752722
rect 676121 752664 676126 752720
rect 676182 752664 676322 752720
rect 676121 752662 676322 752664
rect 676121 752659 676187 752662
rect 673862 752524 673868 752588
rect 673932 752586 673938 752588
rect 673932 752526 676292 752586
rect 673932 752524 673938 752526
rect 676213 752314 676279 752317
rect 676213 752312 676322 752314
rect 676213 752256 676218 752312
rect 676274 752256 676322 752312
rect 676213 752251 676322 752256
rect 676262 752148 676322 752251
rect 676213 751906 676279 751909
rect 676213 751904 676322 751906
rect 676213 751848 676218 751904
rect 676274 751848 676322 751904
rect 676213 751843 676322 751848
rect 676262 751740 676322 751843
rect 683070 751093 683130 751332
rect 683070 751088 683179 751093
rect 683070 751032 683118 751088
rect 683174 751032 683179 751088
rect 683070 751030 683179 751032
rect 683113 751027 683179 751030
rect 683070 750516 683130 750924
rect 40534 750348 40540 750412
rect 40604 750410 40610 750412
rect 41781 750410 41847 750413
rect 40604 750408 41847 750410
rect 40604 750352 41786 750408
rect 41842 750352 41847 750408
rect 40604 750350 41847 750352
rect 40604 750348 40610 750350
rect 41781 750347 41847 750350
rect 683113 750274 683179 750277
rect 683070 750272 683179 750274
rect 683070 750216 683118 750272
rect 683174 750216 683179 750272
rect 683070 750211 683179 750216
rect 651557 750138 651623 750141
rect 650164 750136 651623 750138
rect 650164 750080 651562 750136
rect 651618 750080 651623 750136
rect 683070 750108 683130 750211
rect 650164 750078 651623 750080
rect 651557 750075 651623 750078
rect 42374 749260 42380 749324
rect 42444 749322 42450 749324
rect 42701 749322 42767 749325
rect 42444 749320 42767 749322
rect 42444 749264 42706 749320
rect 42762 749264 42767 749320
rect 42444 749262 42767 749264
rect 42444 749260 42450 749262
rect 42701 749259 42767 749262
rect 41638 746540 41644 746604
rect 41708 746602 41714 746604
rect 42609 746602 42675 746605
rect 41708 746600 42675 746602
rect 41708 746544 42614 746600
rect 42670 746544 42675 746600
rect 41708 746542 42675 746544
rect 41708 746540 41714 746542
rect 42609 746539 42675 746542
rect 41454 742324 41460 742388
rect 41524 742386 41530 742388
rect 41781 742386 41847 742389
rect 41524 742384 41847 742386
rect 41524 742328 41786 742384
rect 41842 742328 41847 742384
rect 41524 742326 41847 742328
rect 41524 742324 41530 742326
rect 41781 742323 41847 742326
rect 675661 741708 675727 741709
rect 675661 741704 675708 741708
rect 675772 741706 675778 741708
rect 675661 741648 675666 741704
rect 675661 741644 675708 741648
rect 675772 741646 675818 741706
rect 675772 741644 675778 741646
rect 675661 741643 675727 741644
rect 62113 741298 62179 741301
rect 62113 741296 64492 741298
rect 62113 741240 62118 741296
rect 62174 741240 64492 741296
rect 62113 741238 64492 741240
rect 62113 741235 62179 741238
rect 651557 736810 651623 736813
rect 650164 736808 651623 736810
rect 650164 736752 651562 736808
rect 651618 736752 651623 736808
rect 650164 736750 651623 736752
rect 651557 736747 651623 736750
rect 674833 736130 674899 736133
rect 675518 736130 675524 736132
rect 674833 736128 675524 736130
rect 674833 736072 674838 736128
rect 674894 736072 675524 736128
rect 674833 736070 675524 736072
rect 674833 736067 674899 736070
rect 675518 736068 675524 736070
rect 675588 736068 675594 736132
rect 675753 734362 675819 734365
rect 676622 734362 676628 734364
rect 675753 734360 676628 734362
rect 675753 734304 675758 734360
rect 675814 734304 676628 734360
rect 675753 734302 676628 734304
rect 675753 734299 675819 734302
rect 676622 734300 676628 734302
rect 676692 734300 676698 734364
rect 675753 733002 675819 733005
rect 677174 733002 677180 733004
rect 675753 733000 677180 733002
rect 675753 732944 675758 733000
rect 675814 732944 677180 733000
rect 675753 732942 677180 732944
rect 675753 732939 675819 732942
rect 677174 732940 677180 732942
rect 677244 732940 677250 733004
rect 31526 731101 31586 731340
rect 31477 731096 31586 731101
rect 31477 731040 31482 731096
rect 31538 731040 31586 731096
rect 31477 731038 31586 731040
rect 31661 731098 31727 731101
rect 31661 731096 31770 731098
rect 31661 731040 31666 731096
rect 31722 731040 31770 731096
rect 31477 731035 31543 731038
rect 31661 731035 31770 731040
rect 31710 730932 31770 731035
rect 31569 730690 31635 730693
rect 31526 730688 31635 730690
rect 31526 730632 31574 730688
rect 31630 730632 31635 730688
rect 31526 730627 31635 730632
rect 31526 730524 31586 730627
rect 31385 730282 31451 730285
rect 31342 730280 31451 730282
rect 31342 730224 31390 730280
rect 31446 730224 31451 730280
rect 31342 730219 31451 730224
rect 31342 730116 31402 730219
rect 40358 729468 40418 729708
rect 40350 729404 40356 729468
rect 40420 729404 40426 729468
rect 42793 729330 42859 729333
rect 41492 729328 42859 729330
rect 41492 729272 42798 729328
rect 42854 729272 42859 729328
rect 41492 729270 42859 729272
rect 42793 729267 42859 729270
rect 44265 728922 44331 728925
rect 41492 728920 44331 728922
rect 41492 728864 44270 728920
rect 44326 728864 44331 728920
rect 41492 728862 44331 728864
rect 44265 728859 44331 728862
rect 39982 728588 39988 728652
rect 40052 728588 40058 728652
rect 39990 728484 40050 728588
rect 675477 728380 675543 728381
rect 675661 728380 675727 728381
rect 675477 728378 675524 728380
rect 675432 728376 675524 728378
rect 675432 728320 675482 728376
rect 675432 728318 675524 728320
rect 675477 728316 675524 728318
rect 675588 728316 675594 728380
rect 675661 728376 675708 728380
rect 675772 728378 675778 728380
rect 675661 728320 675666 728376
rect 675661 728316 675708 728320
rect 675772 728318 675818 728378
rect 675772 728316 675778 728318
rect 675477 728315 675543 728316
rect 675661 728315 675727 728316
rect 62113 728242 62179 728245
rect 62113 728240 64492 728242
rect 62113 728184 62118 728240
rect 62174 728184 64492 728240
rect 62113 728182 64492 728184
rect 62113 728179 62179 728182
rect 40174 727836 40234 728076
rect 40166 727772 40172 727836
rect 40236 727772 40242 727836
rect 44725 727698 44791 727701
rect 41492 727696 44791 727698
rect 41492 727640 44730 727696
rect 44786 727640 44791 727696
rect 41492 727638 44791 727640
rect 44725 727635 44791 727638
rect 44541 727290 44607 727293
rect 41492 727288 44607 727290
rect 41492 727232 44546 727288
rect 44602 727232 44607 727288
rect 41492 727230 44607 727232
rect 44541 727227 44607 727230
rect 674966 727228 674972 727292
rect 675036 727290 675042 727292
rect 678237 727290 678303 727293
rect 675036 727288 678303 727290
rect 675036 727232 678242 727288
rect 678298 727232 678303 727288
rect 675036 727230 678303 727232
rect 675036 727228 675042 727230
rect 678237 727227 678303 727230
rect 30974 726613 31034 726852
rect 30974 726608 31083 726613
rect 30974 726552 31022 726608
rect 31078 726552 31083 726608
rect 30974 726550 31083 726552
rect 31017 726547 31083 726550
rect 675150 726548 675156 726612
rect 675220 726610 675226 726612
rect 680997 726610 681063 726613
rect 675220 726608 681063 726610
rect 675220 726552 681002 726608
rect 681058 726552 681063 726608
rect 675220 726550 681063 726552
rect 675220 726548 675226 726550
rect 680997 726547 681063 726550
rect 40726 726205 40786 726444
rect 40677 726200 40786 726205
rect 40677 726144 40682 726200
rect 40738 726144 40786 726200
rect 40677 726142 40786 726144
rect 40677 726139 40743 726142
rect 39254 725797 39314 726036
rect 39254 725792 39363 725797
rect 39254 725736 39302 725792
rect 39358 725736 39363 725792
rect 39254 725734 39363 725736
rect 39297 725731 39363 725734
rect 41462 725388 41522 725628
rect 41454 725324 41460 725388
rect 41524 725324 41530 725388
rect 42057 725250 42123 725253
rect 41492 725248 42123 725250
rect 41492 725192 42062 725248
rect 42118 725192 42123 725248
rect 41492 725190 42123 725192
rect 42057 725187 42123 725190
rect 40726 724573 40786 724812
rect 40726 724568 40835 724573
rect 40726 724512 40774 724568
rect 40830 724512 40835 724568
rect 40726 724510 40835 724512
rect 40769 724507 40835 724510
rect 44357 724434 44423 724437
rect 41492 724432 44423 724434
rect 41492 724376 44362 724432
rect 44418 724376 44423 724432
rect 41492 724374 44423 724376
rect 44357 724371 44423 724374
rect 676070 724372 676076 724436
rect 676140 724434 676146 724436
rect 679617 724434 679683 724437
rect 676140 724432 679683 724434
rect 676140 724376 679622 724432
rect 679678 724376 679683 724432
rect 676140 724374 679683 724376
rect 676140 724372 676146 724374
rect 679617 724371 679683 724374
rect 35758 723757 35818 723996
rect 35758 723752 35867 723757
rect 35758 723696 35806 723752
rect 35862 723696 35867 723752
rect 35758 723694 35867 723696
rect 35801 723691 35867 723694
rect 35758 723349 35818 723588
rect 652017 723482 652083 723485
rect 650164 723480 652083 723482
rect 650164 723424 652022 723480
rect 652078 723424 652083 723480
rect 650164 723422 652083 723424
rect 652017 723419 652083 723422
rect 35709 723344 35818 723349
rect 35709 723288 35714 723344
rect 35770 723288 35818 723344
rect 35709 723286 35818 723288
rect 40861 723346 40927 723349
rect 40861 723344 40970 723346
rect 40861 723288 40866 723344
rect 40922 723288 40970 723344
rect 35709 723283 35775 723286
rect 40861 723283 40970 723288
rect 40910 723180 40970 723283
rect 42977 722802 43043 722805
rect 41492 722800 43043 722802
rect 41492 722744 42982 722800
rect 43038 722744 43043 722800
rect 41492 722742 43043 722744
rect 42977 722739 43043 722742
rect 44449 722394 44515 722397
rect 41492 722392 44515 722394
rect 41492 722336 44454 722392
rect 44510 722336 44515 722392
rect 41492 722334 44515 722336
rect 44449 722331 44515 722334
rect 44173 721986 44239 721989
rect 41492 721984 44239 721986
rect 41492 721928 44178 721984
rect 44234 721928 44239 721984
rect 41492 721926 44239 721928
rect 44173 721923 44239 721926
rect 675526 721634 676138 721694
rect 675526 721561 675586 721634
rect 675477 721556 675586 721561
rect 40542 721308 40602 721548
rect 675477 721500 675482 721556
rect 675538 721500 675586 721556
rect 675477 721498 675586 721500
rect 675661 721558 675727 721561
rect 676078 721560 676138 721634
rect 675886 721558 675892 721560
rect 675661 721556 675892 721558
rect 675661 721500 675666 721556
rect 675722 721500 675892 721556
rect 675661 721498 675892 721500
rect 675477 721495 675543 721498
rect 675661 721495 675727 721498
rect 675886 721496 675892 721498
rect 675956 721496 675962 721560
rect 676070 721496 676076 721560
rect 676140 721496 676146 721560
rect 40534 721244 40540 721308
rect 40604 721244 40610 721308
rect 41462 720901 41522 721140
rect 41462 720896 41571 720901
rect 41462 720840 41510 720896
rect 41566 720840 41571 720896
rect 41462 720838 41571 720840
rect 41505 720835 41571 720838
rect 27662 720324 27722 720732
rect 41462 719677 41522 719916
rect 41462 719672 41571 719677
rect 41462 719616 41510 719672
rect 41566 719616 41571 719672
rect 41462 719614 41571 719616
rect 41505 719611 41571 719614
rect 676029 716546 676095 716549
rect 676029 716544 676292 716546
rect 676029 716488 676034 716544
rect 676090 716488 676292 716544
rect 676029 716486 676292 716488
rect 676029 716483 676095 716486
rect 39297 716138 39363 716141
rect 41638 716138 41644 716140
rect 39297 716136 41644 716138
rect 39297 716080 39302 716136
rect 39358 716080 41644 716136
rect 39297 716078 41644 716080
rect 39297 716075 39363 716078
rect 41638 716076 41644 716078
rect 41708 716076 41714 716140
rect 676029 716138 676095 716141
rect 676029 716136 676292 716138
rect 676029 716080 676034 716136
rect 676090 716080 676292 716136
rect 676029 716078 676292 716080
rect 676029 716075 676095 716078
rect 676029 715730 676095 715733
rect 676029 715728 676292 715730
rect 676029 715672 676034 715728
rect 676090 715672 676292 715728
rect 676029 715670 676292 715672
rect 676029 715667 676095 715670
rect 31017 715458 31083 715461
rect 41822 715458 41828 715460
rect 31017 715456 41828 715458
rect 31017 715400 31022 715456
rect 31078 715400 41828 715456
rect 31017 715398 41828 715400
rect 31017 715395 31083 715398
rect 41822 715396 41828 715398
rect 41892 715396 41898 715460
rect 62113 715322 62179 715325
rect 674741 715322 674807 715325
rect 62113 715320 64492 715322
rect 62113 715264 62118 715320
rect 62174 715264 64492 715320
rect 62113 715262 64492 715264
rect 674741 715320 676292 715322
rect 674741 715264 674746 715320
rect 674802 715264 676292 715320
rect 674741 715262 676292 715264
rect 62113 715259 62179 715262
rect 674741 715259 674807 715262
rect 674741 714914 674807 714917
rect 674741 714912 676292 714914
rect 674741 714856 674746 714912
rect 674802 714856 676292 714912
rect 674741 714854 676292 714856
rect 674741 714851 674807 714854
rect 676029 714506 676095 714509
rect 676029 714504 676292 714506
rect 676029 714448 676034 714504
rect 676090 714448 676292 714504
rect 676029 714446 676292 714448
rect 676029 714443 676095 714446
rect 676029 714098 676095 714101
rect 676029 714096 676292 714098
rect 676029 714040 676034 714096
rect 676090 714040 676292 714096
rect 676029 714038 676292 714040
rect 676029 714035 676095 714038
rect 42057 713828 42123 713829
rect 42006 713826 42012 713828
rect 41966 713766 42012 713826
rect 42076 713824 42123 713828
rect 42118 713768 42123 713824
rect 42006 713764 42012 713766
rect 42076 713764 42123 713768
rect 42057 713763 42123 713764
rect 676029 713690 676095 713693
rect 676029 713688 676292 713690
rect 676029 713632 676034 713688
rect 676090 713632 676292 713688
rect 676029 713630 676292 713632
rect 676029 713627 676095 713630
rect 676949 713492 677015 713493
rect 676949 713488 676996 713492
rect 677060 713490 677066 713492
rect 676949 713432 676954 713488
rect 676949 713428 676996 713432
rect 677060 713430 677106 713490
rect 677060 713428 677066 713430
rect 676949 713427 677015 713428
rect 42190 713220 42196 713284
rect 42260 713282 42266 713284
rect 42425 713282 42491 713285
rect 42260 713280 42491 713282
rect 42260 713224 42430 713280
rect 42486 713224 42491 713280
rect 42260 713222 42491 713224
rect 42260 713220 42266 713222
rect 42425 713219 42491 713222
rect 676029 713282 676095 713285
rect 676029 713280 676292 713282
rect 676029 713224 676034 713280
rect 676090 713224 676292 713280
rect 676029 713222 676292 713224
rect 676029 713219 676095 713222
rect 676029 712874 676095 712877
rect 676029 712872 676292 712874
rect 676029 712816 676034 712872
rect 676090 712816 676292 712872
rect 676029 712814 676292 712816
rect 676029 712811 676095 712814
rect 676029 712466 676095 712469
rect 676029 712464 676292 712466
rect 676029 712408 676034 712464
rect 676090 712408 676292 712464
rect 676029 712406 676292 712408
rect 676029 712403 676095 712406
rect 678237 712058 678303 712061
rect 678237 712056 678316 712058
rect 678237 712000 678242 712056
rect 678298 712000 678316 712056
rect 678237 711998 678316 712000
rect 678237 711995 678303 711998
rect 676029 711650 676095 711653
rect 676029 711648 676292 711650
rect 676029 711592 676034 711648
rect 676090 711592 676292 711648
rect 676029 711590 676292 711592
rect 676029 711587 676095 711590
rect 679617 711242 679683 711245
rect 679604 711240 679683 711242
rect 679604 711184 679622 711240
rect 679678 711184 679683 711240
rect 679604 711182 679683 711184
rect 679617 711179 679683 711182
rect 40534 710772 40540 710836
rect 40604 710834 40610 710836
rect 42517 710834 42583 710837
rect 40604 710832 42583 710834
rect 40604 710776 42522 710832
rect 42578 710776 42583 710832
rect 40604 710774 42583 710776
rect 40604 710772 40610 710774
rect 42517 710771 42583 710774
rect 680997 710834 681063 710837
rect 680997 710832 681076 710834
rect 680997 710776 681002 710832
rect 681058 710776 681076 710832
rect 680997 710774 681076 710776
rect 680997 710771 681063 710774
rect 676029 710426 676095 710429
rect 676029 710424 676292 710426
rect 676029 710368 676034 710424
rect 676090 710368 676292 710424
rect 676029 710366 676292 710368
rect 676029 710363 676095 710366
rect 651557 710290 651623 710293
rect 650164 710288 651623 710290
rect 650164 710232 651562 710288
rect 651618 710232 651623 710288
rect 650164 710230 651623 710232
rect 651557 710227 651623 710230
rect 676029 710018 676095 710021
rect 676029 710016 676292 710018
rect 676029 709960 676034 710016
rect 676090 709960 676292 710016
rect 676029 709958 676292 709960
rect 676029 709955 676095 709958
rect 676029 709610 676095 709613
rect 676029 709608 676292 709610
rect 676029 709552 676034 709608
rect 676090 709552 676292 709608
rect 676029 709550 676292 709552
rect 676029 709547 676095 709550
rect 676029 709202 676095 709205
rect 676029 709200 676292 709202
rect 676029 709144 676034 709200
rect 676090 709144 676292 709200
rect 676029 709142 676292 709144
rect 676029 709139 676095 709142
rect 676029 708794 676095 708797
rect 676029 708792 676292 708794
rect 676029 708736 676034 708792
rect 676090 708736 676292 708792
rect 676029 708734 676292 708736
rect 676029 708731 676095 708734
rect 42190 708460 42196 708524
rect 42260 708522 42266 708524
rect 42517 708522 42583 708525
rect 42260 708520 42583 708522
rect 42260 708464 42522 708520
rect 42578 708464 42583 708520
rect 42260 708462 42583 708464
rect 42260 708460 42266 708462
rect 42517 708459 42583 708462
rect 676029 708386 676095 708389
rect 676029 708384 676292 708386
rect 676029 708328 676034 708384
rect 676090 708328 676292 708384
rect 676029 708326 676292 708328
rect 676029 708323 676095 708326
rect 676029 707978 676095 707981
rect 676029 707976 676292 707978
rect 676029 707920 676034 707976
rect 676090 707920 676292 707976
rect 676029 707918 676292 707920
rect 676029 707915 676095 707918
rect 676029 707570 676095 707573
rect 676029 707568 676292 707570
rect 676029 707512 676034 707568
rect 676090 707512 676292 707568
rect 676029 707510 676292 707512
rect 676029 707507 676095 707510
rect 676029 707162 676095 707165
rect 676029 707160 676292 707162
rect 676029 707104 676034 707160
rect 676090 707104 676292 707160
rect 676029 707102 676292 707104
rect 676029 707099 676095 707102
rect 42057 706756 42123 706757
rect 42006 706754 42012 706756
rect 41966 706694 42012 706754
rect 42076 706752 42123 706756
rect 42118 706696 42123 706752
rect 42006 706692 42012 706694
rect 42076 706692 42123 706696
rect 42057 706691 42123 706692
rect 675937 706754 676003 706757
rect 675937 706752 676292 706754
rect 675937 706696 675942 706752
rect 675998 706696 676292 706752
rect 675937 706694 676292 706696
rect 675937 706691 676003 706694
rect 676029 706346 676095 706349
rect 676029 706344 676292 706346
rect 676029 706288 676034 706344
rect 676090 706288 676292 706344
rect 676029 706286 676292 706288
rect 676029 706283 676095 706286
rect 676262 705500 676322 705908
rect 42241 705122 42307 705125
rect 42517 705122 42583 705125
rect 42241 705120 42583 705122
rect 42241 705064 42246 705120
rect 42302 705064 42522 705120
rect 42578 705064 42583 705120
rect 42241 705062 42583 705064
rect 42241 705059 42307 705062
rect 42517 705059 42583 705062
rect 676029 705122 676095 705125
rect 676029 705120 676292 705122
rect 676029 705064 676034 705120
rect 676090 705064 676292 705120
rect 676029 705062 676292 705064
rect 676029 705059 676095 705062
rect 41822 703700 41828 703764
rect 41892 703762 41898 703764
rect 42425 703762 42491 703765
rect 41892 703760 42491 703762
rect 41892 703704 42430 703760
rect 42486 703704 42491 703760
rect 41892 703702 42491 703704
rect 41892 703700 41898 703702
rect 42425 703699 42491 703702
rect 41454 702340 41460 702404
rect 41524 702402 41530 702404
rect 41781 702402 41847 702405
rect 41524 702400 41847 702402
rect 41524 702344 41786 702400
rect 41842 702344 41847 702400
rect 41524 702342 41847 702344
rect 41524 702340 41530 702342
rect 41781 702339 41847 702342
rect 62757 702266 62823 702269
rect 62757 702264 64492 702266
rect 62757 702208 62762 702264
rect 62818 702208 64492 702264
rect 62757 702206 64492 702208
rect 62757 702203 62823 702206
rect 41638 699348 41644 699412
rect 41708 699410 41714 699412
rect 41781 699410 41847 699413
rect 41708 699408 41847 699410
rect 41708 699352 41786 699408
rect 41842 699352 41847 699408
rect 41708 699350 41847 699352
rect 41708 699348 41714 699350
rect 41781 699347 41847 699350
rect 652017 696962 652083 696965
rect 675385 696964 675451 696965
rect 675334 696962 675340 696964
rect 650164 696960 652083 696962
rect 650164 696904 652022 696960
rect 652078 696904 652083 696960
rect 650164 696902 652083 696904
rect 675294 696902 675340 696962
rect 675404 696960 675451 696964
rect 675446 696904 675451 696960
rect 652017 696899 652083 696902
rect 675334 696900 675340 696902
rect 675404 696900 675451 696904
rect 675385 696899 675451 696900
rect 675477 694788 675543 694789
rect 675477 694784 675524 694788
rect 675588 694786 675594 694788
rect 675477 694728 675482 694784
rect 675477 694724 675524 694728
rect 675588 694726 675634 694786
rect 675588 694724 675594 694726
rect 675477 694723 675543 694724
rect 675753 694242 675819 694245
rect 676438 694242 676444 694244
rect 675753 694240 676444 694242
rect 675753 694184 675758 694240
rect 675814 694184 676444 694240
rect 675753 694182 676444 694184
rect 675753 694179 675819 694182
rect 676438 694180 676444 694182
rect 676508 694180 676514 694244
rect 62113 689210 62179 689213
rect 62113 689208 64492 689210
rect 62113 689152 62118 689208
rect 62174 689152 64492 689208
rect 62113 689150 64492 689152
rect 62113 689147 62179 689150
rect 35617 688394 35683 688397
rect 35574 688392 35683 688394
rect 35574 688336 35622 688392
rect 35678 688336 35683 688392
rect 35574 688331 35683 688336
rect 35574 688092 35634 688331
rect 35801 687714 35867 687717
rect 35788 687712 35867 687714
rect 35788 687656 35806 687712
rect 35862 687656 35867 687712
rect 35788 687654 35867 687656
rect 35801 687651 35867 687654
rect 675753 687442 675819 687445
rect 676806 687442 676812 687444
rect 675753 687440 676812 687442
rect 675753 687384 675758 687440
rect 675814 687384 676812 687440
rect 675753 687382 676812 687384
rect 675753 687379 675819 687382
rect 676806 687380 676812 687382
rect 676876 687380 676882 687444
rect 30281 687306 30347 687309
rect 30268 687304 30347 687306
rect 30268 687248 30286 687304
rect 30342 687248 30347 687304
rect 30268 687246 30347 687248
rect 30281 687243 30347 687246
rect 40350 687108 40356 687172
rect 40420 687108 40426 687172
rect 40358 686868 40418 687108
rect 44633 686490 44699 686493
rect 41492 686488 44699 686490
rect 41492 686432 44638 686488
rect 44694 686432 44699 686488
rect 41492 686430 44699 686432
rect 44633 686427 44699 686430
rect 675661 686220 675727 686221
rect 675661 686216 675708 686220
rect 675772 686218 675778 686220
rect 675661 686160 675666 686216
rect 675661 686156 675708 686160
rect 675772 686158 675818 686218
rect 675772 686156 675778 686158
rect 675661 686155 675727 686156
rect 44265 686082 44331 686085
rect 41492 686080 44331 686082
rect 41492 686024 44270 686080
rect 44326 686024 44331 686080
rect 41492 686022 44331 686024
rect 44265 686019 44331 686022
rect 44265 685674 44331 685677
rect 41492 685672 44331 685674
rect 41492 685616 44270 685672
rect 44326 685616 44331 685672
rect 41492 685614 44331 685616
rect 44265 685611 44331 685614
rect 40166 685476 40172 685540
rect 40236 685476 40242 685540
rect 40174 685236 40234 685476
rect 39990 684724 40050 684828
rect 39982 684660 39988 684724
rect 40052 684660 40058 684724
rect 44541 684450 44607 684453
rect 41492 684448 44607 684450
rect 41492 684392 44546 684448
rect 44602 684392 44607 684448
rect 41492 684390 44607 684392
rect 44541 684387 44607 684390
rect 44357 684042 44423 684045
rect 41492 684040 44423 684042
rect 41492 683984 44362 684040
rect 44418 683984 44423 684040
rect 41492 683982 44423 683984
rect 44357 683979 44423 683982
rect 39297 683634 39363 683637
rect 651833 683634 651899 683637
rect 39284 683632 39363 683634
rect 39284 683576 39302 683632
rect 39358 683576 39363 683632
rect 39284 683574 39363 683576
rect 650164 683632 651899 683634
rect 650164 683576 651838 683632
rect 651894 683576 651899 683632
rect 650164 683574 651899 683576
rect 39297 683571 39363 683574
rect 651833 683571 651899 683574
rect 675385 683364 675451 683365
rect 675334 683362 675340 683364
rect 675294 683302 675340 683362
rect 675404 683360 675451 683364
rect 675446 683304 675451 683360
rect 675334 683300 675340 683302
rect 675404 683300 675451 683304
rect 675518 683300 675524 683364
rect 675588 683362 675594 683364
rect 675753 683362 675819 683365
rect 675588 683360 675819 683362
rect 675588 683304 675758 683360
rect 675814 683304 675819 683360
rect 675588 683302 675819 683304
rect 675588 683300 675594 683302
rect 675385 683299 675451 683300
rect 675753 683299 675819 683302
rect 675477 683226 675543 683229
rect 675702 683226 675708 683228
rect 675477 683224 675708 683226
rect 41462 683090 41522 683196
rect 675477 683168 675482 683224
rect 675538 683168 675708 683224
rect 675477 683166 675708 683168
rect 675477 683163 675543 683166
rect 675702 683164 675708 683166
rect 675772 683164 675778 683228
rect 676438 683164 676444 683228
rect 676508 683164 676514 683228
rect 676446 683093 676506 683164
rect 41689 683090 41755 683093
rect 41462 683088 41755 683090
rect 41462 683032 41694 683088
rect 41750 683032 41755 683088
rect 41462 683030 41755 683032
rect 676446 683088 676555 683093
rect 676446 683032 676494 683088
rect 676550 683032 676555 683088
rect 676446 683030 676555 683032
rect 41689 683027 41755 683030
rect 676489 683027 676555 683030
rect 32397 682818 32463 682821
rect 32397 682816 32476 682818
rect 32397 682760 32402 682816
rect 32458 682760 32476 682816
rect 32397 682758 32476 682760
rect 32397 682755 32463 682758
rect 41462 682276 41522 682380
rect 41454 682212 41460 682276
rect 41524 682212 41530 682276
rect 41462 681866 41522 681972
rect 41689 681866 41755 681869
rect 41462 681864 41755 681866
rect 41462 681808 41694 681864
rect 41750 681808 41755 681864
rect 41462 681806 41755 681808
rect 41689 681803 41755 681806
rect 675886 681804 675892 681868
rect 675956 681866 675962 681868
rect 679617 681866 679683 681869
rect 675956 681864 679683 681866
rect 675956 681808 679622 681864
rect 679678 681808 679683 681864
rect 675956 681806 679683 681808
rect 675956 681804 675962 681806
rect 679617 681803 679683 681806
rect 31017 681594 31083 681597
rect 31004 681592 31083 681594
rect 31004 681536 31022 681592
rect 31078 681536 31083 681592
rect 31004 681534 31083 681536
rect 31017 681531 31083 681534
rect 42793 681186 42859 681189
rect 41492 681184 42859 681186
rect 41492 681128 42798 681184
rect 42854 681128 42859 681184
rect 41492 681126 42859 681128
rect 42793 681123 42859 681126
rect 41965 680778 42031 680781
rect 41492 680776 42031 680778
rect 41492 680720 41970 680776
rect 42026 680720 42031 680776
rect 41492 680718 42031 680720
rect 41965 680715 42031 680718
rect 35157 680370 35223 680373
rect 35157 680368 35236 680370
rect 35157 680312 35162 680368
rect 35218 680312 35236 680368
rect 35157 680310 35236 680312
rect 35157 680307 35223 680310
rect 44173 679962 44239 679965
rect 41492 679960 44239 679962
rect 41492 679904 44178 679960
rect 44234 679904 44239 679960
rect 41492 679902 44239 679904
rect 44173 679899 44239 679902
rect 40542 679420 40602 679524
rect 40534 679356 40540 679420
rect 40604 679356 40610 679420
rect 42885 679146 42951 679149
rect 41492 679144 42951 679146
rect 41492 679088 42890 679144
rect 42946 679088 42951 679144
rect 41492 679086 42951 679088
rect 42885 679083 42951 679086
rect 44449 678738 44515 678741
rect 41492 678736 44515 678738
rect 41492 678680 44454 678736
rect 44510 678680 44515 678736
rect 41492 678678 44515 678680
rect 44449 678675 44515 678678
rect 40726 678196 40786 678300
rect 676070 678268 676076 678332
rect 676140 678330 676146 678332
rect 679709 678330 679775 678333
rect 676140 678328 679775 678330
rect 676140 678272 679714 678328
rect 679770 678272 679775 678328
rect 676140 678270 679775 678272
rect 676140 678268 676146 678270
rect 679709 678267 679775 678270
rect 40718 678132 40724 678196
rect 40788 678132 40794 678196
rect 30606 677788 30666 677892
rect 30598 677724 30604 677788
rect 30668 677724 30674 677788
rect 27662 677076 27722 677484
rect 30465 676868 30531 676871
rect 30422 676866 30531 676868
rect 30422 676810 30470 676866
rect 30526 676810 30531 676866
rect 30422 676805 30531 676810
rect 30422 676698 30482 676805
rect 30422 676668 30636 676698
rect 30452 676638 30666 676668
rect 30606 676564 30666 676638
rect 30598 676500 30604 676564
rect 30668 676500 30674 676564
rect 675150 676364 675156 676428
rect 675220 676426 675226 676428
rect 675385 676426 675451 676429
rect 675220 676424 675451 676426
rect 675220 676368 675390 676424
rect 675446 676368 675451 676424
rect 675220 676366 675451 676368
rect 675220 676364 675226 676366
rect 675385 676363 675451 676366
rect 675753 676426 675819 676429
rect 675886 676426 675892 676428
rect 675753 676424 675892 676426
rect 675753 676368 675758 676424
rect 675814 676368 675892 676424
rect 675753 676366 675892 676368
rect 675753 676363 675819 676366
rect 675886 676364 675892 676366
rect 675956 676364 675962 676428
rect 676489 676426 676555 676429
rect 676990 676426 676996 676428
rect 676489 676424 676996 676426
rect 676489 676368 676494 676424
rect 676550 676368 676996 676424
rect 676489 676366 676996 676368
rect 676489 676363 676555 676366
rect 676990 676364 676996 676366
rect 677060 676364 677066 676428
rect 62113 676154 62179 676157
rect 62113 676152 64492 676154
rect 62113 676096 62118 676152
rect 62174 676096 64492 676152
rect 62113 676094 64492 676096
rect 62113 676091 62179 676094
rect 32397 671394 32463 671397
rect 41638 671394 41644 671396
rect 32397 671392 41644 671394
rect 32397 671336 32402 671392
rect 32458 671336 41644 671392
rect 32397 671334 41644 671336
rect 32397 671331 32463 671334
rect 41638 671332 41644 671334
rect 41708 671332 41714 671396
rect 676262 671125 676322 671364
rect 676213 671120 676322 671125
rect 676213 671064 676218 671120
rect 676274 671064 676322 671120
rect 676213 671062 676322 671064
rect 676213 671059 676279 671062
rect 39297 670986 39363 670989
rect 42374 670986 42380 670988
rect 39297 670984 42380 670986
rect 39297 670928 39302 670984
rect 39358 670928 42380 670984
rect 39297 670926 42380 670928
rect 39297 670923 39363 670926
rect 42374 670924 42380 670926
rect 42444 670924 42450 670988
rect 676029 670986 676095 670989
rect 676029 670984 676292 670986
rect 676029 670928 676034 670984
rect 676090 670928 676292 670984
rect 676029 670926 676292 670928
rect 676029 670923 676095 670926
rect 41781 670716 41847 670717
rect 42057 670716 42123 670717
rect 41781 670714 41828 670716
rect 41736 670712 41828 670714
rect 41736 670656 41786 670712
rect 41736 670654 41828 670656
rect 41781 670652 41828 670654
rect 41892 670652 41898 670716
rect 42006 670652 42012 670716
rect 42076 670714 42123 670716
rect 42076 670712 42168 670714
rect 42118 670656 42168 670712
rect 42076 670654 42168 670656
rect 42076 670652 42123 670654
rect 41781 670651 41847 670652
rect 42057 670651 42123 670652
rect 651557 670442 651623 670445
rect 650164 670440 651623 670442
rect 650164 670384 651562 670440
rect 651618 670384 651623 670440
rect 650164 670382 651623 670384
rect 651557 670379 651623 670382
rect 676121 670306 676187 670309
rect 676262 670306 676322 670548
rect 676121 670304 676322 670306
rect 676121 670248 676126 670304
rect 676182 670248 676322 670304
rect 676121 670246 676322 670248
rect 676121 670243 676187 670246
rect 42190 670108 42196 670172
rect 42260 670170 42266 670172
rect 42425 670170 42491 670173
rect 42260 670168 42491 670170
rect 42260 670112 42430 670168
rect 42486 670112 42491 670168
rect 42260 670110 42491 670112
rect 42260 670108 42266 670110
rect 42425 670107 42491 670110
rect 674741 670170 674807 670173
rect 674741 670168 676292 670170
rect 674741 670112 674746 670168
rect 674802 670112 676292 670168
rect 674741 670110 676292 670112
rect 674741 670107 674807 670110
rect 676262 669493 676322 669732
rect 676213 669488 676322 669493
rect 676213 669432 676218 669488
rect 676274 669432 676322 669488
rect 676213 669430 676322 669432
rect 676213 669427 676279 669430
rect 676029 669354 676095 669357
rect 676029 669352 676292 669354
rect 676029 669296 676034 669352
rect 676090 669296 676292 669352
rect 676029 669294 676292 669296
rect 676029 669291 676095 669294
rect 672349 669082 672415 669085
rect 672942 669082 672948 669084
rect 672349 669080 672948 669082
rect 672349 669024 672354 669080
rect 672410 669024 672948 669080
rect 672349 669022 672948 669024
rect 672349 669019 672415 669022
rect 672942 669020 672948 669022
rect 673012 669020 673018 669084
rect 676262 668677 676322 668916
rect 676213 668672 676322 668677
rect 676213 668616 676218 668672
rect 676274 668616 676322 668672
rect 676213 668614 676322 668616
rect 676213 668611 676279 668614
rect 41873 668540 41939 668541
rect 41822 668538 41828 668540
rect 41782 668478 41828 668538
rect 41892 668536 41939 668540
rect 41934 668480 41939 668536
rect 41822 668476 41828 668478
rect 41892 668476 41939 668480
rect 41873 668475 41939 668476
rect 676029 668538 676095 668541
rect 676029 668536 676292 668538
rect 676029 668480 676034 668536
rect 676090 668480 676292 668536
rect 676029 668478 676292 668480
rect 676029 668475 676095 668478
rect 41822 668340 41828 668404
rect 41892 668402 41898 668404
rect 42374 668402 42380 668404
rect 41892 668342 42380 668402
rect 41892 668340 41898 668342
rect 42374 668340 42380 668342
rect 42444 668340 42450 668404
rect 674741 668130 674807 668133
rect 674741 668128 676292 668130
rect 674741 668072 674746 668128
rect 674802 668072 676292 668128
rect 674741 668070 676292 668072
rect 674741 668067 674807 668070
rect 676262 667453 676322 667692
rect 676213 667448 676322 667453
rect 676213 667392 676218 667448
rect 676274 667392 676322 667448
rect 676213 667390 676322 667392
rect 676213 667387 676279 667390
rect 676029 667314 676095 667317
rect 676029 667312 676292 667314
rect 676029 667256 676034 667312
rect 676090 667256 676292 667312
rect 676029 667254 676292 667256
rect 676029 667251 676095 667254
rect 679617 667042 679683 667045
rect 679574 667040 679683 667042
rect 679574 666984 679622 667040
rect 679678 666984 679683 667040
rect 679574 666979 679683 666984
rect 679574 666876 679634 666979
rect 676121 666226 676187 666229
rect 676262 666226 676322 666468
rect 676121 666224 676322 666226
rect 676121 666168 676126 666224
rect 676182 666168 676322 666224
rect 676121 666166 676322 666168
rect 676121 666163 676187 666166
rect 676262 665821 676322 666060
rect 676213 665816 676322 665821
rect 676213 665760 676218 665816
rect 676274 665760 676322 665816
rect 676213 665758 676322 665760
rect 679709 665818 679775 665821
rect 679709 665816 679818 665818
rect 679709 665760 679714 665816
rect 679770 665760 679818 665816
rect 676213 665755 676279 665758
rect 679709 665755 679818 665760
rect 679758 665652 679818 665755
rect 40718 665348 40724 665412
rect 40788 665410 40794 665412
rect 41781 665410 41847 665413
rect 40788 665408 41847 665410
rect 40788 665352 41786 665408
rect 41842 665352 41847 665408
rect 40788 665350 41847 665352
rect 40788 665348 40794 665350
rect 41781 665347 41847 665350
rect 676029 665274 676095 665277
rect 676029 665272 676292 665274
rect 676029 665216 676034 665272
rect 676090 665216 676292 665272
rect 676029 665214 676292 665216
rect 676029 665211 676095 665214
rect 676213 665002 676279 665005
rect 676213 665000 676322 665002
rect 676213 664944 676218 665000
rect 676274 664944 676322 665000
rect 676213 664939 676322 664944
rect 676262 664836 676322 664939
rect 40534 664532 40540 664596
rect 40604 664594 40610 664596
rect 41781 664594 41847 664597
rect 40604 664592 41847 664594
rect 40604 664536 41786 664592
rect 41842 664536 41847 664592
rect 40604 664534 41847 664536
rect 40604 664532 40610 664534
rect 41781 664531 41847 664534
rect 676262 664189 676322 664428
rect 676213 664184 676322 664189
rect 676213 664128 676218 664184
rect 676274 664128 676322 664184
rect 676213 664126 676322 664128
rect 676213 664123 676279 664126
rect 676262 663781 676322 664020
rect 676213 663776 676322 663781
rect 676213 663720 676218 663776
rect 676274 663720 676322 663776
rect 676213 663718 676322 663720
rect 676213 663715 676279 663718
rect 676262 663373 676322 663612
rect 42057 663372 42123 663373
rect 42006 663370 42012 663372
rect 41966 663310 42012 663370
rect 42076 663368 42123 663372
rect 42118 663312 42123 663368
rect 42006 663308 42012 663310
rect 42076 663308 42123 663312
rect 42057 663307 42123 663308
rect 676213 663368 676322 663373
rect 676213 663312 676218 663368
rect 676274 663312 676322 663368
rect 676213 663310 676322 663312
rect 676213 663307 676279 663310
rect 677174 663308 677180 663372
rect 677244 663308 677250 663372
rect 677182 663204 677242 663308
rect 62113 663098 62179 663101
rect 62113 663096 64492 663098
rect 62113 663040 62118 663096
rect 62174 663040 64492 663096
rect 62113 663038 64492 663040
rect 62113 663035 62179 663038
rect 676622 662900 676628 662964
rect 676692 662900 676698 662964
rect 676630 662796 676690 662900
rect 676029 662418 676095 662421
rect 676029 662416 676292 662418
rect 676029 662360 676034 662416
rect 676090 662360 676292 662416
rect 676029 662358 676292 662360
rect 676029 662355 676095 662358
rect 676262 661741 676322 661980
rect 676213 661736 676322 661741
rect 676213 661680 676218 661736
rect 676274 661680 676322 661736
rect 676213 661678 676322 661680
rect 676213 661675 676279 661678
rect 41454 661268 41460 661332
rect 41524 661330 41530 661332
rect 42701 661330 42767 661333
rect 41524 661328 42767 661330
rect 41524 661272 42706 661328
rect 42762 661272 42767 661328
rect 41524 661270 42767 661272
rect 41524 661268 41530 661270
rect 42701 661267 42767 661270
rect 676121 661330 676187 661333
rect 676262 661330 676322 661572
rect 676121 661328 676322 661330
rect 676121 661272 676126 661328
rect 676182 661272 676322 661328
rect 676121 661270 676322 661272
rect 676121 661267 676187 661270
rect 683070 660925 683130 661164
rect 683070 660920 683179 660925
rect 683070 660864 683118 660920
rect 683174 660864 683179 660920
rect 683070 660862 683179 660864
rect 683113 660859 683179 660862
rect 42149 660516 42215 660517
rect 42149 660514 42196 660516
rect 42104 660512 42196 660514
rect 42104 660456 42154 660512
rect 42104 660454 42196 660456
rect 42149 660452 42196 660454
rect 42260 660452 42266 660516
rect 42149 660451 42215 660452
rect 41822 660316 41828 660380
rect 41892 660378 41898 660380
rect 42517 660378 42583 660381
rect 41892 660376 42583 660378
rect 41892 660320 42522 660376
rect 42578 660320 42583 660376
rect 685830 660348 685890 660756
rect 41892 660318 42583 660320
rect 41892 660316 41898 660318
rect 42517 660315 42583 660318
rect 683113 660106 683179 660109
rect 683070 660104 683179 660106
rect 683070 660048 683118 660104
rect 683174 660048 683179 660104
rect 683070 660043 683179 660048
rect 683070 659940 683130 660043
rect 41638 658276 41644 658340
rect 41708 658338 41714 658340
rect 42333 658338 42399 658341
rect 41708 658336 42399 658338
rect 41708 658280 42338 658336
rect 42394 658280 42399 658336
rect 41708 658278 42399 658280
rect 41708 658276 41714 658278
rect 42333 658275 42399 658278
rect 651557 657114 651623 657117
rect 650164 657112 651623 657114
rect 650164 657056 651562 657112
rect 651618 657056 651623 657112
rect 650164 657054 651623 657056
rect 651557 657051 651623 657054
rect 62113 650042 62179 650045
rect 62113 650040 64492 650042
rect 62113 649984 62118 650040
rect 62174 649984 64492 650040
rect 62113 649982 64492 649984
rect 62113 649979 62179 649982
rect 675385 649908 675451 649909
rect 675334 649906 675340 649908
rect 675294 649846 675340 649906
rect 675404 649904 675451 649908
rect 675446 649848 675451 649904
rect 675334 649844 675340 649846
rect 675404 649844 675451 649848
rect 675385 649843 675451 649844
rect 675753 648682 675819 648685
rect 676622 648682 676628 648684
rect 675753 648680 676628 648682
rect 675753 648624 675758 648680
rect 675814 648624 676628 648680
rect 675753 648622 676628 648624
rect 675753 648619 675819 648622
rect 676622 648620 676628 648622
rect 676692 648620 676698 648684
rect 675201 645962 675267 645965
rect 675518 645962 675524 645964
rect 675201 645960 675524 645962
rect 675201 645904 675206 645960
rect 675262 645904 675524 645960
rect 675201 645902 675524 645904
rect 675201 645899 675267 645902
rect 675518 645900 675524 645902
rect 675588 645900 675594 645964
rect 35574 644741 35634 644912
rect 35574 644736 35683 644741
rect 35801 644738 35867 644741
rect 35574 644680 35622 644736
rect 35678 644680 35683 644736
rect 35574 644678 35683 644680
rect 35617 644675 35683 644678
rect 35758 644736 35867 644738
rect 35758 644680 35806 644736
rect 35862 644680 35867 644736
rect 35758 644675 35867 644680
rect 675753 644738 675819 644741
rect 677174 644738 677180 644740
rect 675753 644736 677180 644738
rect 675753 644680 675758 644736
rect 675814 644680 677180 644736
rect 675753 644678 677180 644680
rect 675753 644675 675819 644678
rect 677174 644676 677180 644678
rect 677244 644676 677250 644740
rect 35758 644504 35818 644675
rect 677174 644602 677180 644604
rect 675710 644542 677180 644602
rect 41462 643922 41522 644096
rect 41462 643862 45570 643922
rect 44633 643786 44699 643789
rect 41462 643784 44699 643786
rect 41462 643728 44638 643784
rect 44694 643728 44699 643784
rect 41462 643726 44699 643728
rect 41462 643688 41522 643726
rect 44633 643723 44699 643726
rect 45510 643514 45570 643862
rect 651557 643786 651623 643789
rect 650164 643784 651623 643786
rect 650164 643728 651562 643784
rect 651618 643728 651623 643784
rect 650164 643726 651623 643728
rect 651557 643723 651623 643726
rect 62757 643514 62823 643517
rect 45510 643512 62823 643514
rect 45510 643456 62762 643512
rect 62818 643456 62823 643512
rect 45510 643454 62823 643456
rect 62757 643451 62823 643454
rect 41462 643242 41522 643280
rect 44173 643242 44239 643245
rect 41462 643240 44239 643242
rect 41462 643184 44178 643240
rect 44234 643184 44239 643240
rect 41462 643182 44239 643184
rect 44173 643179 44239 643182
rect 675710 643109 675770 644542
rect 677174 644540 677180 644542
rect 677244 644540 677250 644604
rect 44265 643106 44331 643109
rect 41462 643104 44331 643106
rect 41462 643048 44270 643104
rect 44326 643048 44331 643104
rect 41462 643046 44331 643048
rect 41462 642872 41522 643046
rect 44265 643043 44331 643046
rect 675661 643104 675770 643109
rect 675661 643048 675666 643104
rect 675722 643048 675770 643104
rect 675661 643046 675770 643048
rect 675661 643043 675727 643046
rect 39982 642228 39988 642292
rect 40052 642228 40058 642292
rect 41462 642290 41522 642464
rect 44633 642290 44699 642293
rect 41462 642288 44699 642290
rect 41462 642232 44638 642288
rect 44694 642232 44699 642288
rect 41462 642230 44699 642232
rect 39990 642056 40050 642228
rect 44633 642227 44699 642230
rect 39990 641476 40050 641648
rect 39982 641412 39988 641476
rect 40052 641412 40058 641476
rect 44357 641474 44423 641477
rect 41462 641472 44423 641474
rect 41462 641416 44362 641472
rect 44418 641416 44423 641472
rect 41462 641414 44423 641416
rect 41462 641240 41522 641414
rect 44357 641411 44423 641414
rect 41462 640658 41522 640832
rect 44725 640658 44791 640661
rect 41462 640656 44791 640658
rect 41462 640600 44730 640656
rect 44786 640600 44791 640656
rect 41462 640598 44791 640600
rect 44725 640595 44791 640598
rect 35206 640253 35266 640424
rect 35157 640248 35266 640253
rect 35157 640192 35162 640248
rect 35218 640192 35266 640248
rect 35157 640190 35266 640192
rect 35157 640187 35223 640190
rect 39254 639845 39314 640016
rect 39254 639840 39363 639845
rect 39254 639784 39302 639840
rect 39358 639784 39363 639840
rect 39254 639782 39363 639784
rect 39297 639779 39363 639782
rect 41462 639436 41522 639608
rect 41454 639372 41460 639436
rect 41524 639372 41530 639436
rect 40726 639029 40786 639200
rect 40677 639024 40786 639029
rect 40677 638968 40682 639024
rect 40738 638968 40786 639024
rect 40677 638966 40786 638968
rect 40677 638963 40743 638966
rect 41462 638618 41522 638792
rect 675201 638754 675267 638757
rect 675334 638754 675340 638756
rect 675201 638752 675340 638754
rect 675201 638696 675206 638752
rect 675262 638696 675340 638752
rect 675201 638694 675340 638696
rect 675201 638691 675267 638694
rect 675334 638692 675340 638694
rect 675404 638692 675410 638756
rect 42885 638618 42951 638621
rect 41462 638616 42951 638618
rect 41462 638560 42890 638616
rect 42946 638560 42951 638616
rect 41462 638558 42951 638560
rect 42885 638555 42951 638558
rect 32446 638213 32506 638384
rect 32397 638208 32506 638213
rect 675477 638212 675543 638213
rect 675477 638210 675524 638212
rect 32397 638152 32402 638208
rect 32458 638152 32506 638208
rect 32397 638150 32506 638152
rect 675432 638208 675524 638210
rect 675432 638152 675482 638208
rect 675432 638150 675524 638152
rect 32397 638147 32463 638150
rect 675477 638148 675524 638150
rect 675588 638148 675594 638212
rect 675477 638147 675543 638148
rect 33734 637805 33794 637976
rect 676622 637876 676628 637940
rect 676692 637938 676698 637940
rect 676857 637938 676923 637941
rect 676692 637936 676923 637938
rect 676692 637880 676862 637936
rect 676918 637880 676923 637936
rect 676692 637878 676923 637880
rect 676692 637876 676698 637878
rect 676857 637875 676923 637878
rect 676990 637876 676996 637940
rect 677060 637938 677066 637940
rect 677501 637938 677567 637941
rect 677060 637936 677567 637938
rect 677060 637880 677506 637936
rect 677562 637880 677567 637936
rect 677060 637878 677567 637880
rect 677060 637876 677066 637878
rect 677501 637875 677567 637878
rect 33734 637800 33843 637805
rect 33734 637744 33782 637800
rect 33838 637744 33843 637800
rect 33734 637742 33843 637744
rect 33777 637739 33843 637742
rect 40910 637397 40970 637568
rect 675886 637468 675892 637532
rect 675956 637530 675962 637532
rect 680997 637530 681063 637533
rect 675956 637528 681063 637530
rect 675956 637472 681002 637528
rect 681058 637472 681063 637528
rect 675956 637470 681063 637472
rect 675956 637468 675962 637470
rect 680997 637467 681063 637470
rect 40861 637392 40970 637397
rect 40861 637336 40866 637392
rect 40922 637336 40970 637392
rect 40861 637334 40970 637336
rect 40861 637331 40927 637334
rect 675150 637332 675156 637396
rect 675220 637394 675226 637396
rect 679617 637394 679683 637397
rect 675220 637392 679683 637394
rect 675220 637336 679622 637392
rect 679678 637336 679683 637392
rect 675220 637334 679683 637336
rect 675220 637332 675226 637334
rect 679617 637331 679683 637334
rect 41462 636986 41522 637160
rect 62113 637122 62179 637125
rect 62113 637120 64492 637122
rect 62113 637064 62118 637120
rect 62174 637064 64492 637120
rect 62113 637062 64492 637064
rect 62113 637059 62179 637062
rect 44449 636986 44515 636989
rect 41462 636984 44515 636986
rect 41462 636928 44454 636984
rect 44510 636928 44515 636984
rect 41462 636926 44515 636928
rect 44449 636923 44515 636926
rect 40910 636580 40970 636752
rect 40902 636516 40908 636580
rect 40972 636516 40978 636580
rect 40542 636172 40602 636344
rect 40534 636108 40540 636172
rect 40604 636108 40610 636172
rect 41462 635762 41522 635936
rect 42793 635762 42859 635765
rect 41462 635760 42859 635762
rect 41462 635704 42798 635760
rect 42854 635704 42859 635760
rect 41462 635702 42859 635704
rect 42793 635699 42859 635702
rect 41462 635354 41522 635528
rect 44541 635354 44607 635357
rect 41462 635352 44607 635354
rect 41462 635296 44546 635352
rect 44602 635296 44607 635352
rect 41462 635294 44607 635296
rect 44541 635291 44607 635294
rect 40726 634948 40786 635120
rect 40718 634884 40724 634948
rect 40788 634884 40794 634948
rect 41462 634538 41522 634712
rect 41462 634478 41890 634538
rect 30422 633896 30482 634304
rect 41830 633722 41890 634478
rect 41462 633662 41890 633722
rect 41462 633450 41522 633662
rect 54477 633450 54543 633453
rect 41462 633448 54543 633450
rect 41462 633392 54482 633448
rect 54538 633392 54543 633448
rect 41462 633390 54543 633392
rect 54477 633387 54543 633390
rect 675201 631410 675267 631413
rect 676070 631410 676076 631412
rect 675201 631408 676076 631410
rect 675201 631352 675206 631408
rect 675262 631352 676076 631408
rect 675201 631350 676076 631352
rect 675201 631347 675267 631350
rect 676070 631348 676076 631350
rect 676140 631348 676146 631412
rect 676857 631410 676923 631413
rect 676990 631410 676996 631412
rect 676857 631408 676996 631410
rect 676857 631352 676862 631408
rect 676918 631352 676996 631408
rect 676857 631350 676996 631352
rect 676857 631347 676923 631350
rect 676990 631348 676996 631350
rect 677060 631348 677066 631412
rect 651557 630594 651623 630597
rect 650164 630592 651623 630594
rect 650164 630536 651562 630592
rect 651618 630536 651623 630592
rect 650164 630534 651623 630536
rect 651557 630531 651623 630534
rect 33777 629914 33843 629917
rect 41638 629914 41644 629916
rect 33777 629912 41644 629914
rect 33777 629856 33782 629912
rect 33838 629856 41644 629912
rect 33777 629854 41644 629856
rect 33777 629851 33843 629854
rect 41638 629852 41644 629854
rect 41708 629852 41714 629916
rect 40861 629234 40927 629237
rect 42190 629234 42196 629236
rect 40861 629232 42196 629234
rect 40861 629176 40866 629232
rect 40922 629176 42196 629232
rect 40861 629174 42196 629176
rect 40861 629171 40927 629174
rect 42190 629172 42196 629174
rect 42260 629172 42266 629236
rect 40677 629098 40743 629101
rect 42006 629098 42012 629100
rect 40677 629096 42012 629098
rect 40677 629040 40682 629096
rect 40738 629040 42012 629096
rect 40677 629038 42012 629040
rect 40677 629035 40743 629038
rect 42006 629036 42012 629038
rect 42076 629036 42082 629100
rect 35157 628554 35223 628557
rect 41822 628554 41828 628556
rect 35157 628552 41828 628554
rect 35157 628496 35162 628552
rect 35218 628496 41828 628552
rect 35157 628494 41828 628496
rect 35157 628491 35223 628494
rect 41822 628492 41828 628494
rect 41892 628492 41898 628556
rect 676121 626106 676187 626109
rect 676262 626106 676322 626348
rect 676121 626104 676322 626106
rect 676121 626048 676126 626104
rect 676182 626048 676322 626104
rect 676121 626046 676322 626048
rect 676121 626043 676187 626046
rect 676262 625701 676322 625940
rect 676213 625696 676322 625701
rect 676213 625640 676218 625696
rect 676274 625640 676322 625696
rect 676213 625638 676322 625640
rect 676213 625635 676279 625638
rect 676262 625293 676322 625532
rect 40902 625228 40908 625292
rect 40972 625290 40978 625292
rect 40972 625230 42442 625290
rect 40972 625228 40978 625230
rect 42382 625154 42442 625230
rect 676213 625288 676322 625293
rect 676213 625232 676218 625288
rect 676274 625232 676322 625288
rect 676213 625230 676322 625232
rect 676213 625227 676279 625230
rect 42517 625154 42583 625157
rect 42382 625152 42583 625154
rect 42382 625096 42522 625152
rect 42578 625096 42583 625152
rect 42382 625094 42583 625096
rect 42517 625091 42583 625094
rect 676262 624885 676322 625124
rect 676213 624880 676322 624885
rect 676213 624824 676218 624880
rect 676274 624824 676322 624880
rect 676213 624822 676322 624824
rect 676213 624819 676279 624822
rect 676121 624474 676187 624477
rect 676262 624474 676322 624716
rect 676121 624472 676322 624474
rect 676121 624416 676126 624472
rect 676182 624416 676322 624472
rect 676121 624414 676322 624416
rect 676121 624411 676187 624414
rect 676262 624069 676322 624308
rect 62113 624066 62179 624069
rect 62113 624064 64492 624066
rect 62113 624008 62118 624064
rect 62174 624008 64492 624064
rect 62113 624006 64492 624008
rect 676213 624064 676322 624069
rect 676213 624008 676218 624064
rect 676274 624008 676322 624064
rect 676213 624006 676322 624008
rect 62113 624003 62179 624006
rect 676213 624003 676279 624006
rect 676029 623930 676095 623933
rect 676029 623928 676292 623930
rect 676029 623872 676034 623928
rect 676090 623872 676292 623928
rect 676029 623870 676292 623872
rect 676029 623867 676095 623870
rect 40718 623732 40724 623796
rect 40788 623794 40794 623796
rect 42517 623794 42583 623797
rect 40788 623792 42583 623794
rect 40788 623736 42522 623792
rect 42578 623736 42583 623792
rect 40788 623734 42583 623736
rect 40788 623732 40794 623734
rect 42517 623731 42583 623734
rect 676213 623658 676279 623661
rect 676213 623656 676322 623658
rect 676213 623600 676218 623656
rect 676274 623600 676322 623656
rect 676213 623595 676322 623600
rect 676262 623492 676322 623595
rect 676029 623114 676095 623117
rect 676029 623112 676292 623114
rect 676029 623056 676034 623112
rect 676090 623056 676292 623112
rect 676029 623054 676292 623056
rect 676029 623051 676095 623054
rect 676213 622842 676279 622845
rect 676213 622840 676322 622842
rect 676213 622784 676218 622840
rect 676274 622784 676322 622840
rect 676213 622779 676322 622784
rect 676262 622676 676322 622779
rect 676029 622298 676095 622301
rect 676029 622296 676292 622298
rect 676029 622240 676034 622296
rect 676090 622240 676292 622296
rect 676029 622238 676292 622240
rect 676029 622235 676095 622238
rect 679617 622026 679683 622029
rect 679574 622024 679683 622026
rect 679574 621968 679622 622024
rect 679678 621968 679683 622024
rect 679574 621963 679683 621968
rect 679574 621860 679634 621963
rect 681089 621618 681155 621621
rect 681046 621616 681155 621618
rect 681046 621560 681094 621616
rect 681150 621560 681155 621616
rect 681046 621555 681155 621560
rect 40534 621420 40540 621484
rect 40604 621482 40610 621484
rect 41781 621482 41847 621485
rect 40604 621480 41847 621482
rect 40604 621424 41786 621480
rect 41842 621424 41847 621480
rect 681046 621452 681106 621555
rect 40604 621422 41847 621424
rect 40604 621420 40610 621422
rect 41781 621419 41847 621422
rect 676213 621210 676279 621213
rect 676213 621208 676322 621210
rect 676213 621152 676218 621208
rect 676274 621152 676322 621208
rect 676213 621147 676322 621152
rect 676262 621044 676322 621147
rect 680997 620802 681063 620805
rect 680997 620800 681106 620802
rect 680997 620744 681002 620800
rect 681058 620744 681106 620800
rect 680997 620739 681106 620744
rect 681046 620636 681106 620739
rect 676262 619989 676322 620228
rect 676213 619984 676322 619989
rect 676213 619928 676218 619984
rect 676274 619928 676322 619984
rect 676213 619926 676322 619928
rect 676213 619923 676279 619926
rect 676029 619850 676095 619853
rect 676029 619848 676292 619850
rect 676029 619792 676034 619848
rect 676090 619792 676292 619848
rect 676029 619790 676292 619792
rect 676029 619787 676095 619790
rect 676262 619173 676322 619412
rect 676213 619168 676322 619173
rect 676213 619112 676218 619168
rect 676274 619112 676322 619168
rect 676213 619110 676322 619112
rect 676213 619107 676279 619110
rect 42006 618972 42012 619036
rect 42076 619034 42082 619036
rect 42241 619034 42307 619037
rect 42076 619032 42307 619034
rect 42076 618976 42246 619032
rect 42302 618976 42307 619032
rect 42076 618974 42307 618976
rect 42076 618972 42082 618974
rect 42241 618971 42307 618974
rect 676029 619034 676095 619037
rect 676029 619032 676292 619034
rect 676029 618976 676034 619032
rect 676090 618976 676292 619032
rect 676029 618974 676292 618976
rect 676029 618971 676095 618974
rect 677501 618762 677567 618765
rect 677501 618760 677610 618762
rect 677501 618704 677506 618760
rect 677562 618704 677610 618760
rect 677501 618699 677610 618704
rect 677550 618596 677610 618699
rect 676806 618292 676812 618356
rect 676876 618292 676882 618356
rect 676814 618188 676874 618292
rect 676262 617541 676322 617780
rect 676213 617536 676322 617541
rect 676213 617480 676218 617536
rect 676274 617480 676322 617536
rect 676213 617478 676322 617480
rect 676213 617475 676279 617478
rect 676029 617402 676095 617405
rect 676029 617400 676292 617402
rect 676029 617344 676034 617400
rect 676090 617344 676292 617400
rect 676029 617342 676292 617344
rect 676029 617339 676095 617342
rect 652385 617266 652451 617269
rect 650164 617264 652451 617266
rect 650164 617208 652390 617264
rect 652446 617208 652451 617264
rect 650164 617206 652451 617208
rect 652385 617203 652451 617206
rect 676029 616994 676095 616997
rect 676029 616992 676292 616994
rect 676029 616936 676034 616992
rect 676090 616936 676292 616992
rect 676029 616934 676292 616936
rect 676029 616931 676095 616934
rect 41822 616796 41828 616860
rect 41892 616858 41898 616860
rect 42517 616858 42583 616861
rect 41892 616856 42583 616858
rect 41892 616800 42522 616856
rect 42578 616800 42583 616856
rect 41892 616798 42583 616800
rect 41892 616796 41898 616798
rect 42517 616795 42583 616798
rect 42149 616724 42215 616725
rect 42149 616722 42196 616724
rect 42104 616720 42196 616722
rect 42104 616664 42154 616720
rect 42104 616662 42196 616664
rect 42149 616660 42196 616662
rect 42260 616660 42266 616724
rect 676213 616722 676279 616725
rect 676213 616720 676322 616722
rect 676213 616664 676218 616720
rect 676274 616664 676322 616720
rect 42149 616659 42215 616660
rect 676213 616659 676322 616664
rect 676262 616556 676322 616659
rect 683070 615909 683130 616148
rect 683070 615904 683179 615909
rect 683070 615848 683118 615904
rect 683174 615848 683179 615904
rect 683070 615846 683179 615848
rect 683113 615843 683179 615846
rect 683070 615332 683130 615740
rect 683113 615090 683179 615093
rect 683070 615088 683179 615090
rect 683070 615032 683118 615088
rect 683174 615032 683179 615088
rect 683070 615027 683179 615032
rect 683070 614924 683130 615027
rect 41454 614076 41460 614140
rect 41524 614138 41530 614140
rect 42517 614138 42583 614141
rect 41524 614136 42583 614138
rect 41524 614080 42522 614136
rect 42578 614080 42583 614136
rect 41524 614078 42583 614080
rect 41524 614076 41530 614078
rect 42517 614075 42583 614078
rect 41638 613396 41644 613460
rect 41708 613458 41714 613460
rect 41781 613458 41847 613461
rect 41708 613456 41847 613458
rect 41708 613400 41786 613456
rect 41842 613400 41847 613456
rect 41708 613398 41847 613400
rect 41708 613396 41714 613398
rect 41781 613395 41847 613398
rect 62113 611010 62179 611013
rect 62113 611008 64492 611010
rect 62113 610952 62118 611008
rect 62174 610952 64492 611008
rect 62113 610950 64492 610952
rect 62113 610947 62179 610950
rect 675385 606524 675451 606525
rect 675334 606522 675340 606524
rect 675294 606462 675340 606522
rect 675404 606520 675451 606524
rect 675446 606464 675451 606520
rect 675334 606460 675340 606462
rect 675404 606460 675451 606464
rect 675385 606459 675451 606460
rect 651557 603938 651623 603941
rect 650164 603936 651623 603938
rect 650164 603880 651562 603936
rect 651618 603880 651623 603936
rect 650164 603878 651623 603880
rect 651557 603875 651623 603878
rect 35801 601898 35867 601901
rect 35758 601896 35867 601898
rect 35758 601840 35806 601896
rect 35862 601840 35867 601896
rect 35758 601835 35867 601840
rect 35758 601732 35818 601835
rect 35801 601490 35867 601493
rect 35758 601488 35867 601490
rect 35758 601432 35806 601488
rect 35862 601432 35867 601488
rect 35758 601427 35867 601432
rect 35758 601324 35818 601427
rect 35709 601082 35775 601085
rect 35709 601080 35818 601082
rect 35709 601024 35714 601080
rect 35770 601024 35818 601080
rect 35709 601019 35818 601024
rect 35758 600916 35818 601019
rect 675201 600946 675267 600949
rect 675702 600946 675708 600948
rect 675201 600944 675708 600946
rect 675201 600888 675206 600944
rect 675262 600888 675708 600944
rect 675201 600886 675708 600888
rect 675201 600883 675267 600886
rect 675702 600884 675708 600886
rect 675772 600884 675778 600948
rect 35617 600674 35683 600677
rect 35574 600672 35683 600674
rect 35574 600616 35622 600672
rect 35678 600616 35683 600672
rect 35574 600611 35683 600616
rect 35574 600508 35634 600611
rect 44173 600130 44239 600133
rect 41492 600128 44239 600130
rect 41492 600072 44178 600128
rect 44234 600072 44239 600128
rect 41492 600070 44239 600072
rect 44173 600067 44239 600070
rect 44633 599722 44699 599725
rect 41492 599720 44699 599722
rect 41492 599664 44638 599720
rect 44694 599664 44699 599720
rect 41492 599662 44699 599664
rect 44633 599659 44699 599662
rect 42793 599314 42859 599317
rect 41492 599312 42859 599314
rect 41492 599256 42798 599312
rect 42854 599256 42859 599312
rect 41492 599254 42859 599256
rect 42793 599251 42859 599254
rect 39982 598980 39988 599044
rect 40052 598980 40058 599044
rect 675753 599042 675819 599045
rect 676806 599042 676812 599044
rect 675753 599040 676812 599042
rect 675753 598984 675758 599040
rect 675814 598984 676812 599040
rect 675753 598982 676812 598984
rect 39990 598876 40050 598980
rect 675753 598979 675819 598982
rect 676806 598980 676812 598982
rect 676876 598980 676882 599044
rect 39990 598228 40050 598468
rect 39982 598164 39988 598228
rect 40052 598164 40058 598228
rect 44725 598090 44791 598093
rect 41492 598088 44791 598090
rect 41492 598032 44730 598088
rect 44786 598032 44791 598088
rect 41492 598030 44791 598032
rect 44725 598027 44791 598030
rect 62113 597954 62179 597957
rect 62113 597952 64492 597954
rect 62113 597896 62118 597952
rect 62174 597896 64492 597952
rect 62113 597894 64492 597896
rect 62113 597891 62179 597894
rect 44265 597682 44331 597685
rect 41492 597680 44331 597682
rect 41492 597624 44270 597680
rect 44326 597624 44331 597680
rect 41492 597622 44331 597624
rect 44265 597619 44331 597622
rect 39254 597005 39314 597244
rect 39254 597000 39363 597005
rect 39254 596944 39302 597000
rect 39358 596944 39363 597000
rect 39254 596942 39363 596944
rect 39297 596939 39363 596942
rect 40910 596597 40970 596836
rect 40861 596592 40970 596597
rect 40861 596536 40866 596592
rect 40922 596536 40970 596592
rect 40861 596534 40970 596536
rect 40861 596531 40927 596534
rect 40726 596189 40786 596428
rect 40677 596184 40786 596189
rect 40677 596128 40682 596184
rect 40738 596128 40786 596184
rect 40677 596126 40786 596128
rect 40677 596123 40743 596126
rect 42057 596050 42123 596053
rect 41492 596048 42123 596050
rect 41492 595992 42062 596048
rect 42118 595992 42123 596048
rect 41492 595990 42123 595992
rect 42057 595987 42123 595990
rect 44357 595642 44423 595645
rect 41492 595640 44423 595642
rect 41492 595584 44362 595640
rect 44418 595584 44423 595640
rect 41492 595582 44423 595584
rect 44357 595579 44423 595582
rect 675569 595372 675635 595373
rect 675518 595370 675524 595372
rect 675478 595310 675524 595370
rect 675588 595368 675635 595372
rect 675630 595312 675635 595368
rect 675518 595308 675524 595310
rect 675588 595308 675635 595312
rect 675569 595307 675635 595308
rect 33734 594965 33794 595204
rect 31661 594962 31727 594965
rect 31661 594960 31770 594962
rect 31661 594904 31666 594960
rect 31722 594904 31770 594960
rect 31661 594899 31770 594904
rect 33734 594960 33843 594965
rect 33734 594904 33782 594960
rect 33838 594904 33843 594960
rect 33734 594902 33843 594904
rect 33777 594899 33843 594902
rect 31710 594796 31770 594899
rect 42885 594418 42951 594421
rect 41492 594416 42951 594418
rect 41492 594360 42890 594416
rect 42946 594360 42951 594416
rect 41492 594358 42951 594360
rect 42885 594355 42951 594358
rect 42149 594010 42215 594013
rect 41492 594008 42215 594010
rect 41492 593952 42154 594008
rect 42210 593952 42215 594008
rect 41492 593950 42215 593952
rect 42149 593947 42215 593950
rect 32446 593333 32506 593572
rect 32397 593328 32506 593333
rect 32397 593272 32402 593328
rect 32458 593272 32506 593328
rect 32397 593270 32506 593272
rect 32397 593267 32463 593270
rect 44633 593194 44699 593197
rect 675753 593196 675819 593197
rect 675702 593194 675708 593196
rect 41492 593192 44699 593194
rect 41492 593136 44638 593192
rect 44694 593136 44699 593192
rect 41492 593134 44699 593136
rect 675662 593134 675708 593194
rect 675772 593192 675819 593196
rect 675814 593136 675819 593192
rect 44633 593131 44699 593134
rect 675702 593132 675708 593134
rect 675772 593132 675819 593136
rect 675753 593131 675819 593132
rect 675569 593060 675635 593061
rect 675518 592996 675524 593060
rect 675588 593058 675635 593060
rect 675588 593056 675680 593058
rect 675630 593000 675680 593056
rect 675588 592998 675680 593000
rect 675588 592996 675635 592998
rect 675569 592995 675635 592996
rect 44449 592786 44515 592789
rect 41492 592784 44515 592786
rect 41492 592728 44454 592784
rect 44510 592728 44515 592784
rect 41492 592726 44515 592728
rect 44449 592723 44515 592726
rect 40542 592108 40602 592348
rect 40534 592044 40540 592108
rect 40604 592044 40610 592108
rect 675334 592044 675340 592108
rect 675404 592106 675410 592108
rect 675477 592106 675543 592109
rect 675404 592104 675543 592106
rect 675404 592048 675482 592104
rect 675538 592048 675543 592104
rect 675404 592046 675543 592048
rect 675404 592044 675410 592046
rect 675477 592043 675543 592046
rect 676990 592044 676996 592108
rect 677060 592106 677066 592108
rect 677501 592106 677567 592109
rect 677060 592104 677567 592106
rect 677060 592048 677506 592104
rect 677562 592048 677567 592104
rect 677060 592046 677567 592048
rect 677060 592044 677066 592046
rect 677501 592043 677567 592046
rect 40726 591700 40786 591940
rect 40718 591636 40724 591700
rect 40788 591636 40794 591700
rect 41462 591293 41522 591532
rect 676070 591364 676076 591428
rect 676140 591426 676146 591428
rect 682377 591426 682443 591429
rect 676140 591424 682443 591426
rect 676140 591368 682382 591424
rect 682438 591368 682443 591424
rect 676140 591366 682443 591368
rect 676140 591364 676146 591366
rect 682377 591363 682443 591366
rect 41462 591288 41571 591293
rect 41462 591232 41510 591288
rect 41566 591232 41571 591288
rect 41462 591230 41571 591232
rect 41505 591227 41571 591230
rect 30422 590716 30482 591124
rect 651557 590746 651623 590749
rect 650164 590744 651623 590746
rect 650164 590688 651562 590744
rect 651618 590688 651623 590744
rect 650164 590686 651623 590688
rect 651557 590683 651623 590686
rect 41462 590069 41522 590308
rect 41462 590064 41571 590069
rect 41462 590008 41510 590064
rect 41566 590008 41571 590064
rect 41462 590006 41571 590008
rect 41505 590003 41571 590006
rect 31661 587210 31727 587213
rect 41454 587210 41460 587212
rect 31661 587208 41460 587210
rect 31661 587152 31666 587208
rect 31722 587152 41460 587208
rect 31661 587150 41460 587152
rect 31661 587147 31727 587150
rect 41454 587148 41460 587150
rect 41524 587148 41530 587212
rect 675569 586258 675635 586261
rect 675702 586258 675708 586260
rect 675569 586256 675708 586258
rect 675569 586200 675574 586256
rect 675630 586200 675708 586256
rect 675569 586198 675708 586200
rect 675569 586195 675635 586198
rect 675702 586196 675708 586198
rect 675772 586196 675778 586260
rect 675845 586258 675911 586261
rect 676070 586258 676076 586260
rect 675845 586256 676076 586258
rect 675845 586200 675850 586256
rect 675906 586200 676076 586256
rect 675845 586198 676076 586200
rect 675845 586195 675911 586198
rect 676070 586196 676076 586198
rect 676140 586196 676146 586260
rect 40861 585444 40927 585445
rect 40861 585442 40908 585444
rect 40816 585440 40908 585442
rect 40816 585384 40866 585440
rect 40816 585382 40908 585384
rect 40861 585380 40908 585382
rect 40972 585380 40978 585444
rect 40861 585379 40927 585380
rect 39297 585170 39363 585173
rect 42374 585170 42380 585172
rect 39297 585168 42380 585170
rect 39297 585112 39302 585168
rect 39358 585112 42380 585168
rect 39297 585110 42380 585112
rect 39297 585107 39363 585110
rect 42374 585108 42380 585110
rect 42444 585108 42450 585172
rect 62113 584898 62179 584901
rect 62113 584896 64492 584898
rect 62113 584840 62118 584896
rect 62174 584840 64492 584896
rect 62113 584838 64492 584840
rect 62113 584835 62179 584838
rect 40677 584646 40743 584649
rect 42006 584646 42012 584648
rect 40677 584644 42012 584646
rect 40677 584588 40682 584644
rect 40738 584588 42012 584644
rect 40677 584586 42012 584588
rect 40677 584583 40743 584586
rect 42006 584584 42012 584586
rect 42076 584584 42082 584648
rect 675477 584626 675543 584629
rect 675886 584626 675892 584628
rect 675477 584624 675892 584626
rect 675477 584568 675482 584624
rect 675538 584568 675892 584624
rect 675477 584566 675892 584568
rect 675477 584563 675543 584566
rect 675886 584564 675892 584566
rect 675956 584564 675962 584628
rect 41597 584512 41663 584513
rect 41597 584510 41644 584512
rect 41552 584508 41644 584510
rect 41552 584452 41602 584508
rect 41552 584450 41644 584452
rect 41597 584448 41644 584450
rect 41708 584448 41714 584512
rect 41597 584447 41663 584448
rect 42149 584218 42215 584221
rect 42558 584218 42564 584220
rect 42149 584216 42564 584218
rect 42149 584160 42154 584216
rect 42210 584160 42564 584216
rect 42149 584158 42564 584160
rect 42149 584155 42215 584158
rect 42558 584156 42564 584158
rect 42628 584156 42634 584220
rect 40902 581708 40908 581772
rect 40972 581770 40978 581772
rect 41781 581770 41847 581773
rect 40972 581768 41847 581770
rect 40972 581712 41786 581768
rect 41842 581712 41847 581768
rect 40972 581710 41847 581712
rect 40972 581708 40978 581710
rect 41781 581707 41847 581710
rect 676029 581090 676095 581093
rect 676029 581088 676292 581090
rect 676029 581032 676034 581088
rect 676090 581032 676292 581088
rect 676029 581030 676292 581032
rect 676029 581027 676095 581030
rect 676121 580546 676187 580549
rect 676262 580546 676322 580652
rect 676121 580544 676322 580546
rect 676121 580488 676126 580544
rect 676182 580488 676322 580544
rect 676121 580486 676322 580488
rect 676121 580483 676187 580486
rect 41638 580212 41644 580276
rect 41708 580274 41714 580276
rect 41781 580274 41847 580277
rect 41708 580272 41847 580274
rect 41708 580216 41786 580272
rect 41842 580216 41847 580272
rect 41708 580214 41847 580216
rect 41708 580212 41714 580214
rect 41781 580211 41847 580214
rect 676029 580274 676095 580277
rect 676029 580272 676292 580274
rect 676029 580216 676034 580272
rect 676090 580216 676292 580272
rect 676029 580214 676292 580216
rect 676029 580211 676095 580214
rect 676213 580138 676279 580141
rect 676213 580136 676322 580138
rect 676213 580080 676218 580136
rect 676274 580080 676322 580136
rect 676213 580075 676322 580080
rect 676262 579836 676322 580075
rect 676262 579325 676322 579428
rect 676262 579320 676371 579325
rect 676262 579264 676310 579320
rect 676366 579264 676371 579320
rect 676262 579262 676371 579264
rect 676305 579259 676371 579262
rect 40718 578988 40724 579052
rect 40788 579050 40794 579052
rect 41781 579050 41847 579053
rect 40788 579048 41847 579050
rect 40788 578992 41786 579048
rect 41842 578992 41847 579048
rect 40788 578990 41847 578992
rect 40788 578988 40794 578990
rect 41781 578987 41847 578990
rect 676262 578917 676322 579020
rect 676213 578912 676322 578917
rect 676213 578856 676218 578912
rect 676274 578856 676322 578912
rect 676213 578854 676322 578856
rect 676213 578851 676279 578854
rect 676121 578506 676187 578509
rect 676262 578506 676322 578612
rect 676121 578504 676322 578506
rect 676121 578448 676126 578504
rect 676182 578448 676322 578504
rect 676121 578446 676322 578448
rect 676121 578443 676187 578446
rect 676029 578234 676095 578237
rect 676029 578232 676292 578234
rect 676029 578176 676034 578232
rect 676090 578176 676292 578232
rect 676029 578174 676292 578176
rect 676029 578171 676095 578174
rect 676262 577693 676322 577796
rect 676213 577688 676322 577693
rect 676213 577632 676218 577688
rect 676274 577632 676322 577688
rect 676213 577630 676322 577632
rect 676213 577627 676279 577630
rect 40534 577492 40540 577556
rect 40604 577554 40610 577556
rect 41781 577554 41847 577557
rect 40604 577552 41847 577554
rect 40604 577496 41786 577552
rect 41842 577496 41847 577552
rect 40604 577494 41847 577496
rect 40604 577492 40610 577494
rect 41781 577491 41847 577494
rect 651557 577418 651623 577421
rect 650164 577416 651623 577418
rect 650164 577360 651562 577416
rect 651618 577360 651623 577416
rect 650164 577358 651623 577360
rect 651557 577355 651623 577358
rect 676029 577418 676095 577421
rect 676029 577416 676292 577418
rect 676029 577360 676034 577416
rect 676090 577360 676292 577416
rect 676029 577358 676292 577360
rect 676029 577355 676095 577358
rect 676029 577010 676095 577013
rect 676029 577008 676292 577010
rect 676029 576952 676034 577008
rect 676090 576952 676292 577008
rect 676029 576950 676292 576952
rect 676029 576947 676095 576950
rect 676121 576466 676187 576469
rect 676262 576466 676322 576572
rect 676121 576464 676322 576466
rect 676121 576408 676126 576464
rect 676182 576408 676322 576464
rect 676121 576406 676322 576408
rect 676121 576403 676187 576406
rect 676262 576061 676322 576164
rect 676213 576056 676322 576061
rect 676213 576000 676218 576056
rect 676274 576000 676322 576056
rect 676213 575998 676322 576000
rect 676213 575995 676279 575998
rect 676029 575786 676095 575789
rect 676029 575784 676292 575786
rect 676029 575728 676034 575784
rect 676090 575728 676292 575784
rect 676029 575726 676292 575728
rect 676029 575723 676095 575726
rect 682377 575650 682443 575653
rect 682334 575648 682443 575650
rect 682334 575592 682382 575648
rect 682438 575592 682443 575648
rect 682334 575587 682443 575592
rect 682334 575348 682394 575587
rect 676029 574970 676095 574973
rect 676029 574968 676292 574970
rect 676029 574912 676034 574968
rect 676090 574912 676292 574968
rect 676029 574910 676292 574912
rect 676029 574907 676095 574910
rect 676262 574429 676322 574532
rect 676213 574424 676322 574429
rect 676213 574368 676218 574424
rect 676274 574368 676322 574424
rect 676213 574366 676322 574368
rect 676213 574363 676279 574366
rect 676029 574154 676095 574157
rect 676029 574152 676292 574154
rect 676029 574096 676034 574152
rect 676090 574096 676292 574152
rect 676029 574094 676292 574096
rect 676029 574091 676095 574094
rect 42333 574020 42399 574021
rect 42333 574018 42380 574020
rect 42288 574016 42380 574018
rect 42288 573960 42338 574016
rect 42288 573958 42380 573960
rect 42333 573956 42380 573958
rect 42444 573956 42450 574020
rect 42333 573955 42399 573956
rect 42149 573882 42215 573885
rect 42558 573882 42564 573884
rect 42149 573880 42564 573882
rect 42149 573824 42154 573880
rect 42210 573824 42564 573880
rect 42149 573822 42564 573824
rect 42149 573819 42215 573822
rect 42558 573820 42564 573822
rect 42628 573820 42634 573884
rect 676029 573746 676095 573749
rect 676029 573744 676292 573746
rect 676029 573688 676034 573744
rect 676090 573688 676292 573744
rect 676029 573686 676292 573688
rect 676029 573683 676095 573686
rect 677501 573610 677567 573613
rect 677501 573608 677610 573610
rect 677501 573552 677506 573608
rect 677562 573552 677610 573608
rect 677501 573547 677610 573552
rect 677550 573308 677610 573547
rect 677174 573140 677180 573204
rect 677244 573140 677250 573204
rect 677182 572900 677242 573140
rect 677358 572732 677364 572796
rect 677428 572732 677434 572796
rect 677366 572492 677426 572732
rect 676262 571981 676322 572084
rect 676213 571976 676322 571981
rect 676213 571920 676218 571976
rect 676274 571920 676322 571976
rect 676213 571918 676322 571920
rect 676213 571915 676279 571918
rect 62113 571842 62179 571845
rect 62113 571840 64492 571842
rect 62113 571784 62118 571840
rect 62174 571784 64492 571840
rect 62113 571782 64492 571784
rect 62113 571779 62179 571782
rect 676262 571573 676322 571676
rect 42006 571508 42012 571572
rect 42076 571570 42082 571572
rect 42701 571570 42767 571573
rect 42076 571568 42767 571570
rect 42076 571512 42706 571568
rect 42762 571512 42767 571568
rect 42076 571510 42767 571512
rect 42076 571508 42082 571510
rect 42701 571507 42767 571510
rect 676213 571568 676322 571573
rect 676213 571512 676218 571568
rect 676274 571512 676322 571568
rect 676213 571510 676322 571512
rect 676213 571507 676279 571510
rect 676262 571165 676322 571268
rect 676213 571160 676322 571165
rect 676213 571104 676218 571160
rect 676274 571104 676322 571160
rect 676213 571102 676322 571104
rect 676213 571099 676279 571102
rect 683070 570757 683130 570860
rect 683070 570752 683179 570757
rect 683070 570696 683118 570752
rect 683174 570696 683179 570752
rect 683070 570694 683179 570696
rect 683113 570691 683179 570694
rect 41454 570420 41460 570484
rect 41524 570482 41530 570484
rect 42149 570482 42215 570485
rect 41524 570480 42215 570482
rect 41524 570424 42154 570480
rect 42210 570424 42215 570480
rect 41524 570422 42215 570424
rect 41524 570420 41530 570422
rect 42149 570419 42215 570422
rect 685830 570044 685890 570452
rect 683113 569938 683179 569941
rect 683070 569936 683179 569938
rect 683070 569880 683118 569936
rect 683174 569880 683179 569936
rect 683070 569875 683179 569880
rect 683070 569636 683130 569875
rect 652109 564090 652175 564093
rect 650164 564088 652175 564090
rect 650164 564032 652114 564088
rect 652170 564032 652175 564088
rect 650164 564030 652175 564032
rect 652109 564027 652175 564030
rect 675753 562730 675819 562733
rect 676622 562730 676628 562732
rect 675753 562728 676628 562730
rect 675753 562672 675758 562728
rect 675814 562672 676628 562728
rect 675753 562670 676628 562672
rect 675753 562667 675819 562670
rect 676622 562668 676628 562670
rect 676692 562668 676698 562732
rect 675334 561172 675340 561236
rect 675404 561234 675410 561236
rect 675477 561234 675543 561237
rect 675404 561232 675543 561234
rect 675404 561176 675482 561232
rect 675538 561176 675543 561232
rect 675404 561174 675543 561176
rect 675404 561172 675410 561174
rect 675477 561171 675543 561174
rect 675569 559604 675635 559605
rect 675518 559602 675524 559604
rect 675478 559542 675524 559602
rect 675588 559600 675635 559604
rect 675630 559544 675635 559600
rect 675518 559540 675524 559542
rect 675588 559540 675635 559544
rect 675569 559539 675635 559540
rect 677174 559058 677180 559060
rect 675710 558998 677180 559058
rect 675710 558925 675770 558998
rect 677174 558996 677180 558998
rect 677244 558996 677250 559060
rect 675710 558920 675819 558925
rect 675710 558864 675758 558920
rect 675814 558864 675819 558920
rect 675710 558862 675819 558864
rect 675753 558859 675819 558862
rect 62113 558786 62179 558789
rect 62113 558784 64492 558786
rect 62113 558728 62118 558784
rect 62174 558728 64492 558784
rect 62113 558726 64492 558728
rect 62113 558723 62179 558726
rect 35758 558381 35818 558484
rect 35617 558378 35683 558381
rect 35574 558376 35683 558378
rect 35574 558320 35622 558376
rect 35678 558320 35683 558376
rect 35574 558315 35683 558320
rect 35758 558376 35867 558381
rect 35758 558320 35806 558376
rect 35862 558320 35867 558376
rect 35758 558318 35867 558320
rect 35801 558315 35867 558318
rect 35574 558076 35634 558315
rect 35709 557970 35775 557973
rect 35709 557968 35818 557970
rect 35709 557912 35714 557968
rect 35770 557912 35818 557968
rect 35709 557907 35818 557912
rect 35758 557668 35818 557907
rect 44173 557290 44239 557293
rect 41492 557288 44239 557290
rect 41492 557232 44178 557288
rect 44234 557232 44239 557288
rect 41492 557230 44239 557232
rect 44173 557227 44239 557230
rect 44633 556882 44699 556885
rect 41492 556880 44699 556882
rect 41492 556824 44638 556880
rect 44694 556824 44699 556880
rect 41492 556822 44699 556824
rect 44633 556819 44699 556822
rect 42793 556474 42859 556477
rect 41492 556472 42859 556474
rect 41492 556416 42798 556472
rect 42854 556416 42859 556472
rect 41492 556414 42859 556416
rect 42793 556411 42859 556414
rect 42793 556066 42859 556069
rect 41492 556064 42859 556066
rect 41492 556008 42798 556064
rect 42854 556008 42859 556064
rect 41492 556006 42859 556008
rect 42793 556003 42859 556006
rect 39982 555868 39988 555932
rect 40052 555868 40058 555932
rect 39990 555628 40050 555868
rect 44357 555250 44423 555253
rect 41492 555248 44423 555250
rect 41492 555192 44362 555248
rect 44418 555192 44423 555248
rect 41492 555190 44423 555192
rect 44357 555187 44423 555190
rect 44265 554842 44331 554845
rect 41492 554840 44331 554842
rect 41492 554784 44270 554840
rect 44326 554784 44331 554840
rect 41492 554782 44331 554784
rect 44265 554779 44331 554782
rect 674925 554842 674991 554845
rect 675518 554842 675524 554844
rect 674925 554840 675524 554842
rect 674925 554784 674930 554840
rect 674986 554784 675524 554840
rect 674925 554782 675524 554784
rect 674925 554779 674991 554782
rect 675518 554780 675524 554782
rect 675588 554780 675594 554844
rect 44265 554434 44331 554437
rect 41492 554432 44331 554434
rect 41492 554376 44270 554432
rect 44326 554376 44331 554432
rect 41492 554374 44331 554376
rect 44265 554371 44331 554374
rect 675753 554026 675819 554029
rect 677174 554026 677180 554028
rect 675753 554024 677180 554026
rect 40910 553893 40970 553996
rect 675753 553968 675758 554024
rect 675814 553968 677180 554024
rect 675753 553966 677180 553968
rect 675753 553963 675819 553966
rect 677174 553964 677180 553966
rect 677244 553964 677250 554028
rect 40861 553888 40970 553893
rect 40861 553832 40866 553888
rect 40922 553832 40970 553888
rect 40861 553830 40970 553832
rect 40861 553827 40927 553830
rect 40726 553485 40786 553588
rect 40677 553480 40786 553485
rect 40677 553424 40682 553480
rect 40738 553424 40786 553480
rect 40677 553422 40786 553424
rect 40677 553419 40743 553422
rect 40910 553077 40970 553180
rect 40910 553072 41019 553077
rect 40910 553016 40958 553072
rect 41014 553016 41019 553072
rect 40910 553014 41019 553016
rect 40953 553011 41019 553014
rect 32446 552669 32506 552772
rect 32397 552664 32506 552669
rect 32397 552608 32402 552664
rect 32458 552608 32506 552664
rect 32397 552606 32506 552608
rect 32397 552603 32463 552606
rect 40726 552261 40786 552364
rect 40726 552256 40835 552261
rect 40726 552200 40774 552256
rect 40830 552200 40835 552256
rect 40726 552198 40835 552200
rect 40769 552195 40835 552198
rect 675753 551986 675819 551989
rect 676990 551986 676996 551988
rect 675753 551984 676996 551986
rect 30974 551853 31034 551956
rect 675753 551928 675758 551984
rect 675814 551928 676996 551984
rect 675753 551926 676996 551928
rect 675753 551923 675819 551926
rect 676990 551924 676996 551926
rect 677060 551924 677066 551988
rect 30974 551848 31083 551853
rect 30974 551792 31022 551848
rect 31078 551792 31083 551848
rect 30974 551790 31083 551792
rect 31017 551787 31083 551790
rect 42885 551578 42951 551581
rect 41492 551576 42951 551578
rect 41492 551520 42890 551576
rect 42946 551520 42951 551576
rect 41492 551518 42951 551520
rect 42885 551515 42951 551518
rect 44449 551170 44515 551173
rect 41492 551168 44515 551170
rect 41492 551112 44454 551168
rect 44510 551112 44515 551168
rect 41492 551110 44515 551112
rect 44449 551107 44515 551110
rect 651557 550898 651623 550901
rect 650164 550896 651623 550898
rect 650164 550840 651562 550896
rect 651618 550840 651623 550896
rect 650164 550838 651623 550840
rect 651557 550835 651623 550838
rect 40726 550628 40786 550732
rect 40718 550564 40724 550628
rect 40788 550564 40794 550628
rect 44173 550354 44239 550357
rect 41492 550352 44239 550354
rect 41492 550296 44178 550352
rect 44234 550296 44239 550352
rect 41492 550294 44239 550296
rect 44173 550291 44239 550294
rect 675017 550354 675083 550357
rect 675334 550354 675340 550356
rect 675017 550352 675340 550354
rect 675017 550296 675022 550352
rect 675078 550296 675340 550352
rect 675017 550294 675340 550296
rect 675017 550291 675083 550294
rect 675334 550292 675340 550294
rect 675404 550292 675410 550356
rect 43069 549946 43135 549949
rect 41492 549944 43135 549946
rect 41492 549888 43074 549944
rect 43130 549888 43135 549944
rect 41492 549886 43135 549888
rect 43069 549883 43135 549886
rect 40542 549404 40602 549508
rect 40534 549340 40540 549404
rect 40604 549340 40610 549404
rect 40910 548996 40970 549100
rect 40902 548932 40908 548996
rect 40972 548932 40978 548996
rect 44541 548722 44607 548725
rect 41492 548720 44607 548722
rect 41492 548664 44546 548720
rect 44602 548664 44607 548720
rect 41492 548662 44607 548664
rect 44541 548659 44607 548662
rect 31710 548181 31770 548284
rect 31661 548176 31770 548181
rect 31661 548120 31666 548176
rect 31722 548120 31770 548176
rect 31661 548118 31770 548120
rect 31661 548115 31727 548118
rect 674373 548042 674439 548045
rect 674373 548040 674666 548042
rect 674373 547984 674378 548040
rect 674434 547984 674666 548040
rect 674373 547982 674666 547984
rect 674373 547979 674439 547982
rect 674606 547909 674666 547982
rect 674606 547904 674715 547909
rect 27662 547468 27722 547890
rect 674606 547848 674654 547904
rect 674710 547848 674715 547904
rect 674606 547846 674715 547848
rect 674649 547843 674715 547846
rect 35758 546957 35818 547060
rect 35758 546952 35867 546957
rect 35758 546896 35806 546952
rect 35862 546896 35867 546952
rect 35758 546894 35867 546896
rect 35801 546891 35867 546894
rect 675702 546756 675708 546820
rect 675772 546818 675778 546820
rect 678237 546818 678303 546821
rect 675772 546816 678303 546818
rect 675772 546760 678242 546816
rect 678298 546760 678303 546816
rect 675772 546758 678303 546760
rect 675772 546756 675778 546758
rect 678237 546755 678303 546758
rect 675886 546620 675892 546684
rect 675956 546682 675962 546684
rect 679617 546682 679683 546685
rect 675956 546680 679683 546682
rect 675956 546624 679622 546680
rect 679678 546624 679683 546680
rect 675956 546622 679683 546624
rect 675956 546620 675962 546622
rect 679617 546619 679683 546622
rect 676622 546484 676628 546548
rect 676692 546546 676698 546548
rect 677501 546546 677567 546549
rect 676692 546544 677567 546546
rect 676692 546488 677506 546544
rect 677562 546488 677567 546544
rect 676692 546486 677567 546488
rect 676692 546484 676698 546486
rect 677501 546483 677567 546486
rect 62113 545866 62179 545869
rect 62113 545864 64492 545866
rect 62113 545808 62118 545864
rect 62174 545808 64492 545864
rect 62113 545806 64492 545808
rect 62113 545803 62179 545806
rect 40861 545186 40927 545189
rect 41454 545186 41460 545188
rect 40861 545184 41460 545186
rect 40861 545128 40866 545184
rect 40922 545128 41460 545184
rect 40861 545126 41460 545128
rect 40861 545123 40927 545126
rect 41454 545124 41460 545126
rect 41524 545124 41530 545188
rect 676806 543628 676812 543692
rect 676876 543690 676882 543692
rect 683297 543690 683363 543693
rect 676876 543688 683363 543690
rect 676876 543632 683302 543688
rect 683358 543632 683363 543688
rect 676876 543630 683363 543632
rect 676876 543628 676882 543630
rect 683297 543627 683363 543630
rect 40953 543010 41019 543013
rect 41638 543010 41644 543012
rect 40953 543008 41644 543010
rect 40953 542952 40958 543008
rect 41014 542952 41644 543008
rect 40953 542950 41644 542952
rect 40953 542947 41019 542950
rect 41638 542948 41644 542950
rect 41708 542948 41714 543012
rect 676070 542948 676076 543012
rect 676140 543010 676146 543012
rect 678329 543010 678395 543013
rect 676140 543008 678395 543010
rect 676140 542952 678334 543008
rect 678390 542952 678395 543008
rect 676140 542950 678395 542952
rect 676140 542948 676146 542950
rect 678329 542947 678395 542950
rect 32397 542874 32463 542877
rect 41822 542874 41828 542876
rect 32397 542872 41828 542874
rect 32397 542816 32402 542872
rect 32458 542816 41828 542872
rect 32397 542814 41828 542816
rect 32397 542811 32463 542814
rect 41822 542812 41828 542814
rect 41892 542812 41898 542876
rect 40769 542330 40835 542333
rect 42006 542330 42012 542332
rect 40769 542328 42012 542330
rect 40769 542272 40774 542328
rect 40830 542272 42012 542328
rect 40769 542270 42012 542272
rect 40769 542267 40835 542270
rect 42006 542268 42012 542270
rect 42076 542268 42082 542332
rect 651557 537570 651623 537573
rect 650164 537568 651623 537570
rect 650164 537512 651562 537568
rect 651618 537512 651623 537568
rect 650164 537510 651623 537512
rect 651557 537507 651623 537510
rect 676262 535941 676322 536112
rect 42006 535876 42012 535940
rect 42076 535938 42082 535940
rect 42609 535938 42675 535941
rect 42076 535936 42675 535938
rect 42076 535880 42614 535936
rect 42670 535880 42675 535936
rect 42076 535878 42675 535880
rect 42076 535876 42082 535878
rect 42609 535875 42675 535878
rect 676213 535936 676322 535941
rect 676213 535880 676218 535936
rect 676274 535880 676322 535936
rect 676213 535878 676322 535880
rect 676213 535875 676279 535878
rect 676029 535734 676095 535737
rect 676029 535732 676292 535734
rect 676029 535676 676034 535732
rect 676090 535676 676292 535732
rect 676029 535674 676292 535676
rect 676029 535671 676095 535674
rect 676121 535122 676187 535125
rect 676262 535122 676322 535296
rect 676121 535120 676322 535122
rect 676121 535064 676126 535120
rect 676182 535064 676322 535120
rect 676121 535062 676322 535064
rect 676121 535059 676187 535062
rect 676262 534717 676322 534888
rect 676213 534712 676322 534717
rect 676213 534656 676218 534712
rect 676274 534656 676322 534712
rect 676213 534654 676322 534656
rect 676213 534651 676279 534654
rect 40902 534516 40908 534580
rect 40972 534578 40978 534580
rect 41781 534578 41847 534581
rect 40972 534576 41847 534578
rect 40972 534520 41786 534576
rect 41842 534520 41847 534576
rect 40972 534518 41847 534520
rect 40972 534516 40978 534518
rect 41781 534515 41847 534518
rect 675937 534510 676003 534513
rect 675937 534508 676292 534510
rect 675937 534452 675942 534508
rect 675998 534452 676292 534508
rect 675937 534450 676292 534452
rect 675937 534447 676003 534450
rect 676213 534306 676279 534309
rect 676213 534304 676322 534306
rect 676213 534248 676218 534304
rect 676274 534248 676322 534304
rect 676213 534243 676322 534248
rect 40718 534108 40724 534172
rect 40788 534170 40794 534172
rect 40788 534110 42626 534170
rect 40788 534108 40794 534110
rect 42566 533901 42626 534110
rect 676262 534072 676322 534243
rect 42566 533896 42675 533901
rect 42566 533840 42614 533896
rect 42670 533840 42675 533896
rect 42566 533838 42675 533840
rect 42609 533835 42675 533838
rect 683806 533493 683866 533664
rect 683806 533488 683915 533493
rect 683806 533432 683854 533488
rect 683910 533432 683915 533488
rect 683806 533430 683915 533432
rect 683849 533427 683915 533430
rect 676029 533286 676095 533289
rect 676029 533284 676292 533286
rect 676029 533228 676034 533284
rect 676090 533228 676292 533284
rect 676029 533226 676292 533228
rect 676029 533223 676095 533226
rect 676029 532878 676095 532881
rect 676029 532876 676292 532878
rect 676029 532820 676034 532876
rect 676090 532820 676292 532876
rect 676029 532818 676292 532820
rect 676029 532815 676095 532818
rect 62113 532810 62179 532813
rect 62113 532808 64492 532810
rect 62113 532752 62118 532808
rect 62174 532752 64492 532808
rect 62113 532750 64492 532752
rect 62113 532747 62179 532750
rect 41822 532612 41828 532676
rect 41892 532674 41898 532676
rect 42333 532674 42399 532677
rect 41892 532672 42399 532674
rect 41892 532616 42338 532672
rect 42394 532616 42399 532672
rect 41892 532614 42399 532616
rect 41892 532612 41898 532614
rect 42333 532611 42399 532614
rect 676213 532674 676279 532677
rect 676213 532672 676322 532674
rect 676213 532616 676218 532672
rect 676274 532616 676322 532672
rect 676213 532611 676322 532616
rect 676262 532440 676322 532611
rect 677182 531861 677242 532032
rect 677182 531856 677291 531861
rect 679617 531858 679683 531861
rect 677182 531800 677230 531856
rect 677286 531800 677291 531856
rect 677182 531798 677291 531800
rect 677225 531795 677291 531798
rect 679574 531856 679683 531858
rect 679574 531800 679622 531856
rect 679678 531800 679683 531856
rect 679574 531795 679683 531800
rect 679574 531624 679634 531795
rect 40534 531388 40540 531452
rect 40604 531450 40610 531452
rect 41781 531450 41847 531453
rect 40604 531448 41847 531450
rect 40604 531392 41786 531448
rect 41842 531392 41847 531448
rect 40604 531390 41847 531392
rect 40604 531388 40610 531390
rect 41781 531387 41847 531390
rect 678237 531450 678303 531453
rect 678237 531448 678346 531450
rect 678237 531392 678242 531448
rect 678298 531392 678346 531448
rect 678237 531387 678346 531392
rect 678286 531216 678346 531387
rect 676121 530634 676187 530637
rect 676262 530634 676322 530808
rect 678329 530634 678395 530637
rect 676121 530632 676322 530634
rect 676121 530576 676126 530632
rect 676182 530576 676322 530632
rect 676121 530574 676322 530576
rect 678286 530632 678395 530634
rect 678286 530576 678334 530632
rect 678390 530576 678395 530632
rect 676121 530571 676187 530574
rect 678286 530571 678395 530576
rect 678286 530400 678346 530571
rect 676213 530226 676279 530229
rect 676213 530224 676322 530226
rect 676213 530168 676218 530224
rect 676274 530168 676322 530224
rect 676213 530163 676322 530168
rect 676262 529992 676322 530163
rect 41454 529892 41460 529956
rect 41524 529954 41530 529956
rect 41524 529894 42258 529954
rect 41524 529892 41530 529894
rect 42198 529546 42258 529894
rect 42333 529546 42399 529549
rect 42198 529544 42399 529546
rect 42198 529488 42338 529544
rect 42394 529488 42399 529544
rect 42198 529486 42399 529488
rect 42333 529483 42399 529486
rect 41638 529348 41644 529412
rect 41708 529410 41714 529412
rect 42609 529410 42675 529413
rect 41708 529408 42675 529410
rect 41708 529352 42614 529408
rect 42670 529352 42675 529408
rect 41708 529350 42675 529352
rect 41708 529348 41714 529350
rect 42609 529347 42675 529350
rect 676121 529410 676187 529413
rect 676262 529410 676322 529584
rect 676121 529408 676322 529410
rect 676121 529352 676126 529408
rect 676182 529352 676322 529408
rect 676121 529350 676322 529352
rect 676121 529347 676187 529350
rect 676262 529005 676322 529176
rect 676213 529000 676322 529005
rect 676213 528944 676218 529000
rect 676274 528944 676322 529000
rect 676213 528942 676322 528944
rect 676397 529002 676463 529005
rect 676397 529000 676506 529002
rect 676397 528944 676402 529000
rect 676458 528944 676506 529000
rect 676213 528939 676279 528942
rect 676397 528939 676506 528944
rect 676446 528768 676506 528939
rect 675845 528390 675911 528393
rect 675845 528388 676292 528390
rect 675845 528332 675850 528388
rect 675906 528332 676292 528388
rect 675845 528330 676292 528332
rect 675845 528327 675911 528330
rect 676262 527781 676322 527952
rect 676213 527776 676322 527781
rect 683297 527778 683363 527781
rect 676213 527720 676218 527776
rect 676274 527720 676322 527776
rect 676213 527718 676322 527720
rect 683254 527776 683363 527778
rect 683254 527720 683302 527776
rect 683358 527720 683363 527776
rect 676213 527715 676279 527718
rect 683254 527715 683363 527720
rect 683254 527544 683314 527715
rect 675845 527166 675911 527169
rect 675845 527164 676292 527166
rect 675845 527108 675850 527164
rect 675906 527108 676292 527164
rect 675845 527106 676292 527108
rect 675845 527103 675911 527106
rect 676213 526962 676279 526965
rect 676213 526960 676322 526962
rect 676213 526904 676218 526960
rect 676274 526904 676322 526960
rect 676213 526899 676322 526904
rect 676262 526728 676322 526899
rect 676213 526554 676279 526557
rect 676213 526552 676322 526554
rect 676213 526496 676218 526552
rect 676274 526496 676322 526552
rect 676213 526491 676322 526496
rect 676262 526320 676322 526491
rect 683070 525741 683130 525912
rect 683070 525736 683179 525741
rect 683070 525680 683118 525736
rect 683174 525680 683179 525736
rect 683070 525678 683179 525680
rect 683113 525675 683179 525678
rect 685830 525096 685890 525504
rect 683113 524922 683179 524925
rect 683070 524920 683179 524922
rect 683070 524864 683118 524920
rect 683174 524864 683179 524920
rect 683070 524859 683179 524864
rect 683070 524688 683130 524859
rect 651557 524242 651623 524245
rect 650164 524240 651623 524242
rect 650164 524184 651562 524240
rect 651618 524184 651623 524240
rect 650164 524182 651623 524184
rect 651557 524179 651623 524182
rect 62113 519754 62179 519757
rect 62113 519752 64492 519754
rect 62113 519696 62118 519752
rect 62174 519696 64492 519752
rect 62113 519694 64492 519696
rect 62113 519691 62179 519694
rect 651557 511050 651623 511053
rect 650164 511048 651623 511050
rect 650164 510992 651562 511048
rect 651618 510992 651623 511048
rect 650164 510990 651623 510992
rect 651557 510987 651623 510990
rect 62113 506698 62179 506701
rect 62113 506696 64492 506698
rect 62113 506640 62118 506696
rect 62174 506640 64492 506696
rect 62113 506638 64492 506640
rect 62113 506635 62179 506638
rect 651557 497722 651623 497725
rect 650164 497720 651623 497722
rect 650164 497664 651562 497720
rect 651618 497664 651623 497720
rect 650164 497662 651623 497664
rect 651557 497659 651623 497662
rect 62113 493642 62179 493645
rect 62113 493640 64492 493642
rect 62113 493584 62118 493640
rect 62174 493584 64492 493640
rect 62113 493582 64492 493584
rect 62113 493579 62179 493582
rect 677409 492420 677475 492421
rect 677358 492418 677364 492420
rect 677318 492358 677364 492418
rect 677428 492416 677475 492420
rect 677470 492360 677475 492416
rect 677358 492356 677364 492358
rect 677428 492356 677475 492360
rect 677409 492355 677475 492356
rect 675845 492146 675911 492149
rect 675845 492144 676292 492146
rect 675845 492088 675850 492144
rect 675906 492088 676292 492144
rect 675845 492086 676292 492088
rect 675845 492083 675911 492086
rect 675937 491738 676003 491741
rect 675937 491736 676292 491738
rect 675937 491680 675942 491736
rect 675998 491680 676292 491736
rect 675937 491678 676292 491680
rect 675937 491675 676003 491678
rect 675937 491330 676003 491333
rect 675937 491328 676292 491330
rect 675937 491272 675942 491328
rect 675998 491272 676292 491328
rect 675937 491270 676292 491272
rect 675937 491267 676003 491270
rect 675753 490922 675819 490925
rect 675753 490920 676292 490922
rect 675753 490864 675758 490920
rect 675814 490864 676292 490920
rect 675753 490862 676292 490864
rect 675753 490859 675819 490862
rect 675937 490514 676003 490517
rect 675937 490512 676292 490514
rect 675937 490456 675942 490512
rect 675998 490456 676292 490512
rect 675937 490454 676292 490456
rect 675937 490451 676003 490454
rect 677366 489933 677426 490076
rect 677317 489928 677426 489933
rect 677317 489872 677322 489928
rect 677378 489872 677426 489928
rect 677317 489870 677426 489872
rect 677317 489867 677383 489870
rect 675845 489698 675911 489701
rect 675845 489696 676292 489698
rect 675845 489640 675850 489696
rect 675906 489640 676292 489696
rect 675845 489638 676292 489640
rect 675845 489635 675911 489638
rect 676029 489290 676095 489293
rect 676029 489288 676292 489290
rect 676029 489232 676034 489288
rect 676090 489232 676292 489288
rect 676029 489230 676292 489232
rect 676029 489227 676095 489230
rect 676029 488882 676095 488885
rect 676029 488880 676292 488882
rect 676029 488824 676034 488880
rect 676090 488824 676292 488880
rect 676029 488822 676292 488824
rect 676029 488819 676095 488822
rect 676029 488474 676095 488477
rect 676029 488472 676292 488474
rect 676029 488416 676034 488472
rect 676090 488416 676292 488472
rect 676029 488414 676292 488416
rect 676029 488411 676095 488414
rect 676029 488066 676095 488069
rect 676029 488064 676292 488066
rect 676029 488008 676034 488064
rect 676090 488008 676292 488064
rect 676029 488006 676292 488008
rect 676029 488003 676095 488006
rect 680997 487658 681063 487661
rect 680997 487656 681076 487658
rect 680997 487600 681002 487656
rect 681058 487600 681076 487656
rect 680997 487598 681076 487600
rect 680997 487595 681063 487598
rect 679709 487250 679775 487253
rect 679709 487248 679788 487250
rect 679709 487192 679714 487248
rect 679770 487192 679788 487248
rect 679709 487190 679788 487192
rect 679709 487187 679775 487190
rect 676029 486842 676095 486845
rect 676029 486840 676292 486842
rect 676029 486784 676034 486840
rect 676090 486784 676292 486840
rect 676029 486782 676292 486784
rect 676029 486779 676095 486782
rect 679617 486434 679683 486437
rect 679604 486432 679683 486434
rect 679604 486376 679622 486432
rect 679678 486376 679683 486432
rect 679604 486374 679683 486376
rect 679617 486371 679683 486374
rect 676029 486026 676095 486029
rect 676029 486024 676292 486026
rect 676029 485968 676034 486024
rect 676090 485968 676292 486024
rect 676029 485966 676292 485968
rect 676029 485963 676095 485966
rect 674741 485618 674807 485621
rect 674741 485616 676292 485618
rect 674741 485560 674746 485616
rect 674802 485560 676292 485616
rect 674741 485558 676292 485560
rect 674741 485555 674807 485558
rect 675937 485210 676003 485213
rect 675937 485208 676292 485210
rect 675937 485152 675942 485208
rect 675998 485152 676292 485208
rect 675937 485150 676292 485152
rect 675937 485147 676003 485150
rect 675937 484802 676003 484805
rect 675937 484800 676292 484802
rect 675937 484744 675942 484800
rect 675998 484744 676292 484800
rect 675937 484742 676292 484744
rect 675937 484739 676003 484742
rect 651557 484530 651623 484533
rect 650164 484528 651623 484530
rect 650164 484472 651562 484528
rect 651618 484472 651623 484528
rect 650164 484470 651623 484472
rect 651557 484467 651623 484470
rect 677409 484394 677475 484397
rect 677396 484392 677475 484394
rect 677396 484336 677414 484392
rect 677470 484336 677475 484392
rect 677396 484334 677475 484336
rect 677409 484331 677475 484334
rect 676070 484060 676076 484124
rect 676140 484060 676146 484124
rect 676078 483986 676138 484060
rect 676078 483926 676292 483986
rect 676070 483652 676076 483716
rect 676140 483652 676146 483716
rect 676078 483578 676138 483652
rect 676078 483518 676292 483578
rect 675937 483170 676003 483173
rect 675937 483168 676292 483170
rect 675937 483112 675942 483168
rect 675998 483112 676292 483168
rect 675937 483110 676292 483112
rect 675937 483107 676003 483110
rect 675937 482762 676003 482765
rect 675937 482760 676292 482762
rect 675937 482704 675942 482760
rect 675998 482704 676292 482760
rect 675937 482702 676292 482704
rect 675937 482699 676003 482702
rect 674649 482354 674715 482357
rect 674649 482352 676292 482354
rect 674649 482296 674654 482352
rect 674710 482296 676292 482352
rect 674649 482294 676292 482296
rect 674649 482291 674715 482294
rect 676078 481886 676292 481946
rect 676078 480722 676138 481886
rect 685830 481100 685890 481508
rect 678973 480722 679039 480725
rect 676078 480720 679166 480722
rect 676078 480664 678978 480720
rect 679034 480664 679166 480720
rect 676078 480662 679166 480664
rect 678973 480659 679039 480662
rect 62113 480586 62179 480589
rect 62113 480584 64492 480586
rect 62113 480528 62118 480584
rect 62174 480528 64492 480584
rect 62113 480526 64492 480528
rect 62113 480523 62179 480526
rect 672073 474874 672139 474877
rect 672942 474874 672948 474876
rect 672073 474872 672948 474874
rect 672073 474816 672078 474872
rect 672134 474816 672948 474872
rect 672073 474814 672948 474816
rect 672073 474811 672139 474814
rect 672942 474812 672948 474814
rect 673012 474812 673018 474876
rect 651649 471202 651715 471205
rect 650164 471200 651715 471202
rect 650164 471144 651654 471200
rect 651710 471144 651715 471200
rect 650164 471142 651715 471144
rect 651649 471139 651715 471142
rect 62113 467530 62179 467533
rect 62113 467528 64492 467530
rect 62113 467472 62118 467528
rect 62174 467472 64492 467528
rect 62113 467470 64492 467472
rect 62113 467467 62179 467470
rect 651557 457874 651623 457877
rect 650164 457872 651623 457874
rect 650164 457816 651562 457872
rect 651618 457816 651623 457872
rect 650164 457814 651623 457816
rect 651557 457811 651623 457814
rect 62113 454610 62179 454613
rect 62113 454608 64492 454610
rect 62113 454552 62118 454608
rect 62174 454552 64492 454608
rect 62113 454550 64492 454552
rect 62113 454547 62179 454550
rect 651557 444546 651623 444549
rect 650164 444544 651623 444546
rect 650164 444488 651562 444544
rect 651618 444488 651623 444544
rect 650164 444486 651623 444488
rect 651557 444483 651623 444486
rect 62113 441554 62179 441557
rect 62113 441552 64492 441554
rect 62113 441496 62118 441552
rect 62174 441496 64492 441552
rect 62113 441494 64492 441496
rect 62113 441491 62179 441494
rect 651557 431354 651623 431357
rect 650164 431352 651623 431354
rect 650164 431296 651562 431352
rect 651618 431296 651623 431352
rect 650164 431294 651623 431296
rect 651557 431291 651623 431294
rect 43161 430946 43227 430949
rect 41492 430944 43227 430946
rect 41492 430888 43166 430944
rect 43222 430888 43227 430944
rect 41492 430886 43227 430888
rect 43161 430883 43227 430886
rect 41781 430538 41847 430541
rect 41492 430536 41847 430538
rect 41492 430480 41786 430536
rect 41842 430480 41847 430536
rect 41492 430478 41847 430480
rect 41781 430475 41847 430478
rect 43621 430130 43687 430133
rect 41492 430128 43687 430130
rect 41492 430072 43626 430128
rect 43682 430072 43687 430128
rect 41492 430070 43687 430072
rect 43621 430067 43687 430070
rect 44633 429722 44699 429725
rect 41492 429720 44699 429722
rect 41492 429664 44638 429720
rect 44694 429664 44699 429720
rect 41492 429662 44699 429664
rect 44633 429659 44699 429662
rect 44173 429314 44239 429317
rect 41492 429312 44239 429314
rect 41492 429256 44178 429312
rect 44234 429256 44239 429312
rect 41492 429254 44239 429256
rect 44173 429251 44239 429254
rect 42793 428906 42859 428909
rect 41492 428904 42859 428906
rect 41492 428848 42798 428904
rect 42854 428848 42859 428904
rect 41492 428846 42859 428848
rect 42793 428843 42859 428846
rect 42793 428498 42859 428501
rect 41492 428496 42859 428498
rect 41492 428440 42798 428496
rect 42854 428440 42859 428496
rect 41492 428438 42859 428440
rect 42793 428435 42859 428438
rect 62113 428498 62179 428501
rect 62113 428496 64492 428498
rect 62113 428440 62118 428496
rect 62174 428440 64492 428496
rect 62113 428438 64492 428440
rect 62113 428435 62179 428438
rect 44357 428090 44423 428093
rect 41492 428088 44423 428090
rect 41492 428032 44362 428088
rect 44418 428032 44423 428088
rect 41492 428030 44423 428032
rect 44357 428027 44423 428030
rect 44357 427682 44423 427685
rect 41492 427680 44423 427682
rect 41492 427624 44362 427680
rect 44418 427624 44423 427680
rect 41492 427622 44423 427624
rect 44357 427619 44423 427622
rect 44265 427274 44331 427277
rect 41492 427272 44331 427274
rect 41492 427216 44270 427272
rect 44326 427216 44331 427272
rect 41492 427214 44331 427216
rect 44265 427211 44331 427214
rect 44541 426866 44607 426869
rect 41492 426864 44607 426866
rect 41492 426808 44546 426864
rect 44602 426808 44607 426864
rect 41492 426806 44607 426808
rect 44541 426803 44607 426806
rect 41822 426458 41828 426460
rect 41492 426398 41828 426458
rect 41822 426396 41828 426398
rect 41892 426396 41898 426460
rect 32397 426050 32463 426053
rect 32397 426048 32476 426050
rect 32397 425992 32402 426048
rect 32458 425992 32476 426048
rect 32397 425990 32476 425992
rect 32397 425987 32463 425990
rect 41822 425642 41828 425644
rect 41492 425582 41828 425642
rect 41822 425580 41828 425582
rect 41892 425580 41898 425644
rect 35157 425234 35223 425237
rect 35157 425232 35236 425234
rect 35157 425176 35162 425232
rect 35218 425176 35236 425232
rect 35157 425174 35236 425176
rect 35157 425171 35223 425174
rect 42190 424826 42196 424828
rect 41492 424766 42196 424826
rect 42190 424764 42196 424766
rect 42260 424764 42266 424828
rect 32489 424418 32555 424421
rect 32476 424416 32555 424418
rect 32476 424360 32494 424416
rect 32550 424360 32555 424416
rect 32476 424358 32555 424360
rect 32489 424355 32555 424358
rect 41822 424010 41828 424012
rect 41492 423950 41828 424010
rect 41822 423948 41828 423950
rect 41892 423948 41898 424012
rect 42006 423602 42012 423604
rect 41492 423542 42012 423602
rect 42006 423540 42012 423542
rect 42076 423540 42082 423604
rect 42885 423194 42951 423197
rect 41492 423192 42951 423194
rect 41492 423136 42890 423192
rect 42946 423136 42951 423192
rect 41492 423134 42951 423136
rect 42885 423131 42951 423134
rect 41822 422786 41828 422788
rect 41492 422726 41828 422786
rect 41822 422724 41828 422726
rect 41892 422724 41898 422788
rect 31017 422378 31083 422381
rect 31004 422376 31083 422378
rect 31004 422320 31022 422376
rect 31078 422320 31083 422376
rect 31004 422318 31083 422320
rect 31017 422315 31083 422318
rect 44449 421970 44515 421973
rect 41492 421968 44515 421970
rect 41492 421912 44454 421968
rect 44510 421912 44515 421968
rect 41492 421910 44515 421912
rect 44449 421907 44515 421910
rect 42977 421562 43043 421565
rect 41492 421560 43043 421562
rect 41492 421504 42982 421560
rect 43038 421504 43043 421560
rect 41492 421502 43043 421504
rect 42977 421499 43043 421502
rect 44633 421154 44699 421157
rect 41492 421152 44699 421154
rect 41492 421096 44638 421152
rect 44694 421096 44699 421152
rect 41492 421094 44699 421096
rect 44633 421091 44699 421094
rect 40049 420678 40055 420742
rect 40119 420740 40125 420742
rect 40119 420680 40158 420740
rect 40119 420678 40125 420680
rect 21774 419900 21834 420308
rect 41781 419522 41847 419525
rect 41492 419520 41847 419522
rect 40049 419450 40055 419514
rect 40119 419450 40125 419514
rect 41492 419464 41786 419520
rect 41842 419464 41847 419520
rect 41492 419462 41847 419464
rect 41781 419459 41847 419462
rect 651557 418026 651623 418029
rect 650164 418024 651623 418026
rect 650164 417968 651562 418024
rect 651618 417968 651623 418024
rect 650164 417966 651623 417968
rect 651557 417963 651623 417966
rect 62113 415442 62179 415445
rect 62113 415440 64492 415442
rect 62113 415384 62118 415440
rect 62174 415384 64492 415440
rect 62113 415382 64492 415384
rect 62113 415379 62179 415382
rect 41822 415244 41828 415308
rect 41892 415244 41898 415308
rect 41830 415034 41890 415244
rect 42006 415034 42012 415036
rect 41830 414974 42012 415034
rect 42006 414972 42012 414974
rect 42076 414972 42082 415036
rect 35157 414762 35223 414765
rect 41454 414762 41460 414764
rect 35157 414760 41460 414762
rect 35157 414704 35162 414760
rect 35218 414704 41460 414760
rect 35157 414702 41460 414704
rect 35157 414699 35223 414702
rect 41454 414700 41460 414702
rect 41524 414700 41530 414764
rect 32397 414626 32463 414629
rect 41822 414626 41828 414628
rect 32397 414624 41828 414626
rect 32397 414568 32402 414624
rect 32458 414568 41828 414624
rect 32397 414566 41828 414568
rect 32397 414563 32463 414566
rect 41822 414564 41828 414566
rect 41892 414564 41898 414628
rect 41873 411228 41939 411229
rect 41822 411226 41828 411228
rect 41782 411166 41828 411226
rect 41892 411224 41939 411228
rect 41934 411168 41939 411224
rect 41822 411164 41828 411166
rect 41892 411164 41939 411168
rect 41873 411163 41939 411164
rect 41086 409396 41092 409460
rect 41156 409458 41162 409460
rect 41781 409458 41847 409461
rect 41156 409456 41847 409458
rect 41156 409400 41786 409456
rect 41842 409400 41847 409456
rect 41156 409398 41847 409400
rect 41156 409396 41162 409398
rect 41781 409395 41847 409398
rect 41638 406268 41644 406332
rect 41708 406330 41714 406332
rect 41781 406330 41847 406333
rect 41708 406328 41847 406330
rect 41708 406272 41786 406328
rect 41842 406272 41847 406328
rect 41708 406270 41847 406272
rect 41708 406268 41714 406270
rect 41781 406267 41847 406270
rect 652017 404698 652083 404701
rect 650164 404696 652083 404698
rect 650164 404640 652022 404696
rect 652078 404640 652083 404696
rect 650164 404638 652083 404640
rect 652017 404635 652083 404638
rect 676262 403749 676322 403852
rect 676262 403744 676371 403749
rect 676262 403688 676310 403744
rect 676366 403688 676371 403744
rect 676262 403686 676371 403688
rect 676305 403683 676371 403686
rect 676262 403341 676322 403444
rect 676213 403336 676322 403341
rect 676213 403280 676218 403336
rect 676274 403280 676322 403336
rect 676213 403278 676322 403280
rect 676397 403338 676463 403341
rect 676397 403336 676506 403338
rect 676397 403280 676402 403336
rect 676458 403280 676506 403336
rect 676213 403275 676279 403278
rect 676397 403275 676506 403280
rect 676446 403036 676506 403275
rect 676121 402930 676187 402933
rect 676121 402928 676322 402930
rect 676121 402872 676126 402928
rect 676182 402872 676322 402928
rect 676121 402870 676322 402872
rect 676121 402867 676187 402870
rect 676262 402628 676322 402870
rect 42057 402524 42123 402525
rect 42006 402522 42012 402524
rect 41966 402462 42012 402522
rect 42076 402520 42123 402524
rect 42118 402464 42123 402520
rect 42006 402460 42012 402462
rect 42076 402460 42123 402464
rect 42057 402459 42123 402460
rect 62113 402386 62179 402389
rect 62113 402384 64492 402386
rect 62113 402328 62118 402384
rect 62174 402328 64492 402384
rect 62113 402326 64492 402328
rect 62113 402323 62179 402326
rect 676262 402117 676322 402220
rect 676213 402112 676322 402117
rect 676213 402056 676218 402112
rect 676274 402056 676322 402112
rect 676213 402054 676322 402056
rect 676213 402051 676279 402054
rect 41454 401780 41460 401844
rect 41524 401842 41530 401844
rect 41781 401842 41847 401845
rect 41524 401840 41847 401842
rect 41524 401784 41786 401840
rect 41842 401784 41847 401840
rect 41524 401782 41847 401784
rect 41524 401780 41530 401782
rect 41781 401779 41847 401782
rect 676029 401842 676095 401845
rect 676029 401840 676292 401842
rect 676029 401784 676034 401840
rect 676090 401784 676292 401840
rect 676029 401782 676292 401784
rect 676029 401779 676095 401782
rect 676262 401301 676322 401404
rect 676213 401296 676322 401301
rect 676213 401240 676218 401296
rect 676274 401240 676322 401296
rect 676213 401238 676322 401240
rect 677317 401298 677383 401301
rect 677317 401296 677426 401298
rect 677317 401240 677322 401296
rect 677378 401240 677426 401296
rect 676213 401235 676279 401238
rect 677317 401235 677426 401240
rect 677366 400996 677426 401235
rect 674741 400618 674807 400621
rect 674741 400616 676292 400618
rect 674741 400560 674746 400616
rect 674802 400560 676292 400616
rect 674741 400558 676292 400560
rect 674741 400555 674807 400558
rect 677225 400482 677291 400485
rect 677182 400480 677291 400482
rect 677182 400424 677230 400480
rect 677286 400424 677291 400480
rect 677182 400419 677291 400424
rect 677182 400180 677242 400419
rect 40534 400012 40540 400076
rect 40604 400074 40610 400076
rect 41781 400074 41847 400077
rect 40604 400072 41847 400074
rect 40604 400016 41786 400072
rect 41842 400016 41847 400072
rect 40604 400014 41847 400016
rect 40604 400012 40610 400014
rect 41781 400011 41847 400014
rect 676262 399669 676322 399772
rect 40902 399604 40908 399668
rect 40972 399666 40978 399668
rect 41781 399666 41847 399669
rect 40972 399664 41847 399666
rect 40972 399608 41786 399664
rect 41842 399608 41847 399664
rect 40972 399606 41847 399608
rect 40972 399604 40978 399606
rect 41781 399603 41847 399606
rect 676213 399664 676322 399669
rect 676213 399608 676218 399664
rect 676274 399608 676322 399664
rect 676213 399606 676322 399608
rect 676213 399603 676279 399606
rect 675886 399332 675892 399396
rect 675956 399394 675962 399396
rect 675956 399334 676292 399394
rect 675956 399332 675962 399334
rect 40718 398788 40724 398852
rect 40788 398850 40794 398852
rect 41781 398850 41847 398853
rect 676262 398852 676322 398956
rect 40788 398848 41847 398850
rect 40788 398792 41786 398848
rect 41842 398792 41847 398848
rect 40788 398790 41847 398792
rect 40788 398788 40794 398790
rect 41781 398787 41847 398790
rect 676254 398788 676260 398852
rect 676324 398788 676330 398852
rect 676029 398578 676095 398581
rect 676029 398576 676292 398578
rect 676029 398520 676034 398576
rect 676090 398520 676292 398576
rect 676029 398518 676292 398520
rect 676029 398515 676095 398518
rect 676029 398170 676095 398173
rect 676029 398168 676292 398170
rect 676029 398112 676034 398168
rect 676090 398112 676292 398168
rect 676029 398110 676292 398112
rect 676029 398107 676095 398110
rect 676814 397629 676874 397732
rect 676814 397624 676923 397629
rect 676814 397568 676862 397624
rect 676918 397568 676923 397624
rect 676814 397566 676923 397568
rect 676857 397563 676923 397566
rect 676446 397220 676506 397324
rect 676438 397156 676444 397220
rect 676508 397156 676514 397220
rect 676998 396813 677058 396916
rect 676949 396808 677058 396813
rect 676949 396752 676954 396808
rect 677010 396752 677058 396808
rect 676949 396750 677058 396752
rect 676949 396747 677015 396750
rect 678286 396405 678346 396508
rect 678286 396400 678395 396405
rect 678286 396344 678334 396400
rect 678390 396344 678395 396400
rect 678286 396342 678395 396344
rect 678329 396339 678395 396342
rect 678286 395997 678346 396100
rect 678237 395992 678346 395997
rect 678237 395936 678242 395992
rect 678298 395936 678346 395992
rect 678237 395934 678346 395936
rect 678237 395931 678303 395934
rect 676446 395589 676506 395692
rect 676397 395584 676506 395589
rect 676397 395528 676402 395584
rect 676458 395528 676506 395584
rect 676397 395526 676506 395528
rect 676397 395523 676463 395526
rect 676070 395116 676076 395180
rect 676140 395178 676146 395180
rect 676262 395178 676322 395284
rect 676140 395118 676322 395178
rect 676140 395116 676146 395118
rect 676446 394773 676506 394876
rect 676446 394768 676555 394773
rect 676446 394712 676494 394768
rect 676550 394712 676555 394768
rect 676446 394710 676555 394712
rect 676489 394707 676555 394710
rect 676262 394365 676322 394468
rect 676213 394360 676322 394365
rect 676213 394304 676218 394360
rect 676274 394304 676322 394360
rect 676213 394302 676322 394304
rect 676213 394299 676279 394302
rect 676262 393957 676322 394060
rect 676213 393952 676322 393957
rect 676213 393896 676218 393952
rect 676274 393896 676322 393952
rect 676213 393894 676322 393896
rect 676213 393891 676279 393894
rect 683070 393549 683130 393652
rect 683070 393544 683179 393549
rect 683070 393488 683118 393544
rect 683174 393488 683179 393544
rect 683070 393486 683179 393488
rect 683113 393483 683179 393486
rect 685830 392836 685890 393244
rect 683070 392325 683130 392428
rect 683070 392320 683179 392325
rect 683070 392264 683118 392320
rect 683174 392264 683179 392320
rect 683070 392262 683179 392264
rect 683113 392259 683179 392262
rect 651557 391506 651623 391509
rect 650164 391504 651623 391506
rect 650164 391448 651562 391504
rect 651618 391448 651623 391504
rect 650164 391446 651623 391448
rect 651557 391443 651623 391446
rect 62113 389330 62179 389333
rect 62113 389328 64492 389330
rect 62113 389272 62118 389328
rect 62174 389272 64492 389328
rect 62113 389270 64492 389272
rect 62113 389267 62179 389270
rect 675518 388452 675524 388516
rect 675588 388514 675594 388516
rect 676857 388514 676923 388517
rect 675588 388512 676923 388514
rect 675588 388456 676862 388512
rect 676918 388456 676923 388512
rect 675588 388454 676923 388456
rect 675588 388452 675594 388454
rect 676857 388451 676923 388454
rect 35758 387565 35818 387668
rect 675702 387636 675708 387700
rect 675772 387698 675778 387700
rect 676397 387698 676463 387701
rect 675772 387696 676463 387698
rect 675772 387640 676402 387696
rect 676458 387640 676463 387696
rect 675772 387638 676463 387640
rect 675772 387636 675778 387638
rect 676397 387635 676463 387638
rect 35758 387560 35867 387565
rect 35758 387504 35806 387560
rect 35862 387504 35867 387560
rect 35758 387502 35867 387504
rect 35801 387499 35867 387502
rect 675334 387500 675340 387564
rect 675404 387562 675410 387564
rect 678329 387562 678395 387565
rect 675404 387560 678395 387562
rect 675404 387504 678334 387560
rect 678390 387504 678395 387560
rect 675404 387502 678395 387504
rect 675404 387500 675410 387502
rect 678329 387499 678395 387502
rect 35758 387157 35818 387260
rect 35617 387154 35683 387157
rect 35574 387152 35683 387154
rect 35574 387096 35622 387152
rect 35678 387096 35683 387152
rect 35574 387091 35683 387096
rect 35758 387152 35867 387157
rect 35758 387096 35806 387152
rect 35862 387096 35867 387152
rect 35758 387094 35867 387096
rect 35801 387091 35867 387094
rect 35574 386852 35634 387091
rect 35709 386746 35775 386749
rect 35709 386744 35818 386746
rect 35709 386688 35714 386744
rect 35770 386688 35818 386744
rect 35709 386683 35818 386688
rect 35758 386444 35818 386683
rect 44633 386066 44699 386069
rect 41492 386064 44699 386066
rect 41492 386008 44638 386064
rect 44694 386008 44699 386064
rect 41492 386006 44699 386008
rect 44633 386003 44699 386006
rect 42793 385658 42859 385661
rect 41492 385656 42859 385658
rect 41492 385600 42798 385656
rect 42854 385600 42859 385656
rect 41492 385598 42859 385600
rect 42793 385595 42859 385598
rect 44173 385250 44239 385253
rect 41492 385248 44239 385250
rect 41492 385192 44178 385248
rect 44234 385192 44239 385248
rect 41492 385190 44239 385192
rect 44173 385187 44239 385190
rect 675753 384978 675819 384981
rect 675886 384978 675892 384980
rect 675753 384976 675892 384978
rect 675753 384920 675758 384976
rect 675814 384920 675892 384976
rect 675753 384918 675892 384920
rect 675753 384915 675819 384918
rect 675886 384916 675892 384918
rect 675956 384916 675962 384980
rect 44357 384842 44423 384845
rect 41492 384840 44423 384842
rect 41492 384784 44362 384840
rect 44418 384784 44423 384840
rect 41492 384782 44423 384784
rect 44357 384779 44423 384782
rect 44725 384434 44791 384437
rect 41492 384432 44791 384434
rect 41492 384376 44730 384432
rect 44786 384376 44791 384432
rect 41492 384374 44791 384376
rect 44725 384371 44791 384374
rect 44541 384026 44607 384029
rect 41492 384024 44607 384026
rect 41492 383968 44546 384024
rect 44602 383968 44607 384024
rect 41492 383966 44607 383968
rect 44541 383963 44607 383966
rect 42793 383618 42859 383621
rect 41492 383616 42859 383618
rect 41492 383560 42798 383616
rect 42854 383560 42859 383616
rect 41492 383558 42859 383560
rect 42793 383555 42859 383558
rect 40726 383076 40786 383180
rect 40718 383012 40724 383076
rect 40788 383012 40794 383076
rect 40910 382669 40970 382772
rect 40861 382664 40970 382669
rect 40861 382608 40866 382664
rect 40922 382608 40970 382664
rect 40861 382606 40970 382608
rect 40861 382603 40927 382606
rect 40542 382260 40602 382364
rect 675385 382260 675451 382261
rect 40534 382196 40540 382260
rect 40604 382196 40610 382260
rect 675334 382258 675340 382260
rect 675294 382198 675340 382258
rect 675404 382256 675451 382260
rect 675446 382200 675451 382256
rect 675334 382196 675340 382198
rect 675404 382196 675451 382200
rect 675385 382195 675451 382196
rect 41462 381852 41522 381956
rect 41454 381788 41460 381852
rect 41524 381788 41530 381852
rect 37966 381445 38026 381548
rect 37917 381440 38026 381445
rect 37917 381384 37922 381440
rect 37978 381384 38026 381440
rect 37917 381382 38026 381384
rect 37917 381379 37983 381382
rect 30974 381037 31034 381140
rect 30974 381032 31083 381037
rect 30974 380976 31022 381032
rect 31078 380976 31083 381032
rect 30974 380974 31083 380976
rect 31017 380971 31083 380974
rect 43161 380762 43227 380765
rect 41492 380760 43227 380762
rect 41492 380704 43166 380760
rect 43222 380704 43227 380760
rect 41492 380702 43227 380704
rect 43161 380699 43227 380702
rect 42977 380354 43043 380357
rect 41492 380352 43043 380354
rect 41492 380296 42982 380352
rect 43038 380296 43043 380352
rect 41492 380294 43043 380296
rect 42977 380291 43043 380294
rect 40910 379812 40970 379916
rect 40902 379748 40908 379812
rect 40972 379748 40978 379812
rect 40726 379405 40786 379508
rect 40677 379400 40786 379405
rect 40677 379344 40682 379400
rect 40738 379344 40786 379400
rect 40677 379342 40786 379344
rect 40677 379339 40743 379342
rect 44449 379130 44515 379133
rect 41492 379128 44515 379130
rect 41492 379072 44454 379128
rect 44510 379072 44515 379128
rect 41492 379070 44515 379072
rect 44449 379067 44515 379070
rect 43069 378722 43135 378725
rect 41492 378720 43135 378722
rect 41492 378664 43074 378720
rect 43130 378664 43135 378720
rect 41492 378662 43135 378664
rect 43069 378659 43135 378662
rect 675477 378724 675543 378725
rect 675477 378720 675524 378724
rect 675588 378722 675594 378724
rect 675477 378664 675482 378720
rect 675477 378660 675524 378664
rect 675588 378662 675634 378722
rect 675588 378660 675594 378662
rect 675477 378659 675543 378660
rect 33734 378181 33794 378284
rect 33734 378176 33843 378181
rect 651557 378178 651623 378181
rect 33734 378120 33782 378176
rect 33838 378120 33843 378176
rect 33734 378118 33843 378120
rect 650164 378176 651623 378178
rect 650164 378120 651562 378176
rect 651618 378120 651623 378176
rect 650164 378118 651623 378120
rect 33777 378115 33843 378118
rect 651557 378115 651623 378118
rect 44541 377906 44607 377909
rect 41492 377904 44607 377906
rect 41492 377848 44546 377904
rect 44602 377848 44607 377904
rect 41492 377846 44607 377848
rect 44541 377843 44607 377846
rect 675753 377634 675819 377637
rect 676070 377634 676076 377636
rect 675753 377632 676076 377634
rect 675753 377576 675758 377632
rect 675814 377576 676076 377632
rect 675753 377574 676076 377576
rect 675753 377571 675819 377574
rect 676070 377572 676076 377574
rect 676140 377572 676146 377636
rect 35758 377365 35818 377468
rect 35758 377360 35867 377365
rect 35758 377304 35806 377360
rect 35862 377304 35867 377360
rect 35758 377302 35867 377304
rect 35801 377299 35867 377302
rect 27662 376652 27722 377060
rect 62113 376274 62179 376277
rect 62113 376272 64492 376274
rect 41462 376141 41522 376244
rect 62113 376216 62118 376272
rect 62174 376216 64492 376272
rect 62113 376214 64492 376216
rect 62113 376211 62179 376214
rect 41462 376136 41571 376141
rect 41462 376080 41510 376136
rect 41566 376080 41571 376136
rect 41462 376078 41571 376080
rect 41505 376075 41571 376078
rect 675753 375460 675819 375461
rect 675702 375458 675708 375460
rect 675662 375398 675708 375458
rect 675772 375456 675819 375460
rect 675814 375400 675819 375456
rect 675702 375396 675708 375398
rect 675772 375396 675819 375400
rect 675753 375395 675819 375396
rect 675753 373690 675819 373693
rect 676254 373690 676260 373692
rect 675753 373688 676260 373690
rect 675753 373632 675758 373688
rect 675814 373632 676260 373688
rect 675753 373630 676260 373632
rect 675753 373627 675819 373630
rect 676254 373628 676260 373630
rect 676324 373628 676330 373692
rect 675753 372058 675819 372061
rect 676438 372058 676444 372060
rect 675753 372056 676444 372058
rect 675753 372000 675758 372056
rect 675814 372000 676444 372056
rect 675753 371998 676444 372000
rect 675753 371995 675819 371998
rect 676438 371996 676444 371998
rect 676508 371996 676514 372060
rect 33777 371922 33843 371925
rect 42006 371922 42012 371924
rect 33777 371920 42012 371922
rect 33777 371864 33782 371920
rect 33838 371864 42012 371920
rect 33777 371862 42012 371864
rect 33777 371859 33843 371862
rect 42006 371860 42012 371862
rect 42076 371860 42082 371924
rect 37917 371378 37983 371381
rect 41638 371378 41644 371380
rect 37917 371376 41644 371378
rect 37917 371320 37922 371376
rect 37978 371320 41644 371376
rect 37917 371318 41644 371320
rect 37917 371315 37983 371318
rect 41638 371316 41644 371318
rect 41708 371316 41714 371380
rect 41781 370292 41847 370293
rect 41781 370290 41828 370292
rect 41736 370288 41828 370290
rect 41736 370232 41786 370288
rect 41736 370230 41828 370232
rect 41781 370228 41828 370230
rect 41892 370228 41898 370292
rect 41781 370227 41847 370228
rect 41873 366348 41939 366349
rect 41822 366346 41828 366348
rect 41782 366286 41828 366346
rect 41892 366344 41939 366348
rect 41934 366288 41939 366344
rect 41822 366284 41828 366286
rect 41892 366284 41939 366288
rect 41873 366283 41939 366284
rect 652017 364850 652083 364853
rect 650164 364848 652083 364850
rect 650164 364792 652022 364848
rect 652078 364792 652083 364848
rect 650164 364790 652083 364792
rect 652017 364787 652083 364790
rect 41965 363764 42031 363765
rect 41965 363760 42012 363764
rect 42076 363762 42082 363764
rect 41965 363704 41970 363760
rect 41965 363700 42012 363704
rect 42076 363702 42122 363762
rect 42076 363700 42082 363702
rect 41965 363699 42031 363700
rect 62113 363354 62179 363357
rect 62113 363352 64492 363354
rect 62113 363296 62118 363352
rect 62174 363296 64492 363352
rect 62113 363294 64492 363296
rect 62113 363291 62179 363294
rect 41638 362884 41644 362948
rect 41708 362946 41714 362948
rect 41781 362946 41847 362949
rect 41708 362944 41847 362946
rect 41708 362888 41786 362944
rect 41842 362888 41847 362944
rect 41708 362886 41847 362888
rect 41708 362884 41714 362886
rect 41781 362883 41847 362886
rect 40902 360164 40908 360228
rect 40972 360226 40978 360228
rect 40972 360166 41706 360226
rect 40972 360164 40978 360166
rect 41646 360090 41706 360166
rect 41781 360090 41847 360093
rect 41646 360088 41847 360090
rect 41646 360032 41786 360088
rect 41842 360032 41847 360088
rect 41646 360030 41847 360032
rect 41781 360027 41847 360030
rect 41454 358668 41460 358732
rect 41524 358730 41530 358732
rect 41781 358730 41847 358733
rect 41524 358728 41847 358730
rect 41524 358672 41786 358728
rect 41842 358672 41847 358728
rect 41524 358670 41847 358672
rect 41524 358668 41530 358670
rect 41781 358667 41847 358670
rect 675845 358730 675911 358733
rect 675845 358728 676292 358730
rect 675845 358672 675850 358728
rect 675906 358672 676292 358728
rect 675845 358670 676292 358672
rect 675845 358667 675911 358670
rect 675937 358322 676003 358325
rect 675937 358320 676292 358322
rect 675937 358264 675942 358320
rect 675998 358264 676292 358320
rect 675937 358262 676292 358264
rect 675937 358259 676003 358262
rect 676029 357914 676095 357917
rect 676029 357912 676292 357914
rect 676029 357856 676034 357912
rect 676090 357856 676292 357912
rect 676029 357854 676292 357856
rect 676029 357851 676095 357854
rect 676029 357506 676095 357509
rect 676029 357504 676292 357506
rect 676029 357448 676034 357504
rect 676090 357448 676292 357504
rect 676029 357446 676292 357448
rect 676029 357443 676095 357446
rect 676029 357098 676095 357101
rect 676029 357096 676292 357098
rect 676029 357040 676034 357096
rect 676090 357040 676292 357096
rect 676029 357038 676292 357040
rect 676029 357035 676095 357038
rect 40718 356900 40724 356964
rect 40788 356962 40794 356964
rect 41781 356962 41847 356965
rect 40788 356960 41847 356962
rect 40788 356904 41786 356960
rect 41842 356904 41847 356960
rect 40788 356902 41847 356904
rect 40788 356900 40794 356902
rect 41781 356899 41847 356902
rect 676029 356690 676095 356693
rect 676029 356688 676292 356690
rect 676029 356632 676034 356688
rect 676090 356632 676292 356688
rect 676029 356630 676292 356632
rect 676029 356627 676095 356630
rect 676029 356282 676095 356285
rect 676029 356280 676292 356282
rect 676029 356224 676034 356280
rect 676090 356224 676292 356280
rect 676029 356222 676292 356224
rect 676029 356219 676095 356222
rect 674741 355874 674807 355877
rect 674741 355872 676292 355874
rect 674741 355816 674746 355872
rect 674802 355816 676292 355872
rect 674741 355814 676292 355816
rect 674741 355811 674807 355814
rect 40534 355676 40540 355740
rect 40604 355738 40610 355740
rect 41781 355738 41847 355741
rect 40604 355736 41847 355738
rect 40604 355680 41786 355736
rect 41842 355680 41847 355736
rect 40604 355678 41847 355680
rect 40604 355676 40610 355678
rect 41781 355675 41847 355678
rect 674741 355466 674807 355469
rect 674741 355464 676292 355466
rect 674741 355408 674746 355464
rect 674802 355408 676292 355464
rect 674741 355406 676292 355408
rect 674741 355403 674807 355406
rect 676029 355058 676095 355061
rect 676029 355056 676292 355058
rect 676029 355000 676034 355056
rect 676090 355000 676292 355056
rect 676029 354998 676292 355000
rect 676029 354995 676095 354998
rect 676029 354650 676095 354653
rect 676029 354648 676292 354650
rect 676029 354592 676034 354648
rect 676090 354592 676292 354648
rect 676029 354590 676292 354592
rect 676029 354587 676095 354590
rect 675518 354180 675524 354244
rect 675588 354242 675594 354244
rect 675588 354182 676292 354242
rect 675588 354180 675594 354182
rect 676078 353774 676292 353834
rect 676078 353700 676138 353774
rect 676070 353636 676076 353700
rect 676140 353636 676146 353700
rect 675334 353364 675340 353428
rect 675404 353426 675410 353428
rect 675404 353366 676292 353426
rect 675404 353364 675410 353366
rect 675886 352956 675892 353020
rect 675956 353018 675962 353020
rect 675956 352958 676292 353018
rect 675956 352956 675962 352958
rect 678237 352610 678303 352613
rect 678237 352608 678316 352610
rect 678237 352552 678242 352608
rect 678298 352552 678316 352608
rect 678237 352550 678316 352552
rect 678237 352547 678303 352550
rect 676078 352142 676292 352202
rect 676078 352068 676138 352142
rect 676070 352004 676076 352068
rect 676140 352004 676146 352068
rect 676029 351794 676095 351797
rect 676029 351792 676292 351794
rect 676029 351736 676034 351792
rect 676090 351736 676292 351792
rect 676029 351734 676292 351736
rect 676029 351731 676095 351734
rect 651557 351658 651623 351661
rect 650164 351656 651623 351658
rect 650164 351600 651562 351656
rect 651618 351600 651623 351656
rect 650164 351598 651623 351600
rect 651557 351595 651623 351598
rect 676814 351150 676874 351356
rect 676806 351086 676812 351150
rect 676876 351086 676882 351150
rect 676029 350978 676095 350981
rect 676029 350976 676292 350978
rect 676029 350920 676034 350976
rect 676090 350920 676292 350976
rect 676029 350918 676292 350920
rect 676029 350915 676095 350918
rect 676029 350570 676095 350573
rect 676029 350568 676292 350570
rect 676029 350512 676034 350568
rect 676090 350512 676292 350568
rect 676029 350510 676292 350512
rect 676029 350507 676095 350510
rect 62113 350298 62179 350301
rect 62113 350296 64492 350298
rect 62113 350240 62118 350296
rect 62174 350240 64492 350296
rect 62113 350238 64492 350240
rect 62113 350235 62179 350238
rect 675937 350162 676003 350165
rect 675937 350160 676292 350162
rect 675937 350104 675942 350160
rect 675998 350104 676292 350160
rect 675937 350102 676292 350104
rect 675937 350099 676003 350102
rect 676029 349754 676095 349757
rect 676029 349752 676292 349754
rect 676029 349696 676034 349752
rect 676090 349696 676292 349752
rect 676029 349694 676292 349696
rect 676029 349691 676095 349694
rect 676029 349346 676095 349349
rect 676029 349344 676292 349346
rect 676029 349288 676034 349344
rect 676090 349288 676292 349344
rect 676029 349286 676292 349288
rect 676029 349283 676095 349286
rect 676029 348938 676095 348941
rect 676029 348936 676292 348938
rect 676029 348880 676034 348936
rect 676090 348880 676292 348936
rect 676029 348878 676292 348880
rect 676029 348875 676095 348878
rect 676029 348530 676095 348533
rect 676029 348528 676292 348530
rect 676029 348472 676034 348528
rect 676090 348472 676292 348528
rect 676029 348470 676292 348472
rect 676029 348467 676095 348470
rect 676262 347684 676322 348092
rect 676029 347306 676095 347309
rect 676029 347304 676292 347306
rect 676029 347248 676034 347304
rect 676090 347248 676292 347304
rect 676029 347246 676292 347248
rect 676029 347243 676095 347246
rect 675937 346626 676003 346629
rect 676622 346626 676628 346628
rect 675937 346624 676628 346626
rect 675937 346568 675942 346624
rect 675998 346568 676628 346624
rect 675937 346566 676628 346568
rect 675937 346563 676003 346566
rect 676622 346564 676628 346566
rect 676692 346564 676698 346628
rect 676121 346490 676187 346493
rect 677174 346490 677180 346492
rect 676121 346488 677180 346490
rect 676121 346432 676126 346488
rect 676182 346432 677180 346488
rect 676121 346430 677180 346432
rect 676121 346427 676187 346430
rect 677174 346428 677180 346430
rect 677244 346428 677250 346492
rect 27613 344722 27679 344725
rect 27613 344720 27722 344722
rect 27613 344664 27618 344720
rect 27674 344664 27722 344720
rect 27613 344659 27722 344664
rect 27662 344556 27722 344659
rect 35801 344314 35867 344317
rect 35758 344312 35867 344314
rect 35758 344256 35806 344312
rect 35862 344256 35867 344312
rect 35758 344251 35867 344256
rect 35758 344148 35818 344251
rect 35709 343906 35775 343909
rect 35709 343904 35818 343906
rect 35709 343848 35714 343904
rect 35770 343848 35818 343904
rect 35709 343843 35818 343848
rect 35758 343740 35818 343843
rect 675518 343572 675524 343636
rect 675588 343634 675594 343636
rect 678237 343634 678303 343637
rect 675588 343632 678303 343634
rect 675588 343576 678242 343632
rect 678298 343576 678303 343632
rect 675588 343574 678303 343576
rect 675588 343572 675594 343574
rect 678237 343571 678303 343574
rect 44633 343362 44699 343365
rect 41492 343360 44699 343362
rect 41492 343304 44638 343360
rect 44694 343304 44699 343360
rect 41492 343302 44699 343304
rect 44633 343299 44699 343302
rect 44265 342954 44331 342957
rect 41492 342952 44331 342954
rect 41492 342896 44270 342952
rect 44326 342896 44331 342952
rect 41492 342894 44331 342896
rect 44265 342891 44331 342894
rect 44173 342546 44239 342549
rect 41492 342544 44239 342546
rect 41492 342488 44178 342544
rect 44234 342488 44239 342544
rect 41492 342486 44239 342488
rect 44173 342483 44239 342486
rect 675293 342274 675359 342277
rect 676857 342274 676923 342277
rect 675293 342272 676923 342274
rect 675293 342216 675298 342272
rect 675354 342216 676862 342272
rect 676918 342216 676923 342272
rect 675293 342214 676923 342216
rect 675293 342211 675359 342214
rect 676857 342211 676923 342214
rect 44541 342138 44607 342141
rect 41492 342136 44607 342138
rect 41492 342080 44546 342136
rect 44602 342080 44607 342136
rect 41492 342078 44607 342080
rect 44541 342075 44607 342078
rect 44725 341730 44791 341733
rect 41492 341728 44791 341730
rect 41492 341672 44730 341728
rect 44786 341672 44791 341728
rect 41492 341670 44791 341672
rect 44725 341667 44791 341670
rect 42885 341322 42951 341325
rect 41492 341320 42951 341322
rect 41492 341264 42890 341320
rect 42946 341264 42951 341320
rect 41492 341262 42951 341264
rect 42885 341259 42951 341262
rect 42793 340914 42859 340917
rect 41492 340912 42859 340914
rect 41492 340856 42798 340912
rect 42854 340856 42859 340912
rect 41492 340854 42859 340856
rect 42793 340851 42859 340854
rect 675661 340780 675727 340781
rect 675661 340776 675708 340780
rect 675772 340778 675778 340780
rect 675661 340720 675666 340776
rect 675661 340716 675708 340720
rect 675772 340718 675818 340778
rect 675772 340716 675778 340718
rect 675661 340715 675727 340716
rect 42793 340506 42859 340509
rect 41492 340504 42859 340506
rect 41492 340448 42798 340504
rect 42854 340448 42859 340504
rect 41492 340446 42859 340448
rect 42793 340443 42859 340446
rect 40726 339828 40786 340068
rect 40718 339764 40724 339828
rect 40788 339764 40794 339828
rect 30974 339421 31034 339660
rect 30974 339416 31083 339421
rect 30974 339360 31022 339416
rect 31078 339360 31083 339416
rect 30974 339358 31083 339360
rect 31017 339355 31083 339358
rect 675753 339418 675819 339421
rect 675886 339418 675892 339420
rect 675753 339416 675892 339418
rect 675753 339360 675758 339416
rect 675814 339360 675892 339416
rect 675753 339358 675892 339360
rect 675753 339355 675819 339358
rect 675886 339356 675892 339358
rect 675956 339356 675962 339420
rect 40542 339012 40602 339252
rect 40534 338948 40540 339012
rect 40604 338948 40610 339012
rect 42006 338874 42012 338876
rect 41492 338814 42012 338874
rect 42006 338812 42012 338814
rect 42076 338812 42082 338876
rect 32446 338197 32506 338436
rect 651649 338330 651715 338333
rect 650164 338328 651715 338330
rect 650164 338272 651654 338328
rect 651710 338272 651715 338328
rect 650164 338270 651715 338272
rect 651649 338267 651715 338270
rect 32397 338192 32506 338197
rect 32397 338136 32402 338192
rect 32458 338136 32506 338192
rect 32397 338134 32506 338136
rect 32397 338131 32463 338134
rect 44173 338058 44239 338061
rect 41492 338056 44239 338058
rect 41492 338000 44178 338056
rect 44234 338000 44239 338056
rect 41492 337998 44239 338000
rect 44173 337995 44239 337998
rect 675753 337922 675819 337925
rect 676070 337922 676076 337924
rect 675753 337920 676076 337922
rect 675753 337864 675758 337920
rect 675814 337864 676076 337920
rect 675753 337862 676076 337864
rect 675753 337859 675819 337862
rect 676070 337860 676076 337862
rect 676140 337860 676146 337924
rect 40910 337380 40970 337620
rect 40902 337316 40908 337380
rect 40972 337316 40978 337380
rect 62113 337242 62179 337245
rect 62113 337240 64492 337242
rect 41462 336970 41522 337212
rect 62113 337184 62118 337240
rect 62174 337184 64492 337240
rect 62113 337182 64492 337184
rect 62113 337179 62179 337182
rect 41638 336970 41644 336972
rect 41462 336910 41644 336970
rect 41638 336908 41644 336910
rect 41708 336908 41714 336972
rect 42977 336834 43043 336837
rect 41492 336832 43043 336834
rect 41492 336776 42982 336832
rect 43038 336776 43043 336832
rect 41492 336774 43043 336776
rect 42977 336771 43043 336774
rect 44357 336426 44423 336429
rect 41492 336424 44423 336426
rect 41492 336368 44362 336424
rect 44418 336368 44423 336424
rect 41492 336366 44423 336368
rect 44357 336363 44423 336366
rect 41278 335748 41338 335988
rect 675753 335882 675819 335885
rect 676990 335882 676996 335884
rect 675753 335880 676996 335882
rect 675753 335824 675758 335880
rect 675814 335824 676996 335880
rect 675753 335822 676996 335824
rect 675753 335819 675819 335822
rect 676990 335820 676996 335822
rect 677060 335820 677066 335884
rect 41270 335684 41276 335748
rect 41340 335684 41346 335748
rect 41094 335340 41154 335580
rect 41086 335276 41092 335340
rect 41156 335276 41162 335340
rect 674833 335338 674899 335341
rect 676806 335338 676812 335340
rect 674833 335336 676812 335338
rect 674833 335280 674838 335336
rect 674894 335280 676812 335336
rect 674833 335278 676812 335280
rect 674833 335275 674899 335278
rect 676806 335276 676812 335278
rect 676876 335276 676882 335340
rect 43069 335202 43135 335205
rect 41492 335200 43135 335202
rect 41492 335144 43074 335200
rect 43130 335144 43135 335200
rect 41492 335142 43135 335144
rect 43069 335139 43135 335142
rect 44449 334794 44515 334797
rect 41492 334792 44515 334794
rect 41492 334736 44454 334792
rect 44510 334736 44515 334792
rect 41492 334734 44515 334736
rect 44449 334731 44515 334734
rect 30422 334117 30482 334356
rect 30373 334112 30482 334117
rect 30373 334056 30378 334112
rect 30434 334056 30482 334112
rect 30373 334054 30482 334056
rect 30373 334051 30439 334054
rect 30422 333540 30482 333948
rect 675477 333572 675543 333573
rect 675477 333568 675524 333572
rect 675588 333570 675594 333572
rect 675477 333512 675482 333568
rect 675477 333508 675524 333512
rect 675588 333510 675634 333570
rect 675588 333508 675594 333510
rect 675477 333507 675543 333508
rect 30373 333298 30439 333301
rect 30373 333296 30482 333298
rect 30373 333240 30378 333296
rect 30434 333240 30482 333296
rect 30373 333235 30482 333240
rect 30422 333132 30482 333235
rect 676622 332618 676628 332620
rect 675710 332558 676628 332618
rect 675710 332213 675770 332558
rect 676622 332556 676628 332558
rect 676692 332556 676698 332620
rect 675710 332208 675819 332213
rect 675710 332152 675758 332208
rect 675814 332152 675819 332208
rect 675710 332150 675819 332152
rect 675753 332147 675819 332150
rect 32397 327858 32463 327861
rect 41454 327858 41460 327860
rect 32397 327856 41460 327858
rect 32397 327800 32402 327856
rect 32458 327800 41460 327856
rect 32397 327798 41460 327800
rect 32397 327795 32463 327798
rect 41454 327796 41460 327798
rect 41524 327796 41530 327860
rect 31017 327722 31083 327725
rect 41822 327722 41828 327724
rect 31017 327720 41828 327722
rect 31017 327664 31022 327720
rect 31078 327664 41828 327720
rect 31017 327662 41828 327664
rect 31017 327659 31083 327662
rect 41822 327660 41828 327662
rect 41892 327660 41898 327724
rect 675109 325682 675175 325685
rect 676438 325682 676444 325684
rect 675109 325680 676444 325682
rect 675109 325624 675114 325680
rect 675170 325624 676444 325680
rect 675109 325622 676444 325624
rect 675109 325619 675175 325622
rect 676438 325620 676444 325622
rect 676508 325620 676514 325684
rect 675753 325546 675819 325549
rect 676254 325546 676260 325548
rect 675753 325544 676260 325546
rect 675753 325488 675758 325544
rect 675814 325488 676260 325544
rect 675753 325486 676260 325488
rect 675753 325483 675819 325486
rect 676254 325484 676260 325486
rect 676324 325484 676330 325548
rect 651557 325002 651623 325005
rect 650164 325000 651623 325002
rect 650164 324944 651562 325000
rect 651618 324944 651623 325000
rect 650164 324942 651623 324944
rect 651557 324939 651623 324942
rect 41781 324868 41847 324869
rect 41781 324864 41828 324868
rect 41892 324866 41898 324868
rect 41781 324808 41786 324864
rect 41781 324804 41828 324808
rect 41892 324806 41938 324866
rect 41892 324804 41898 324806
rect 41781 324803 41847 324804
rect 62113 324186 62179 324189
rect 62113 324184 64492 324186
rect 62113 324128 62118 324184
rect 62174 324128 64492 324184
rect 62113 324126 64492 324128
rect 62113 324123 62179 324126
rect 41270 321132 41276 321196
rect 41340 321194 41346 321196
rect 41781 321194 41847 321197
rect 41340 321192 41847 321194
rect 41340 321136 41786 321192
rect 41842 321136 41847 321192
rect 41340 321134 41847 321136
rect 41340 321132 41346 321134
rect 41781 321131 41847 321134
rect 41454 319908 41460 319972
rect 41524 319970 41530 319972
rect 41781 319970 41847 319973
rect 41524 319968 41847 319970
rect 41524 319912 41786 319968
rect 41842 319912 41847 319968
rect 41524 319910 41847 319912
rect 41524 319908 41530 319910
rect 41781 319907 41847 319910
rect 41086 317324 41092 317388
rect 41156 317386 41162 317388
rect 41781 317386 41847 317389
rect 41156 317384 41847 317386
rect 41156 317328 41786 317384
rect 41842 317328 41847 317384
rect 41156 317326 41847 317328
rect 41156 317324 41162 317326
rect 41781 317323 41847 317326
rect 41638 315828 41644 315892
rect 41708 315890 41714 315892
rect 41781 315890 41847 315893
rect 41708 315888 41847 315890
rect 41708 315832 41786 315888
rect 41842 315832 41847 315888
rect 41708 315830 41847 315832
rect 41708 315828 41714 315830
rect 41781 315827 41847 315830
rect 41965 315484 42031 315485
rect 41965 315480 42012 315484
rect 42076 315482 42082 315484
rect 41965 315424 41970 315480
rect 41965 315420 42012 315424
rect 42076 315422 42122 315482
rect 42076 315420 42082 315422
rect 41965 315419 42031 315420
rect 40718 313788 40724 313852
rect 40788 313850 40794 313852
rect 41873 313850 41939 313853
rect 40788 313848 41939 313850
rect 40788 313792 41878 313848
rect 41934 313792 41939 313848
rect 40788 313790 41939 313792
rect 40788 313788 40794 313790
rect 41873 313787 41939 313790
rect 676029 313714 676095 313717
rect 676029 313712 676292 313714
rect 676029 313656 676034 313712
rect 676090 313656 676292 313712
rect 676029 313654 676292 313656
rect 676029 313651 676095 313654
rect 676213 313578 676279 313581
rect 676213 313576 676322 313578
rect 676213 313520 676218 313576
rect 676274 313520 676322 313576
rect 676213 313515 676322 313520
rect 676262 313276 676322 313515
rect 40902 313108 40908 313172
rect 40972 313170 40978 313172
rect 41781 313170 41847 313173
rect 40972 313168 41847 313170
rect 40972 313112 41786 313168
rect 41842 313112 41847 313168
rect 40972 313110 41847 313112
rect 40972 313108 40978 313110
rect 41781 313107 41847 313110
rect 676121 312762 676187 312765
rect 676262 312762 676322 312868
rect 676121 312760 676322 312762
rect 676121 312704 676126 312760
rect 676182 312704 676322 312760
rect 676121 312702 676322 312704
rect 676121 312699 676187 312702
rect 676262 312357 676322 312460
rect 40534 312292 40540 312356
rect 40604 312354 40610 312356
rect 41781 312354 41847 312357
rect 40604 312352 41847 312354
rect 40604 312296 41786 312352
rect 41842 312296 41847 312352
rect 40604 312294 41847 312296
rect 40604 312292 40610 312294
rect 41781 312291 41847 312294
rect 676213 312352 676322 312357
rect 676213 312296 676218 312352
rect 676274 312296 676322 312352
rect 676213 312294 676322 312296
rect 676213 312291 676279 312294
rect 676262 311949 676322 312052
rect 676213 311944 676322 311949
rect 676213 311888 676218 311944
rect 676274 311888 676322 311944
rect 676213 311886 676322 311888
rect 676213 311883 676279 311886
rect 651557 311810 651623 311813
rect 650164 311808 651623 311810
rect 650164 311752 651562 311808
rect 651618 311752 651623 311808
rect 650164 311750 651623 311752
rect 651557 311747 651623 311750
rect 676262 311541 676322 311644
rect 676213 311536 676322 311541
rect 676213 311480 676218 311536
rect 676274 311480 676322 311536
rect 676213 311478 676322 311480
rect 676213 311475 676279 311478
rect 62113 311130 62179 311133
rect 676121 311130 676187 311133
rect 676262 311130 676322 311236
rect 62113 311128 64492 311130
rect 62113 311072 62118 311128
rect 62174 311072 64492 311128
rect 62113 311070 64492 311072
rect 676121 311128 676322 311130
rect 676121 311072 676126 311128
rect 676182 311072 676322 311128
rect 676121 311070 676322 311072
rect 62113 311067 62179 311070
rect 676121 311067 676187 311070
rect 674741 310858 674807 310861
rect 674741 310856 676292 310858
rect 674741 310800 674746 310856
rect 674802 310800 676292 310856
rect 674741 310798 676292 310800
rect 674741 310795 674807 310798
rect 676262 310317 676322 310420
rect 676213 310312 676322 310317
rect 676213 310256 676218 310312
rect 676274 310256 676322 310312
rect 676213 310254 676322 310256
rect 676213 310251 676279 310254
rect 676029 310042 676095 310045
rect 676029 310040 676292 310042
rect 676029 309984 676034 310040
rect 676090 309984 676292 310040
rect 676029 309982 676292 309984
rect 676029 309979 676095 309982
rect 676262 309501 676322 309604
rect 676213 309496 676322 309501
rect 676213 309440 676218 309496
rect 676274 309440 676322 309496
rect 676213 309438 676322 309440
rect 676213 309435 676279 309438
rect 679574 309093 679634 309196
rect 679574 309088 679683 309093
rect 679574 309032 679622 309088
rect 679678 309032 679683 309088
rect 679574 309030 679683 309032
rect 679617 309027 679683 309030
rect 676446 308684 676506 308788
rect 676438 308620 676444 308684
rect 676508 308620 676514 308684
rect 678286 308277 678346 308380
rect 678237 308272 678346 308277
rect 678237 308216 678242 308272
rect 678298 308216 678346 308272
rect 678237 308214 678346 308216
rect 678237 308211 678303 308214
rect 675886 307940 675892 308004
rect 675956 308002 675962 308004
rect 675956 307942 676292 308002
rect 675956 307940 675962 307942
rect 679758 307461 679818 307564
rect 679709 307456 679818 307461
rect 679709 307400 679714 307456
rect 679770 307400 679818 307456
rect 679709 307398 679818 307400
rect 679709 307395 679775 307398
rect 676262 307052 676322 307156
rect 676254 306988 676260 307052
rect 676324 306988 676330 307052
rect 676814 306645 676874 306748
rect 676814 306640 676923 306645
rect 676814 306584 676862 306640
rect 676918 306584 676923 306640
rect 676814 306582 676923 306584
rect 676857 306579 676923 306582
rect 676446 306237 676506 306340
rect 676397 306232 676506 306237
rect 676397 306176 676402 306232
rect 676458 306176 676506 306232
rect 676397 306174 676506 306176
rect 676397 306171 676463 306174
rect 676446 305829 676506 305932
rect 676446 305824 676555 305829
rect 676446 305768 676494 305824
rect 676550 305768 676555 305824
rect 676446 305766 676555 305768
rect 676489 305763 676555 305766
rect 676070 305356 676076 305420
rect 676140 305418 676146 305420
rect 676262 305418 676322 305524
rect 676140 305358 676322 305418
rect 676140 305356 676146 305358
rect 676630 305012 676690 305116
rect 676622 304948 676628 305012
rect 676692 304948 676698 305012
rect 676262 304605 676322 304708
rect 676262 304600 676371 304605
rect 676262 304544 676310 304600
rect 676366 304544 676371 304600
rect 676262 304542 676371 304544
rect 676305 304539 676371 304542
rect 676121 304194 676187 304197
rect 676262 304194 676322 304300
rect 676121 304192 676322 304194
rect 676121 304136 676126 304192
rect 676182 304136 676322 304192
rect 676121 304134 676322 304136
rect 676121 304131 676187 304134
rect 676262 303789 676322 303892
rect 676213 303784 676322 303789
rect 676213 303728 676218 303784
rect 676274 303728 676322 303784
rect 676213 303726 676322 303728
rect 676213 303723 676279 303726
rect 683070 303381 683130 303484
rect 683070 303376 683179 303381
rect 683070 303320 683118 303376
rect 683174 303320 683179 303376
rect 683070 303318 683179 303320
rect 683113 303315 683179 303318
rect 685830 302668 685890 303076
rect 683113 302562 683179 302565
rect 683070 302560 683179 302562
rect 683070 302504 683118 302560
rect 683174 302504 683179 302560
rect 683070 302499 683179 302504
rect 683070 302260 683130 302499
rect 35801 301610 35867 301613
rect 35758 301608 35867 301610
rect 35758 301552 35806 301608
rect 35862 301552 35867 301608
rect 35758 301547 35867 301552
rect 35758 301308 35818 301547
rect 35801 300930 35867 300933
rect 35788 300928 35867 300930
rect 35788 300872 35806 300928
rect 35862 300872 35867 300928
rect 35788 300870 35867 300872
rect 35801 300867 35867 300870
rect 45001 300522 45067 300525
rect 41492 300520 45067 300522
rect 41492 300464 45006 300520
rect 45062 300464 45067 300520
rect 41492 300462 45067 300464
rect 45001 300459 45067 300462
rect 44265 300114 44331 300117
rect 41492 300112 44331 300114
rect 41492 300056 44270 300112
rect 44326 300056 44331 300112
rect 41492 300054 44331 300056
rect 44265 300051 44331 300054
rect 44357 299706 44423 299709
rect 41492 299704 44423 299706
rect 41492 299648 44362 299704
rect 44418 299648 44423 299704
rect 41492 299646 44423 299648
rect 44357 299643 44423 299646
rect 675702 299372 675708 299436
rect 675772 299434 675778 299436
rect 679617 299434 679683 299437
rect 675772 299432 679683 299434
rect 675772 299376 679622 299432
rect 679678 299376 679683 299432
rect 675772 299374 679683 299376
rect 675772 299372 675778 299374
rect 679617 299371 679683 299374
rect 44541 299298 44607 299301
rect 41492 299296 44607 299298
rect 41492 299240 44546 299296
rect 44602 299240 44607 299296
rect 41492 299238 44607 299240
rect 44541 299235 44607 299238
rect 44265 298890 44331 298893
rect 41492 298888 44331 298890
rect 41492 298832 44270 298888
rect 44326 298832 44331 298888
rect 41492 298830 44331 298832
rect 44265 298827 44331 298830
rect 42885 298482 42951 298485
rect 652017 298482 652083 298485
rect 41492 298480 42951 298482
rect 41492 298424 42890 298480
rect 42946 298424 42951 298480
rect 41492 298422 42951 298424
rect 650164 298480 652083 298482
rect 650164 298424 652022 298480
rect 652078 298424 652083 298480
rect 650164 298422 652083 298424
rect 42885 298419 42951 298422
rect 652017 298419 652083 298422
rect 62113 298210 62179 298213
rect 62113 298208 64492 298210
rect 62113 298152 62118 298208
rect 62174 298152 64492 298208
rect 62113 298150 64492 298152
rect 62113 298147 62179 298150
rect 44173 298074 44239 298077
rect 41492 298072 44239 298074
rect 41492 298016 44178 298072
rect 44234 298016 44239 298072
rect 41492 298014 44239 298016
rect 44173 298011 44239 298014
rect 675886 297876 675892 297940
rect 675956 297938 675962 297940
rect 679709 297938 679775 297941
rect 675956 297936 679775 297938
rect 675956 297880 679714 297936
rect 679770 297880 679775 297936
rect 675956 297878 679775 297880
rect 675956 297876 675962 297878
rect 679709 297875 679775 297878
rect 42793 297666 42859 297669
rect 41492 297664 42859 297666
rect 41492 297608 42798 297664
rect 42854 297608 42859 297664
rect 41492 297606 42859 297608
rect 42793 297603 42859 297606
rect 675334 297332 675340 297396
rect 675404 297394 675410 297396
rect 676397 297394 676463 297397
rect 675404 297392 676463 297394
rect 675404 297336 676402 297392
rect 676458 297336 676463 297392
rect 675404 297334 676463 297336
rect 675404 297332 675410 297334
rect 676397 297331 676463 297334
rect 42793 297258 42859 297261
rect 41492 297256 42859 297258
rect 41492 297200 42798 297256
rect 42854 297200 42859 297256
rect 41492 297198 42859 297200
rect 42793 297195 42859 297198
rect 42742 296850 42748 296852
rect 41492 296790 42748 296850
rect 42742 296788 42748 296790
rect 42812 296788 42818 296852
rect 35157 296442 35223 296445
rect 35157 296440 35236 296442
rect 35157 296384 35162 296440
rect 35218 296384 35236 296440
rect 35157 296382 35236 296384
rect 35157 296379 35223 296382
rect 41822 296034 41828 296036
rect 41492 295974 41828 296034
rect 41822 295972 41828 295974
rect 41892 295972 41898 296036
rect 42006 295626 42012 295628
rect 41492 295566 42012 295626
rect 42006 295564 42012 295566
rect 42076 295564 42082 295628
rect 42885 295218 42951 295221
rect 41492 295216 42951 295218
rect 41492 295160 42890 295216
rect 42946 295160 42951 295216
rect 41492 295158 42951 295160
rect 42885 295155 42951 295158
rect 32397 294810 32463 294813
rect 675753 294812 675819 294813
rect 32397 294808 32476 294810
rect 32397 294752 32402 294808
rect 32458 294752 32476 294808
rect 32397 294750 32476 294752
rect 32397 294747 32463 294750
rect 675702 294748 675708 294812
rect 675772 294810 675819 294812
rect 675772 294808 675864 294810
rect 675814 294752 675864 294808
rect 675772 294750 675864 294752
rect 675772 294748 675819 294750
rect 675753 294747 675819 294748
rect 41822 294402 41828 294404
rect 41492 294342 41828 294402
rect 41822 294340 41828 294342
rect 41892 294340 41898 294404
rect 42558 293994 42564 293996
rect 41492 293934 42564 293994
rect 42558 293932 42564 293934
rect 42628 293932 42634 293996
rect 44449 293586 44515 293589
rect 41492 293584 44515 293586
rect 41492 293528 44454 293584
rect 44510 293528 44515 293584
rect 41492 293526 44515 293528
rect 44449 293523 44515 293526
rect 41822 293178 41828 293180
rect 41492 293118 41828 293178
rect 41822 293116 41828 293118
rect 41892 293116 41898 293180
rect 41822 292770 41828 292772
rect 41492 292710 41828 292770
rect 41822 292708 41828 292710
rect 41892 292708 41898 292772
rect 675477 292636 675543 292637
rect 675477 292634 675524 292636
rect 675432 292632 675524 292634
rect 675432 292576 675482 292632
rect 675432 292574 675524 292576
rect 675477 292572 675524 292574
rect 675588 292572 675594 292636
rect 675477 292571 675543 292572
rect 42977 292362 43043 292365
rect 41492 292360 43043 292362
rect 41492 292304 42982 292360
rect 43038 292304 43043 292360
rect 41492 292302 43043 292304
rect 42977 292299 43043 292302
rect 675385 292092 675451 292093
rect 675334 292090 675340 292092
rect 675294 292030 675340 292090
rect 675404 292088 675451 292092
rect 675446 292032 675451 292088
rect 675334 292028 675340 292030
rect 675404 292028 675451 292032
rect 675385 292027 675451 292028
rect 43161 291954 43227 291957
rect 41492 291952 43227 291954
rect 41492 291896 43166 291952
rect 43222 291896 43227 291952
rect 41492 291894 43227 291896
rect 43161 291891 43227 291894
rect 44541 291546 44607 291549
rect 41492 291544 44607 291546
rect 41492 291488 44546 291544
rect 44602 291488 44607 291544
rect 41492 291486 44607 291488
rect 44541 291483 44607 291486
rect 45001 291138 45067 291141
rect 41492 291136 45067 291138
rect 41492 291080 45006 291136
rect 45062 291080 45067 291136
rect 41492 291078 45067 291080
rect 45001 291075 45067 291078
rect 43897 290730 43963 290733
rect 41492 290728 43963 290730
rect 41492 290672 43902 290728
rect 43958 290672 43963 290728
rect 41492 290670 43963 290672
rect 43897 290667 43963 290670
rect 51809 289914 51875 289917
rect 41492 289912 51875 289914
rect 41492 289856 51814 289912
rect 51870 289856 51875 289912
rect 41492 289854 51875 289856
rect 51809 289851 51875 289854
rect 675661 288420 675727 288421
rect 675661 288416 675708 288420
rect 675772 288418 675778 288420
rect 675661 288360 675666 288416
rect 675661 288356 675708 288360
rect 675772 288358 675818 288418
rect 675772 288356 675778 288358
rect 675661 288355 675727 288356
rect 675753 287330 675819 287333
rect 676622 287330 676628 287332
rect 675753 287328 676628 287330
rect 675753 287272 675758 287328
rect 675814 287272 676628 287328
rect 675753 287270 676628 287272
rect 675753 287267 675819 287270
rect 676622 287268 676628 287270
rect 676692 287268 676698 287332
rect 675753 285562 675819 285565
rect 676070 285562 676076 285564
rect 675753 285560 676076 285562
rect 675753 285504 675758 285560
rect 675814 285504 676076 285560
rect 675753 285502 676076 285504
rect 675753 285499 675819 285502
rect 676070 285500 676076 285502
rect 676140 285500 676146 285564
rect 651557 285290 651623 285293
rect 650164 285288 651623 285290
rect 650164 285232 651562 285288
rect 651618 285232 651623 285288
rect 650164 285230 651623 285232
rect 651557 285227 651623 285230
rect 62113 285154 62179 285157
rect 62113 285152 64492 285154
rect 62113 285096 62118 285152
rect 62174 285096 64492 285152
rect 62113 285094 64492 285096
rect 62113 285091 62179 285094
rect 35157 284882 35223 284885
rect 41454 284882 41460 284884
rect 35157 284880 41460 284882
rect 35157 284824 35162 284880
rect 35218 284824 41460 284880
rect 35157 284822 41460 284824
rect 35157 284819 35223 284822
rect 41454 284820 41460 284822
rect 41524 284820 41530 284884
rect 675753 283658 675819 283661
rect 676438 283658 676444 283660
rect 675753 283656 676444 283658
rect 675753 283600 675758 283656
rect 675814 283600 676444 283656
rect 675753 283598 676444 283600
rect 675753 283595 675819 283598
rect 676438 283596 676444 283598
rect 676508 283596 676514 283660
rect 41454 281420 41460 281484
rect 41524 281482 41530 281484
rect 41781 281482 41847 281485
rect 41524 281480 41847 281482
rect 41524 281424 41786 281480
rect 41842 281424 41847 281480
rect 41524 281422 41847 281424
rect 41524 281420 41530 281422
rect 41781 281419 41847 281422
rect 675753 281482 675819 281485
rect 676254 281482 676260 281484
rect 675753 281480 676260 281482
rect 675753 281424 675758 281480
rect 675814 281424 676260 281480
rect 675753 281422 676260 281424
rect 675753 281419 675819 281422
rect 676254 281420 676260 281422
rect 676324 281420 676330 281484
rect 40902 279788 40908 279852
rect 40972 279850 40978 279852
rect 41781 279850 41847 279853
rect 40972 279848 41847 279850
rect 40972 279792 41786 279848
rect 41842 279792 41847 279848
rect 40972 279790 41847 279792
rect 40972 279788 40978 279790
rect 41781 279787 41847 279790
rect 41086 278020 41092 278084
rect 41156 278082 41162 278084
rect 41781 278082 41847 278085
rect 41156 278080 41847 278082
rect 41156 278024 41786 278080
rect 41842 278024 41847 278080
rect 41156 278022 41847 278024
rect 41156 278020 41162 278022
rect 41781 278019 41847 278022
rect 391933 275498 391999 275501
rect 544653 275498 544719 275501
rect 391933 275496 544719 275498
rect 391933 275440 391938 275496
rect 391994 275440 544658 275496
rect 544714 275440 544719 275496
rect 391933 275438 544719 275440
rect 391933 275435 391999 275438
rect 544653 275435 544719 275438
rect 371233 275362 371299 275365
rect 537569 275362 537635 275365
rect 371233 275360 537635 275362
rect 371233 275304 371238 275360
rect 371294 275304 537574 275360
rect 537630 275304 537635 275360
rect 371233 275302 537635 275304
rect 371233 275299 371299 275302
rect 537569 275299 537635 275302
rect 409689 275226 409755 275229
rect 640425 275226 640491 275229
rect 409689 275224 640491 275226
rect 409689 275168 409694 275224
rect 409750 275168 640430 275224
rect 640486 275168 640491 275224
rect 409689 275166 640491 275168
rect 409689 275163 409755 275166
rect 640425 275163 640491 275166
rect 382181 274138 382247 274141
rect 569493 274138 569559 274141
rect 382181 274136 569559 274138
rect 382181 274080 382186 274136
rect 382242 274080 569498 274136
rect 569554 274080 569559 274136
rect 382181 274078 569559 274080
rect 382181 274075 382247 274078
rect 569493 274075 569559 274078
rect 401041 274002 401107 274005
rect 619081 274002 619147 274005
rect 401041 274000 619147 274002
rect 401041 273944 401046 274000
rect 401102 273944 619086 274000
rect 619142 273944 619147 274000
rect 401041 273942 619147 273944
rect 401041 273939 401107 273942
rect 619081 273939 619147 273942
rect 411897 273866 411963 273869
rect 629753 273866 629819 273869
rect 411897 273864 629819 273866
rect 411897 273808 411902 273864
rect 411958 273808 629758 273864
rect 629814 273808 629819 273864
rect 411897 273806 629819 273808
rect 411897 273803 411963 273806
rect 629753 273803 629819 273806
rect 41781 273052 41847 273053
rect 41781 273048 41828 273052
rect 41892 273050 41898 273052
rect 41781 272992 41786 273048
rect 41781 272988 41828 272992
rect 41892 272990 41938 273050
rect 41892 272988 41898 272990
rect 41781 272987 41847 272988
rect 383377 272778 383443 272781
rect 572989 272778 573055 272781
rect 383377 272776 573055 272778
rect 383377 272720 383382 272776
rect 383438 272720 572994 272776
rect 573050 272720 573055 272776
rect 383377 272718 573055 272720
rect 383377 272715 383443 272718
rect 572989 272715 573055 272718
rect 404169 272642 404235 272645
rect 628557 272642 628623 272645
rect 404169 272640 628623 272642
rect 404169 272584 404174 272640
rect 404230 272584 628562 272640
rect 628618 272584 628623 272640
rect 404169 272582 628623 272584
rect 404169 272579 404235 272582
rect 628557 272579 628623 272582
rect 406929 272506 406995 272509
rect 635641 272506 635707 272509
rect 406929 272504 635707 272506
rect 406929 272448 406934 272504
rect 406990 272448 635646 272504
rect 635702 272448 635707 272504
rect 406929 272446 635707 272448
rect 406929 272443 406995 272446
rect 635641 272443 635707 272446
rect 41638 272172 41644 272236
rect 41708 272234 41714 272236
rect 41781 272234 41847 272237
rect 41708 272232 41847 272234
rect 41708 272176 41786 272232
rect 41842 272176 41847 272232
rect 41708 272174 41847 272176
rect 41708 272172 41714 272174
rect 41781 272171 41847 272174
rect 406101 271418 406167 271421
rect 448973 271418 449039 271421
rect 406101 271416 449039 271418
rect 406101 271360 406106 271416
rect 406162 271360 448978 271416
rect 449034 271360 449039 271416
rect 406101 271358 449039 271360
rect 406101 271355 406167 271358
rect 448973 271355 449039 271358
rect 379329 271282 379395 271285
rect 562409 271282 562475 271285
rect 379329 271280 562475 271282
rect 379329 271224 379334 271280
rect 379390 271224 562414 271280
rect 562470 271224 562475 271280
rect 379329 271222 562475 271224
rect 379329 271219 379395 271222
rect 562409 271219 562475 271222
rect 395705 271146 395771 271149
rect 604913 271146 604979 271149
rect 395705 271144 604979 271146
rect 395705 271088 395710 271144
rect 395766 271088 604918 271144
rect 604974 271088 604979 271144
rect 395705 271086 604979 271088
rect 395705 271083 395771 271086
rect 604913 271083 604979 271086
rect 41965 270468 42031 270469
rect 41965 270464 42012 270468
rect 42076 270466 42082 270468
rect 41965 270408 41970 270464
rect 41965 270404 42012 270408
rect 42076 270406 42122 270466
rect 42076 270404 42082 270406
rect 41965 270403 42031 270404
rect 376477 270058 376543 270061
rect 554773 270058 554839 270061
rect 376477 270056 554839 270058
rect 376477 270000 376482 270056
rect 376538 270000 554778 270056
rect 554834 270000 554839 270056
rect 376477 269998 554839 270000
rect 376477 269995 376543 269998
rect 554773 269995 554839 269998
rect 386045 269922 386111 269925
rect 579613 269922 579679 269925
rect 386045 269920 579679 269922
rect 386045 269864 386050 269920
rect 386106 269864 579618 269920
rect 579674 269864 579679 269920
rect 386045 269862 579679 269864
rect 386045 269859 386111 269862
rect 579613 269859 579679 269862
rect 40718 269724 40724 269788
rect 40788 269786 40794 269788
rect 41781 269786 41847 269789
rect 40788 269784 41847 269786
rect 40788 269728 41786 269784
rect 41842 269728 41847 269784
rect 40788 269726 41847 269728
rect 40788 269724 40794 269726
rect 41781 269723 41847 269726
rect 394969 269786 395035 269789
rect 603073 269786 603139 269789
rect 394969 269784 603139 269786
rect 394969 269728 394974 269784
rect 395030 269728 603078 269784
rect 603134 269728 603139 269784
rect 394969 269726 603139 269728
rect 394969 269723 395035 269726
rect 603073 269723 603139 269726
rect 40534 269044 40540 269108
rect 40604 269106 40610 269108
rect 41781 269106 41847 269109
rect 40604 269104 41847 269106
rect 40604 269048 41786 269104
rect 41842 269048 41847 269104
rect 40604 269046 41847 269048
rect 40604 269044 40610 269046
rect 41781 269043 41847 269046
rect 398465 268698 398531 268701
rect 612733 268698 612799 268701
rect 398465 268696 612799 268698
rect 398465 268640 398470 268696
rect 398526 268640 612738 268696
rect 612794 268640 612799 268696
rect 398465 268638 612799 268640
rect 398465 268635 398531 268638
rect 612733 268635 612799 268638
rect 676262 268565 676322 268668
rect 405733 268562 405799 268565
rect 622393 268562 622459 268565
rect 405733 268560 622459 268562
rect 405733 268504 405738 268560
rect 405794 268504 622398 268560
rect 622454 268504 622459 268560
rect 405733 268502 622459 268504
rect 405733 268499 405799 268502
rect 622393 268499 622459 268502
rect 676213 268560 676322 268565
rect 676213 268504 676218 268560
rect 676274 268504 676322 268560
rect 676213 268502 676322 268504
rect 676213 268499 676279 268502
rect 402513 268426 402579 268429
rect 623773 268426 623839 268429
rect 402513 268424 623839 268426
rect 402513 268368 402518 268424
rect 402574 268368 623778 268424
rect 623834 268368 623839 268424
rect 402513 268366 623839 268368
rect 402513 268363 402579 268366
rect 623773 268363 623839 268366
rect 676121 268154 676187 268157
rect 676262 268154 676322 268260
rect 676121 268152 676322 268154
rect 676121 268096 676126 268152
rect 676182 268096 676322 268152
rect 676121 268094 676322 268096
rect 676121 268091 676187 268094
rect 676262 267749 676322 267852
rect 676213 267744 676322 267749
rect 676213 267688 676218 267744
rect 676274 267688 676322 267744
rect 676213 267686 676322 267688
rect 676213 267683 676279 267686
rect 676262 267341 676322 267444
rect 407389 267338 407455 267341
rect 457989 267338 458055 267341
rect 407389 267336 458055 267338
rect 407389 267280 407394 267336
rect 407450 267280 457994 267336
rect 458050 267280 458055 267336
rect 407389 267278 458055 267280
rect 407389 267275 407455 267278
rect 457989 267275 458055 267278
rect 676213 267336 676322 267341
rect 676213 267280 676218 267336
rect 676274 267280 676322 267336
rect 676213 267278 676322 267280
rect 676213 267275 676279 267278
rect 410977 267202 411043 267205
rect 645853 267202 645919 267205
rect 410977 267200 645919 267202
rect 410977 267144 410982 267200
rect 411038 267144 645858 267200
rect 645914 267144 645919 267200
rect 410977 267142 645919 267144
rect 410977 267139 411043 267142
rect 645853 267139 645919 267142
rect 389173 267066 389239 267069
rect 404353 267066 404419 267069
rect 389173 267064 404419 267066
rect 389173 267008 389178 267064
rect 389234 267008 404358 267064
rect 404414 267008 404419 267064
rect 389173 267006 404419 267008
rect 389173 267003 389239 267006
rect 404353 267003 404419 267006
rect 412265 267066 412331 267069
rect 648613 267066 648679 267069
rect 412265 267064 648679 267066
rect 412265 267008 412270 267064
rect 412326 267008 648618 267064
rect 648674 267008 648679 267064
rect 412265 267006 648679 267008
rect 412265 267003 412331 267006
rect 648613 267003 648679 267006
rect 676029 267066 676095 267069
rect 676029 267064 676292 267066
rect 676029 267008 676034 267064
rect 676090 267008 676292 267064
rect 676029 267006 676292 267008
rect 676029 267003 676095 267006
rect 676262 266525 676322 266628
rect 402053 266522 402119 266525
rect 405733 266522 405799 266525
rect 402053 266520 405799 266522
rect 402053 266464 402058 266520
rect 402114 266464 405738 266520
rect 405794 266464 405799 266520
rect 402053 266462 405799 266464
rect 402053 266459 402119 266462
rect 405733 266459 405799 266462
rect 676213 266520 676322 266525
rect 676213 266464 676218 266520
rect 676274 266464 676322 266520
rect 676213 266462 676322 266464
rect 676213 266459 676279 266462
rect 404721 266386 404787 266389
rect 411897 266386 411963 266389
rect 404721 266384 411963 266386
rect 404721 266328 404726 266384
rect 404782 266328 411902 266384
rect 411958 266328 411963 266384
rect 404721 266326 411963 266328
rect 404721 266323 404787 266326
rect 411897 266323 411963 266326
rect 676262 266117 676322 266220
rect 676213 266112 676322 266117
rect 676213 266056 676218 266112
rect 676274 266056 676322 266112
rect 676213 266054 676322 266056
rect 676213 266051 676279 266054
rect 388253 265842 388319 265845
rect 585133 265842 585199 265845
rect 388253 265840 585199 265842
rect 388253 265784 388258 265840
rect 388314 265784 585138 265840
rect 585194 265784 585199 265840
rect 388253 265782 585199 265784
rect 388253 265779 388319 265782
rect 585133 265779 585199 265782
rect 676029 265842 676095 265845
rect 676029 265840 676292 265842
rect 676029 265784 676034 265840
rect 676090 265784 676292 265840
rect 676029 265782 676292 265784
rect 676029 265779 676095 265782
rect 405181 265706 405247 265709
rect 630673 265706 630739 265709
rect 405181 265704 630739 265706
rect 405181 265648 405186 265704
rect 405242 265648 630678 265704
rect 630734 265648 630739 265704
rect 405181 265646 630739 265648
rect 405181 265643 405247 265646
rect 630673 265643 630739 265646
rect 407849 265570 407915 265573
rect 637573 265570 637639 265573
rect 407849 265568 637639 265570
rect 407849 265512 407854 265568
rect 407910 265512 637578 265568
rect 637634 265512 637639 265568
rect 407849 265510 637639 265512
rect 407849 265507 407915 265510
rect 637573 265507 637639 265510
rect 676262 265301 676322 265404
rect 676213 265296 676322 265301
rect 676213 265240 676218 265296
rect 676274 265240 676322 265296
rect 676213 265238 676322 265240
rect 676213 265235 676279 265238
rect 674741 265026 674807 265029
rect 674741 265024 676292 265026
rect 674741 264968 674746 265024
rect 674802 264968 676292 265024
rect 674741 264966 676292 264968
rect 674741 264963 674807 264966
rect 676262 264485 676322 264588
rect 676213 264480 676322 264485
rect 676213 264424 676218 264480
rect 676274 264424 676322 264480
rect 676213 264422 676322 264424
rect 676213 264419 676279 264422
rect 396993 264210 397059 264213
rect 401225 264210 401291 264213
rect 396993 264208 401291 264210
rect 396993 264152 396998 264208
rect 397054 264152 401230 264208
rect 401286 264152 401291 264208
rect 396993 264150 401291 264152
rect 396993 264147 397059 264150
rect 401225 264147 401291 264150
rect 676262 264077 676322 264180
rect 676262 264072 676371 264077
rect 676262 264016 676310 264072
rect 676366 264016 676371 264072
rect 676262 264014 676371 264016
rect 676305 264011 676371 264014
rect 676814 263669 676874 263772
rect 676814 263664 676923 263669
rect 676814 263608 676862 263664
rect 676918 263608 676923 263664
rect 676814 263606 676923 263608
rect 676857 263603 676923 263606
rect 675385 263394 675451 263397
rect 675385 263392 676292 263394
rect 675385 263336 675390 263392
rect 675446 263336 676292 263392
rect 675385 263334 676292 263336
rect 675385 263331 675451 263334
rect 676029 262986 676095 262989
rect 676029 262984 676292 262986
rect 676029 262928 676034 262984
rect 676090 262928 676292 262984
rect 676029 262926 676292 262928
rect 676029 262923 676095 262926
rect 676029 262578 676095 262581
rect 676029 262576 676292 262578
rect 676029 262520 676034 262576
rect 676090 262520 676292 262576
rect 676029 262518 676292 262520
rect 676029 262515 676095 262518
rect 415301 262306 415367 262309
rect 412436 262304 415367 262306
rect 412436 262248 415306 262304
rect 415362 262248 415367 262304
rect 412436 262246 415367 262248
rect 415301 262243 415367 262246
rect 676262 262037 676322 262140
rect 676213 262032 676322 262037
rect 676213 261976 676218 262032
rect 676274 261976 676322 262032
rect 676213 261974 676322 261976
rect 676213 261971 676279 261974
rect 676262 261629 676322 261732
rect 676213 261624 676322 261629
rect 676213 261568 676218 261624
rect 676274 261568 676322 261624
rect 676213 261566 676322 261568
rect 676213 261563 676279 261566
rect 676262 261221 676322 261324
rect 676213 261216 676322 261221
rect 676213 261160 676218 261216
rect 676274 261160 676322 261216
rect 676213 261158 676322 261160
rect 676213 261155 676279 261158
rect 677182 260812 677242 260916
rect 677174 260748 677180 260812
rect 677244 260748 677250 260812
rect 676998 260404 677058 260508
rect 676990 260340 676996 260404
rect 677060 260340 677066 260404
rect 676262 259997 676322 260100
rect 676213 259992 676322 259997
rect 676213 259936 676218 259992
rect 676274 259936 676322 259992
rect 676213 259934 676322 259936
rect 676213 259931 676279 259934
rect 676814 259588 676874 259692
rect 676806 259524 676812 259588
rect 676876 259524 676882 259588
rect 414197 259178 414263 259181
rect 412436 259176 414263 259178
rect 412436 259120 414202 259176
rect 414258 259120 414263 259176
rect 412436 259118 414263 259120
rect 414197 259115 414263 259118
rect 676121 259178 676187 259181
rect 676262 259178 676322 259284
rect 676121 259176 676322 259178
rect 676121 259120 676126 259176
rect 676182 259120 676322 259176
rect 676121 259118 676322 259120
rect 676121 259115 676187 259118
rect 676262 258773 676322 258876
rect 676213 258768 676322 258773
rect 676213 258712 676218 258768
rect 676274 258712 676322 258768
rect 676213 258710 676322 258712
rect 676213 258707 676279 258710
rect 189073 258634 189139 258637
rect 189073 258632 191820 258634
rect 189073 258576 189078 258632
rect 189134 258576 191820 258632
rect 189073 258574 191820 258576
rect 189073 258571 189139 258574
rect 683070 258365 683130 258468
rect 28349 258362 28415 258365
rect 28349 258360 28458 258362
rect 28349 258304 28354 258360
rect 28410 258304 28458 258360
rect 28349 258299 28458 258304
rect 683070 258360 683179 258365
rect 683070 258304 683118 258360
rect 683174 258304 683179 258360
rect 683070 258302 683179 258304
rect 683113 258299 683179 258302
rect 28398 258060 28458 258299
rect 683070 257652 683130 258060
rect 31710 257549 31770 257652
rect 31477 257546 31543 257549
rect 31477 257544 31586 257546
rect 31477 257488 31482 257544
rect 31538 257488 31586 257544
rect 31477 257483 31586 257488
rect 31661 257544 31770 257549
rect 683113 257546 683179 257549
rect 31661 257488 31666 257544
rect 31722 257488 31770 257544
rect 31661 257486 31770 257488
rect 683070 257544 683179 257546
rect 683070 257488 683118 257544
rect 683174 257488 683179 257544
rect 31661 257483 31727 257486
rect 683070 257483 683179 257488
rect 31526 257244 31586 257483
rect 683070 257244 683130 257483
rect 31569 257138 31635 257141
rect 31526 257136 31635 257138
rect 31526 257080 31574 257136
rect 31630 257080 31635 257136
rect 31526 257075 31635 257080
rect 31526 256836 31586 257075
rect 42885 256458 42951 256461
rect 41492 256456 42951 256458
rect 41492 256400 42890 256456
rect 42946 256400 42951 256456
rect 41492 256398 42951 256400
rect 42885 256395 42951 256398
rect 44265 256050 44331 256053
rect 41492 256048 44331 256050
rect 41492 255992 44270 256048
rect 44326 255992 44331 256048
rect 41492 255990 44331 255992
rect 44265 255987 44331 255990
rect 415301 255914 415367 255917
rect 412436 255912 415367 255914
rect 412436 255856 415306 255912
rect 415362 255856 415367 255912
rect 412436 255854 415367 255856
rect 415301 255851 415367 255854
rect 43345 255642 43411 255645
rect 41492 255640 43411 255642
rect 41492 255584 43350 255640
rect 43406 255584 43411 255640
rect 41492 255582 43411 255584
rect 43345 255579 43411 255582
rect 44173 255234 44239 255237
rect 41492 255232 44239 255234
rect 41492 255176 44178 255232
rect 44234 255176 44239 255232
rect 41492 255174 44239 255176
rect 44173 255171 44239 255174
rect 44265 254826 44331 254829
rect 41492 254824 44331 254826
rect 41492 254768 44270 254824
rect 44326 254768 44331 254824
rect 41492 254766 44331 254768
rect 44265 254763 44331 254766
rect 42793 254418 42859 254421
rect 41492 254416 42859 254418
rect 41492 254360 42798 254416
rect 42854 254360 42859 254416
rect 41492 254358 42859 254360
rect 42793 254355 42859 254358
rect 44725 254010 44791 254013
rect 41492 254008 44791 254010
rect 41492 253952 44730 254008
rect 44786 253952 44791 254008
rect 41492 253950 44791 253952
rect 44725 253947 44791 253950
rect 30974 253469 31034 253572
rect 30974 253464 31083 253469
rect 30974 253408 31022 253464
rect 31078 253408 31083 253464
rect 30974 253406 31083 253408
rect 31017 253403 31083 253406
rect 32446 253061 32506 253164
rect 175038 253132 175044 253196
rect 175108 253194 175114 253196
rect 185209 253194 185275 253197
rect 175108 253192 185275 253194
rect 175108 253136 185214 253192
rect 185270 253136 185275 253192
rect 175108 253134 185275 253136
rect 175108 253132 175114 253134
rect 185209 253131 185275 253134
rect 32397 253056 32506 253061
rect 32397 253000 32402 253056
rect 32458 253000 32506 253056
rect 32397 252998 32506 253000
rect 32397 252995 32463 252998
rect 42977 252786 43043 252789
rect 414381 252786 414447 252789
rect 41492 252784 43043 252786
rect 41492 252728 42982 252784
rect 43038 252728 43043 252784
rect 41492 252726 43043 252728
rect 412436 252784 414447 252786
rect 412436 252728 414386 252784
rect 414442 252728 414447 252784
rect 412436 252726 414447 252728
rect 42977 252723 43043 252726
rect 414381 252723 414447 252726
rect 31158 252245 31218 252348
rect 31109 252240 31218 252245
rect 31109 252184 31114 252240
rect 31170 252184 31218 252240
rect 31109 252182 31218 252184
rect 31109 252179 31175 252182
rect 43161 251970 43227 251973
rect 41492 251968 43227 251970
rect 41492 251912 43166 251968
rect 43222 251912 43227 251968
rect 41492 251910 43227 251912
rect 43161 251907 43227 251910
rect 44173 251562 44239 251565
rect 41492 251560 44239 251562
rect 41492 251504 44178 251560
rect 44234 251504 44239 251560
rect 41492 251502 44239 251504
rect 44173 251499 44239 251502
rect 675150 251500 675156 251564
rect 675220 251562 675226 251564
rect 676857 251562 676923 251565
rect 675220 251560 676923 251562
rect 675220 251504 676862 251560
rect 676918 251504 676923 251560
rect 675220 251502 676923 251504
rect 675220 251500 675226 251502
rect 676857 251499 676923 251502
rect 44357 251154 44423 251157
rect 41492 251152 44423 251154
rect 41492 251096 44362 251152
rect 44418 251096 44423 251152
rect 41492 251094 44423 251096
rect 44357 251091 44423 251094
rect 43069 250746 43135 250749
rect 41492 250744 43135 250746
rect 41492 250688 43074 250744
rect 43130 250688 43135 250744
rect 41492 250686 43135 250688
rect 43069 250683 43135 250686
rect 40542 250204 40602 250308
rect 40534 250140 40540 250204
rect 40604 250140 40610 250204
rect 40726 249796 40786 249900
rect 40718 249732 40724 249796
rect 40788 249732 40794 249796
rect 675150 249596 675156 249660
rect 675220 249596 675226 249660
rect 44541 249522 44607 249525
rect 414197 249522 414263 249525
rect 41492 249520 44607 249522
rect 41492 249464 44546 249520
rect 44602 249464 44607 249520
rect 41492 249462 44607 249464
rect 412436 249520 414263 249522
rect 412436 249464 414202 249520
rect 414258 249464 414263 249520
rect 412436 249462 414263 249464
rect 44541 249459 44607 249462
rect 414197 249459 414263 249462
rect 43253 249114 43319 249117
rect 41492 249112 43319 249114
rect 41492 249056 43258 249112
rect 43314 249056 43319 249112
rect 41492 249054 43319 249056
rect 43253 249051 43319 249054
rect 44909 248706 44975 248709
rect 41492 248704 44975 248706
rect 41492 248648 44914 248704
rect 44970 248648 44975 248704
rect 41492 248646 44975 248648
rect 44909 248643 44975 248646
rect 675158 248301 675218 249596
rect 44633 248298 44699 248301
rect 41492 248296 44699 248298
rect 41492 248240 44638 248296
rect 44694 248240 44699 248296
rect 41492 248238 44699 248240
rect 44633 248235 44699 248238
rect 675109 248296 675218 248301
rect 675109 248240 675114 248296
rect 675170 248240 675218 248296
rect 675109 248238 675218 248240
rect 675109 248235 675175 248238
rect 190361 248026 190427 248029
rect 190361 248024 191820 248026
rect 190361 247968 190366 248024
rect 190422 247968 191820 248024
rect 190361 247966 191820 247968
rect 190361 247963 190427 247966
rect 41462 247754 41522 247860
rect 41462 247694 55230 247754
rect 41462 247346 41522 247452
rect 55170 247346 55230 247694
rect 191097 247346 191163 247349
rect 41462 247286 45570 247346
rect 55170 247344 191163 247346
rect 55170 247288 191102 247344
rect 191158 247288 191163 247344
rect 55170 247286 191163 247288
rect 45510 247210 45570 247286
rect 191097 247283 191163 247286
rect 189717 247210 189783 247213
rect 45510 247208 189783 247210
rect 45510 247152 189722 247208
rect 189778 247152 189783 247208
rect 45510 247150 189783 247152
rect 189717 247147 189783 247150
rect 675753 246666 675819 246669
rect 677174 246666 677180 246668
rect 675753 246664 677180 246666
rect 35758 246533 35818 246636
rect 675753 246608 675758 246664
rect 675814 246608 677180 246664
rect 675753 246606 677180 246608
rect 675753 246603 675819 246606
rect 677174 246604 677180 246606
rect 677244 246604 677250 246668
rect 35758 246528 35867 246533
rect 35758 246472 35806 246528
rect 35862 246472 35867 246528
rect 35758 246470 35867 246472
rect 35801 246467 35867 246470
rect 415301 246394 415367 246397
rect 412436 246392 415367 246394
rect 412436 246336 415306 246392
rect 415362 246336 415367 246392
rect 412436 246334 415367 246336
rect 415301 246331 415367 246334
rect 674465 245714 674531 245717
rect 675702 245714 675708 245716
rect 674465 245712 675708 245714
rect 674465 245656 674470 245712
rect 674526 245656 675708 245712
rect 674465 245654 675708 245656
rect 674465 245651 674531 245654
rect 675702 245652 675708 245654
rect 675772 245652 675778 245716
rect 675753 245442 675819 245445
rect 676806 245442 676812 245444
rect 675753 245440 676812 245442
rect 675753 245384 675758 245440
rect 675814 245384 676812 245440
rect 675753 245382 676812 245384
rect 675753 245379 675819 245382
rect 676806 245380 676812 245382
rect 676876 245380 676882 245444
rect 414381 243130 414447 243133
rect 412436 243128 414447 243130
rect 412436 243072 414386 243128
rect 414442 243072 414447 243128
rect 412436 243070 414447 243072
rect 414381 243067 414447 243070
rect 174997 241636 175063 241637
rect 174997 241634 175044 241636
rect 174952 241632 175044 241634
rect 174952 241576 175002 241632
rect 174952 241574 175044 241576
rect 174997 241572 175044 241574
rect 175108 241572 175114 241636
rect 174997 241571 175063 241572
rect 41965 240682 42031 240685
rect 41965 240680 42074 240682
rect 41965 240624 41970 240680
rect 42026 240624 42074 240680
rect 41965 240619 42074 240624
rect 42014 238509 42074 240619
rect 414933 240002 414999 240005
rect 412436 240000 414999 240002
rect 412436 239944 414938 240000
rect 414994 239944 414999 240000
rect 412436 239942 414999 239944
rect 414933 239939 414999 239942
rect 42701 238778 42767 238781
rect 42701 238776 42810 238778
rect 42701 238720 42706 238776
rect 42762 238720 42810 238776
rect 42701 238715 42810 238720
rect 41965 238504 42074 238509
rect 41965 238448 41970 238504
rect 42026 238448 42074 238504
rect 41965 238446 42074 238448
rect 41965 238443 42031 238446
rect 42006 238036 42012 238100
rect 42076 238098 42082 238100
rect 42750 238098 42810 238715
rect 675293 238642 675359 238645
rect 676990 238642 676996 238644
rect 675293 238640 676996 238642
rect 675293 238584 675298 238640
rect 675354 238584 676996 238640
rect 675293 238582 676996 238584
rect 675293 238579 675359 238582
rect 676990 238580 676996 238582
rect 677060 238580 677066 238644
rect 42076 238038 42810 238098
rect 42076 238036 42082 238038
rect 42190 237356 42196 237420
rect 42260 237418 42266 237420
rect 42701 237418 42767 237421
rect 42260 237416 42767 237418
rect 42260 237360 42706 237416
rect 42762 237360 42767 237416
rect 42260 237358 42767 237360
rect 42260 237356 42266 237358
rect 42701 237355 42767 237358
rect 189073 237418 189139 237421
rect 189073 237416 191820 237418
rect 189073 237360 189078 237416
rect 189134 237360 191820 237416
rect 189073 237358 191820 237360
rect 189073 237355 189139 237358
rect 675753 236876 675819 236877
rect 675702 236874 675708 236876
rect 675662 236814 675708 236874
rect 675772 236872 675819 236876
rect 675814 236816 675819 236872
rect 675702 236812 675708 236814
rect 675772 236812 675819 236816
rect 675753 236811 675819 236812
rect 40718 236676 40724 236740
rect 40788 236738 40794 236740
rect 41781 236738 41847 236741
rect 414197 236738 414263 236741
rect 40788 236736 41847 236738
rect 40788 236680 41786 236736
rect 41842 236680 41847 236736
rect 40788 236678 41847 236680
rect 412436 236736 414263 236738
rect 412436 236680 414202 236736
rect 414258 236680 414263 236736
rect 412436 236678 414263 236680
rect 40788 236676 40794 236678
rect 41781 236675 41847 236678
rect 414197 236675 414263 236678
rect 415301 233610 415367 233613
rect 412436 233608 415367 233610
rect 412436 233552 415306 233608
rect 415362 233552 415367 233608
rect 412436 233550 415367 233552
rect 415301 233547 415367 233550
rect 40534 232868 40540 232932
rect 40604 232930 40610 232932
rect 42425 232930 42491 232933
rect 40604 232928 42491 232930
rect 40604 232872 42430 232928
rect 42486 232872 42491 232928
rect 40604 232870 42491 232872
rect 40604 232868 40610 232870
rect 42425 232867 42491 232870
rect 43529 231162 43595 231165
rect 647366 231162 647372 231164
rect 43529 231160 647372 231162
rect 43529 231104 43534 231160
rect 43590 231104 647372 231160
rect 43529 231102 647372 231104
rect 43529 231099 43595 231102
rect 647366 231100 647372 231102
rect 647436 231100 647442 231164
rect 196617 230346 196683 230349
rect 199009 230346 199075 230349
rect 196617 230344 199075 230346
rect 196617 230288 196622 230344
rect 196678 230288 199014 230344
rect 199070 230288 199075 230344
rect 196617 230286 199075 230288
rect 196617 230283 196683 230286
rect 199009 230283 199075 230286
rect 376937 230346 377003 230349
rect 428641 230346 428707 230349
rect 376937 230344 428707 230346
rect 376937 230288 376942 230344
rect 376998 230288 428646 230344
rect 428702 230288 428707 230344
rect 376937 230286 428707 230288
rect 376937 230283 377003 230286
rect 428641 230283 428707 230286
rect 381537 230210 381603 230213
rect 478137 230210 478203 230213
rect 381537 230208 478203 230210
rect 381537 230152 381542 230208
rect 381598 230152 478142 230208
rect 478198 230152 478203 230208
rect 381537 230150 478203 230152
rect 381537 230147 381603 230150
rect 478137 230147 478203 230150
rect 375833 230074 375899 230077
rect 486417 230074 486483 230077
rect 375833 230072 486483 230074
rect 375833 230016 375838 230072
rect 375894 230016 486422 230072
rect 486478 230016 486483 230072
rect 375833 230014 486483 230016
rect 375833 230011 375899 230014
rect 486417 230011 486483 230014
rect 64137 229938 64203 229941
rect 196157 229938 196223 229941
rect 64137 229936 196223 229938
rect 64137 229880 64142 229936
rect 64198 229880 196162 229936
rect 196218 229880 196223 229936
rect 64137 229878 196223 229880
rect 64137 229875 64203 229878
rect 196157 229875 196223 229878
rect 378685 229938 378751 229941
rect 493317 229938 493383 229941
rect 378685 229936 493383 229938
rect 378685 229880 378690 229936
rect 378746 229880 493322 229936
rect 493378 229880 493383 229936
rect 378685 229878 493383 229880
rect 378685 229875 378751 229878
rect 493317 229875 493383 229878
rect 57881 229802 57947 229805
rect 194777 229802 194843 229805
rect 57881 229800 194843 229802
rect 57881 229744 57886 229800
rect 57942 229744 194782 229800
rect 194838 229744 194843 229800
rect 57881 229742 194843 229744
rect 57881 229739 57947 229742
rect 194777 229739 194843 229742
rect 380157 229802 380223 229805
rect 496077 229802 496143 229805
rect 380157 229800 496143 229802
rect 380157 229744 380162 229800
rect 380218 229744 496082 229800
rect 496138 229744 496143 229800
rect 380157 229742 496143 229744
rect 380157 229739 380223 229742
rect 496077 229739 496143 229742
rect 646129 229666 646195 229669
rect 646446 229666 646452 229668
rect 646129 229664 646452 229666
rect 646129 229608 646134 229664
rect 646190 229608 646452 229664
rect 646129 229606 646452 229608
rect 646129 229603 646195 229606
rect 646446 229604 646452 229606
rect 646516 229604 646522 229668
rect 42149 228988 42215 228989
rect 42149 228986 42196 228988
rect 42104 228984 42196 228986
rect 42104 228928 42154 228984
rect 42104 228926 42196 228928
rect 42149 228924 42196 228926
rect 42260 228924 42266 228988
rect 42149 228923 42215 228924
rect 387241 228714 387307 228717
rect 513373 228714 513439 228717
rect 387241 228712 513439 228714
rect 387241 228656 387246 228712
rect 387302 228656 513378 228712
rect 513434 228656 513439 228712
rect 387241 228654 513439 228656
rect 387241 228651 387307 228654
rect 513373 228651 513439 228654
rect 399385 228578 399451 228581
rect 541525 228578 541591 228581
rect 399385 228576 541591 228578
rect 399385 228520 399390 228576
rect 399446 228520 541530 228576
rect 541586 228520 541591 228576
rect 399385 228518 541591 228520
rect 399385 228515 399451 228518
rect 541525 228515 541591 228518
rect 90541 228442 90607 228445
rect 207933 228442 207999 228445
rect 90541 228440 207999 228442
rect 90541 228384 90546 228440
rect 90602 228384 207938 228440
rect 207994 228384 207999 228440
rect 90541 228382 207999 228384
rect 90541 228379 90607 228382
rect 207933 228379 207999 228382
rect 402605 228442 402671 228445
rect 549253 228442 549319 228445
rect 402605 228440 549319 228442
rect 402605 228384 402610 228440
rect 402666 228384 549258 228440
rect 549314 228384 549319 228440
rect 402605 228382 549319 228384
rect 402605 228379 402671 228382
rect 549253 228379 549319 228382
rect 86861 228306 86927 228309
rect 206553 228306 206619 228309
rect 86861 228304 206619 228306
rect 86861 228248 86866 228304
rect 86922 228248 206558 228304
rect 206614 228248 206619 228304
rect 86861 228246 206619 228248
rect 86861 228243 86927 228246
rect 206553 228243 206619 228246
rect 411069 228306 411135 228309
rect 564433 228306 564499 228309
rect 411069 228304 564499 228306
rect 411069 228248 411074 228304
rect 411130 228248 564438 228304
rect 564494 228248 564499 228304
rect 411069 228246 564499 228248
rect 411069 228243 411135 228246
rect 564433 228243 564499 228246
rect 41965 227356 42031 227357
rect 41965 227352 42012 227356
rect 42076 227354 42082 227356
rect 380525 227354 380591 227357
rect 496905 227354 496971 227357
rect 41965 227296 41970 227352
rect 41965 227292 42012 227296
rect 42076 227294 42122 227354
rect 380525 227352 496971 227354
rect 380525 227296 380530 227352
rect 380586 227296 496910 227352
rect 496966 227296 496971 227352
rect 380525 227294 496971 227296
rect 42076 227292 42082 227294
rect 41965 227291 42031 227292
rect 380525 227291 380591 227294
rect 496905 227291 496971 227294
rect 72969 227218 73035 227221
rect 201493 227218 201559 227221
rect 72969 227216 201559 227218
rect 72969 227160 72974 227216
rect 73030 227160 201498 227216
rect 201554 227160 201559 227216
rect 72969 227158 201559 227160
rect 72969 227155 73035 227158
rect 201493 227155 201559 227158
rect 383009 227218 383075 227221
rect 502517 227218 502583 227221
rect 383009 227216 502583 227218
rect 383009 227160 383014 227216
rect 383070 227160 502522 227216
rect 502578 227160 502583 227216
rect 383009 227158 502583 227160
rect 383009 227155 383075 227158
rect 502517 227155 502583 227158
rect 62757 227082 62823 227085
rect 197261 227082 197327 227085
rect 62757 227080 197327 227082
rect 62757 227024 62762 227080
rect 62818 227024 197266 227080
rect 197322 227024 197327 227080
rect 62757 227022 197327 227024
rect 62757 227019 62823 227022
rect 197261 227019 197327 227022
rect 388345 227082 388411 227085
rect 515489 227082 515555 227085
rect 388345 227080 515555 227082
rect 388345 227024 388350 227080
rect 388406 227024 515494 227080
rect 515550 227024 515555 227080
rect 388345 227022 515555 227024
rect 388345 227019 388411 227022
rect 515489 227019 515555 227022
rect 59261 226946 59327 226949
rect 195789 226946 195855 226949
rect 59261 226944 195855 226946
rect 59261 226888 59266 226944
rect 59322 226888 195794 226944
rect 195850 226888 195855 226944
rect 59261 226886 195855 226888
rect 59261 226883 59327 226886
rect 195789 226883 195855 226886
rect 407941 226946 408007 226949
rect 561673 226946 561739 226949
rect 407941 226944 561739 226946
rect 407941 226888 407946 226944
rect 408002 226888 561678 226944
rect 561734 226888 561739 226944
rect 407941 226886 561739 226888
rect 407941 226883 408007 226886
rect 561673 226883 561739 226886
rect 386229 225994 386295 225997
rect 510705 225994 510771 225997
rect 386229 225992 510771 225994
rect 386229 225936 386234 225992
rect 386290 225936 510710 225992
rect 510766 225936 510771 225992
rect 386229 225934 510771 225936
rect 386229 225931 386295 225934
rect 510705 225931 510771 225934
rect 394049 225858 394115 225861
rect 528921 225858 528987 225861
rect 394049 225856 528987 225858
rect 394049 225800 394054 225856
rect 394110 225800 528926 225856
rect 528982 225800 528987 225856
rect 394049 225798 528987 225800
rect 394049 225795 394115 225798
rect 528921 225795 528987 225798
rect 93025 225722 93091 225725
rect 210049 225722 210115 225725
rect 93025 225720 210115 225722
rect 93025 225664 93030 225720
rect 93086 225664 210054 225720
rect 210110 225664 210115 225720
rect 93025 225662 210115 225664
rect 93025 225659 93091 225662
rect 210049 225659 210115 225662
rect 396441 225722 396507 225725
rect 534073 225722 534139 225725
rect 396441 225720 534139 225722
rect 396441 225664 396446 225720
rect 396502 225664 534078 225720
rect 534134 225664 534139 225720
rect 396441 225662 534139 225664
rect 396441 225659 396507 225662
rect 534073 225659 534139 225662
rect 89529 225586 89595 225589
rect 208669 225586 208735 225589
rect 89529 225584 208735 225586
rect 89529 225528 89534 225584
rect 89590 225528 208674 225584
rect 208730 225528 208735 225584
rect 89529 225526 208735 225528
rect 89529 225523 89595 225526
rect 208669 225523 208735 225526
rect 400489 225586 400555 225589
rect 544009 225586 544075 225589
rect 400489 225584 544075 225586
rect 400489 225528 400494 225584
rect 400550 225528 544014 225584
rect 544070 225528 544075 225584
rect 400489 225526 544075 225528
rect 400489 225523 400555 225526
rect 544009 225523 544075 225526
rect 377673 224770 377739 224773
rect 490189 224770 490255 224773
rect 377673 224768 490255 224770
rect 377673 224712 377678 224768
rect 377734 224712 490194 224768
rect 490250 224712 490255 224768
rect 377673 224710 490255 224712
rect 377673 224707 377739 224710
rect 490189 224707 490255 224710
rect 78489 224634 78555 224637
rect 202597 224634 202663 224637
rect 78489 224632 202663 224634
rect 78489 224576 78494 224632
rect 78550 224576 202602 224632
rect 202658 224576 202663 224632
rect 78489 224574 202663 224576
rect 78489 224571 78555 224574
rect 202597 224571 202663 224574
rect 381905 224634 381971 224637
rect 499573 224634 499639 224637
rect 381905 224632 499639 224634
rect 381905 224576 381910 224632
rect 381966 224576 499578 224632
rect 499634 224576 499639 224632
rect 381905 224574 499639 224576
rect 381905 224571 381971 224574
rect 499573 224571 499639 224574
rect 72049 224498 72115 224501
rect 199745 224498 199811 224501
rect 72049 224496 199811 224498
rect 72049 224440 72054 224496
rect 72110 224440 199750 224496
rect 199806 224440 199811 224496
rect 72049 224438 199811 224440
rect 72049 224435 72115 224438
rect 199745 224435 199811 224438
rect 384021 224498 384087 224501
rect 505369 224498 505435 224501
rect 384021 224496 505435 224498
rect 384021 224440 384026 224496
rect 384082 224440 505374 224496
rect 505430 224440 505435 224496
rect 384021 224438 505435 224440
rect 384021 224435 384087 224438
rect 505369 224435 505435 224438
rect 69473 224362 69539 224365
rect 200113 224362 200179 224365
rect 69473 224360 200179 224362
rect 69473 224304 69478 224360
rect 69534 224304 200118 224360
rect 200174 224304 200179 224360
rect 69473 224302 200179 224304
rect 69473 224299 69539 224302
rect 200113 224299 200179 224302
rect 401133 224362 401199 224365
rect 545757 224362 545823 224365
rect 401133 224360 545823 224362
rect 401133 224304 401138 224360
rect 401194 224304 545762 224360
rect 545818 224304 545823 224360
rect 401133 224302 545823 224304
rect 401133 224299 401199 224302
rect 545757 224299 545823 224302
rect 61929 224226 61995 224229
rect 195421 224226 195487 224229
rect 61929 224224 195487 224226
rect 61929 224168 61934 224224
rect 61990 224168 195426 224224
rect 195482 224168 195487 224224
rect 61929 224166 195487 224168
rect 61929 224163 61995 224166
rect 195421 224163 195487 224166
rect 406101 224226 406167 224229
rect 556705 224226 556771 224229
rect 406101 224224 556771 224226
rect 406101 224168 406106 224224
rect 406162 224168 556710 224224
rect 556766 224168 556771 224224
rect 406101 224166 556771 224168
rect 406101 224163 406167 224166
rect 556705 224163 556771 224166
rect 675937 223546 676003 223549
rect 675937 223544 676292 223546
rect 675937 223488 675942 223544
rect 675998 223488 676292 223544
rect 675937 223486 676292 223488
rect 675937 223483 676003 223486
rect 99005 223274 99071 223277
rect 211153 223274 211219 223277
rect 99005 223272 211219 223274
rect 99005 223216 99010 223272
rect 99066 223216 211158 223272
rect 211214 223216 211219 223272
rect 99005 223214 211219 223216
rect 99005 223211 99071 223214
rect 211153 223211 211219 223214
rect 376201 223274 376267 223277
rect 487797 223274 487863 223277
rect 376201 223272 487863 223274
rect 376201 223216 376206 223272
rect 376262 223216 487802 223272
rect 487858 223216 487863 223272
rect 376201 223214 487863 223216
rect 376201 223211 376267 223214
rect 487797 223211 487863 223214
rect 92289 223138 92355 223141
rect 208025 223138 208091 223141
rect 92289 223136 208091 223138
rect 92289 223080 92294 223136
rect 92350 223080 208030 223136
rect 208086 223080 208091 223136
rect 92289 223078 208091 223080
rect 92289 223075 92355 223078
rect 208025 223075 208091 223078
rect 379053 223138 379119 223141
rect 494145 223138 494211 223141
rect 379053 223136 494211 223138
rect 379053 223080 379058 223136
rect 379114 223080 494150 223136
rect 494206 223080 494211 223136
rect 379053 223078 494211 223080
rect 379053 223075 379119 223078
rect 494145 223075 494211 223078
rect 676029 223138 676095 223141
rect 676029 223136 676292 223138
rect 676029 223080 676034 223136
rect 676090 223080 676292 223136
rect 676029 223078 676292 223080
rect 676029 223075 676095 223078
rect 58617 223002 58683 223005
rect 194041 223002 194107 223005
rect 58617 223000 194107 223002
rect 58617 222944 58622 223000
rect 58678 222944 194046 223000
rect 194102 222944 194107 223000
rect 58617 222942 194107 222944
rect 58617 222939 58683 222942
rect 194041 222939 194107 222942
rect 389357 223002 389423 223005
rect 517973 223002 518039 223005
rect 389357 223000 518039 223002
rect 389357 222944 389362 223000
rect 389418 222944 517978 223000
rect 518034 222944 518039 223000
rect 389357 222942 518039 222944
rect 389357 222939 389423 222942
rect 517973 222939 518039 222942
rect 55121 222866 55187 222869
rect 192385 222866 192451 222869
rect 55121 222864 192451 222866
rect 55121 222808 55126 222864
rect 55182 222808 192390 222864
rect 192446 222808 192451 222864
rect 55121 222806 192451 222808
rect 55121 222803 55187 222806
rect 192385 222803 192451 222806
rect 390461 222866 390527 222869
rect 520457 222866 520523 222869
rect 390461 222864 520523 222866
rect 390461 222808 390466 222864
rect 390522 222808 520462 222864
rect 520518 222808 520523 222864
rect 390461 222806 520523 222808
rect 390461 222803 390527 222806
rect 520457 222803 520523 222806
rect 675845 222730 675911 222733
rect 675845 222728 676292 222730
rect 675845 222672 675850 222728
rect 675906 222672 676292 222728
rect 675845 222670 676292 222672
rect 675845 222667 675911 222670
rect 676029 222322 676095 222325
rect 676029 222320 676292 222322
rect 676029 222264 676034 222320
rect 676090 222264 676292 222320
rect 676029 222262 676292 222264
rect 676029 222259 676095 222262
rect 73705 221914 73771 221917
rect 200573 221914 200639 221917
rect 73705 221912 200639 221914
rect 73705 221856 73710 221912
rect 73766 221856 200578 221912
rect 200634 221856 200639 221912
rect 73705 221854 200639 221856
rect 73705 221851 73771 221854
rect 200573 221851 200639 221854
rect 400673 221914 400739 221917
rect 528093 221914 528159 221917
rect 400673 221912 528159 221914
rect 400673 221856 400678 221912
rect 400734 221856 528098 221912
rect 528154 221856 528159 221912
rect 400673 221854 528159 221856
rect 400673 221851 400739 221854
rect 528093 221851 528159 221854
rect 676029 221914 676095 221917
rect 676029 221912 676292 221914
rect 676029 221856 676034 221912
rect 676090 221856 676292 221912
rect 676029 221854 676292 221856
rect 676029 221851 676095 221854
rect 70209 221778 70275 221781
rect 199101 221778 199167 221781
rect 70209 221776 199167 221778
rect 70209 221720 70214 221776
rect 70270 221720 199106 221776
rect 199162 221720 199167 221776
rect 70209 221718 199167 221720
rect 70209 221715 70275 221718
rect 199101 221715 199167 221718
rect 392853 221778 392919 221781
rect 525885 221778 525951 221781
rect 392853 221776 525951 221778
rect 392853 221720 392858 221776
rect 392914 221720 525890 221776
rect 525946 221720 525951 221776
rect 392853 221718 525951 221720
rect 392853 221715 392919 221718
rect 525885 221715 525951 221718
rect 66989 221642 67055 221645
rect 197721 221642 197787 221645
rect 66989 221640 197787 221642
rect 66989 221584 66994 221640
rect 67050 221584 197726 221640
rect 197782 221584 197787 221640
rect 66989 221582 197787 221584
rect 66989 221579 67055 221582
rect 197721 221579 197787 221582
rect 397177 221642 397243 221645
rect 536005 221642 536071 221645
rect 397177 221640 536071 221642
rect 397177 221584 397182 221640
rect 397238 221584 536010 221640
rect 536066 221584 536071 221640
rect 397177 221582 536071 221584
rect 397177 221579 397243 221582
rect 536005 221579 536071 221582
rect 56869 221506 56935 221509
rect 193397 221506 193463 221509
rect 56869 221504 193463 221506
rect 56869 221448 56874 221504
rect 56930 221448 193402 221504
rect 193458 221448 193463 221504
rect 56869 221446 193463 221448
rect 56869 221443 56935 221446
rect 193397 221443 193463 221446
rect 404997 221506 405063 221509
rect 546677 221506 546743 221509
rect 404997 221504 546743 221506
rect 404997 221448 405002 221504
rect 405058 221448 546682 221504
rect 546738 221448 546743 221504
rect 404997 221446 546743 221448
rect 404997 221443 405063 221446
rect 546677 221443 546743 221446
rect 676029 221506 676095 221509
rect 676029 221504 676292 221506
rect 676029 221448 676034 221504
rect 676090 221448 676292 221504
rect 676029 221446 676292 221448
rect 676029 221443 676095 221446
rect 674741 221098 674807 221101
rect 674741 221096 676292 221098
rect 674741 221040 674746 221096
rect 674802 221040 676292 221096
rect 674741 221038 676292 221040
rect 674741 221035 674807 221038
rect 676029 220690 676095 220693
rect 676029 220688 676292 220690
rect 676029 220632 676034 220688
rect 676090 220632 676292 220688
rect 676029 220630 676292 220632
rect 676029 220627 676095 220630
rect 389173 220554 389239 220557
rect 495617 220554 495683 220557
rect 389173 220552 495683 220554
rect 389173 220496 389178 220552
rect 389234 220496 495622 220552
rect 495678 220496 495683 220552
rect 389173 220494 495683 220496
rect 389173 220491 389239 220494
rect 495617 220491 495683 220494
rect 380341 220418 380407 220421
rect 489453 220418 489519 220421
rect 380341 220416 489519 220418
rect 380341 220360 380346 220416
rect 380402 220360 489458 220416
rect 489514 220360 489519 220416
rect 380341 220358 489519 220360
rect 380341 220355 380407 220358
rect 489453 220355 489519 220358
rect 74441 220282 74507 220285
rect 201585 220282 201651 220285
rect 74441 220280 201651 220282
rect 74441 220224 74446 220280
rect 74502 220224 201590 220280
rect 201646 220224 201651 220280
rect 74441 220222 201651 220224
rect 74441 220219 74507 220222
rect 201585 220219 201651 220222
rect 382181 220282 382247 220285
rect 498653 220282 498719 220285
rect 382181 220280 498719 220282
rect 382181 220224 382186 220280
rect 382242 220224 498658 220280
rect 498714 220224 498719 220280
rect 382181 220222 498719 220224
rect 382181 220219 382247 220222
rect 498653 220219 498719 220222
rect 676029 220282 676095 220285
rect 676029 220280 676292 220282
rect 676029 220224 676034 220280
rect 676090 220224 676292 220280
rect 676029 220222 676292 220224
rect 676029 220219 676095 220222
rect 67541 220146 67607 220149
rect 196617 220146 196683 220149
rect 67541 220144 196683 220146
rect 67541 220088 67546 220144
rect 67602 220088 196622 220144
rect 196678 220088 196683 220144
rect 67541 220086 196683 220088
rect 67541 220083 67607 220086
rect 196617 220083 196683 220086
rect 384849 220146 384915 220149
rect 507209 220146 507275 220149
rect 384849 220144 507275 220146
rect 384849 220088 384854 220144
rect 384910 220088 507214 220144
rect 507270 220088 507275 220144
rect 384849 220086 507275 220088
rect 384849 220083 384915 220086
rect 507209 220083 507275 220086
rect 676029 219874 676095 219877
rect 676029 219872 676292 219874
rect 676029 219816 676034 219872
rect 676090 219816 676292 219872
rect 676029 219814 676292 219816
rect 676029 219811 676095 219814
rect 507209 219466 507275 219469
rect 623957 219466 624023 219469
rect 507209 219464 624023 219466
rect 507209 219408 507214 219464
rect 507270 219408 623962 219464
rect 624018 219408 624023 219464
rect 507209 219406 624023 219408
rect 507209 219403 507275 219406
rect 623957 219403 624023 219406
rect 676029 219466 676095 219469
rect 676029 219464 676292 219466
rect 676029 219408 676034 219464
rect 676090 219408 676292 219464
rect 676029 219406 676292 219408
rect 676029 219403 676095 219406
rect 676029 219058 676095 219061
rect 676029 219056 676292 219058
rect 676029 219000 676034 219056
rect 676090 219000 676292 219056
rect 676029 218998 676292 219000
rect 676029 218995 676095 218998
rect 117957 218650 118023 218653
rect 663885 218650 663951 218653
rect 117957 218648 663951 218650
rect 117957 218592 117962 218648
rect 118018 218592 663890 218648
rect 663946 218592 663951 218648
rect 117957 218590 663951 218592
rect 117957 218587 118023 218590
rect 663885 218587 663951 218590
rect 675886 218588 675892 218652
rect 675956 218650 675962 218652
rect 675956 218590 676292 218650
rect 675956 218588 675962 218590
rect 675702 218180 675708 218244
rect 675772 218242 675778 218244
rect 675772 218182 676292 218242
rect 675772 218180 675778 218182
rect 675518 217772 675524 217836
rect 675588 217834 675594 217836
rect 675588 217774 676292 217834
rect 675588 217772 675594 217774
rect 679617 217426 679683 217429
rect 679604 217424 679683 217426
rect 679604 217368 679622 217424
rect 679678 217368 679683 217424
rect 679604 217366 679683 217368
rect 679617 217363 679683 217366
rect 532969 217018 533035 217021
rect 628925 217018 628991 217021
rect 532969 217016 628991 217018
rect 532969 216960 532974 217016
rect 533030 216960 628930 217016
rect 628986 216960 628991 217016
rect 532969 216958 628991 216960
rect 532969 216955 533035 216958
rect 628925 216955 628991 216958
rect 675845 217018 675911 217021
rect 675845 217016 676292 217018
rect 675845 216960 675850 217016
rect 675906 216960 676292 217016
rect 675845 216958 676292 216960
rect 675845 216955 675911 216958
rect 492581 216882 492647 216885
rect 622025 216882 622091 216885
rect 492581 216880 622091 216882
rect 492581 216824 492586 216880
rect 492642 216824 622030 216880
rect 622086 216824 622091 216880
rect 492581 216822 622091 216824
rect 492581 216819 492647 216822
rect 622025 216819 622091 216822
rect 489085 216746 489151 216749
rect 620921 216746 620987 216749
rect 489085 216744 620987 216746
rect 489085 216688 489090 216744
rect 489146 216688 620926 216744
rect 620982 216688 620987 216744
rect 489085 216686 620987 216688
rect 489085 216683 489151 216686
rect 620921 216683 620987 216686
rect 676029 216610 676095 216613
rect 676029 216608 676292 216610
rect 676029 216552 676034 216608
rect 676090 216552 676292 216608
rect 676029 216550 676292 216552
rect 676029 216547 676095 216550
rect 578877 216202 578943 216205
rect 576380 216200 578943 216202
rect 576380 216144 578882 216200
rect 578938 216144 578943 216200
rect 576380 216142 578943 216144
rect 578877 216139 578943 216142
rect 676029 216202 676095 216205
rect 676029 216200 676292 216202
rect 676029 216144 676034 216200
rect 676090 216144 676292 216200
rect 676029 216142 676292 216144
rect 676029 216139 676095 216142
rect 676029 215794 676095 215797
rect 676029 215792 676292 215794
rect 676029 215736 676034 215792
rect 676090 215736 676292 215792
rect 676029 215734 676292 215736
rect 676029 215731 676095 215734
rect 676622 215494 676628 215558
rect 676692 215494 676698 215558
rect 676630 215356 676690 215494
rect 28717 215114 28783 215117
rect 28717 215112 28826 215114
rect 28717 215056 28722 215112
rect 28778 215056 28826 215112
rect 28717 215051 28826 215056
rect 28766 214948 28826 215051
rect 675937 214978 676003 214981
rect 675937 214976 676292 214978
rect 675937 214920 675942 214976
rect 675998 214920 676292 214976
rect 675937 214918 676292 214920
rect 675937 214915 676003 214918
rect 35801 214706 35867 214709
rect 579245 214706 579311 214709
rect 35758 214704 35867 214706
rect 35758 214648 35806 214704
rect 35862 214648 35867 214704
rect 35758 214643 35867 214648
rect 576380 214704 579311 214706
rect 576380 214648 579250 214704
rect 579306 214648 579311 214704
rect 576380 214646 579311 214648
rect 579245 214643 579311 214646
rect 35758 214540 35818 214643
rect 676998 214334 677058 214540
rect 35801 214298 35867 214301
rect 35758 214296 35867 214298
rect 35758 214240 35806 214296
rect 35862 214240 35867 214296
rect 676990 214270 676996 214334
rect 677060 214270 677066 214334
rect 35758 214235 35867 214240
rect 35758 214132 35818 214235
rect 676029 214162 676095 214165
rect 676029 214160 676292 214162
rect 676029 214104 676034 214160
rect 676090 214104 676292 214160
rect 676029 214102 676292 214104
rect 676029 214099 676095 214102
rect 676029 214028 676095 214029
rect 676029 214026 676076 214028
rect 675984 214024 676076 214026
rect 675984 213968 676034 214024
rect 675984 213966 676076 213968
rect 676029 213964 676076 213966
rect 676140 213964 676146 214028
rect 676029 213963 676095 213964
rect 42885 213754 42951 213757
rect 41492 213752 42951 213754
rect 41492 213696 42890 213752
rect 42946 213696 42951 213752
rect 41492 213694 42951 213696
rect 42885 213691 42951 213694
rect 676029 213754 676095 213757
rect 676029 213752 676292 213754
rect 676029 213696 676034 213752
rect 676090 213696 676292 213752
rect 676029 213694 676292 213696
rect 676029 213691 676095 213694
rect 41505 213482 41571 213485
rect 41462 213480 41571 213482
rect 41462 213424 41510 213480
rect 41566 213424 41571 213480
rect 41462 213419 41571 213424
rect 41462 213316 41522 213419
rect 676029 213346 676095 213349
rect 676029 213344 676292 213346
rect 676029 213288 676034 213344
rect 676090 213288 676292 213344
rect 676029 213286 676292 213288
rect 676029 213283 676095 213286
rect 578969 213210 579035 213213
rect 576380 213208 579035 213210
rect 576380 213152 578974 213208
rect 579030 213152 579035 213208
rect 576380 213150 579035 213152
rect 578969 213147 579035 213150
rect 646446 213012 646452 213076
rect 646516 213074 646522 213076
rect 647141 213074 647207 213077
rect 646516 213072 647207 213074
rect 646516 213016 647146 213072
rect 647202 213016 647207 213072
rect 646516 213014 647207 213016
rect 646516 213012 646522 213014
rect 647141 213011 647207 213014
rect 647366 213012 647372 213076
rect 647436 213074 647442 213076
rect 648521 213074 648587 213077
rect 647436 213072 648587 213074
rect 647436 213016 648526 213072
rect 648582 213016 648587 213072
rect 647436 213014 648587 213016
rect 647436 213012 647442 213014
rect 648521 213011 648587 213014
rect 43345 212938 43411 212941
rect 41492 212936 43411 212938
rect 41492 212880 43350 212936
rect 43406 212880 43411 212936
rect 41492 212878 43411 212880
rect 43345 212875 43411 212878
rect 47209 212530 47275 212533
rect 41492 212528 47275 212530
rect 41492 212472 47214 212528
rect 47270 212472 47275 212528
rect 676262 212500 676322 212908
rect 41492 212470 47275 212472
rect 47209 212467 47275 212470
rect 44265 212122 44331 212125
rect 41492 212120 44331 212122
rect 41492 212064 44270 212120
rect 44326 212064 44331 212120
rect 41492 212062 44331 212064
rect 44265 212059 44331 212062
rect 676029 212122 676095 212125
rect 676029 212120 676292 212122
rect 676029 212064 676034 212120
rect 676090 212064 676292 212120
rect 676029 212062 676292 212064
rect 676029 212059 676095 212062
rect 41321 211850 41387 211853
rect 41278 211848 41387 211850
rect 41278 211792 41326 211848
rect 41382 211792 41387 211848
rect 41278 211787 41387 211792
rect 41278 211684 41338 211787
rect 578417 211714 578483 211717
rect 576380 211712 578483 211714
rect 576380 211656 578422 211712
rect 578478 211656 578483 211712
rect 576380 211654 578483 211656
rect 578417 211651 578483 211654
rect 675937 211442 676003 211445
rect 676806 211442 676812 211444
rect 675937 211440 676812 211442
rect 675937 211384 675942 211440
rect 675998 211384 676812 211440
rect 675937 211382 676812 211384
rect 675937 211379 676003 211382
rect 676806 211380 676812 211382
rect 676876 211380 676882 211444
rect 44725 211306 44791 211309
rect 41492 211304 44791 211306
rect 41492 211248 44730 211304
rect 44786 211248 44791 211304
rect 41492 211246 44791 211248
rect 44725 211243 44791 211246
rect 675845 211306 675911 211309
rect 676438 211306 676444 211308
rect 675845 211304 676444 211306
rect 675845 211248 675850 211304
rect 675906 211248 676444 211304
rect 675845 211246 676444 211248
rect 675845 211243 675911 211246
rect 676438 211244 676444 211246
rect 676508 211244 676514 211308
rect 41462 210626 41522 210868
rect 50061 210626 50127 210629
rect 41462 210624 50127 210626
rect 41462 210568 50066 210624
rect 50122 210568 50127 210624
rect 41462 210566 50127 210568
rect 50061 210563 50127 210566
rect 30974 210221 31034 210460
rect 30974 210216 31083 210221
rect 578509 210218 578575 210221
rect 30974 210160 31022 210216
rect 31078 210160 31083 210216
rect 30974 210158 31083 210160
rect 576380 210216 578575 210218
rect 576380 210160 578514 210216
rect 578570 210160 578575 210216
rect 576380 210158 578575 210160
rect 31017 210155 31083 210158
rect 578509 210155 578575 210158
rect 41462 209810 41522 210052
rect 675702 209884 675708 209948
rect 675772 209884 675778 209948
rect 41638 209810 41644 209812
rect 41462 209750 41644 209810
rect 41638 209748 41644 209750
rect 41708 209748 41714 209812
rect 665449 209810 665515 209813
rect 665449 209808 666570 209810
rect 665449 209752 665454 209808
rect 665510 209752 666570 209808
rect 665449 209750 666570 209752
rect 665449 209747 665515 209750
rect 40542 209404 40602 209644
rect 603073 209538 603139 209541
rect 666510 209538 666570 209750
rect 675710 209674 675770 209884
rect 675886 209674 675892 209676
rect 675710 209614 675892 209674
rect 675886 209612 675892 209614
rect 675956 209612 675962 209676
rect 603073 209536 606556 209538
rect 603073 209480 603078 209536
rect 603134 209480 606556 209536
rect 603073 209478 606556 209480
rect 666510 209478 666754 209538
rect 603073 209475 603139 209478
rect 40534 209340 40540 209404
rect 40604 209340 40610 209404
rect 42793 209266 42859 209269
rect 666694 209266 666754 209478
rect 667933 209266 667999 209269
rect 41492 209264 42859 209266
rect 41492 209208 42798 209264
rect 42854 209208 42859 209264
rect 41492 209206 42859 209208
rect 666356 209264 667999 209266
rect 666356 209208 667938 209264
rect 667994 209208 667999 209264
rect 666356 209206 667999 209208
rect 42793 209203 42859 209206
rect 667933 209203 667999 209206
rect 39297 208586 39363 208589
rect 41462 208588 41522 208828
rect 579521 208722 579587 208725
rect 576380 208720 579587 208722
rect 576380 208664 579526 208720
rect 579582 208664 579587 208720
rect 576380 208662 579587 208664
rect 579521 208659 579587 208662
rect 39254 208584 39363 208586
rect 39254 208528 39302 208584
rect 39358 208528 39363 208584
rect 39254 208523 39363 208528
rect 41454 208524 41460 208588
rect 41524 208524 41530 208588
rect 603165 208586 603231 208589
rect 603165 208584 606556 208586
rect 603165 208528 603170 208584
rect 603226 208528 606556 208584
rect 603165 208526 606556 208528
rect 603165 208523 603231 208526
rect 39254 208420 39314 208523
rect 676070 208252 676076 208316
rect 676140 208314 676146 208316
rect 676857 208314 676923 208317
rect 676140 208312 676923 208314
rect 676140 208256 676862 208312
rect 676918 208256 676923 208312
rect 676140 208254 676923 208256
rect 676140 208252 676146 208254
rect 676857 208251 676923 208254
rect 44173 208042 44239 208045
rect 41492 208040 44239 208042
rect 41492 207984 44178 208040
rect 44234 207984 44239 208040
rect 41492 207982 44239 207984
rect 44173 207979 44239 207982
rect 42885 207634 42951 207637
rect 41492 207632 42951 207634
rect 41492 207576 42890 207632
rect 42946 207576 42951 207632
rect 41492 207574 42951 207576
rect 42885 207571 42951 207574
rect 603073 207498 603139 207501
rect 603073 207496 606556 207498
rect 603073 207440 603078 207496
rect 603134 207440 606556 207496
rect 603073 207438 606556 207440
rect 603073 207435 603139 207438
rect 578785 207226 578851 207229
rect 576380 207224 578851 207226
rect 40726 206956 40786 207196
rect 576380 207168 578790 207224
rect 578846 207168 578851 207224
rect 576380 207166 578851 207168
rect 578785 207163 578851 207166
rect 675334 207164 675340 207228
rect 675404 207226 675410 207228
rect 679617 207226 679683 207229
rect 675404 207224 679683 207226
rect 675404 207168 679622 207224
rect 679678 207168 679683 207224
rect 675404 207166 679683 207168
rect 675404 207164 675410 207166
rect 679617 207163 679683 207166
rect 40718 206892 40724 206956
rect 40788 206892 40794 206956
rect 43345 206818 43411 206821
rect 41492 206816 43411 206818
rect 41492 206760 43350 206816
rect 43406 206760 43411 206816
rect 41492 206758 43411 206760
rect 43345 206755 43411 206758
rect 603073 206546 603139 206549
rect 603073 206544 606556 206546
rect 603073 206488 603078 206544
rect 603134 206488 606556 206544
rect 603073 206486 606556 206488
rect 603073 206483 603139 206486
rect 43161 206410 43227 206413
rect 41492 206408 43227 206410
rect 41492 206352 43166 206408
rect 43222 206352 43227 206408
rect 41492 206350 43227 206352
rect 43161 206347 43227 206350
rect 42977 206002 43043 206005
rect 41492 206000 43043 206002
rect 41492 205944 42982 206000
rect 43038 205944 43043 206000
rect 41492 205942 43043 205944
rect 42977 205939 43043 205942
rect 667933 205866 667999 205869
rect 666356 205864 667999 205866
rect 666356 205808 667938 205864
rect 667994 205808 667999 205864
rect 666356 205806 667999 205808
rect 667933 205803 667999 205806
rect 579429 205730 579495 205733
rect 576380 205728 579495 205730
rect 576380 205672 579434 205728
rect 579490 205672 579495 205728
rect 576380 205670 579495 205672
rect 579429 205667 579495 205670
rect 43437 205594 43503 205597
rect 41492 205592 43503 205594
rect 41492 205536 43442 205592
rect 43498 205536 43503 205592
rect 41492 205534 43503 205536
rect 43437 205531 43503 205534
rect 675753 205594 675819 205597
rect 675886 205594 675892 205596
rect 675753 205592 675892 205594
rect 675753 205536 675758 205592
rect 675814 205536 675892 205592
rect 675753 205534 675892 205536
rect 675753 205531 675819 205534
rect 675886 205532 675892 205534
rect 675956 205532 675962 205596
rect 603073 205458 603139 205461
rect 603073 205456 606556 205458
rect 603073 205400 603078 205456
rect 603134 205400 606556 205456
rect 603073 205398 606556 205400
rect 603073 205395 603139 205398
rect 43253 205186 43319 205189
rect 41492 205184 43319 205186
rect 41492 205128 43258 205184
rect 43314 205128 43319 205184
rect 41492 205126 43319 205128
rect 43253 205123 43319 205126
rect 675753 205050 675819 205053
rect 676070 205050 676076 205052
rect 675753 205048 676076 205050
rect 675753 204992 675758 205048
rect 675814 204992 676076 205048
rect 675753 204990 676076 204992
rect 675753 204987 675819 204990
rect 676070 204988 676076 204990
rect 676140 204988 676146 205052
rect 31293 204914 31359 204917
rect 31293 204912 31402 204914
rect 31293 204856 31298 204912
rect 31354 204856 31402 204912
rect 31293 204851 31402 204856
rect 31342 204748 31402 204851
rect 31109 204506 31175 204509
rect 603165 204506 603231 204509
rect 31109 204504 31218 204506
rect 31109 204448 31114 204504
rect 31170 204448 31218 204504
rect 31109 204443 31218 204448
rect 603165 204504 606556 204506
rect 603165 204448 603170 204504
rect 603226 204448 606556 204504
rect 603165 204446 606556 204448
rect 603165 204443 603231 204446
rect 31158 204340 31218 204443
rect 578877 204234 578943 204237
rect 666829 204234 666895 204237
rect 675753 204236 675819 204237
rect 675702 204234 675708 204236
rect 576380 204232 578943 204234
rect 576380 204176 578882 204232
rect 578938 204176 578943 204232
rect 576380 204174 578943 204176
rect 666356 204232 666895 204234
rect 666356 204176 666834 204232
rect 666890 204176 666895 204232
rect 666356 204174 666895 204176
rect 675662 204174 675708 204234
rect 675772 204232 675819 204236
rect 675814 204176 675819 204232
rect 578877 204171 578943 204174
rect 666829 204171 666895 204174
rect 675702 204172 675708 204174
rect 675772 204172 675819 204176
rect 675753 204171 675819 204172
rect 35758 203285 35818 203524
rect 603073 203418 603139 203421
rect 603073 203416 606556 203418
rect 603073 203360 603078 203416
rect 603134 203360 606556 203416
rect 603073 203358 606556 203360
rect 603073 203355 603139 203358
rect 35758 203280 35867 203285
rect 35758 203224 35806 203280
rect 35862 203224 35867 203280
rect 35758 203222 35867 203224
rect 35801 203219 35867 203222
rect 675109 202874 675175 202877
rect 676990 202874 676996 202876
rect 675109 202872 676996 202874
rect 675109 202816 675114 202872
rect 675170 202816 676996 202872
rect 675109 202814 676996 202816
rect 675109 202811 675175 202814
rect 676990 202812 676996 202814
rect 677060 202812 677066 202876
rect 579245 202738 579311 202741
rect 576380 202736 579311 202738
rect 576380 202680 579250 202736
rect 579306 202680 579311 202736
rect 576380 202678 579311 202680
rect 579245 202675 579311 202678
rect 675477 202740 675543 202741
rect 675477 202736 675524 202740
rect 675588 202738 675594 202740
rect 675477 202680 675482 202736
rect 675477 202676 675524 202680
rect 675588 202678 675634 202738
rect 675588 202676 675594 202678
rect 675477 202675 675543 202676
rect 603073 202466 603139 202469
rect 603073 202464 606556 202466
rect 603073 202408 603078 202464
rect 603134 202408 606556 202464
rect 603073 202406 606556 202408
rect 603073 202403 603139 202406
rect 603073 201378 603139 201381
rect 674833 201378 674899 201381
rect 676806 201378 676812 201380
rect 603073 201376 606556 201378
rect 603073 201320 603078 201376
rect 603134 201320 606556 201376
rect 603073 201318 606556 201320
rect 674833 201376 676812 201378
rect 674833 201320 674838 201376
rect 674894 201320 676812 201376
rect 674833 201318 676812 201320
rect 603073 201315 603139 201318
rect 674833 201315 674899 201318
rect 676806 201316 676812 201318
rect 676876 201316 676882 201380
rect 578233 201242 578299 201245
rect 576380 201240 578299 201242
rect 576380 201184 578238 201240
rect 578294 201184 578299 201240
rect 576380 201182 578299 201184
rect 578233 201179 578299 201182
rect 666829 200834 666895 200837
rect 666356 200832 666895 200834
rect 666356 200776 666834 200832
rect 666890 200776 666895 200832
rect 666356 200774 666895 200776
rect 666829 200771 666895 200774
rect 603165 200426 603231 200429
rect 603165 200424 606556 200426
rect 603165 200368 603170 200424
rect 603226 200368 606556 200424
rect 603165 200366 606556 200368
rect 603165 200363 603231 200366
rect 578417 199746 578483 199749
rect 576380 199744 578483 199746
rect 576380 199688 578422 199744
rect 578478 199688 578483 199744
rect 576380 199686 578483 199688
rect 578417 199683 578483 199686
rect 31017 199338 31083 199341
rect 41822 199338 41828 199340
rect 31017 199336 41828 199338
rect 31017 199280 31022 199336
rect 31078 199280 41828 199336
rect 31017 199278 41828 199280
rect 31017 199275 31083 199278
rect 41822 199276 41828 199278
rect 41892 199276 41898 199340
rect 603073 199338 603139 199341
rect 603073 199336 606556 199338
rect 603073 199280 603078 199336
rect 603134 199280 606556 199336
rect 603073 199278 606556 199280
rect 603073 199275 603139 199278
rect 666737 199066 666803 199069
rect 667933 199066 667999 199069
rect 666356 199064 667999 199066
rect 666356 199008 666742 199064
rect 666798 199008 667938 199064
rect 667994 199008 667999 199064
rect 666356 199006 667999 199008
rect 666737 199003 666803 199006
rect 667933 199003 667999 199006
rect 603073 198386 603139 198389
rect 675753 198386 675819 198389
rect 676070 198386 676076 198388
rect 603073 198384 606556 198386
rect 603073 198328 603078 198384
rect 603134 198328 606556 198384
rect 603073 198326 606556 198328
rect 675753 198384 676076 198386
rect 675753 198328 675758 198384
rect 675814 198328 676076 198384
rect 675753 198326 676076 198328
rect 603073 198323 603139 198326
rect 675753 198323 675819 198326
rect 676070 198324 676076 198326
rect 676140 198324 676146 198388
rect 579061 198250 579127 198253
rect 576380 198248 579127 198250
rect 576380 198192 579066 198248
rect 579122 198192 579127 198248
rect 576380 198190 579127 198192
rect 579061 198187 579127 198190
rect 39297 197706 39363 197709
rect 39297 197704 41890 197706
rect 39297 197648 39302 197704
rect 39358 197648 41890 197704
rect 39297 197646 41890 197648
rect 39297 197643 39363 197646
rect 41830 197165 41890 197646
rect 603073 197298 603139 197301
rect 603073 197296 606556 197298
rect 603073 197240 603078 197296
rect 603134 197240 606556 197296
rect 603073 197238 606556 197240
rect 603073 197235 603139 197238
rect 41830 197160 41939 197165
rect 41830 197104 41878 197160
rect 41934 197104 41939 197160
rect 41830 197102 41939 197104
rect 41873 197099 41939 197102
rect 579521 196754 579587 196757
rect 576380 196752 579587 196754
rect 576380 196696 579526 196752
rect 579582 196696 579587 196752
rect 576380 196694 579587 196696
rect 579521 196691 579587 196694
rect 603165 196346 603231 196349
rect 603165 196344 606556 196346
rect 603165 196288 603170 196344
rect 603226 196288 606556 196344
rect 603165 196286 606556 196288
rect 603165 196283 603231 196286
rect 667933 195666 667999 195669
rect 666356 195664 667999 195666
rect 666356 195608 667938 195664
rect 667994 195608 667999 195664
rect 666356 195606 667999 195608
rect 667933 195603 667999 195606
rect 40718 195332 40724 195396
rect 40788 195394 40794 195396
rect 42190 195394 42196 195396
rect 40788 195334 42196 195394
rect 40788 195332 40794 195334
rect 42190 195332 42196 195334
rect 42260 195332 42266 195396
rect 675753 195394 675819 195397
rect 676622 195394 676628 195396
rect 675753 195392 676628 195394
rect 675753 195336 675758 195392
rect 675814 195336 676628 195392
rect 675753 195334 676628 195336
rect 675753 195331 675819 195334
rect 676622 195332 676628 195334
rect 676692 195332 676698 195396
rect 41638 195196 41644 195260
rect 41708 195258 41714 195260
rect 41781 195258 41847 195261
rect 579521 195258 579587 195261
rect 41708 195256 41847 195258
rect 41708 195200 41786 195256
rect 41842 195200 41847 195256
rect 41708 195198 41847 195200
rect 576380 195256 579587 195258
rect 576380 195200 579526 195256
rect 579582 195200 579587 195256
rect 576380 195198 579587 195200
rect 41708 195196 41714 195198
rect 41781 195195 41847 195198
rect 579521 195195 579587 195198
rect 603073 195258 603139 195261
rect 603073 195256 606556 195258
rect 603073 195200 603078 195256
rect 603134 195200 606556 195256
rect 603073 195198 606556 195200
rect 603073 195195 603139 195198
rect 603073 194306 603139 194309
rect 603073 194304 606556 194306
rect 603073 194248 603078 194304
rect 603134 194248 606556 194304
rect 603073 194246 606556 194248
rect 603073 194243 603139 194246
rect 666553 194034 666619 194037
rect 666356 194032 666619 194034
rect 666356 193976 666558 194032
rect 666614 193976 666619 194032
rect 666356 193974 666619 193976
rect 666553 193971 666619 193974
rect 579521 193626 579587 193629
rect 576380 193624 579587 193626
rect 576380 193568 579526 193624
rect 579582 193568 579587 193624
rect 576380 193566 579587 193568
rect 579521 193563 579587 193566
rect 603073 193218 603139 193221
rect 603073 193216 606556 193218
rect 603073 193160 603078 193216
rect 603134 193160 606556 193216
rect 603073 193158 606556 193160
rect 603073 193155 603139 193158
rect 603073 192266 603139 192269
rect 603073 192264 606556 192266
rect 603073 192208 603078 192264
rect 603134 192208 606556 192264
rect 603073 192206 606556 192208
rect 603073 192203 603139 192206
rect 579521 192130 579587 192133
rect 576380 192128 579587 192130
rect 576380 192072 579526 192128
rect 579582 192072 579587 192128
rect 576380 192070 579587 192072
rect 579521 192067 579587 192070
rect 603073 191178 603139 191181
rect 603073 191176 606556 191178
rect 603073 191120 603078 191176
rect 603134 191120 606556 191176
rect 603073 191118 606556 191120
rect 603073 191115 603139 191118
rect 579245 190634 579311 190637
rect 666553 190634 666619 190637
rect 576380 190632 579311 190634
rect 576380 190576 579250 190632
rect 579306 190576 579311 190632
rect 576380 190574 579311 190576
rect 666356 190632 666619 190634
rect 666356 190576 666558 190632
rect 666614 190576 666619 190632
rect 666356 190574 666619 190576
rect 579245 190571 579311 190574
rect 666553 190571 666619 190574
rect 675753 190362 675819 190365
rect 676438 190362 676444 190364
rect 675753 190360 676444 190362
rect 675753 190304 675758 190360
rect 675814 190304 676444 190360
rect 675753 190302 676444 190304
rect 675753 190299 675819 190302
rect 676438 190300 676444 190302
rect 676508 190300 676514 190364
rect 41454 190164 41460 190228
rect 41524 190226 41530 190228
rect 41781 190226 41847 190229
rect 41524 190224 41847 190226
rect 41524 190168 41786 190224
rect 41842 190168 41847 190224
rect 41524 190166 41847 190168
rect 41524 190164 41530 190166
rect 41781 190163 41847 190166
rect 603165 190226 603231 190229
rect 674833 190226 674899 190229
rect 676254 190226 676260 190228
rect 603165 190224 606556 190226
rect 603165 190168 603170 190224
rect 603226 190168 606556 190224
rect 603165 190166 606556 190168
rect 674833 190224 676260 190226
rect 674833 190168 674838 190224
rect 674894 190168 676260 190224
rect 674833 190166 676260 190168
rect 603165 190163 603231 190166
rect 674833 190163 674899 190166
rect 676254 190164 676260 190166
rect 676324 190164 676330 190228
rect 578233 189138 578299 189141
rect 576380 189136 578299 189138
rect 576380 189080 578238 189136
rect 578294 189080 578299 189136
rect 576380 189078 578299 189080
rect 578233 189075 578299 189078
rect 603073 189138 603139 189141
rect 603073 189136 606556 189138
rect 603073 189080 603078 189136
rect 603134 189080 606556 189136
rect 603073 189078 606556 189080
rect 603073 189075 603139 189078
rect 666553 189002 666619 189005
rect 666356 189000 666619 189002
rect 666356 188944 666558 189000
rect 666614 188944 666619 189000
rect 666356 188942 666619 188944
rect 666553 188939 666619 188942
rect 603073 188186 603139 188189
rect 603073 188184 606556 188186
rect 603073 188128 603078 188184
rect 603134 188128 606556 188184
rect 603073 188126 606556 188128
rect 603073 188123 603139 188126
rect 579245 187642 579311 187645
rect 576380 187640 579311 187642
rect 576380 187584 579250 187640
rect 579306 187584 579311 187640
rect 576380 187582 579311 187584
rect 579245 187579 579311 187582
rect 42149 187372 42215 187373
rect 42149 187370 42196 187372
rect 42104 187368 42196 187370
rect 42104 187312 42154 187368
rect 42104 187310 42196 187312
rect 42149 187308 42196 187310
rect 42260 187308 42266 187372
rect 42149 187307 42215 187308
rect 603073 187098 603139 187101
rect 603073 187096 606556 187098
rect 603073 187040 603078 187096
rect 603134 187040 606556 187096
rect 603073 187038 606556 187040
rect 603073 187035 603139 187038
rect 579521 186146 579587 186149
rect 576380 186144 579587 186146
rect 576380 186088 579526 186144
rect 579582 186088 579587 186144
rect 576380 186086 579587 186088
rect 579521 186083 579587 186086
rect 603165 186146 603231 186149
rect 603165 186144 606556 186146
rect 603165 186088 603170 186144
rect 603226 186088 606556 186144
rect 603165 186086 606556 186088
rect 603165 186083 603231 186086
rect 666553 185602 666619 185605
rect 666356 185600 666619 185602
rect 666356 185544 666558 185600
rect 666614 185544 666619 185600
rect 666356 185542 666619 185544
rect 666553 185539 666619 185542
rect 603073 185058 603139 185061
rect 603073 185056 606556 185058
rect 603073 185000 603078 185056
rect 603134 185000 606556 185056
rect 603073 184998 606556 185000
rect 603073 184995 603139 184998
rect 578877 184650 578943 184653
rect 576380 184648 578943 184650
rect 576380 184592 578882 184648
rect 578938 184592 578943 184648
rect 576380 184590 578943 184592
rect 578877 184587 578943 184590
rect 41873 184244 41939 184245
rect 41822 184242 41828 184244
rect 41782 184182 41828 184242
rect 41892 184240 41939 184244
rect 41934 184184 41939 184240
rect 41822 184180 41828 184182
rect 41892 184180 41939 184184
rect 41873 184179 41939 184180
rect 603073 184106 603139 184109
rect 603073 184104 606556 184106
rect 603073 184048 603078 184104
rect 603134 184048 606556 184104
rect 603073 184046 606556 184048
rect 603073 184043 603139 184046
rect 667933 183834 667999 183837
rect 666356 183832 667999 183834
rect 666356 183776 667938 183832
rect 667994 183776 667999 183832
rect 666356 183774 667999 183776
rect 667933 183771 667999 183774
rect 579429 183154 579495 183157
rect 576380 183152 579495 183154
rect 576380 183096 579434 183152
rect 579490 183096 579495 183152
rect 576380 183094 579495 183096
rect 579429 183091 579495 183094
rect 40534 182956 40540 183020
rect 40604 183018 40610 183020
rect 41781 183018 41847 183021
rect 40604 183016 41847 183018
rect 40604 182960 41786 183016
rect 41842 182960 41847 183016
rect 40604 182958 41847 182960
rect 40604 182956 40610 182958
rect 41781 182955 41847 182958
rect 603073 183018 603139 183021
rect 603073 183016 606556 183018
rect 603073 182960 603078 183016
rect 603134 182960 606556 183016
rect 603073 182958 606556 182960
rect 603073 182955 603139 182958
rect 603165 182066 603231 182069
rect 603165 182064 606556 182066
rect 603165 182008 603170 182064
rect 603226 182008 606556 182064
rect 603165 182006 606556 182008
rect 603165 182003 603231 182006
rect 579521 181658 579587 181661
rect 576380 181656 579587 181658
rect 576380 181600 579526 181656
rect 579582 181600 579587 181656
rect 576380 181598 579587 181600
rect 579521 181595 579587 181598
rect 603073 180978 603139 180981
rect 603073 180976 606556 180978
rect 603073 180920 603078 180976
rect 603134 180920 606556 180976
rect 603073 180918 606556 180920
rect 603073 180915 603139 180918
rect 668025 180434 668091 180437
rect 666356 180432 668091 180434
rect 666356 180376 668030 180432
rect 668086 180376 668091 180432
rect 666356 180374 668091 180376
rect 668025 180371 668091 180374
rect 578877 180162 578943 180165
rect 576380 180160 578943 180162
rect 576380 180104 578882 180160
rect 578938 180104 578943 180160
rect 576380 180102 578943 180104
rect 578877 180099 578943 180102
rect 603073 180026 603139 180029
rect 603073 180024 606556 180026
rect 603073 179968 603078 180024
rect 603134 179968 606556 180024
rect 603073 179966 606556 179968
rect 603073 179963 603139 179966
rect 603073 178938 603139 178941
rect 603073 178936 606556 178938
rect 603073 178880 603078 178936
rect 603134 178880 606556 178936
rect 603073 178878 606556 178880
rect 603073 178875 603139 178878
rect 667933 178802 667999 178805
rect 666356 178800 667999 178802
rect 666356 178744 667938 178800
rect 667994 178744 667999 178800
rect 666356 178742 667999 178744
rect 667933 178739 667999 178742
rect 579337 178666 579403 178669
rect 576380 178664 579403 178666
rect 576380 178608 579342 178664
rect 579398 178608 579403 178664
rect 576380 178606 579403 178608
rect 579337 178603 579403 178606
rect 675937 178530 676003 178533
rect 675937 178528 676292 178530
rect 675937 178472 675942 178528
rect 675998 178472 676292 178528
rect 675937 178470 676292 178472
rect 675937 178467 676003 178470
rect 676029 178122 676095 178125
rect 676029 178120 676292 178122
rect 676029 178064 676034 178120
rect 676090 178064 676292 178120
rect 676029 178062 676292 178064
rect 676029 178059 676095 178062
rect 603165 177986 603231 177989
rect 603165 177984 606556 177986
rect 603165 177928 603170 177984
rect 603226 177928 606556 177984
rect 603165 177926 606556 177928
rect 603165 177923 603231 177926
rect 675937 177714 676003 177717
rect 675937 177712 676292 177714
rect 675937 177656 675942 177712
rect 675998 177656 676292 177712
rect 675937 177654 676292 177656
rect 675937 177651 676003 177654
rect 676029 177306 676095 177309
rect 676029 177304 676292 177306
rect 676029 177248 676034 177304
rect 676090 177248 676292 177304
rect 676029 177246 676292 177248
rect 676029 177243 676095 177246
rect 578233 177170 578299 177173
rect 576380 177168 578299 177170
rect 576380 177112 578238 177168
rect 578294 177112 578299 177168
rect 576380 177110 578299 177112
rect 578233 177107 578299 177110
rect 603073 176898 603139 176901
rect 676029 176898 676095 176901
rect 603073 176896 606556 176898
rect 603073 176840 603078 176896
rect 603134 176840 606556 176896
rect 603073 176838 606556 176840
rect 676029 176896 676292 176898
rect 676029 176840 676034 176896
rect 676090 176840 676292 176896
rect 676029 176838 676292 176840
rect 603073 176835 603139 176838
rect 676029 176835 676095 176838
rect 674741 176490 674807 176493
rect 674741 176488 676292 176490
rect 674741 176432 674746 176488
rect 674802 176432 676292 176488
rect 674741 176430 676292 176432
rect 674741 176427 674807 176430
rect 676029 176082 676095 176085
rect 676029 176080 676292 176082
rect 676029 176024 676034 176080
rect 676090 176024 676292 176080
rect 676029 176022 676292 176024
rect 676029 176019 676095 176022
rect 603073 175946 603139 175949
rect 603073 175944 606556 175946
rect 603073 175888 603078 175944
rect 603134 175888 606556 175944
rect 603073 175886 606556 175888
rect 603073 175883 603139 175886
rect 578325 175674 578391 175677
rect 576380 175672 578391 175674
rect 576380 175616 578330 175672
rect 578386 175616 578391 175672
rect 576380 175614 578391 175616
rect 578325 175611 578391 175614
rect 676029 175674 676095 175677
rect 676029 175672 676292 175674
rect 676029 175616 676034 175672
rect 676090 175616 676292 175672
rect 676029 175614 676292 175616
rect 676029 175611 676095 175614
rect 667933 175402 667999 175405
rect 666356 175400 667999 175402
rect 666356 175344 667938 175400
rect 667994 175344 667999 175400
rect 666356 175342 667999 175344
rect 667933 175339 667999 175342
rect 676029 175266 676095 175269
rect 676029 175264 676292 175266
rect 676029 175208 676034 175264
rect 676090 175208 676292 175264
rect 676029 175206 676292 175208
rect 676029 175203 676095 175206
rect 603073 174858 603139 174861
rect 676029 174858 676095 174861
rect 603073 174856 606556 174858
rect 603073 174800 603078 174856
rect 603134 174800 606556 174856
rect 603073 174798 606556 174800
rect 676029 174856 676292 174858
rect 676029 174800 676034 174856
rect 676090 174800 676292 174856
rect 676029 174798 676292 174800
rect 603073 174795 603139 174798
rect 676029 174795 676095 174798
rect 674741 174450 674807 174453
rect 674741 174448 676292 174450
rect 674741 174392 674746 174448
rect 674802 174392 676292 174448
rect 674741 174390 676292 174392
rect 674741 174387 674807 174390
rect 578417 174178 578483 174181
rect 576380 174176 578483 174178
rect 576380 174120 578422 174176
rect 578478 174120 578483 174176
rect 576380 174118 578483 174120
rect 578417 174115 578483 174118
rect 675334 173980 675340 174044
rect 675404 174042 675410 174044
rect 675404 173982 676292 174042
rect 675404 173980 675410 173982
rect 603717 173906 603783 173909
rect 603717 173904 606556 173906
rect 603717 173848 603722 173904
rect 603778 173848 606556 173904
rect 603717 173846 606556 173848
rect 603717 173843 603783 173846
rect 667933 173634 667999 173637
rect 668301 173634 668367 173637
rect 666356 173632 668367 173634
rect 666356 173576 667938 173632
rect 667994 173576 668306 173632
rect 668362 173576 668367 173632
rect 666356 173574 668367 173576
rect 667933 173571 667999 173574
rect 668301 173571 668367 173574
rect 676078 173574 676292 173634
rect 676078 173500 676138 173574
rect 676070 173436 676076 173500
rect 676140 173436 676146 173500
rect 678237 173226 678303 173229
rect 678237 173224 678316 173226
rect 678237 173168 678242 173224
rect 678298 173168 678316 173224
rect 678237 173166 678316 173168
rect 678237 173163 678303 173166
rect 603073 172818 603139 172821
rect 676029 172818 676095 172821
rect 603073 172816 606556 172818
rect 603073 172760 603078 172816
rect 603134 172760 606556 172816
rect 603073 172758 606556 172760
rect 676029 172816 676292 172818
rect 676029 172760 676034 172816
rect 676090 172760 676292 172816
rect 676029 172758 676292 172760
rect 603073 172755 603139 172758
rect 676029 172755 676095 172758
rect 578785 172682 578851 172685
rect 576380 172680 578851 172682
rect 576380 172624 578790 172680
rect 578846 172624 578851 172680
rect 576380 172622 578851 172624
rect 578785 172619 578851 172622
rect 676029 172410 676095 172413
rect 676029 172408 676292 172410
rect 676029 172352 676034 172408
rect 676090 172352 676292 172408
rect 676029 172350 676292 172352
rect 676029 172347 676095 172350
rect 676078 171942 676292 172002
rect 603073 171866 603139 171869
rect 676078 171868 676138 171942
rect 603073 171864 606556 171866
rect 603073 171808 603078 171864
rect 603134 171808 606556 171864
rect 603073 171806 606556 171808
rect 603073 171803 603139 171806
rect 676070 171804 676076 171868
rect 676140 171804 676146 171868
rect 676765 171594 676831 171597
rect 676765 171592 676844 171594
rect 676765 171536 676770 171592
rect 676826 171536 676844 171592
rect 676765 171534 676844 171536
rect 676765 171531 676831 171534
rect 578693 171186 578759 171189
rect 667933 171186 667999 171189
rect 576380 171184 578759 171186
rect 576380 171128 578698 171184
rect 578754 171128 578759 171184
rect 576380 171126 578759 171128
rect 578693 171123 578759 171126
rect 666510 171184 667999 171186
rect 666510 171128 667938 171184
rect 667994 171128 667999 171184
rect 666510 171126 667999 171128
rect 603165 170778 603231 170781
rect 603165 170776 606556 170778
rect 603165 170720 603170 170776
rect 603226 170720 606556 170776
rect 603165 170718 606556 170720
rect 603165 170715 603231 170718
rect 666510 170506 666570 171126
rect 667933 171123 667999 171126
rect 676029 171186 676095 171189
rect 676029 171184 676292 171186
rect 676029 171128 676034 171184
rect 676090 171128 676292 171184
rect 676029 171126 676292 171128
rect 676029 171123 676095 171126
rect 675886 170716 675892 170780
rect 675956 170778 675962 170780
rect 675956 170718 676292 170778
rect 675956 170716 675962 170718
rect 666510 170446 666754 170506
rect 666694 170234 666754 170446
rect 676029 170370 676095 170373
rect 676029 170368 676292 170370
rect 676029 170312 676034 170368
rect 676090 170312 676292 170368
rect 676029 170310 676292 170312
rect 676029 170307 676095 170310
rect 666356 170174 666754 170234
rect 676581 169962 676647 169965
rect 676581 169960 676660 169962
rect 676581 169904 676586 169960
rect 676642 169904 676660 169960
rect 676581 169902 676660 169904
rect 676581 169899 676647 169902
rect 603073 169826 603139 169829
rect 603073 169824 606556 169826
rect 603073 169768 603078 169824
rect 603134 169768 606556 169824
rect 603073 169766 606556 169768
rect 603073 169763 603139 169766
rect 675702 169628 675708 169692
rect 675772 169690 675778 169692
rect 676029 169690 676095 169693
rect 675772 169688 676095 169690
rect 675772 169632 676034 169688
rect 676090 169632 676095 169688
rect 675772 169630 676095 169632
rect 675772 169628 675778 169630
rect 676029 169627 676095 169630
rect 579429 169554 579495 169557
rect 576380 169552 579495 169554
rect 576380 169496 579434 169552
rect 579490 169496 579495 169552
rect 576380 169494 579495 169496
rect 579429 169491 579495 169494
rect 676029 169554 676095 169557
rect 676029 169552 676292 169554
rect 676029 169496 676034 169552
rect 676090 169496 676292 169552
rect 676029 169494 676292 169496
rect 676029 169491 676095 169494
rect 676029 169146 676095 169149
rect 676029 169144 676292 169146
rect 676029 169088 676034 169144
rect 676090 169088 676292 169144
rect 676029 169086 676292 169088
rect 676029 169083 676095 169086
rect 603073 168738 603139 168741
rect 676029 168738 676095 168741
rect 603073 168736 606556 168738
rect 603073 168680 603078 168736
rect 603134 168680 606556 168736
rect 603073 168678 606556 168680
rect 676029 168736 676292 168738
rect 676029 168680 676034 168736
rect 676090 168680 676292 168736
rect 676029 168678 676292 168680
rect 603073 168675 603139 168678
rect 676029 168675 676095 168678
rect 668301 168602 668367 168605
rect 666356 168600 668367 168602
rect 666356 168544 668306 168600
rect 668362 168544 668367 168600
rect 666356 168542 668367 168544
rect 668301 168539 668367 168542
rect 676029 168330 676095 168333
rect 676029 168328 676292 168330
rect 676029 168272 676034 168328
rect 676090 168272 676292 168328
rect 676029 168270 676292 168272
rect 676029 168267 676095 168270
rect 579337 168058 579403 168061
rect 576380 168056 579403 168058
rect 576380 168000 579342 168056
rect 579398 168000 579403 168056
rect 576380 167998 579403 168000
rect 579337 167995 579403 167998
rect 676029 167922 676095 167925
rect 676029 167920 676292 167922
rect 676029 167864 676034 167920
rect 676090 167864 676292 167920
rect 676029 167862 676292 167864
rect 676029 167859 676095 167862
rect 603073 167786 603139 167789
rect 603073 167784 606556 167786
rect 603073 167728 603078 167784
rect 603134 167728 606556 167784
rect 603073 167726 606556 167728
rect 603073 167723 603139 167726
rect 676029 167106 676095 167109
rect 676029 167104 676292 167106
rect 676029 167048 676034 167104
rect 676090 167048 676292 167104
rect 676029 167046 676292 167048
rect 676029 167043 676095 167046
rect 603809 166698 603875 166701
rect 603809 166696 606556 166698
rect 603809 166640 603814 166696
rect 603870 166640 606556 166696
rect 603809 166638 606556 166640
rect 603809 166635 603875 166638
rect 578601 166562 578667 166565
rect 576380 166560 578667 166562
rect 576380 166504 578606 166560
rect 578662 166504 578667 166560
rect 576380 166502 578667 166504
rect 578601 166499 578667 166502
rect 676581 166428 676647 166429
rect 676765 166428 676831 166429
rect 676581 166426 676628 166428
rect 676536 166424 676628 166426
rect 676536 166368 676586 166424
rect 676536 166366 676628 166368
rect 676581 166364 676628 166366
rect 676692 166364 676698 166428
rect 676765 166424 676812 166428
rect 676876 166426 676882 166428
rect 676765 166368 676770 166424
rect 676765 166364 676812 166368
rect 676876 166366 676922 166426
rect 676876 166364 676882 166366
rect 676581 166363 676647 166364
rect 676765 166363 676831 166364
rect 603073 165746 603139 165749
rect 603073 165744 606556 165746
rect 603073 165688 603078 165744
rect 603134 165688 606556 165744
rect 603073 165686 606556 165688
rect 603073 165683 603139 165686
rect 668301 165202 668367 165205
rect 666356 165200 668367 165202
rect 666356 165144 668306 165200
rect 668362 165144 668367 165200
rect 666356 165142 668367 165144
rect 668301 165139 668367 165142
rect 576350 164386 576410 165036
rect 603073 164658 603139 164661
rect 603073 164656 606556 164658
rect 603073 164600 603078 164656
rect 603134 164600 606556 164656
rect 603073 164598 606556 164600
rect 603073 164595 603139 164598
rect 578233 164386 578299 164389
rect 576350 164384 578299 164386
rect 576350 164328 578238 164384
rect 578294 164328 578299 164384
rect 576350 164326 578299 164328
rect 578233 164323 578299 164326
rect 603073 163706 603139 163709
rect 603073 163704 606556 163706
rect 603073 163648 603078 163704
rect 603134 163648 606556 163704
rect 603073 163646 606556 163648
rect 603073 163643 603139 163646
rect 579521 163570 579587 163573
rect 667933 163570 667999 163573
rect 576380 163568 579587 163570
rect 576380 163512 579526 163568
rect 579582 163512 579587 163568
rect 576380 163510 579587 163512
rect 666356 163568 667999 163570
rect 666356 163512 667938 163568
rect 667994 163512 667999 163568
rect 666356 163510 667999 163512
rect 579521 163507 579587 163510
rect 667933 163507 667999 163510
rect 676070 162692 676076 162756
rect 676140 162754 676146 162756
rect 677041 162754 677107 162757
rect 676140 162752 677107 162754
rect 676140 162696 677046 162752
rect 677102 162696 677107 162752
rect 676140 162694 677107 162696
rect 676140 162692 676146 162694
rect 677041 162691 677107 162694
rect 603073 162618 603139 162621
rect 603073 162616 606556 162618
rect 603073 162560 603078 162616
rect 603134 162560 606556 162616
rect 603073 162558 606556 162560
rect 603073 162555 603139 162558
rect 675518 162556 675524 162620
rect 675588 162618 675594 162620
rect 676857 162618 676923 162621
rect 675588 162616 676923 162618
rect 675588 162560 676862 162616
rect 676918 162560 676923 162616
rect 675588 162558 676923 162560
rect 675588 162556 675594 162558
rect 676857 162555 676923 162558
rect 579153 162074 579219 162077
rect 576380 162072 579219 162074
rect 576380 162016 579158 162072
rect 579214 162016 579219 162072
rect 576380 162014 579219 162016
rect 579153 162011 579219 162014
rect 603717 161666 603783 161669
rect 603717 161664 606556 161666
rect 603717 161608 603722 161664
rect 603778 161608 606556 161664
rect 603717 161606 606556 161608
rect 603717 161603 603783 161606
rect 667933 161530 667999 161533
rect 666510 161528 667999 161530
rect 666510 161472 667938 161528
rect 667994 161472 667999 161528
rect 666510 161470 667999 161472
rect 579245 160578 579311 160581
rect 576380 160576 579311 160578
rect 576380 160520 579250 160576
rect 579306 160520 579311 160576
rect 576380 160518 579311 160520
rect 579245 160515 579311 160518
rect 603073 160578 603139 160581
rect 603073 160576 606556 160578
rect 603073 160520 603078 160576
rect 603134 160520 606556 160576
rect 603073 160518 606556 160520
rect 603073 160515 603139 160518
rect 666510 160442 666570 161470
rect 667933 161467 667999 161470
rect 666510 160382 666754 160442
rect 666694 160170 666754 160382
rect 666356 160110 666754 160170
rect 675753 160034 675819 160037
rect 676806 160034 676812 160036
rect 675753 160032 676812 160034
rect 675753 159976 675758 160032
rect 675814 159976 676812 160032
rect 675753 159974 676812 159976
rect 675753 159971 675819 159974
rect 676806 159972 676812 159974
rect 676876 159972 676882 160036
rect 603073 159626 603139 159629
rect 603073 159624 606556 159626
rect 603073 159568 603078 159624
rect 603134 159568 606556 159624
rect 603073 159566 606556 159568
rect 603073 159563 603139 159566
rect 675334 159428 675340 159492
rect 675404 159490 675410 159492
rect 675477 159490 675543 159493
rect 675404 159488 675543 159490
rect 675404 159432 675482 159488
rect 675538 159432 675543 159488
rect 675404 159430 675543 159432
rect 675404 159428 675410 159430
rect 675477 159427 675543 159430
rect 579061 159082 579127 159085
rect 576380 159080 579127 159082
rect 576380 159024 579066 159080
rect 579122 159024 579127 159080
rect 576380 159022 579127 159024
rect 579061 159019 579127 159022
rect 603165 158538 603231 158541
rect 603165 158536 606556 158538
rect 603165 158480 603170 158536
rect 603226 158480 606556 158536
rect 603165 158478 606556 158480
rect 603165 158475 603231 158478
rect 667933 158402 667999 158405
rect 668669 158402 668735 158405
rect 666356 158400 668735 158402
rect 666356 158344 667938 158400
rect 667994 158344 668674 158400
rect 668730 158344 668735 158400
rect 666356 158342 668735 158344
rect 667933 158339 667999 158342
rect 668669 158339 668735 158342
rect 578877 157586 578943 157589
rect 576380 157584 578943 157586
rect 576380 157528 578882 157584
rect 578938 157528 578943 157584
rect 576380 157526 578943 157528
rect 578877 157523 578943 157526
rect 603073 157586 603139 157589
rect 603073 157584 606556 157586
rect 603073 157528 603078 157584
rect 603134 157528 606556 157584
rect 603073 157526 606556 157528
rect 603073 157523 603139 157526
rect 675661 157452 675727 157453
rect 675661 157448 675708 157452
rect 675772 157450 675778 157452
rect 675661 157392 675666 157448
rect 675661 157388 675708 157392
rect 675772 157390 675818 157450
rect 675772 157388 675778 157390
rect 675661 157387 675727 157388
rect 675477 157044 675543 157045
rect 675477 157040 675524 157044
rect 675588 157042 675594 157044
rect 675477 156984 675482 157040
rect 675477 156980 675524 156984
rect 675588 156982 675634 157042
rect 675588 156980 675594 156982
rect 675477 156979 675543 156980
rect 603073 156498 603139 156501
rect 603073 156496 606556 156498
rect 603073 156440 603078 156496
rect 603134 156440 606556 156496
rect 603073 156438 606556 156440
rect 603073 156435 603139 156438
rect 675753 156362 675819 156365
rect 675886 156362 675892 156364
rect 675753 156360 675892 156362
rect 675753 156304 675758 156360
rect 675814 156304 675892 156360
rect 675753 156302 675892 156304
rect 675753 156299 675819 156302
rect 675886 156300 675892 156302
rect 675956 156300 675962 156364
rect 578969 156090 579035 156093
rect 576380 156088 579035 156090
rect 576380 156032 578974 156088
rect 579030 156032 579035 156088
rect 576380 156030 579035 156032
rect 578969 156027 579035 156030
rect 603073 155546 603139 155549
rect 603073 155544 606556 155546
rect 603073 155488 603078 155544
rect 603134 155488 606556 155544
rect 603073 155486 606556 155488
rect 603073 155483 603139 155486
rect 667933 155002 667999 155005
rect 666356 155000 667999 155002
rect 666356 154944 667938 155000
rect 667994 154944 667999 155000
rect 666356 154942 667999 154944
rect 667933 154939 667999 154942
rect 578325 154594 578391 154597
rect 576380 154592 578391 154594
rect 576380 154536 578330 154592
rect 578386 154536 578391 154592
rect 576380 154534 578391 154536
rect 578325 154531 578391 154534
rect 603165 154458 603231 154461
rect 603165 154456 606556 154458
rect 603165 154400 603170 154456
rect 603226 154400 606556 154456
rect 603165 154398 606556 154400
rect 603165 154395 603231 154398
rect 603073 153506 603139 153509
rect 603073 153504 606556 153506
rect 603073 153448 603078 153504
rect 603134 153448 606556 153504
rect 603073 153446 606556 153448
rect 603073 153443 603139 153446
rect 666553 153370 666619 153373
rect 668577 153370 668643 153373
rect 666356 153368 668643 153370
rect 666356 153312 666558 153368
rect 666614 153312 668582 153368
rect 668638 153312 668643 153368
rect 666356 153310 668643 153312
rect 666553 153307 666619 153310
rect 668577 153307 668643 153310
rect 579521 153098 579587 153101
rect 576380 153096 579587 153098
rect 576380 153040 579526 153096
rect 579582 153040 579587 153096
rect 576380 153038 579587 153040
rect 579521 153035 579587 153038
rect 675753 153098 675819 153101
rect 676070 153098 676076 153100
rect 675753 153096 676076 153098
rect 675753 153040 675758 153096
rect 675814 153040 676076 153096
rect 675753 153038 676076 153040
rect 675753 153035 675819 153038
rect 676070 153036 676076 153038
rect 676140 153036 676146 153100
rect 603073 152418 603139 152421
rect 603073 152416 606556 152418
rect 603073 152360 603078 152416
rect 603134 152360 606556 152416
rect 603073 152358 606556 152360
rect 603073 152355 603139 152358
rect 666553 151874 666619 151877
rect 666510 151872 666619 151874
rect 666510 151816 666558 151872
rect 666614 151816 666619 151872
rect 666510 151811 666619 151816
rect 666510 151770 666616 151811
rect 666556 151605 666616 151770
rect 579429 151602 579495 151605
rect 576380 151600 579495 151602
rect 576380 151544 579434 151600
rect 579490 151544 579495 151600
rect 576380 151542 579495 151544
rect 579429 151539 579495 151542
rect 666553 151600 666619 151605
rect 666553 151544 666558 151600
rect 666614 151544 666619 151600
rect 666553 151539 666619 151544
rect 675753 151602 675819 151605
rect 676622 151602 676628 151604
rect 675753 151600 676628 151602
rect 675753 151544 675758 151600
rect 675814 151544 676628 151600
rect 675753 151542 676628 151544
rect 675753 151539 675819 151542
rect 676622 151540 676628 151542
rect 676692 151540 676698 151604
rect 603073 151466 603139 151469
rect 603073 151464 606556 151466
rect 603073 151408 603078 151464
rect 603134 151408 606556 151464
rect 603073 151406 606556 151408
rect 603073 151403 603139 151406
rect 603073 150378 603139 150381
rect 603073 150376 606556 150378
rect 603073 150320 603078 150376
rect 603134 150320 606556 150376
rect 603073 150318 606556 150320
rect 603073 150315 603139 150318
rect 579429 150106 579495 150109
rect 576380 150104 579495 150106
rect 576380 150048 579434 150104
rect 579490 150048 579495 150104
rect 576380 150046 579495 150048
rect 579429 150043 579495 150046
rect 666553 149970 666619 149973
rect 666356 149968 666619 149970
rect 666356 149912 666558 149968
rect 666614 149912 666619 149968
rect 666356 149910 666619 149912
rect 666553 149907 666619 149910
rect 603901 149426 603967 149429
rect 603901 149424 606556 149426
rect 603901 149368 603906 149424
rect 603962 149368 606556 149424
rect 603901 149366 606556 149368
rect 603901 149363 603967 149366
rect 578509 148610 578575 148613
rect 576380 148608 578575 148610
rect 576380 148552 578514 148608
rect 578570 148552 578575 148608
rect 576380 148550 578575 148552
rect 578509 148547 578575 148550
rect 675753 148474 675819 148477
rect 676438 148474 676444 148476
rect 675753 148472 676444 148474
rect 675753 148416 675758 148472
rect 675814 148416 676444 148472
rect 675753 148414 676444 148416
rect 675753 148411 675819 148414
rect 676438 148412 676444 148414
rect 676508 148412 676514 148476
rect 603073 148338 603139 148341
rect 603073 148336 606556 148338
rect 603073 148280 603078 148336
rect 603134 148280 606556 148336
rect 603073 148278 606556 148280
rect 603073 148275 603139 148278
rect 668301 148202 668367 148205
rect 666356 148200 668367 148202
rect 666356 148144 668306 148200
rect 668362 148144 668367 148200
rect 666356 148142 668367 148144
rect 668301 148139 668367 148142
rect 603073 147386 603139 147389
rect 603073 147384 606556 147386
rect 603073 147328 603078 147384
rect 603134 147328 606556 147384
rect 603073 147326 606556 147328
rect 603073 147323 603139 147326
rect 579521 146978 579587 146981
rect 576380 146976 579587 146978
rect 576380 146920 579526 146976
rect 579582 146920 579587 146976
rect 576380 146918 579587 146920
rect 579521 146915 579587 146918
rect 603165 146298 603231 146301
rect 675753 146298 675819 146301
rect 676254 146298 676260 146300
rect 603165 146296 606556 146298
rect 603165 146240 603170 146296
rect 603226 146240 606556 146296
rect 603165 146238 606556 146240
rect 675753 146296 676260 146298
rect 675753 146240 675758 146296
rect 675814 146240 676260 146296
rect 675753 146238 676260 146240
rect 603165 146235 603231 146238
rect 675753 146235 675819 146238
rect 676254 146236 676260 146238
rect 676324 146236 676330 146300
rect 578693 145482 578759 145485
rect 576380 145480 578759 145482
rect 576380 145424 578698 145480
rect 578754 145424 578759 145480
rect 576380 145422 578759 145424
rect 578693 145419 578759 145422
rect 603717 145346 603783 145349
rect 603717 145344 606556 145346
rect 603717 145288 603722 145344
rect 603778 145288 606556 145344
rect 603717 145286 606556 145288
rect 603717 145283 603783 145286
rect 668301 144938 668367 144941
rect 666356 144936 668367 144938
rect 666356 144880 668306 144936
rect 668362 144880 668367 144936
rect 666356 144878 668367 144880
rect 668301 144875 668367 144878
rect 603073 144258 603139 144261
rect 603073 144256 606556 144258
rect 603073 144200 603078 144256
rect 603134 144200 606556 144256
rect 603073 144198 606556 144200
rect 603073 144195 603139 144198
rect 579521 143986 579587 143989
rect 576380 143984 579587 143986
rect 576380 143928 579526 143984
rect 579582 143928 579587 143984
rect 576380 143926 579587 143928
rect 579521 143923 579587 143926
rect 603809 143306 603875 143309
rect 603809 143304 606556 143306
rect 603809 143248 603814 143304
rect 603870 143248 606556 143304
rect 603809 143246 606556 143248
rect 603809 143243 603875 143246
rect 667933 143170 667999 143173
rect 666356 143168 667999 143170
rect 666356 143112 667938 143168
rect 667994 143112 667999 143168
rect 666356 143110 667999 143112
rect 578693 142490 578759 142493
rect 576380 142488 578759 142490
rect 576380 142432 578698 142488
rect 578754 142432 578759 142488
rect 576380 142430 578759 142432
rect 578693 142427 578759 142430
rect 603073 142218 603139 142221
rect 603073 142216 606556 142218
rect 603073 142160 603078 142216
rect 603134 142160 606556 142216
rect 603073 142158 606556 142160
rect 603073 142155 603139 142158
rect 666510 142085 666570 143110
rect 667933 143107 667999 143110
rect 666510 142080 666619 142085
rect 666510 142024 666558 142080
rect 666614 142024 666619 142080
rect 666510 142022 666619 142024
rect 666553 142019 666619 142022
rect 603073 141266 603139 141269
rect 603073 141264 606556 141266
rect 603073 141208 603078 141264
rect 603134 141208 606556 141264
rect 603073 141206 606556 141208
rect 603073 141203 603139 141206
rect 579337 140994 579403 140997
rect 576380 140992 579403 140994
rect 576380 140936 579342 140992
rect 579398 140936 579403 140992
rect 576380 140934 579403 140936
rect 579337 140931 579403 140934
rect 603073 140178 603139 140181
rect 603073 140176 606556 140178
rect 603073 140120 603078 140176
rect 603134 140120 606556 140176
rect 603073 140118 606556 140120
rect 603073 140115 603139 140118
rect 666553 139770 666619 139773
rect 666356 139768 666619 139770
rect 666356 139712 666558 139768
rect 666614 139712 666619 139768
rect 666356 139710 666619 139712
rect 666553 139707 666619 139710
rect 579153 139498 579219 139501
rect 576380 139496 579219 139498
rect 576380 139440 579158 139496
rect 579214 139440 579219 139496
rect 576380 139438 579219 139440
rect 579153 139435 579219 139438
rect 603165 139226 603231 139229
rect 603165 139224 606556 139226
rect 603165 139168 603170 139224
rect 603226 139168 606556 139224
rect 603165 139166 606556 139168
rect 603165 139163 603231 139166
rect 603073 138138 603139 138141
rect 667933 138138 667999 138141
rect 603073 138136 606556 138138
rect 603073 138080 603078 138136
rect 603134 138080 606556 138136
rect 603073 138078 606556 138080
rect 666356 138136 667999 138138
rect 666356 138080 667938 138136
rect 667994 138080 667999 138136
rect 666356 138078 667999 138080
rect 603073 138075 603139 138078
rect 667933 138075 667999 138078
rect 579521 138002 579587 138005
rect 576380 138000 579587 138002
rect 576380 137944 579526 138000
rect 579582 137944 579587 138000
rect 576380 137942 579587 137944
rect 579521 137939 579587 137942
rect 603073 137186 603139 137189
rect 603073 137184 606556 137186
rect 603073 137128 603078 137184
rect 603134 137128 606556 137184
rect 603073 137126 606556 137128
rect 603073 137123 603139 137126
rect 579521 136506 579587 136509
rect 576380 136504 579587 136506
rect 576380 136448 579526 136504
rect 579582 136448 579587 136504
rect 576380 136446 579587 136448
rect 579521 136443 579587 136446
rect 603073 136098 603139 136101
rect 603073 136096 606556 136098
rect 603073 136040 603078 136096
rect 603134 136040 606556 136096
rect 603073 136038 606556 136040
rect 603073 136035 603139 136038
rect 603165 135146 603231 135149
rect 603165 135144 606556 135146
rect 603165 135088 603170 135144
rect 603226 135088 606556 135144
rect 603165 135086 606556 135088
rect 603165 135083 603231 135086
rect 579245 135010 579311 135013
rect 576380 135008 579311 135010
rect 576380 134952 579250 135008
rect 579306 134952 579311 135008
rect 576380 134950 579311 134952
rect 579245 134947 579311 134950
rect 667933 134738 667999 134741
rect 666356 134736 667999 134738
rect 666356 134680 667938 134736
rect 667994 134680 667999 134736
rect 666356 134678 667999 134680
rect 667933 134675 667999 134678
rect 603073 134058 603139 134061
rect 603073 134056 606556 134058
rect 603073 134000 603078 134056
rect 603134 134000 606556 134056
rect 603073 133998 606556 134000
rect 603073 133995 603139 133998
rect 579061 133514 579127 133517
rect 576380 133512 579127 133514
rect 576380 133456 579066 133512
rect 579122 133456 579127 133512
rect 576380 133454 579127 133456
rect 579061 133451 579127 133454
rect 603073 133106 603139 133109
rect 676121 133106 676187 133109
rect 676262 133106 676322 133348
rect 603073 133104 606556 133106
rect 603073 133048 603078 133104
rect 603134 133048 606556 133104
rect 603073 133046 606556 133048
rect 676121 133104 676322 133106
rect 676121 133048 676126 133104
rect 676182 133048 676322 133104
rect 676121 133046 676322 133048
rect 603073 133043 603139 133046
rect 676121 133043 676187 133046
rect 668577 132970 668643 132973
rect 666356 132968 668643 132970
rect 666356 132912 668582 132968
rect 668638 132912 668643 132968
rect 666356 132910 668643 132912
rect 666510 132429 666570 132910
rect 668577 132907 668643 132910
rect 676029 132970 676095 132973
rect 676029 132968 676292 132970
rect 676029 132912 676034 132968
rect 676090 132912 676292 132968
rect 676029 132910 676292 132912
rect 676029 132907 676095 132910
rect 676213 132698 676279 132701
rect 676213 132696 676322 132698
rect 676213 132640 676218 132696
rect 676274 132640 676322 132696
rect 676213 132635 676322 132640
rect 676262 132532 676322 132635
rect 666510 132424 666619 132429
rect 666510 132368 666558 132424
rect 666614 132368 666619 132424
rect 666510 132366 666619 132368
rect 666553 132363 666619 132366
rect 578877 132018 578943 132021
rect 576380 132016 578943 132018
rect 576380 131960 578882 132016
rect 578938 131960 578943 132016
rect 576380 131958 578943 131960
rect 578877 131955 578943 131958
rect 603073 132018 603139 132021
rect 603073 132016 606556 132018
rect 603073 131960 603078 132016
rect 603134 131960 606556 132016
rect 603073 131958 606556 131960
rect 603073 131955 603139 131958
rect 676262 131885 676322 132124
rect 676213 131880 676322 131885
rect 676213 131824 676218 131880
rect 676274 131824 676322 131880
rect 676213 131822 676322 131824
rect 676213 131819 676279 131822
rect 676121 131474 676187 131477
rect 676262 131474 676322 131716
rect 676121 131472 676322 131474
rect 676121 131416 676126 131472
rect 676182 131416 676322 131472
rect 676121 131414 676322 131416
rect 676121 131411 676187 131414
rect 676029 131338 676095 131341
rect 676029 131336 676292 131338
rect 676029 131280 676034 131336
rect 676090 131280 676292 131336
rect 676029 131278 676292 131280
rect 676029 131275 676095 131278
rect 603165 131066 603231 131069
rect 603165 131064 606556 131066
rect 603165 131008 603170 131064
rect 603226 131008 606556 131064
rect 603165 131006 606556 131008
rect 603165 131003 603231 131006
rect 676121 130658 676187 130661
rect 676262 130658 676322 130900
rect 676121 130656 676322 130658
rect 676121 130600 676126 130656
rect 676182 130600 676322 130656
rect 676121 130598 676322 130600
rect 676121 130595 676187 130598
rect 578325 130522 578391 130525
rect 576380 130520 578391 130522
rect 576380 130464 578330 130520
rect 578386 130464 578391 130520
rect 576380 130462 578391 130464
rect 578325 130459 578391 130462
rect 676262 130253 676322 130492
rect 676213 130248 676322 130253
rect 676213 130192 676218 130248
rect 676274 130192 676322 130248
rect 676213 130190 676322 130192
rect 676213 130187 676279 130190
rect 603073 129978 603139 129981
rect 603073 129976 606556 129978
rect 603073 129920 603078 129976
rect 603134 129920 606556 129976
rect 603073 129918 606556 129920
rect 603073 129915 603139 129918
rect 676262 129845 676322 130084
rect 676213 129840 676322 129845
rect 676213 129784 676218 129840
rect 676274 129784 676322 129840
rect 676213 129782 676322 129784
rect 676213 129779 676279 129782
rect 674741 129706 674807 129709
rect 674741 129704 676292 129706
rect 674741 129648 674746 129704
rect 674802 129648 676292 129704
rect 674741 129646 676292 129648
rect 674741 129643 674807 129646
rect 666553 129570 666619 129573
rect 666356 129568 666619 129570
rect 666356 129512 666558 129568
rect 666614 129512 666619 129568
rect 666356 129510 666619 129512
rect 666553 129507 666619 129510
rect 676262 129029 676322 129268
rect 578969 129026 579035 129029
rect 576380 129024 579035 129026
rect 576380 128968 578974 129024
rect 579030 128968 579035 129024
rect 576380 128966 579035 128968
rect 578969 128963 579035 128966
rect 603073 129026 603139 129029
rect 603073 129024 606556 129026
rect 603073 128968 603078 129024
rect 603134 128968 606556 129024
rect 603073 128966 606556 128968
rect 676213 129024 676322 129029
rect 676213 128968 676218 129024
rect 676274 128968 676322 129024
rect 676213 128966 676322 128968
rect 603073 128963 603139 128966
rect 676213 128963 676279 128966
rect 675334 128828 675340 128892
rect 675404 128890 675410 128892
rect 675404 128830 676292 128890
rect 675404 128828 675410 128830
rect 683622 128213 683682 128452
rect 683622 128208 683731 128213
rect 683622 128152 683670 128208
rect 683726 128152 683731 128208
rect 683622 128150 683731 128152
rect 683665 128147 683731 128150
rect 676029 128074 676095 128077
rect 676029 128072 676292 128074
rect 676029 128016 676034 128072
rect 676090 128016 676292 128072
rect 676029 128014 676292 128016
rect 676029 128011 676095 128014
rect 603073 127938 603139 127941
rect 667933 127938 667999 127941
rect 603073 127936 606556 127938
rect 603073 127880 603078 127936
rect 603134 127880 606556 127936
rect 603073 127878 606556 127880
rect 666356 127936 667999 127938
rect 666356 127880 667938 127936
rect 667994 127880 667999 127936
rect 666356 127878 667999 127880
rect 603073 127875 603139 127878
rect 667933 127875 667999 127878
rect 579521 127530 579587 127533
rect 576380 127528 579587 127530
rect 576380 127472 579526 127528
rect 579582 127472 579587 127528
rect 576380 127470 579587 127472
rect 579521 127467 579587 127470
rect 683070 127397 683130 127636
rect 683070 127392 683179 127397
rect 683070 127336 683118 127392
rect 683174 127336 683179 127392
rect 683070 127334 683179 127336
rect 683113 127331 683179 127334
rect 676814 126989 676874 127228
rect 603165 126986 603231 126989
rect 603165 126984 606556 126986
rect 603165 126928 603170 126984
rect 603226 126928 606556 126984
rect 603165 126926 606556 126928
rect 676814 126984 676923 126989
rect 676814 126928 676862 126984
rect 676918 126928 676923 126984
rect 676814 126926 676923 126928
rect 603165 126923 603231 126926
rect 676857 126923 676923 126926
rect 676262 126580 676322 126820
rect 676254 126516 676260 126580
rect 676324 126516 676330 126580
rect 683254 126173 683314 126412
rect 683254 126168 683363 126173
rect 683254 126112 683302 126168
rect 683358 126112 683363 126168
rect 683254 126110 683363 126112
rect 683297 126107 683363 126110
rect 578693 126034 578759 126037
rect 576380 126032 578759 126034
rect 576380 125976 578698 126032
rect 578754 125976 578759 126032
rect 576380 125974 578759 125976
rect 578693 125971 578759 125974
rect 603073 125898 603139 125901
rect 603073 125896 606556 125898
rect 603073 125840 603078 125896
rect 603134 125840 606556 125896
rect 603073 125838 606556 125840
rect 603073 125835 603139 125838
rect 679574 125765 679634 126004
rect 679574 125760 679683 125765
rect 679574 125704 679622 125760
rect 679678 125704 679683 125760
rect 679574 125702 679683 125704
rect 679617 125699 679683 125702
rect 678286 125357 678346 125596
rect 676397 125354 676463 125357
rect 676397 125352 676506 125354
rect 676397 125296 676402 125352
rect 676458 125296 676506 125352
rect 676397 125291 676506 125296
rect 678237 125352 678346 125357
rect 678237 125296 678242 125352
rect 678298 125296 678346 125352
rect 678237 125294 678346 125296
rect 678237 125291 678303 125294
rect 676446 125188 676506 125291
rect 603073 124946 603139 124949
rect 603073 124944 606556 124946
rect 603073 124888 603078 124944
rect 603134 124888 606556 124944
rect 603073 124886 606556 124888
rect 603073 124883 603139 124886
rect 675702 124884 675708 124948
rect 675772 124946 675778 124948
rect 683113 124946 683179 124949
rect 675772 124944 683179 124946
rect 675772 124888 683118 124944
rect 683174 124888 683179 124944
rect 675772 124886 683179 124888
rect 675772 124884 675778 124886
rect 683113 124883 683179 124886
rect 578417 124538 578483 124541
rect 667933 124538 667999 124541
rect 676446 124540 676506 124780
rect 576380 124536 578483 124538
rect 576380 124480 578422 124536
rect 578478 124480 578483 124536
rect 576380 124478 578483 124480
rect 666356 124536 667999 124538
rect 666356 124480 667938 124536
rect 667994 124480 667999 124536
rect 666356 124478 667999 124480
rect 578417 124475 578483 124478
rect 667933 124475 667999 124478
rect 676438 124476 676444 124540
rect 676508 124476 676514 124540
rect 677550 124133 677610 124372
rect 677550 124128 677659 124133
rect 677550 124072 677598 124128
rect 677654 124072 677659 124128
rect 677550 124070 677659 124072
rect 677593 124067 677659 124070
rect 676029 123994 676095 123997
rect 676029 123992 676292 123994
rect 676029 123936 676034 123992
rect 676090 123936 676292 123992
rect 676029 123934 676292 123936
rect 676029 123931 676095 123934
rect 603073 123858 603139 123861
rect 603073 123856 606556 123858
rect 603073 123800 603078 123856
rect 603134 123800 606556 123856
rect 603073 123798 606556 123800
rect 603073 123795 603139 123798
rect 674741 123586 674807 123589
rect 674741 123584 676292 123586
rect 674741 123528 674746 123584
rect 674802 123528 676292 123584
rect 674741 123526 676292 123528
rect 674741 123523 674807 123526
rect 676262 122909 676322 123148
rect 579245 122906 579311 122909
rect 576380 122904 579311 122906
rect 576380 122848 579250 122904
rect 579306 122848 579311 122904
rect 576380 122846 579311 122848
rect 579245 122843 579311 122846
rect 603165 122906 603231 122909
rect 667933 122906 667999 122909
rect 603165 122904 606556 122906
rect 603165 122848 603170 122904
rect 603226 122848 606556 122904
rect 603165 122846 606556 122848
rect 666356 122904 667999 122906
rect 666356 122848 667938 122904
rect 667994 122848 667999 122904
rect 666356 122846 667999 122848
rect 603165 122843 603231 122846
rect 666510 122773 666570 122846
rect 667933 122843 667999 122846
rect 676213 122904 676322 122909
rect 676213 122848 676218 122904
rect 676274 122848 676322 122904
rect 676213 122846 676322 122848
rect 676213 122843 676279 122846
rect 666510 122768 666619 122773
rect 666510 122712 666558 122768
rect 666614 122712 666619 122768
rect 666510 122710 666619 122712
rect 666553 122707 666619 122710
rect 676121 122498 676187 122501
rect 676262 122498 676322 122740
rect 676121 122496 676322 122498
rect 676121 122440 676126 122496
rect 676182 122440 676322 122496
rect 676121 122438 676322 122440
rect 676121 122435 676187 122438
rect 603073 121818 603139 121821
rect 603073 121816 606556 121818
rect 603073 121760 603078 121816
rect 603134 121760 606556 121816
rect 603073 121758 606556 121760
rect 603073 121755 603139 121758
rect 676262 121685 676322 121924
rect 676213 121680 676322 121685
rect 676213 121624 676218 121680
rect 676274 121624 676322 121680
rect 676213 121622 676322 121624
rect 676213 121619 676279 121622
rect 676806 121620 676812 121684
rect 676876 121682 676882 121684
rect 683665 121682 683731 121685
rect 676876 121680 683731 121682
rect 676876 121624 683670 121680
rect 683726 121624 683731 121680
rect 676876 121622 683731 121624
rect 676876 121620 676882 121622
rect 683665 121619 683731 121622
rect 579521 121410 579587 121413
rect 576380 121408 579587 121410
rect 576380 121352 579526 121408
rect 579582 121352 579587 121408
rect 576380 121350 579587 121352
rect 579521 121347 579587 121350
rect 603073 120866 603139 120869
rect 603073 120864 606556 120866
rect 603073 120808 603078 120864
rect 603134 120808 606556 120864
rect 603073 120806 606556 120808
rect 603073 120803 603139 120806
rect 579245 119914 579311 119917
rect 576380 119912 579311 119914
rect 576380 119856 579250 119912
rect 579306 119856 579311 119912
rect 576380 119854 579311 119856
rect 579245 119851 579311 119854
rect 603073 119778 603139 119781
rect 603073 119776 606556 119778
rect 603073 119720 603078 119776
rect 603134 119720 606556 119776
rect 603073 119718 606556 119720
rect 603073 119715 603139 119718
rect 666553 119506 666619 119509
rect 666356 119504 666619 119506
rect 666356 119448 666558 119504
rect 666614 119448 666619 119504
rect 666356 119446 666619 119448
rect 666553 119443 666619 119446
rect 603717 118826 603783 118829
rect 603717 118824 606556 118826
rect 603717 118768 603722 118824
rect 603778 118768 606556 118824
rect 603717 118766 606556 118768
rect 603717 118763 603783 118766
rect 578509 118418 578575 118421
rect 576380 118416 578575 118418
rect 576380 118360 578514 118416
rect 578570 118360 578575 118416
rect 576380 118358 578575 118360
rect 578509 118355 578575 118358
rect 676070 117948 676076 118012
rect 676140 118010 676146 118012
rect 676857 118010 676923 118013
rect 676140 118008 676923 118010
rect 676140 117952 676862 118008
rect 676918 117952 676923 118008
rect 676140 117950 676923 117952
rect 676140 117948 676146 117950
rect 676857 117947 676923 117950
rect 603073 117738 603139 117741
rect 667933 117738 667999 117741
rect 603073 117736 606556 117738
rect 603073 117680 603078 117736
rect 603134 117680 606556 117736
rect 603073 117678 606556 117680
rect 666356 117736 667999 117738
rect 666356 117680 667938 117736
rect 667994 117680 667999 117736
rect 666356 117678 667999 117680
rect 603073 117675 603139 117678
rect 667933 117675 667999 117678
rect 675886 117268 675892 117332
rect 675956 117330 675962 117332
rect 676397 117330 676463 117333
rect 675956 117328 676463 117330
rect 675956 117272 676402 117328
rect 676458 117272 676463 117328
rect 675956 117270 676463 117272
rect 675956 117268 675962 117270
rect 676397 117267 676463 117270
rect 675518 117132 675524 117196
rect 675588 117194 675594 117196
rect 679617 117194 679683 117197
rect 675588 117192 679683 117194
rect 675588 117136 679622 117192
rect 679678 117136 679683 117192
rect 675588 117134 679683 117136
rect 675588 117132 675594 117134
rect 679617 117131 679683 117134
rect 579521 116922 579587 116925
rect 576380 116920 579587 116922
rect 576380 116864 579526 116920
rect 579582 116864 579587 116920
rect 576380 116862 579587 116864
rect 579521 116859 579587 116862
rect 602337 116786 602403 116789
rect 602337 116784 606556 116786
rect 602337 116728 602342 116784
rect 602398 116728 606556 116784
rect 602337 116726 606556 116728
rect 602337 116723 602403 116726
rect 668393 116106 668459 116109
rect 666356 116104 668459 116106
rect 666356 116048 668398 116104
rect 668454 116048 668459 116104
rect 666356 116046 668459 116048
rect 668393 116043 668459 116046
rect 603073 115698 603139 115701
rect 603073 115696 606556 115698
rect 603073 115640 603078 115696
rect 603134 115640 606556 115696
rect 603073 115638 606556 115640
rect 603073 115635 603139 115638
rect 579429 115426 579495 115429
rect 576380 115424 579495 115426
rect 576380 115368 579434 115424
rect 579490 115368 579495 115424
rect 576380 115366 579495 115368
rect 579429 115363 579495 115366
rect 603165 114746 603231 114749
rect 603165 114744 606556 114746
rect 603165 114688 603170 114744
rect 603226 114688 606556 114744
rect 603165 114686 606556 114688
rect 603165 114683 603231 114686
rect 669221 114338 669287 114341
rect 666356 114336 669287 114338
rect 666356 114280 669226 114336
rect 669282 114280 669287 114336
rect 666356 114278 669287 114280
rect 669221 114275 669287 114278
rect 675385 114204 675451 114205
rect 675334 114202 675340 114204
rect 675294 114142 675340 114202
rect 675404 114200 675451 114204
rect 675446 114144 675451 114200
rect 675334 114140 675340 114142
rect 675404 114140 675451 114144
rect 675385 114139 675451 114140
rect 579245 113930 579311 113933
rect 576380 113928 579311 113930
rect 576380 113872 579250 113928
rect 579306 113872 579311 113928
rect 576380 113870 579311 113872
rect 579245 113867 579311 113870
rect 603073 113658 603139 113661
rect 603073 113656 606556 113658
rect 603073 113600 603078 113656
rect 603134 113600 606556 113656
rect 603073 113598 606556 113600
rect 603073 113595 603139 113598
rect 603073 112706 603139 112709
rect 668853 112706 668919 112709
rect 603073 112704 606556 112706
rect 603073 112648 603078 112704
rect 603134 112648 606556 112704
rect 603073 112646 606556 112648
rect 666356 112704 668919 112706
rect 666356 112648 668858 112704
rect 668914 112648 668919 112704
rect 666356 112646 668919 112648
rect 603073 112643 603139 112646
rect 668853 112643 668919 112646
rect 675661 112572 675727 112573
rect 675661 112568 675708 112572
rect 675772 112570 675778 112572
rect 675661 112512 675666 112568
rect 675661 112508 675708 112512
rect 675772 112510 675818 112570
rect 675772 112508 675778 112510
rect 675661 112507 675727 112508
rect 579521 112434 579587 112437
rect 576380 112432 579587 112434
rect 576380 112376 579526 112432
rect 579582 112376 579587 112432
rect 576380 112374 579587 112376
rect 579521 112371 579587 112374
rect 675477 111756 675543 111757
rect 675477 111752 675524 111756
rect 675588 111754 675594 111756
rect 675477 111696 675482 111752
rect 675477 111692 675524 111696
rect 675588 111694 675634 111754
rect 675588 111692 675594 111694
rect 675477 111691 675543 111692
rect 603809 111618 603875 111621
rect 603809 111616 606556 111618
rect 603809 111560 603814 111616
rect 603870 111560 606556 111616
rect 603809 111558 606556 111560
rect 603809 111555 603875 111558
rect 578693 110938 578759 110941
rect 668301 110938 668367 110941
rect 576380 110936 578759 110938
rect 576380 110880 578698 110936
rect 578754 110880 578759 110936
rect 576380 110878 578759 110880
rect 666356 110936 668367 110938
rect 666356 110880 668306 110936
rect 668362 110880 668367 110936
rect 666356 110878 668367 110880
rect 578693 110875 578759 110878
rect 668301 110875 668367 110878
rect 603073 110666 603139 110669
rect 603073 110664 606556 110666
rect 603073 110608 603078 110664
rect 603134 110608 606556 110664
rect 603073 110606 606556 110608
rect 603073 110603 603139 110606
rect 603073 109578 603139 109581
rect 603073 109576 606556 109578
rect 603073 109520 603078 109576
rect 603134 109520 606556 109576
rect 603073 109518 606556 109520
rect 603073 109515 603139 109518
rect 579521 109442 579587 109445
rect 576380 109440 579587 109442
rect 576380 109384 579526 109440
rect 579582 109384 579587 109440
rect 576380 109382 579587 109384
rect 579521 109379 579587 109382
rect 667933 109306 667999 109309
rect 666356 109304 667999 109306
rect 666356 109248 667938 109304
rect 667994 109248 667999 109304
rect 666356 109246 667999 109248
rect 667933 109243 667999 109246
rect 675109 109034 675175 109037
rect 676438 109034 676444 109036
rect 675109 109032 676444 109034
rect 675109 108976 675114 109032
rect 675170 108976 676444 109032
rect 675109 108974 676444 108976
rect 675109 108971 675175 108974
rect 676438 108972 676444 108974
rect 676508 108972 676514 109036
rect 603073 108626 603139 108629
rect 603073 108624 606556 108626
rect 603073 108568 603078 108624
rect 603134 108568 606556 108624
rect 603073 108566 606556 108568
rect 603073 108563 603139 108566
rect 675753 108218 675819 108221
rect 676070 108218 676076 108220
rect 675753 108216 676076 108218
rect 675753 108160 675758 108216
rect 675814 108160 676076 108216
rect 675753 108158 676076 108160
rect 675753 108155 675819 108158
rect 676070 108156 676076 108158
rect 676140 108156 676146 108220
rect 578785 107946 578851 107949
rect 576380 107944 578851 107946
rect 576380 107888 578790 107944
rect 578846 107888 578851 107944
rect 576380 107886 578851 107888
rect 578785 107883 578851 107886
rect 603165 107538 603231 107541
rect 668117 107538 668183 107541
rect 603165 107536 606556 107538
rect 603165 107480 603170 107536
rect 603226 107480 606556 107536
rect 603165 107478 606556 107480
rect 666356 107536 668183 107538
rect 666356 107480 668122 107536
rect 668178 107480 668183 107536
rect 666356 107478 668183 107480
rect 603165 107475 603231 107478
rect 668117 107475 668183 107478
rect 603073 106586 603139 106589
rect 603073 106584 606556 106586
rect 603073 106528 603078 106584
rect 603134 106528 606556 106584
rect 603073 106526 606556 106528
rect 603073 106523 603139 106526
rect 579429 106450 579495 106453
rect 576380 106448 579495 106450
rect 576380 106392 579434 106448
rect 579490 106392 579495 106448
rect 576380 106390 579495 106392
rect 579429 106387 579495 106390
rect 669221 105906 669287 105909
rect 666356 105904 669287 105906
rect 666356 105848 669226 105904
rect 669282 105848 669287 105904
rect 666356 105846 669287 105848
rect 669221 105843 669287 105846
rect 603073 105498 603139 105501
rect 603073 105496 606556 105498
rect 603073 105440 603078 105496
rect 603134 105440 606556 105496
rect 603073 105438 606556 105440
rect 603073 105435 603139 105438
rect 578233 104954 578299 104957
rect 576380 104952 578299 104954
rect 576380 104896 578238 104952
rect 578294 104896 578299 104952
rect 576380 104894 578299 104896
rect 578233 104891 578299 104894
rect 675753 104818 675819 104821
rect 675886 104818 675892 104820
rect 675753 104816 675892 104818
rect 675753 104760 675758 104816
rect 675814 104760 675892 104816
rect 675753 104758 675892 104760
rect 675753 104755 675819 104758
rect 675886 104756 675892 104758
rect 675956 104756 675962 104820
rect 603073 104546 603139 104549
rect 603073 104544 606556 104546
rect 603073 104488 603078 104544
rect 603134 104488 606556 104544
rect 603073 104486 606556 104488
rect 603073 104483 603139 104486
rect 668669 104138 668735 104141
rect 666356 104136 668735 104138
rect 666356 104080 668674 104136
rect 668730 104080 668735 104136
rect 666356 104078 668735 104080
rect 668669 104075 668735 104078
rect 579337 103458 579403 103461
rect 576380 103456 579403 103458
rect 576380 103400 579342 103456
rect 579398 103400 579403 103456
rect 576380 103398 579403 103400
rect 579337 103395 579403 103398
rect 603165 103458 603231 103461
rect 603165 103456 606556 103458
rect 603165 103400 603170 103456
rect 603226 103400 606556 103456
rect 603165 103398 606556 103400
rect 603165 103395 603231 103398
rect 675753 103186 675819 103189
rect 676806 103186 676812 103188
rect 675753 103184 676812 103186
rect 675753 103128 675758 103184
rect 675814 103128 676812 103184
rect 675753 103126 676812 103128
rect 675753 103123 675819 103126
rect 676806 103124 676812 103126
rect 676876 103124 676882 103188
rect 603073 102506 603139 102509
rect 668761 102506 668827 102509
rect 603073 102504 606556 102506
rect 603073 102448 603078 102504
rect 603134 102448 606556 102504
rect 603073 102446 606556 102448
rect 666356 102504 668827 102506
rect 666356 102448 668766 102504
rect 668822 102448 668827 102504
rect 666356 102446 668827 102448
rect 603073 102443 603139 102446
rect 668761 102443 668827 102446
rect 578325 101962 578391 101965
rect 576380 101960 578391 101962
rect 576380 101904 578330 101960
rect 578386 101904 578391 101960
rect 576380 101902 578391 101904
rect 578325 101899 578391 101902
rect 603073 101418 603139 101421
rect 675753 101418 675819 101421
rect 676254 101418 676260 101420
rect 603073 101416 606556 101418
rect 603073 101360 603078 101416
rect 603134 101360 606556 101416
rect 603073 101358 606556 101360
rect 675753 101416 676260 101418
rect 675753 101360 675758 101416
rect 675814 101360 676260 101416
rect 675753 101358 676260 101360
rect 603073 101355 603139 101358
rect 675753 101355 675819 101358
rect 676254 101356 676260 101358
rect 676324 101356 676330 101420
rect 668577 100874 668643 100877
rect 666356 100872 668643 100874
rect 666356 100816 668582 100872
rect 668638 100816 668643 100872
rect 666356 100814 668643 100816
rect 668577 100811 668643 100814
rect 603441 100466 603507 100469
rect 603441 100464 606556 100466
rect 603441 100408 603446 100464
rect 603502 100408 606556 100464
rect 603441 100406 606556 100408
rect 603441 100403 603507 100406
rect 578693 100330 578759 100333
rect 576380 100328 578759 100330
rect 576380 100272 578698 100328
rect 578754 100272 578759 100328
rect 576380 100270 578759 100272
rect 578693 100267 578759 100270
rect 579521 98834 579587 98837
rect 576380 98832 579587 98834
rect 576380 98776 579526 98832
rect 579582 98776 579587 98832
rect 576380 98774 579587 98776
rect 579521 98771 579587 98774
rect 578693 97338 578759 97341
rect 576380 97336 578759 97338
rect 576380 97280 578698 97336
rect 578754 97280 578759 97336
rect 576380 97278 578759 97280
rect 578693 97275 578759 97278
rect 639822 96460 639828 96524
rect 639892 96522 639898 96524
rect 642265 96522 642331 96525
rect 639892 96520 642331 96522
rect 639892 96464 642270 96520
rect 642326 96464 642331 96520
rect 639892 96462 642331 96464
rect 639892 96460 639898 96462
rect 642265 96459 642331 96462
rect 628281 95978 628347 95981
rect 628238 95976 628347 95978
rect 628238 95920 628286 95976
rect 628342 95920 628347 95976
rect 628238 95915 628347 95920
rect 578509 95842 578575 95845
rect 576380 95840 578575 95842
rect 576380 95784 578514 95840
rect 578570 95784 578575 95840
rect 576380 95782 578575 95784
rect 578509 95779 578575 95782
rect 628238 95404 628298 95915
rect 634670 95780 634676 95844
rect 634740 95842 634746 95844
rect 641713 95842 641779 95845
rect 634740 95840 641779 95842
rect 634740 95784 641718 95840
rect 641774 95784 641779 95840
rect 634740 95782 641779 95784
rect 634740 95780 634746 95782
rect 641713 95779 641779 95782
rect 657353 94754 657419 94757
rect 657310 94752 657419 94754
rect 657310 94696 657358 94752
rect 657414 94696 657419 94752
rect 657310 94691 657419 94696
rect 644657 94618 644723 94621
rect 642988 94616 644723 94618
rect 642988 94560 644662 94616
rect 644718 94560 644723 94616
rect 642988 94558 644723 94560
rect 644657 94555 644723 94558
rect 627821 94482 627887 94485
rect 627821 94480 628268 94482
rect 627821 94424 627826 94480
rect 627882 94424 628268 94480
rect 627821 94422 628268 94424
rect 627821 94419 627887 94422
rect 578601 94346 578667 94349
rect 576380 94344 578667 94346
rect 576380 94288 578606 94344
rect 578662 94288 578667 94344
rect 576380 94286 578667 94288
rect 578601 94283 578667 94286
rect 657310 94180 657370 94691
rect 626533 93530 626599 93533
rect 626533 93528 628268 93530
rect 626533 93472 626538 93528
rect 626594 93472 628268 93528
rect 626533 93470 628268 93472
rect 626533 93467 626599 93470
rect 655329 93394 655395 93397
rect 665357 93394 665423 93397
rect 655329 93392 656788 93394
rect 655329 93336 655334 93392
rect 655390 93336 656788 93392
rect 655329 93334 656788 93336
rect 663596 93392 665423 93394
rect 663596 93336 665362 93392
rect 665418 93336 665423 93392
rect 663596 93334 665423 93336
rect 655329 93331 655395 93334
rect 665357 93331 665423 93334
rect 579521 92850 579587 92853
rect 576380 92848 579587 92850
rect 576380 92792 579526 92848
rect 579582 92792 579587 92848
rect 576380 92790 579587 92792
rect 579521 92787 579587 92790
rect 626349 92578 626415 92581
rect 654777 92578 654843 92581
rect 663793 92578 663859 92581
rect 626349 92576 628268 92578
rect 626349 92520 626354 92576
rect 626410 92520 628268 92576
rect 626349 92518 628268 92520
rect 654777 92576 656788 92578
rect 654777 92520 654782 92576
rect 654838 92520 656788 92576
rect 654777 92518 656788 92520
rect 663596 92576 663859 92578
rect 663596 92520 663798 92576
rect 663854 92520 663859 92576
rect 663596 92518 663859 92520
rect 626349 92515 626415 92518
rect 654777 92515 654843 92518
rect 663793 92515 663859 92518
rect 644749 92170 644815 92173
rect 642988 92168 644815 92170
rect 642988 92112 644754 92168
rect 644810 92112 644815 92168
rect 642988 92110 644815 92112
rect 644749 92107 644815 92110
rect 665173 91762 665239 91765
rect 663596 91760 665239 91762
rect 663596 91704 665178 91760
rect 665234 91704 665239 91760
rect 663596 91702 665239 91704
rect 665173 91699 665239 91702
rect 626441 91626 626507 91629
rect 626441 91624 628268 91626
rect 626441 91568 626446 91624
rect 626502 91568 628268 91624
rect 626441 91566 628268 91568
rect 626441 91563 626507 91566
rect 654317 91490 654383 91493
rect 654317 91488 656788 91490
rect 654317 91432 654322 91488
rect 654378 91432 656788 91488
rect 654317 91430 656788 91432
rect 654317 91427 654383 91430
rect 579521 91354 579587 91357
rect 576380 91352 579587 91354
rect 576380 91296 579526 91352
rect 579582 91296 579587 91352
rect 576380 91294 579587 91296
rect 579521 91291 579587 91294
rect 654317 90674 654383 90677
rect 663885 90674 663951 90677
rect 654317 90672 656788 90674
rect 625061 89994 625127 89997
rect 628238 89994 628298 90644
rect 654317 90616 654322 90672
rect 654378 90616 656788 90672
rect 654317 90614 656788 90616
rect 663596 90672 663951 90674
rect 663596 90616 663890 90672
rect 663946 90616 663951 90672
rect 663596 90614 663951 90616
rect 654317 90611 654383 90614
rect 663885 90611 663951 90614
rect 625061 89992 628298 89994
rect 625061 89936 625066 89992
rect 625122 89936 628298 89992
rect 625061 89934 628298 89936
rect 625061 89931 625127 89934
rect 579521 89858 579587 89861
rect 576380 89856 579587 89858
rect 576380 89800 579526 89856
rect 579582 89800 579587 89856
rect 576380 89798 579587 89800
rect 579521 89795 579587 89798
rect 655421 89858 655487 89861
rect 665265 89858 665331 89861
rect 655421 89856 656788 89858
rect 655421 89800 655426 89856
rect 655482 89800 656788 89856
rect 655421 89798 656788 89800
rect 663596 89856 665331 89858
rect 663596 89800 665270 89856
rect 665326 89800 665331 89856
rect 663596 89798 665331 89800
rect 655421 89795 655487 89798
rect 665265 89795 665331 89798
rect 625797 89722 625863 89725
rect 644473 89722 644539 89725
rect 625797 89720 628268 89722
rect 625797 89664 625802 89720
rect 625858 89664 628268 89720
rect 625797 89662 628268 89664
rect 642988 89720 644539 89722
rect 642988 89664 644478 89720
rect 644534 89664 644539 89720
rect 642988 89662 644539 89664
rect 625797 89659 625863 89662
rect 644473 89659 644539 89662
rect 664069 89042 664135 89045
rect 663596 89040 664135 89042
rect 663596 88984 664074 89040
rect 664130 88984 664135 89040
rect 663596 88982 664135 88984
rect 664069 88979 664135 88982
rect 626441 88906 626507 88909
rect 626441 88904 628268 88906
rect 626441 88848 626446 88904
rect 626502 88848 628268 88904
rect 626441 88846 628268 88848
rect 626441 88843 626507 88846
rect 579521 88362 579587 88365
rect 576380 88360 579587 88362
rect 576380 88304 579526 88360
rect 579582 88304 579587 88360
rect 576380 88302 579587 88304
rect 579521 88299 579587 88302
rect 626441 87954 626507 87957
rect 626441 87952 628268 87954
rect 626441 87896 626446 87952
rect 626502 87896 628268 87952
rect 626441 87894 628268 87896
rect 626441 87891 626507 87894
rect 643093 87682 643159 87685
rect 642958 87680 643159 87682
rect 642958 87624 643098 87680
rect 643154 87624 643159 87680
rect 642958 87622 643159 87624
rect 642958 87108 643018 87622
rect 643093 87619 643159 87622
rect 626349 87002 626415 87005
rect 626349 87000 628268 87002
rect 626349 86944 626354 87000
rect 626410 86944 628268 87000
rect 626349 86942 628268 86944
rect 626349 86939 626415 86942
rect 579521 86866 579587 86869
rect 576380 86864 579587 86866
rect 576380 86808 579526 86864
rect 579582 86808 579587 86864
rect 576380 86806 579587 86808
rect 579521 86803 579587 86806
rect 626441 86050 626507 86053
rect 626441 86048 628268 86050
rect 626441 85992 626446 86048
rect 626502 85992 628268 86048
rect 626441 85990 628268 85992
rect 626441 85987 626507 85990
rect 579521 85370 579587 85373
rect 576380 85368 579587 85370
rect 576380 85312 579526 85368
rect 579582 85312 579587 85368
rect 576380 85310 579587 85312
rect 579521 85307 579587 85310
rect 626441 85098 626507 85101
rect 626441 85096 628268 85098
rect 626441 85040 626446 85096
rect 626502 85040 628268 85096
rect 626441 85038 628268 85040
rect 626441 85035 626507 85038
rect 644565 84690 644631 84693
rect 642988 84688 644631 84690
rect 642988 84632 644570 84688
rect 644626 84632 644631 84688
rect 642988 84630 644631 84632
rect 644565 84627 644631 84630
rect 625613 84146 625679 84149
rect 625613 84144 628268 84146
rect 625613 84088 625618 84144
rect 625674 84088 628268 84144
rect 625613 84086 628268 84088
rect 625613 84083 625679 84086
rect 579521 83874 579587 83877
rect 576380 83872 579587 83874
rect 576380 83816 579526 83872
rect 579582 83816 579587 83872
rect 576380 83814 579587 83816
rect 579521 83811 579587 83814
rect 626073 83194 626139 83197
rect 626073 83192 628268 83194
rect 626073 83136 626078 83192
rect 626134 83136 628268 83192
rect 626073 83134 628268 83136
rect 626073 83131 626139 83134
rect 579153 82378 579219 82381
rect 576380 82376 579219 82378
rect 576380 82320 579158 82376
rect 579214 82320 579219 82376
rect 576380 82318 579219 82320
rect 579153 82315 579219 82318
rect 626441 82242 626507 82245
rect 643277 82242 643343 82245
rect 626441 82240 628268 82242
rect 626441 82184 626446 82240
rect 626502 82184 628268 82240
rect 626441 82182 628268 82184
rect 642988 82240 643343 82242
rect 642988 82184 643282 82240
rect 643338 82184 643343 82240
rect 642988 82182 643343 82184
rect 626441 82179 626507 82182
rect 643277 82179 643343 82182
rect 579521 80882 579587 80885
rect 576380 80880 579587 80882
rect 576380 80824 579526 80880
rect 579582 80824 579587 80880
rect 576380 80822 579587 80824
rect 628790 80882 628850 81396
rect 629201 80882 629267 80885
rect 628790 80880 629267 80882
rect 628790 80824 629206 80880
rect 629262 80824 629267 80880
rect 628790 80822 629267 80824
rect 579521 80819 579587 80822
rect 629201 80819 629267 80822
rect 579061 79386 579127 79389
rect 576380 79384 579127 79386
rect 576380 79328 579066 79384
rect 579122 79328 579127 79384
rect 576380 79326 579127 79328
rect 579061 79323 579127 79326
rect 579521 77890 579587 77893
rect 576380 77888 579587 77890
rect 576380 77832 579526 77888
rect 579582 77832 579587 77888
rect 576380 77830 579587 77832
rect 579521 77827 579587 77830
rect 633893 77754 633959 77757
rect 634670 77754 634676 77756
rect 633893 77752 634676 77754
rect 633893 77696 633898 77752
rect 633954 77696 634676 77752
rect 633893 77694 634676 77696
rect 633893 77691 633959 77694
rect 634670 77692 634676 77694
rect 634740 77692 634746 77756
rect 639597 77754 639663 77757
rect 639822 77754 639828 77756
rect 639597 77752 639828 77754
rect 639597 77696 639602 77752
rect 639658 77696 639828 77752
rect 639597 77694 639828 77696
rect 639597 77691 639663 77694
rect 639822 77692 639828 77694
rect 639892 77692 639898 77756
rect 578969 76258 579035 76261
rect 576380 76256 579035 76258
rect 576380 76200 578974 76256
rect 579030 76200 579035 76256
rect 576380 76198 579035 76200
rect 578969 76195 579035 76198
rect 631133 75986 631199 75989
rect 633893 75986 633959 75989
rect 631133 75984 633959 75986
rect 631133 75928 631138 75984
rect 631194 75928 633898 75984
rect 633954 75928 633959 75984
rect 631133 75926 633959 75928
rect 631133 75923 631199 75926
rect 633893 75923 633959 75926
rect 638902 75108 638908 75172
rect 638972 75170 638978 75172
rect 639229 75170 639295 75173
rect 638972 75168 639295 75170
rect 638972 75112 639234 75168
rect 639290 75112 639295 75168
rect 638972 75110 639295 75112
rect 638972 75108 638978 75110
rect 639229 75107 639295 75110
rect 579521 74762 579587 74765
rect 576380 74760 579587 74762
rect 576380 74704 579526 74760
rect 579582 74704 579587 74760
rect 576380 74702 579587 74704
rect 579521 74699 579587 74702
rect 646865 74490 646931 74493
rect 646668 74488 646931 74490
rect 646668 74432 646870 74488
rect 646926 74432 646931 74488
rect 646668 74430 646931 74432
rect 646865 74427 646931 74430
rect 578877 73266 578943 73269
rect 576380 73264 578943 73266
rect 576380 73208 578882 73264
rect 578938 73208 578943 73264
rect 576380 73206 578943 73208
rect 578877 73203 578943 73206
rect 648705 72994 648771 72997
rect 646668 72992 648771 72994
rect 646668 72936 648710 72992
rect 648766 72936 648771 72992
rect 646668 72934 648771 72936
rect 648705 72931 648771 72934
rect 579521 71770 579587 71773
rect 576380 71768 579587 71770
rect 576380 71712 579526 71768
rect 579582 71712 579587 71768
rect 576380 71710 579587 71712
rect 579521 71707 579587 71710
rect 647325 71498 647391 71501
rect 646668 71496 647391 71498
rect 646668 71440 647330 71496
rect 647386 71440 647391 71496
rect 646668 71438 647391 71440
rect 647325 71435 647391 71438
rect 646129 70410 646195 70413
rect 646086 70408 646195 70410
rect 646086 70352 646134 70408
rect 646190 70352 646195 70408
rect 646086 70347 646195 70352
rect 579245 70274 579311 70277
rect 576380 70272 579311 70274
rect 576380 70216 579250 70272
rect 579306 70216 579311 70272
rect 576380 70214 579311 70216
rect 579245 70211 579311 70214
rect 646086 69972 646146 70347
rect 578693 68778 578759 68781
rect 576380 68776 578759 68778
rect 576380 68720 578698 68776
rect 578754 68720 578759 68776
rect 576380 68718 578759 68720
rect 578693 68715 578759 68718
rect 648797 68506 648863 68509
rect 646668 68504 648863 68506
rect 646668 68448 648802 68504
rect 648858 68448 648863 68504
rect 646668 68446 648863 68448
rect 648797 68443 648863 68446
rect 579521 67282 579587 67285
rect 576380 67280 579587 67282
rect 576380 67224 579526 67280
rect 579582 67224 579587 67280
rect 576380 67222 579587 67224
rect 579521 67219 579587 67222
rect 647417 67010 647483 67013
rect 646668 67008 647483 67010
rect 646668 66952 647422 67008
rect 647478 66952 647483 67008
rect 646668 66950 647483 66952
rect 647417 66947 647483 66950
rect 646129 66058 646195 66061
rect 646086 66056 646195 66058
rect 646086 66000 646134 66056
rect 646190 66000 646195 66056
rect 646086 65995 646195 66000
rect 579521 65786 579587 65789
rect 576380 65784 579587 65786
rect 576380 65728 579526 65784
rect 579582 65728 579587 65784
rect 576380 65726 579587 65728
rect 579521 65723 579587 65726
rect 646086 65484 646146 65995
rect 646129 64426 646195 64429
rect 646086 64424 646195 64426
rect 646086 64368 646134 64424
rect 646190 64368 646195 64424
rect 646086 64363 646195 64368
rect 578693 64290 578759 64293
rect 576380 64288 578759 64290
rect 576380 64232 578698 64288
rect 578754 64232 578759 64288
rect 576380 64230 578759 64232
rect 578693 64227 578759 64230
rect 646086 63988 646146 64363
rect 579521 62794 579587 62797
rect 576380 62792 579587 62794
rect 576380 62736 579526 62792
rect 579582 62736 579587 62792
rect 576380 62734 579587 62736
rect 579521 62731 579587 62734
rect 578693 61298 578759 61301
rect 576380 61296 578759 61298
rect 576380 61240 578698 61296
rect 578754 61240 578759 61296
rect 576380 61238 578759 61240
rect 578693 61235 578759 61238
rect 578877 59802 578943 59805
rect 576380 59800 578943 59802
rect 576380 59744 578882 59800
rect 578938 59744 578943 59800
rect 576380 59742 578943 59744
rect 578877 59739 578943 59742
rect 578877 58306 578943 58309
rect 576380 58304 578943 58306
rect 576380 58248 578882 58304
rect 578938 58248 578943 58304
rect 576380 58246 578943 58248
rect 578877 58243 578943 58246
rect 578877 56810 578943 56813
rect 576380 56808 578943 56810
rect 576380 56752 578882 56808
rect 578938 56752 578943 56808
rect 576380 56750 578943 56752
rect 578877 56747 578943 56750
rect 578233 55314 578299 55317
rect 576380 55312 578299 55314
rect 576380 55256 578238 55312
rect 578294 55256 578299 55312
rect 576380 55254 578299 55256
rect 578233 55251 578299 55254
rect 578325 53818 578391 53821
rect 576380 53816 578391 53818
rect 576380 53760 578330 53816
rect 578386 53760 578391 53816
rect 576380 53758 578391 53760
rect 578325 53755 578391 53758
rect 52177 52458 52243 52461
rect 150295 52458 150361 52461
rect 638902 52458 638908 52460
rect 52177 52456 638908 52458
rect 52177 52400 52182 52456
rect 52238 52400 150300 52456
rect 150356 52400 638908 52456
rect 52177 52398 638908 52400
rect 52177 52395 52243 52398
rect 150295 52395 150361 52398
rect 638902 52396 638908 52398
rect 638972 52396 638978 52460
rect 281441 50554 281507 50557
rect 520222 50554 520228 50556
rect 281441 50552 520228 50554
rect 281441 50496 281446 50552
rect 281502 50496 520228 50552
rect 281441 50494 520228 50496
rect 281441 50491 281507 50494
rect 520222 50492 520228 50494
rect 520292 50492 520298 50556
rect 216121 50418 216187 50421
rect 521694 50418 521700 50420
rect 216121 50416 521700 50418
rect 216121 50360 216126 50416
rect 216182 50360 521700 50416
rect 216121 50358 521700 50360
rect 216121 50355 216187 50358
rect 521694 50356 521700 50358
rect 521764 50356 521770 50420
rect 85113 50282 85179 50285
rect 514702 50282 514708 50284
rect 85113 50280 514708 50282
rect 85113 50224 85118 50280
rect 85174 50224 514708 50280
rect 85113 50222 514708 50224
rect 85113 50219 85179 50222
rect 514702 50220 514708 50222
rect 514772 50220 514778 50284
rect 529790 50220 529796 50284
rect 529860 50282 529866 50284
rect 542997 50282 543063 50285
rect 529860 50280 543063 50282
rect 529860 50224 543002 50280
rect 543058 50224 543063 50280
rect 529860 50222 543063 50224
rect 529860 50220 529866 50222
rect 542997 50219 543063 50222
rect 664253 48514 664319 48517
rect 662094 48512 664319 48514
rect 661480 48456 664258 48512
rect 664314 48456 664319 48512
rect 661480 48454 664319 48456
rect 661480 48452 662154 48454
rect 664253 48451 664319 48454
rect 473169 47698 473235 47701
rect 612825 47698 612891 47701
rect 473169 47696 612891 47698
rect 473169 47640 473174 47696
rect 473230 47640 612830 47696
rect 612886 47640 612891 47696
rect 473169 47638 612891 47640
rect 473169 47635 473235 47638
rect 612825 47635 612891 47638
rect 661174 47565 661234 47761
rect 187550 47500 187556 47564
rect 187620 47562 187626 47564
rect 576117 47562 576183 47565
rect 187620 47560 576183 47562
rect 187620 47504 576122 47560
rect 576178 47504 576183 47560
rect 187620 47502 576183 47504
rect 187620 47500 187626 47502
rect 576117 47499 576183 47502
rect 661125 47560 661234 47565
rect 661125 47504 661130 47560
rect 661186 47504 661234 47560
rect 661125 47502 661234 47504
rect 661125 47499 661191 47502
rect 662413 47426 662479 47429
rect 661388 47424 662479 47426
rect 661388 47368 662418 47424
rect 662474 47368 662479 47424
rect 661388 47366 662479 47368
rect 662413 47363 662479 47366
rect 412449 46746 412515 46749
rect 518566 46746 518572 46748
rect 412449 46744 518572 46746
rect 412449 46688 412454 46744
rect 412510 46688 518572 46744
rect 412449 46686 518572 46688
rect 412449 46683 412515 46686
rect 518566 46684 518572 46686
rect 518636 46684 518642 46748
rect 471646 46548 471652 46612
rect 471716 46610 471722 46612
rect 611353 46610 611419 46613
rect 471716 46608 611419 46610
rect 471716 46552 611358 46608
rect 611414 46552 611419 46608
rect 471716 46550 611419 46552
rect 471716 46548 471722 46550
rect 611353 46547 611419 46550
rect 470133 46474 470199 46477
rect 612733 46474 612799 46477
rect 470133 46472 612799 46474
rect 470133 46416 470138 46472
rect 470194 46416 612738 46472
rect 612794 46416 612799 46472
rect 470133 46414 612799 46416
rect 470133 46411 470199 46414
rect 612733 46411 612799 46414
rect 460606 46276 460612 46340
rect 460676 46338 460682 46340
rect 611445 46338 611511 46341
rect 460676 46336 611511 46338
rect 460676 46280 611450 46336
rect 611506 46280 611511 46336
rect 460676 46278 611511 46280
rect 460676 46276 460682 46278
rect 611445 46275 611511 46278
rect 415117 46202 415183 46205
rect 610157 46202 610223 46205
rect 415117 46200 610223 46202
rect 415117 46144 415122 46200
rect 415178 46144 610162 46200
rect 610218 46144 610223 46200
rect 415117 46142 610223 46144
rect 415117 46139 415183 46142
rect 610157 46139 610223 46142
rect 419717 45250 419783 45253
rect 610065 45250 610131 45253
rect 419717 45248 610131 45250
rect 419717 45192 419722 45248
rect 419778 45192 610070 45248
rect 610126 45192 610131 45248
rect 419717 45190 610131 45192
rect 419717 45187 419783 45190
rect 610065 45187 610131 45190
rect 365110 45052 365116 45116
rect 365180 45114 365186 45116
rect 607305 45114 607371 45117
rect 365180 45112 607371 45114
rect 365180 45056 607310 45112
rect 607366 45056 607371 45112
rect 365180 45054 607371 45056
rect 365180 45052 365186 45054
rect 607305 45051 607371 45054
rect 361982 44916 361988 44980
rect 362052 44978 362058 44980
rect 605833 44978 605899 44981
rect 362052 44976 605899 44978
rect 362052 44920 605838 44976
rect 605894 44920 605899 44976
rect 362052 44918 605899 44920
rect 362052 44916 362058 44918
rect 605833 44915 605899 44918
rect 310094 44780 310100 44844
rect 310164 44842 310170 44844
rect 608593 44842 608659 44845
rect 310164 44840 608659 44842
rect 310164 44784 608598 44840
rect 608654 44784 608659 44840
rect 310164 44782 608659 44784
rect 310164 44780 310170 44782
rect 608593 44779 608659 44782
rect 142337 44298 142403 44301
rect 142110 44296 142403 44298
rect 142110 44240 142342 44296
rect 142398 44240 142403 44296
rect 142110 44238 142403 44240
rect 141918 43964 141924 44028
rect 141988 44026 141994 44028
rect 142110 44026 142170 44238
rect 142337 44235 142403 44238
rect 141988 43966 142170 44026
rect 141988 43964 141994 43966
rect 307293 43482 307359 43485
rect 607213 43482 607279 43485
rect 307293 43480 607279 43482
rect 307293 43424 307298 43480
rect 307354 43424 607218 43480
rect 607274 43424 607279 43480
rect 307293 43422 607279 43424
rect 307293 43419 307359 43422
rect 607213 43419 607279 43422
rect 310099 42396 310165 42397
rect 518617 42396 518683 42397
rect 310094 42394 310100 42396
rect 310008 42334 310100 42394
rect 310094 42332 310100 42334
rect 310164 42332 310170 42396
rect 518566 42332 518572 42396
rect 518636 42394 518683 42396
rect 518636 42392 518728 42394
rect 518678 42336 518728 42392
rect 518636 42334 518728 42336
rect 518636 42332 518683 42334
rect 310099 42331 310165 42332
rect 518617 42331 518683 42332
rect 187509 42124 187575 42125
rect 361941 42124 362007 42125
rect 365069 42124 365135 42125
rect 460565 42124 460631 42125
rect 471605 42124 471671 42125
rect 187509 42122 187556 42124
rect 187464 42120 187556 42122
rect 187464 42064 187514 42120
rect 187464 42062 187556 42064
rect 187509 42060 187556 42062
rect 187620 42060 187626 42124
rect 361941 42122 361988 42124
rect 361896 42120 361988 42122
rect 361896 42064 361946 42120
rect 361896 42062 361988 42064
rect 361941 42060 361988 42062
rect 362052 42060 362058 42124
rect 365069 42122 365116 42124
rect 365024 42120 365116 42122
rect 365024 42064 365074 42120
rect 365024 42062 365116 42064
rect 365069 42060 365116 42062
rect 365180 42060 365186 42124
rect 460565 42122 460612 42124
rect 460520 42120 460612 42122
rect 460520 42064 460570 42120
rect 460520 42062 460612 42064
rect 460565 42060 460612 42062
rect 460676 42060 460682 42124
rect 471605 42122 471652 42124
rect 471560 42120 471652 42122
rect 471560 42064 471610 42120
rect 471560 42062 471652 42064
rect 471605 42060 471652 42062
rect 471716 42060 471722 42124
rect 514702 42060 514708 42124
rect 514772 42122 514778 42124
rect 514845 42122 514911 42125
rect 514772 42120 514911 42122
rect 514772 42064 514850 42120
rect 514906 42064 514911 42120
rect 514772 42062 514911 42064
rect 514772 42060 514778 42062
rect 187509 42059 187575 42060
rect 361941 42059 362007 42060
rect 365069 42059 365135 42060
rect 460565 42059 460631 42060
rect 471605 42059 471671 42060
rect 514845 42059 514911 42062
rect 520222 42060 520228 42124
rect 520292 42122 520298 42124
rect 520365 42122 520431 42125
rect 521745 42124 521811 42125
rect 520292 42120 520431 42122
rect 520292 42064 520370 42120
rect 520426 42064 520431 42120
rect 520292 42062 520431 42064
rect 520292 42060 520298 42062
rect 520365 42059 520431 42062
rect 521694 42060 521700 42124
rect 521764 42122 521811 42124
rect 529657 42122 529723 42125
rect 529790 42122 529796 42124
rect 521764 42120 521856 42122
rect 521806 42064 521856 42120
rect 521764 42062 521856 42064
rect 529657 42120 529796 42122
rect 529657 42064 529662 42120
rect 529718 42064 529796 42120
rect 529657 42062 529796 42064
rect 521764 42060 521811 42062
rect 521745 42059 521811 42060
rect 529657 42059 529723 42062
rect 529790 42060 529796 42062
rect 529860 42060 529866 42124
rect 416681 41850 416747 41853
rect 525885 41850 525951 41853
rect 416681 41848 422310 41850
rect 416681 41792 416686 41848
rect 416742 41792 422310 41848
rect 416681 41790 422310 41792
rect 416681 41787 416747 41790
rect 422250 41442 422310 41790
rect 509190 41848 525951 41850
rect 509190 41792 525890 41848
rect 525946 41792 525951 41848
rect 509190 41790 525951 41792
rect 478781 41578 478847 41581
rect 509190 41578 509250 41790
rect 525885 41787 525951 41790
rect 478781 41576 509250 41578
rect 478781 41520 478786 41576
rect 478842 41520 509250 41576
rect 478781 41518 509250 41520
rect 478781 41515 478847 41518
rect 609973 41442 610039 41445
rect 422250 41440 610039 41442
rect 422250 41384 609978 41440
rect 610034 41384 610039 41440
rect 422250 41382 610039 41384
rect 609973 41379 610039 41382
rect 141693 40354 141759 40357
rect 141918 40354 141924 40356
rect 141693 40352 141924 40354
rect 141693 40296 141698 40352
rect 141754 40296 141924 40352
rect 141693 40294 141924 40296
rect 141693 40291 141759 40294
rect 141918 40292 141924 40294
rect 141988 40292 141994 40356
<< via3 >>
rect 246436 997324 246500 997388
rect 238524 997188 238588 997252
rect 480668 997188 480732 997252
rect 532004 997188 532068 997252
rect 627868 996644 627932 996708
rect 86540 996508 86604 996572
rect 89668 996372 89732 996436
rect 135300 996236 135364 996300
rect 86540 995752 86604 995756
rect 86540 995696 86554 995752
rect 86554 995696 86604 995752
rect 86540 995692 86604 995696
rect 89668 995752 89732 995756
rect 89668 995696 89682 995752
rect 89682 995696 89732 995752
rect 89668 995692 89732 995696
rect 135300 995692 135364 995756
rect 238524 995752 238588 995756
rect 238524 995696 238574 995752
rect 238574 995696 238588 995752
rect 238524 995692 238588 995696
rect 240364 995692 240428 995756
rect 439820 995752 439884 995756
rect 439820 995696 439834 995752
rect 439834 995696 439884 995752
rect 439820 995692 439884 995696
rect 630260 996508 630324 996572
rect 554636 995828 554700 995892
rect 480668 995692 480732 995756
rect 485636 995752 485700 995756
rect 485636 995696 485650 995752
rect 485650 995696 485700 995752
rect 485636 995692 485700 995696
rect 532004 995692 532068 995756
rect 536604 995752 536668 995756
rect 536604 995696 536618 995752
rect 536618 995696 536668 995752
rect 536604 995692 536668 995696
rect 573220 995692 573284 995756
rect 627868 995752 627932 995756
rect 627868 995696 627918 995752
rect 627918 995696 627932 995752
rect 627868 995692 627932 995696
rect 630260 995752 630324 995756
rect 630260 995696 630310 995752
rect 630310 995696 630324 995752
rect 630260 995692 630324 995696
rect 505140 992292 505204 992356
rect 439820 991476 439884 991540
rect 573220 990932 573284 990996
rect 40540 968764 40604 968828
rect 40724 967268 40788 967332
rect 676812 966452 676876 966516
rect 676444 966180 676508 966244
rect 42012 965152 42076 965156
rect 42012 965096 42062 965152
rect 42062 965096 42076 965152
rect 42012 965092 42076 965096
rect 677180 964956 677244 965020
rect 40356 963324 40420 963388
rect 675340 963384 675404 963388
rect 675340 963328 675390 963384
rect 675390 963328 675404 963384
rect 675340 963324 675404 963328
rect 41460 962100 41524 962164
rect 675892 961284 675956 961348
rect 675708 959168 675772 959172
rect 675708 959112 675722 959168
rect 675722 959112 675772 959168
rect 675708 959108 675772 959112
rect 676996 958972 677060 959036
rect 41644 958292 41708 958356
rect 42196 957748 42260 957812
rect 675524 957808 675588 957812
rect 675524 957752 675538 957808
rect 675538 957752 675588 957808
rect 675524 957748 675588 957752
rect 676628 957612 676692 957676
rect 676076 953940 676140 954004
rect 41644 952172 41708 952236
rect 42196 951764 42260 951828
rect 41460 951628 41524 951692
rect 42012 951628 42076 951692
rect 676444 950948 676508 951012
rect 676812 950812 676876 950876
rect 675340 949724 675404 949788
rect 675524 949588 675588 949652
rect 675892 949452 675956 949516
rect 675708 948772 675772 948836
rect 676076 947956 676140 948020
rect 41828 938572 41892 938636
rect 41828 936940 41892 937004
rect 677180 935580 677244 935644
rect 41828 934900 41892 934964
rect 676996 932724 677060 932788
rect 676628 932316 676692 932380
rect 676628 876556 676692 876620
rect 676812 876420 676876 876484
rect 676076 874108 676140 874172
rect 677180 872748 677244 872812
rect 673868 872204 673932 872268
rect 675892 864724 675956 864788
rect 41828 816036 41892 816100
rect 41690 814268 41754 814332
rect 41828 813180 41892 813244
rect 40540 804748 40604 804812
rect 42196 802708 42260 802772
rect 41644 802572 41708 802636
rect 42012 802436 42076 802500
rect 41828 800940 41892 801004
rect 40540 796724 40604 796788
rect 42012 791964 42076 792028
rect 42196 788760 42260 788764
rect 42196 788704 42210 788760
rect 42210 788704 42260 788760
rect 42196 788700 42260 788704
rect 41828 788156 41892 788220
rect 41644 788020 41708 788084
rect 675340 788080 675404 788084
rect 675340 788024 675390 788080
rect 675390 788024 675404 788080
rect 675340 788020 675404 788024
rect 41460 786932 41524 786996
rect 675708 786720 675772 786724
rect 675708 786664 675758 786720
rect 675758 786664 675772 786720
rect 675708 786660 675772 786664
rect 675524 784816 675588 784820
rect 675524 784760 675538 784816
rect 675538 784760 675588 784816
rect 675524 784756 675588 784760
rect 676996 784076 677060 784140
rect 675892 774828 675956 774892
rect 677180 774828 677244 774892
rect 675340 773876 675404 773940
rect 40172 773468 40236 773532
rect 675524 773392 675588 773396
rect 675524 773336 675538 773392
rect 675538 773336 675588 773392
rect 675524 773332 675588 773336
rect 675708 773392 675772 773396
rect 675708 773336 675722 773392
rect 675722 773336 675772 773392
rect 675708 773332 675772 773336
rect 676812 773060 676876 773124
rect 676628 772924 676692 772988
rect 676076 772652 676140 772716
rect 39988 771836 40052 771900
rect 39988 771020 40052 771084
rect 675156 766532 675220 766596
rect 676076 766532 676140 766596
rect 40908 766124 40972 766188
rect 674972 765036 675036 765100
rect 40540 764900 40604 764964
rect 40724 764492 40788 764556
rect 674788 759052 674852 759116
rect 41644 758236 41708 758300
rect 674788 757828 674852 757892
rect 41460 757692 41524 757756
rect 41828 757072 41892 757076
rect 41828 757016 41842 757072
rect 41842 757016 41892 757072
rect 41828 757012 41892 757016
rect 42380 757072 42444 757076
rect 42380 757016 42430 757072
rect 42430 757016 42444 757072
rect 42380 757012 42444 757016
rect 677180 756740 677244 756804
rect 41828 754896 41892 754900
rect 41828 754840 41878 754896
rect 41878 754840 41892 754896
rect 41828 754836 41892 754840
rect 40724 754156 40788 754220
rect 677364 753884 677428 753948
rect 40908 753068 40972 753132
rect 673868 752524 673932 752588
rect 40540 750348 40604 750412
rect 42380 749260 42444 749324
rect 41644 746540 41708 746604
rect 41460 742324 41524 742388
rect 675708 741704 675772 741708
rect 675708 741648 675722 741704
rect 675722 741648 675772 741704
rect 675708 741644 675772 741648
rect 675524 736068 675588 736132
rect 676628 734300 676692 734364
rect 677180 732940 677244 733004
rect 40356 729404 40420 729468
rect 39988 728588 40052 728652
rect 675524 728376 675588 728380
rect 675524 728320 675538 728376
rect 675538 728320 675588 728376
rect 675524 728316 675588 728320
rect 675708 728376 675772 728380
rect 675708 728320 675722 728376
rect 675722 728320 675772 728376
rect 675708 728316 675772 728320
rect 40172 727772 40236 727836
rect 674972 727228 675036 727292
rect 675156 726548 675220 726612
rect 41460 725324 41524 725388
rect 676076 724372 676140 724436
rect 675892 721496 675956 721560
rect 676076 721496 676140 721560
rect 40540 721244 40604 721308
rect 41644 716076 41708 716140
rect 41828 715396 41892 715460
rect 42012 713824 42076 713828
rect 42012 713768 42062 713824
rect 42062 713768 42076 713824
rect 42012 713764 42076 713768
rect 676996 713488 677060 713492
rect 676996 713432 677010 713488
rect 677010 713432 677060 713488
rect 676996 713428 677060 713432
rect 42196 713220 42260 713284
rect 40540 710772 40604 710836
rect 42196 708460 42260 708524
rect 42012 706752 42076 706756
rect 42012 706696 42062 706752
rect 42062 706696 42076 706752
rect 42012 706692 42076 706696
rect 41828 703700 41892 703764
rect 41460 702340 41524 702404
rect 41644 699348 41708 699412
rect 675340 696960 675404 696964
rect 675340 696904 675390 696960
rect 675390 696904 675404 696960
rect 675340 696900 675404 696904
rect 675524 694784 675588 694788
rect 675524 694728 675538 694784
rect 675538 694728 675588 694784
rect 675524 694724 675588 694728
rect 676444 694180 676508 694244
rect 676812 687380 676876 687444
rect 40356 687108 40420 687172
rect 675708 686216 675772 686220
rect 675708 686160 675722 686216
rect 675722 686160 675772 686216
rect 675708 686156 675772 686160
rect 40172 685476 40236 685540
rect 39988 684660 40052 684724
rect 675340 683360 675404 683364
rect 675340 683304 675390 683360
rect 675390 683304 675404 683360
rect 675340 683300 675404 683304
rect 675524 683300 675588 683364
rect 675708 683164 675772 683228
rect 676444 683164 676508 683228
rect 41460 682212 41524 682276
rect 675892 681804 675956 681868
rect 40540 679356 40604 679420
rect 676076 678268 676140 678332
rect 40724 678132 40788 678196
rect 30604 677724 30668 677788
rect 30604 676500 30668 676564
rect 675156 676364 675220 676428
rect 675892 676364 675956 676428
rect 676996 676364 677060 676428
rect 41644 671332 41708 671396
rect 42380 670924 42444 670988
rect 41828 670712 41892 670716
rect 41828 670656 41842 670712
rect 41842 670656 41892 670712
rect 41828 670652 41892 670656
rect 42012 670712 42076 670716
rect 42012 670656 42062 670712
rect 42062 670656 42076 670712
rect 42012 670652 42076 670656
rect 42196 670108 42260 670172
rect 672948 669020 673012 669084
rect 41828 668536 41892 668540
rect 41828 668480 41878 668536
rect 41878 668480 41892 668536
rect 41828 668476 41892 668480
rect 41828 668340 41892 668404
rect 42380 668340 42444 668404
rect 40724 665348 40788 665412
rect 40540 664532 40604 664596
rect 42012 663368 42076 663372
rect 42012 663312 42062 663368
rect 42062 663312 42076 663368
rect 42012 663308 42076 663312
rect 677180 663308 677244 663372
rect 676628 662900 676692 662964
rect 41460 661268 41524 661332
rect 42196 660512 42260 660516
rect 42196 660456 42210 660512
rect 42210 660456 42260 660512
rect 42196 660452 42260 660456
rect 41828 660316 41892 660380
rect 41644 658276 41708 658340
rect 675340 649904 675404 649908
rect 675340 649848 675390 649904
rect 675390 649848 675404 649904
rect 675340 649844 675404 649848
rect 676628 648620 676692 648684
rect 675524 645900 675588 645964
rect 677180 644676 677244 644740
rect 677180 644540 677244 644604
rect 39988 642228 40052 642292
rect 39988 641412 40052 641476
rect 41460 639372 41524 639436
rect 675340 638692 675404 638756
rect 675524 638208 675588 638212
rect 675524 638152 675538 638208
rect 675538 638152 675588 638208
rect 675524 638148 675588 638152
rect 676628 637876 676692 637940
rect 676996 637876 677060 637940
rect 675892 637468 675956 637532
rect 675156 637332 675220 637396
rect 40908 636516 40972 636580
rect 40540 636108 40604 636172
rect 40724 634884 40788 634948
rect 676076 631348 676140 631412
rect 676996 631348 677060 631412
rect 41644 629852 41708 629916
rect 42196 629172 42260 629236
rect 42012 629036 42076 629100
rect 41828 628492 41892 628556
rect 40908 625228 40972 625292
rect 40724 623732 40788 623796
rect 40540 621420 40604 621484
rect 42012 618972 42076 619036
rect 676812 618292 676876 618356
rect 41828 616796 41892 616860
rect 42196 616720 42260 616724
rect 42196 616664 42210 616720
rect 42210 616664 42260 616720
rect 42196 616660 42260 616664
rect 41460 614076 41524 614140
rect 41644 613396 41708 613460
rect 675340 606520 675404 606524
rect 675340 606464 675390 606520
rect 675390 606464 675404 606520
rect 675340 606460 675404 606464
rect 675708 600884 675772 600948
rect 39988 598980 40052 599044
rect 676812 598980 676876 599044
rect 39988 598164 40052 598228
rect 675524 595368 675588 595372
rect 675524 595312 675574 595368
rect 675574 595312 675588 595368
rect 675524 595308 675588 595312
rect 675708 593192 675772 593196
rect 675708 593136 675758 593192
rect 675758 593136 675772 593192
rect 675708 593132 675772 593136
rect 675524 593056 675588 593060
rect 675524 593000 675574 593056
rect 675574 593000 675588 593056
rect 675524 592996 675588 593000
rect 40540 592044 40604 592108
rect 675340 592044 675404 592108
rect 676996 592044 677060 592108
rect 40724 591636 40788 591700
rect 676076 591364 676140 591428
rect 41460 587148 41524 587212
rect 675708 586196 675772 586260
rect 676076 586196 676140 586260
rect 40908 585440 40972 585444
rect 40908 585384 40922 585440
rect 40922 585384 40972 585440
rect 40908 585380 40972 585384
rect 42380 585108 42444 585172
rect 42012 584584 42076 584648
rect 675892 584564 675956 584628
rect 41644 584508 41708 584512
rect 41644 584452 41658 584508
rect 41658 584452 41708 584508
rect 41644 584448 41708 584452
rect 42564 584156 42628 584220
rect 40908 581708 40972 581772
rect 41644 580212 41708 580276
rect 40724 578988 40788 579052
rect 40540 577492 40604 577556
rect 42380 574016 42444 574020
rect 42380 573960 42394 574016
rect 42394 573960 42444 574016
rect 42380 573956 42444 573960
rect 42564 573820 42628 573884
rect 677180 573140 677244 573204
rect 677364 572732 677428 572796
rect 42012 571508 42076 571572
rect 41460 570420 41524 570484
rect 676628 562668 676692 562732
rect 675340 561172 675404 561236
rect 675524 559600 675588 559604
rect 675524 559544 675574 559600
rect 675574 559544 675588 559600
rect 675524 559540 675588 559544
rect 677180 558996 677244 559060
rect 39988 555868 40052 555932
rect 675524 554780 675588 554844
rect 677180 553964 677244 554028
rect 676996 551924 677060 551988
rect 40724 550564 40788 550628
rect 675340 550292 675404 550356
rect 40540 549340 40604 549404
rect 40908 548932 40972 548996
rect 675708 546756 675772 546820
rect 675892 546620 675956 546684
rect 676628 546484 676692 546548
rect 41460 545124 41524 545188
rect 676812 543628 676876 543692
rect 41644 542948 41708 543012
rect 676076 542948 676140 543012
rect 41828 542812 41892 542876
rect 42012 542268 42076 542332
rect 42012 535876 42076 535940
rect 40908 534516 40972 534580
rect 40724 534108 40788 534172
rect 41828 532612 41892 532676
rect 40540 531388 40604 531452
rect 41460 529892 41524 529956
rect 41644 529348 41708 529412
rect 677364 492416 677428 492420
rect 677364 492360 677414 492416
rect 677414 492360 677428 492416
rect 677364 492356 677428 492360
rect 676076 484060 676140 484124
rect 676076 483652 676140 483716
rect 672948 474812 673012 474876
rect 41828 426396 41892 426460
rect 41828 425580 41892 425644
rect 42196 424764 42260 424828
rect 41828 423948 41892 424012
rect 42012 423540 42076 423604
rect 41828 422724 41892 422788
rect 40055 420678 40119 420742
rect 40055 419450 40119 419514
rect 41828 415244 41892 415308
rect 42012 414972 42076 415036
rect 41460 414700 41524 414764
rect 41828 414564 41892 414628
rect 41828 411224 41892 411228
rect 41828 411168 41878 411224
rect 41878 411168 41892 411224
rect 41828 411164 41892 411168
rect 41092 409396 41156 409460
rect 41644 406268 41708 406332
rect 42012 402520 42076 402524
rect 42012 402464 42062 402520
rect 42062 402464 42076 402520
rect 42012 402460 42076 402464
rect 41460 401780 41524 401844
rect 40540 400012 40604 400076
rect 40908 399604 40972 399668
rect 675892 399332 675956 399396
rect 40724 398788 40788 398852
rect 676260 398788 676324 398852
rect 676444 397156 676508 397220
rect 676076 395116 676140 395180
rect 675524 388452 675588 388516
rect 675708 387636 675772 387700
rect 675340 387500 675404 387564
rect 675892 384916 675956 384980
rect 40724 383012 40788 383076
rect 40540 382196 40604 382260
rect 675340 382256 675404 382260
rect 675340 382200 675390 382256
rect 675390 382200 675404 382256
rect 675340 382196 675404 382200
rect 41460 381788 41524 381852
rect 40908 379748 40972 379812
rect 675524 378720 675588 378724
rect 675524 378664 675538 378720
rect 675538 378664 675588 378720
rect 675524 378660 675588 378664
rect 676076 377572 676140 377636
rect 675708 375456 675772 375460
rect 675708 375400 675758 375456
rect 675758 375400 675772 375456
rect 675708 375396 675772 375400
rect 676260 373628 676324 373692
rect 676444 371996 676508 372060
rect 42012 371860 42076 371924
rect 41644 371316 41708 371380
rect 41828 370288 41892 370292
rect 41828 370232 41842 370288
rect 41842 370232 41892 370288
rect 41828 370228 41892 370232
rect 41828 366344 41892 366348
rect 41828 366288 41878 366344
rect 41878 366288 41892 366344
rect 41828 366284 41892 366288
rect 42012 363760 42076 363764
rect 42012 363704 42026 363760
rect 42026 363704 42076 363760
rect 42012 363700 42076 363704
rect 41644 362884 41708 362948
rect 40908 360164 40972 360228
rect 41460 358668 41524 358732
rect 40724 356900 40788 356964
rect 40540 355676 40604 355740
rect 675524 354180 675588 354244
rect 676076 353636 676140 353700
rect 675340 353364 675404 353428
rect 675892 352956 675956 353020
rect 676076 352004 676140 352068
rect 676812 351086 676876 351150
rect 676628 346564 676692 346628
rect 677180 346428 677244 346492
rect 675524 343572 675588 343636
rect 675708 340776 675772 340780
rect 675708 340720 675722 340776
rect 675722 340720 675772 340776
rect 675708 340716 675772 340720
rect 40724 339764 40788 339828
rect 675892 339356 675956 339420
rect 40540 338948 40604 339012
rect 42012 338812 42076 338876
rect 676076 337860 676140 337924
rect 40908 337316 40972 337380
rect 41644 336908 41708 336972
rect 676996 335820 677060 335884
rect 41276 335684 41340 335748
rect 41092 335276 41156 335340
rect 676812 335276 676876 335340
rect 675524 333568 675588 333572
rect 675524 333512 675538 333568
rect 675538 333512 675588 333568
rect 675524 333508 675588 333512
rect 676628 332556 676692 332620
rect 41460 327796 41524 327860
rect 41828 327660 41892 327724
rect 676444 325620 676508 325684
rect 676260 325484 676324 325548
rect 41828 324864 41892 324868
rect 41828 324808 41842 324864
rect 41842 324808 41892 324864
rect 41828 324804 41892 324808
rect 41276 321132 41340 321196
rect 41460 319908 41524 319972
rect 41092 317324 41156 317388
rect 41644 315828 41708 315892
rect 42012 315480 42076 315484
rect 42012 315424 42026 315480
rect 42026 315424 42076 315480
rect 42012 315420 42076 315424
rect 40724 313788 40788 313852
rect 40908 313108 40972 313172
rect 40540 312292 40604 312356
rect 676444 308620 676508 308684
rect 675892 307940 675956 308004
rect 676260 306988 676324 307052
rect 676076 305356 676140 305420
rect 676628 304948 676692 305012
rect 675708 299372 675772 299436
rect 675892 297876 675956 297940
rect 675340 297332 675404 297396
rect 42748 296788 42812 296852
rect 41828 295972 41892 296036
rect 42012 295564 42076 295628
rect 675708 294808 675772 294812
rect 675708 294752 675758 294808
rect 675758 294752 675772 294808
rect 675708 294748 675772 294752
rect 41828 294340 41892 294404
rect 42564 293932 42628 293996
rect 41828 293116 41892 293180
rect 41828 292708 41892 292772
rect 675524 292632 675588 292636
rect 675524 292576 675538 292632
rect 675538 292576 675588 292632
rect 675524 292572 675588 292576
rect 675340 292088 675404 292092
rect 675340 292032 675390 292088
rect 675390 292032 675404 292088
rect 675340 292028 675404 292032
rect 675708 288416 675772 288420
rect 675708 288360 675722 288416
rect 675722 288360 675772 288416
rect 675708 288356 675772 288360
rect 676628 287268 676692 287332
rect 676076 285500 676140 285564
rect 41460 284820 41524 284884
rect 676444 283596 676508 283660
rect 41460 281420 41524 281484
rect 676260 281420 676324 281484
rect 40908 279788 40972 279852
rect 41092 278020 41156 278084
rect 41828 273048 41892 273052
rect 41828 272992 41842 273048
rect 41842 272992 41892 273048
rect 41828 272988 41892 272992
rect 41644 272172 41708 272236
rect 42012 270464 42076 270468
rect 42012 270408 42026 270464
rect 42026 270408 42076 270464
rect 42012 270404 42076 270408
rect 40724 269724 40788 269788
rect 40540 269044 40604 269108
rect 677180 260748 677244 260812
rect 676996 260340 677060 260404
rect 676812 259524 676876 259588
rect 175044 253132 175108 253196
rect 675156 251500 675220 251564
rect 40540 250140 40604 250204
rect 40724 249732 40788 249796
rect 675156 249596 675220 249660
rect 677180 246604 677244 246668
rect 675708 245652 675772 245716
rect 676812 245380 676876 245444
rect 175044 241632 175108 241636
rect 175044 241576 175058 241632
rect 175058 241576 175108 241632
rect 175044 241572 175108 241576
rect 42012 238036 42076 238100
rect 676996 238580 677060 238644
rect 42196 237356 42260 237420
rect 675708 236872 675772 236876
rect 675708 236816 675758 236872
rect 675758 236816 675772 236872
rect 675708 236812 675772 236816
rect 40724 236676 40788 236740
rect 40540 232868 40604 232932
rect 647372 231100 647436 231164
rect 646452 229604 646516 229668
rect 42196 228984 42260 228988
rect 42196 228928 42210 228984
rect 42210 228928 42260 228984
rect 42196 228924 42260 228928
rect 42012 227352 42076 227356
rect 42012 227296 42026 227352
rect 42026 227296 42076 227352
rect 42012 227292 42076 227296
rect 675892 218588 675956 218652
rect 675708 218180 675772 218244
rect 675524 217772 675588 217836
rect 676628 215494 676692 215558
rect 676996 214270 677060 214334
rect 676076 214024 676140 214028
rect 676076 213968 676090 214024
rect 676090 213968 676140 214024
rect 676076 213964 676140 213968
rect 646452 213012 646516 213076
rect 647372 213012 647436 213076
rect 676812 211380 676876 211444
rect 676444 211244 676508 211308
rect 675708 209884 675772 209948
rect 41644 209748 41708 209812
rect 675892 209612 675956 209676
rect 40540 209340 40604 209404
rect 41460 208524 41524 208588
rect 676076 208252 676140 208316
rect 675340 207164 675404 207228
rect 40724 206892 40788 206956
rect 675892 205532 675956 205596
rect 676076 204988 676140 205052
rect 675708 204232 675772 204236
rect 675708 204176 675758 204232
rect 675758 204176 675772 204232
rect 675708 204172 675772 204176
rect 676996 202812 677060 202876
rect 675524 202736 675588 202740
rect 675524 202680 675538 202736
rect 675538 202680 675588 202736
rect 675524 202676 675588 202680
rect 676812 201316 676876 201380
rect 41828 199276 41892 199340
rect 676076 198324 676140 198388
rect 40724 195332 40788 195396
rect 42196 195332 42260 195396
rect 676628 195332 676692 195396
rect 41644 195196 41708 195260
rect 676444 190300 676508 190364
rect 41460 190164 41524 190228
rect 676260 190164 676324 190228
rect 42196 187368 42260 187372
rect 42196 187312 42210 187368
rect 42210 187312 42260 187368
rect 42196 187308 42260 187312
rect 41828 184240 41892 184244
rect 41828 184184 41878 184240
rect 41878 184184 41892 184240
rect 41828 184180 41892 184184
rect 40540 182956 40604 183020
rect 675340 173980 675404 174044
rect 676076 173436 676140 173500
rect 676076 171804 676140 171868
rect 675892 170716 675956 170780
rect 675708 169628 675772 169692
rect 676628 166424 676692 166428
rect 676628 166368 676642 166424
rect 676642 166368 676692 166424
rect 676628 166364 676692 166368
rect 676812 166424 676876 166428
rect 676812 166368 676826 166424
rect 676826 166368 676876 166424
rect 676812 166364 676876 166368
rect 676076 162692 676140 162756
rect 675524 162556 675588 162620
rect 676812 159972 676876 160036
rect 675340 159428 675404 159492
rect 675708 157448 675772 157452
rect 675708 157392 675722 157448
rect 675722 157392 675772 157448
rect 675708 157388 675772 157392
rect 675524 157040 675588 157044
rect 675524 156984 675538 157040
rect 675538 156984 675588 157040
rect 675524 156980 675588 156984
rect 675892 156300 675956 156364
rect 676076 153036 676140 153100
rect 676628 151540 676692 151604
rect 676444 148412 676508 148476
rect 676260 146236 676324 146300
rect 675340 128828 675404 128892
rect 676260 126516 676324 126580
rect 675708 124884 675772 124948
rect 676444 124476 676508 124540
rect 676812 121620 676876 121684
rect 676076 117948 676140 118012
rect 675892 117268 675956 117332
rect 675524 117132 675588 117196
rect 675340 114200 675404 114204
rect 675340 114144 675390 114200
rect 675390 114144 675404 114200
rect 675340 114140 675404 114144
rect 675708 112568 675772 112572
rect 675708 112512 675722 112568
rect 675722 112512 675772 112568
rect 675708 112508 675772 112512
rect 675524 111752 675588 111756
rect 675524 111696 675538 111752
rect 675538 111696 675588 111752
rect 675524 111692 675588 111696
rect 676444 108972 676508 109036
rect 676076 108156 676140 108220
rect 675892 104756 675956 104820
rect 676812 103124 676876 103188
rect 676260 101356 676324 101420
rect 639828 96460 639892 96524
rect 634676 95780 634740 95844
rect 634676 77692 634740 77756
rect 639828 77692 639892 77756
rect 638908 75108 638972 75172
rect 638908 52396 638972 52460
rect 520228 50492 520292 50556
rect 521700 50356 521764 50420
rect 514708 50220 514772 50284
rect 529796 50220 529860 50284
rect 187556 47500 187620 47564
rect 518572 46684 518636 46748
rect 471652 46548 471716 46612
rect 460612 46276 460676 46340
rect 365116 45052 365180 45116
rect 361988 44916 362052 44980
rect 310100 44780 310164 44844
rect 141924 43964 141988 44028
rect 310100 42392 310164 42396
rect 310100 42336 310104 42392
rect 310104 42336 310160 42392
rect 310160 42336 310164 42392
rect 310100 42332 310164 42336
rect 518572 42392 518636 42396
rect 518572 42336 518622 42392
rect 518622 42336 518636 42392
rect 518572 42332 518636 42336
rect 187556 42120 187620 42124
rect 187556 42064 187570 42120
rect 187570 42064 187620 42120
rect 187556 42060 187620 42064
rect 361988 42120 362052 42124
rect 361988 42064 362002 42120
rect 362002 42064 362052 42120
rect 361988 42060 362052 42064
rect 365116 42120 365180 42124
rect 365116 42064 365130 42120
rect 365130 42064 365180 42120
rect 365116 42060 365180 42064
rect 460612 42120 460676 42124
rect 460612 42064 460626 42120
rect 460626 42064 460676 42120
rect 460612 42060 460676 42064
rect 471652 42120 471716 42124
rect 471652 42064 471666 42120
rect 471666 42064 471716 42120
rect 471652 42060 471716 42064
rect 514708 42060 514772 42124
rect 520228 42060 520292 42124
rect 521700 42120 521764 42124
rect 521700 42064 521750 42120
rect 521750 42064 521764 42120
rect 521700 42060 521764 42064
rect 529796 42060 529860 42124
rect 141924 40292 141988 40356
<< metal4 >>
rect 246435 997388 246501 997389
rect 246435 997338 246436 997388
rect 246500 997338 246501 997388
rect 238523 997252 238589 997253
rect 238523 997188 238524 997252
rect 238588 997188 238589 997252
rect 238523 997187 238589 997188
rect 86539 996572 86605 996573
rect 86539 996508 86540 996572
rect 86604 996508 86605 996572
rect 86539 996507 86605 996508
rect 86542 995757 86602 996507
rect 89667 996436 89733 996437
rect 89667 996372 89668 996436
rect 89732 996372 89733 996436
rect 89667 996371 89733 996372
rect 89670 995757 89730 996371
rect 135299 996300 135365 996301
rect 135299 996236 135300 996300
rect 135364 996236 135365 996300
rect 135299 996235 135365 996236
rect 135302 995757 135362 996235
rect 238526 995757 238586 997187
rect 480667 997252 480733 997253
rect 480667 997188 480668 997252
rect 480732 997188 480733 997252
rect 480667 997187 480733 997188
rect 240366 995757 240426 997102
rect 480670 995757 480730 997187
rect 532003 997252 532069 997253
rect 532003 997188 532004 997252
rect 532068 997188 532069 997252
rect 532003 997187 532069 997188
rect 485638 995757 485698 997102
rect 86539 995756 86605 995757
rect 86539 995692 86540 995756
rect 86604 995692 86605 995756
rect 86539 995691 86605 995692
rect 89667 995756 89733 995757
rect 89667 995692 89668 995756
rect 89732 995692 89733 995756
rect 89667 995691 89733 995692
rect 135299 995756 135365 995757
rect 135299 995692 135300 995756
rect 135364 995692 135365 995756
rect 135299 995691 135365 995692
rect 238523 995756 238589 995757
rect 238523 995692 238524 995756
rect 238588 995692 238589 995756
rect 238523 995691 238589 995692
rect 240363 995756 240429 995757
rect 240363 995692 240364 995756
rect 240428 995692 240429 995756
rect 240363 995691 240429 995692
rect 439819 995756 439885 995757
rect 439819 995692 439820 995756
rect 439884 995692 439885 995756
rect 439819 995691 439885 995692
rect 480667 995756 480733 995757
rect 480667 995692 480668 995756
rect 480732 995692 480733 995756
rect 480667 995691 480733 995692
rect 485635 995756 485701 995757
rect 485635 995692 485636 995756
rect 485700 995692 485701 995756
rect 485635 995691 485701 995692
rect 439822 991541 439882 995691
rect 505142 992357 505202 997102
rect 532006 995757 532066 997187
rect 536606 995757 536666 997102
rect 554638 995893 554698 997102
rect 627867 996708 627933 996709
rect 627867 996644 627868 996708
rect 627932 996644 627933 996708
rect 627867 996643 627933 996644
rect 554635 995892 554701 995893
rect 554635 995828 554636 995892
rect 554700 995828 554701 995892
rect 554635 995827 554701 995828
rect 627870 995757 627930 996643
rect 630259 996572 630325 996573
rect 630259 996508 630260 996572
rect 630324 996508 630325 996572
rect 630259 996507 630325 996508
rect 630262 995757 630322 996507
rect 532003 995756 532069 995757
rect 532003 995692 532004 995756
rect 532068 995692 532069 995756
rect 532003 995691 532069 995692
rect 536603 995756 536669 995757
rect 536603 995692 536604 995756
rect 536668 995692 536669 995756
rect 536603 995691 536669 995692
rect 573219 995756 573285 995757
rect 573219 995692 573220 995756
rect 573284 995692 573285 995756
rect 573219 995691 573285 995692
rect 627867 995756 627933 995757
rect 627867 995692 627868 995756
rect 627932 995692 627933 995756
rect 627867 995691 627933 995692
rect 630259 995756 630325 995757
rect 630259 995692 630260 995756
rect 630324 995692 630325 995756
rect 630259 995691 630325 995692
rect 505139 992356 505205 992357
rect 505139 992292 505140 992356
rect 505204 992292 505205 992356
rect 505139 992291 505205 992292
rect 439819 991540 439885 991541
rect 439819 991476 439820 991540
rect 439884 991476 439885 991540
rect 439819 991475 439885 991476
rect 573222 990997 573282 995691
rect 573219 990996 573285 990997
rect 573219 990932 573220 990996
rect 573284 990932 573285 990996
rect 573219 990931 573285 990932
rect 40539 968828 40605 968829
rect 40539 968764 40540 968828
rect 40604 968764 40605 968828
rect 40539 968763 40605 968764
rect 40355 963388 40421 963389
rect 40355 963324 40356 963388
rect 40420 963324 40421 963388
rect 40355 963323 40421 963324
rect 40358 936050 40418 963323
rect 40542 937410 40602 968763
rect 40723 967332 40789 967333
rect 40723 967268 40724 967332
rect 40788 967268 40789 967332
rect 40723 967267 40789 967268
rect 40726 938770 40786 967267
rect 676811 966516 676877 966517
rect 676811 966452 676812 966516
rect 676876 966452 676877 966516
rect 676811 966451 676877 966452
rect 676443 966244 676509 966245
rect 676443 966180 676444 966244
rect 676508 966180 676509 966244
rect 676443 966179 676509 966180
rect 42011 965156 42077 965157
rect 42011 965092 42012 965156
rect 42076 965092 42077 965156
rect 42011 965091 42077 965092
rect 41459 962164 41525 962165
rect 41459 962100 41460 962164
rect 41524 962100 41525 962164
rect 41459 962099 41525 962100
rect 41462 951693 41522 962099
rect 41643 958356 41709 958357
rect 41643 958292 41644 958356
rect 41708 958292 41709 958356
rect 41643 958291 41709 958292
rect 41646 952237 41706 958291
rect 41643 952236 41709 952237
rect 41643 952172 41644 952236
rect 41708 952172 41709 952236
rect 41643 952171 41709 952172
rect 42014 951693 42074 965091
rect 675339 963388 675405 963389
rect 675339 963324 675340 963388
rect 675404 963324 675405 963388
rect 675339 963323 675405 963324
rect 42195 957812 42261 957813
rect 42195 957748 42196 957812
rect 42260 957748 42261 957812
rect 42195 957747 42261 957748
rect 42198 951829 42258 957747
rect 42195 951828 42261 951829
rect 42195 951764 42196 951828
rect 42260 951764 42261 951828
rect 42195 951763 42261 951764
rect 41459 951692 41525 951693
rect 41459 951628 41460 951692
rect 41524 951628 41525 951692
rect 41459 951627 41525 951628
rect 42011 951692 42077 951693
rect 42011 951628 42012 951692
rect 42076 951628 42077 951692
rect 42011 951627 42077 951628
rect 675342 949789 675402 963323
rect 675891 961348 675957 961349
rect 675891 961284 675892 961348
rect 675956 961284 675957 961348
rect 675891 961283 675957 961284
rect 675707 959172 675773 959173
rect 675707 959108 675708 959172
rect 675772 959108 675773 959172
rect 675707 959107 675773 959108
rect 675523 957812 675589 957813
rect 675523 957748 675524 957812
rect 675588 957748 675589 957812
rect 675523 957747 675589 957748
rect 675339 949788 675405 949789
rect 675339 949724 675340 949788
rect 675404 949724 675405 949788
rect 675339 949723 675405 949724
rect 675526 949653 675586 957747
rect 675523 949652 675589 949653
rect 675523 949588 675524 949652
rect 675588 949588 675589 949652
rect 675523 949587 675589 949588
rect 675710 948837 675770 959107
rect 675894 949517 675954 961283
rect 676075 954004 676141 954005
rect 676075 953940 676076 954004
rect 676140 953940 676141 954004
rect 676075 953939 676141 953940
rect 675891 949516 675957 949517
rect 675891 949452 675892 949516
rect 675956 949452 675957 949516
rect 675891 949451 675957 949452
rect 675707 948836 675773 948837
rect 675707 948772 675708 948836
rect 675772 948772 675773 948836
rect 675707 948771 675773 948772
rect 676078 948021 676138 953939
rect 676446 951013 676506 966179
rect 676627 957676 676693 957677
rect 676627 957612 676628 957676
rect 676692 957612 676693 957676
rect 676627 957611 676693 957612
rect 676443 951012 676509 951013
rect 676443 950948 676444 951012
rect 676508 950948 676509 951012
rect 676443 950947 676509 950948
rect 676075 948020 676141 948021
rect 676075 947956 676076 948020
rect 676140 947956 676141 948020
rect 676075 947955 676141 947956
rect 40726 938710 41890 938770
rect 41830 938637 41890 938710
rect 41827 938636 41893 938637
rect 41827 938572 41828 938636
rect 41892 938572 41893 938636
rect 41827 938571 41893 938572
rect 40542 937350 41890 937410
rect 41830 937005 41890 937350
rect 41827 937004 41893 937005
rect 41827 936940 41828 937004
rect 41892 936940 41893 937004
rect 41827 936939 41893 936940
rect 40358 935990 41890 936050
rect 41830 934965 41890 935990
rect 41827 934964 41893 934965
rect 41827 934900 41828 934964
rect 41892 934900 41893 934964
rect 41827 934899 41893 934900
rect 676630 932381 676690 957611
rect 676814 950877 676874 966451
rect 677179 965020 677245 965021
rect 677179 964956 677180 965020
rect 677244 964956 677245 965020
rect 677179 964955 677245 964956
rect 676995 959036 677061 959037
rect 676995 958972 676996 959036
rect 677060 958972 677061 959036
rect 676995 958971 677061 958972
rect 676811 950876 676877 950877
rect 676811 950812 676812 950876
rect 676876 950812 676877 950876
rect 676811 950811 676877 950812
rect 676998 932789 677058 958971
rect 677182 935645 677242 964955
rect 677179 935644 677245 935645
rect 677179 935580 677180 935644
rect 677244 935580 677245 935644
rect 677179 935579 677245 935580
rect 676995 932788 677061 932789
rect 676995 932724 676996 932788
rect 677060 932724 677061 932788
rect 676995 932723 677061 932724
rect 676627 932380 676693 932381
rect 676627 932316 676628 932380
rect 676692 932316 676693 932380
rect 676627 932315 676693 932316
rect 676627 876620 676693 876621
rect 676627 876556 676628 876620
rect 676692 876556 676693 876620
rect 676627 876555 676693 876556
rect 676075 874172 676141 874173
rect 676075 874108 676076 874172
rect 676140 874108 676141 874172
rect 676075 874107 676141 874108
rect 673867 872268 673933 872269
rect 673867 872204 673868 872268
rect 673932 872204 673933 872268
rect 673867 872203 673933 872204
rect 41827 816100 41893 816101
rect 41827 816036 41828 816100
rect 41892 816036 41893 816100
rect 41827 816035 41893 816036
rect 41689 814332 41755 814333
rect 41689 814330 41690 814332
rect 39990 814270 41690 814330
rect 39990 771901 40050 814270
rect 41689 814268 41690 814270
rect 41754 814268 41755 814332
rect 41689 814267 41755 814268
rect 41830 813650 41890 816035
rect 40174 813590 41890 813650
rect 40174 773533 40234 813590
rect 41827 813244 41893 813245
rect 41827 813180 41828 813244
rect 41892 813180 41893 813244
rect 41827 813179 41893 813180
rect 40539 804812 40605 804813
rect 40539 804748 40540 804812
rect 40604 804748 40605 804812
rect 40539 804747 40605 804748
rect 40542 796789 40602 804747
rect 41830 804570 41890 813179
rect 41462 804510 41890 804570
rect 40539 796788 40605 796789
rect 40539 796724 40540 796788
rect 40604 796724 40605 796788
rect 40539 796723 40605 796724
rect 41462 786997 41522 804510
rect 42195 802772 42261 802773
rect 42195 802708 42196 802772
rect 42260 802708 42261 802772
rect 42195 802707 42261 802708
rect 41643 802636 41709 802637
rect 41643 802572 41644 802636
rect 41708 802572 41709 802636
rect 41643 802571 41709 802572
rect 41646 788085 41706 802571
rect 42011 802500 42077 802501
rect 42011 802436 42012 802500
rect 42076 802436 42077 802500
rect 42011 802435 42077 802436
rect 41827 801004 41893 801005
rect 41827 800940 41828 801004
rect 41892 800940 41893 801004
rect 41827 800939 41893 800940
rect 41830 788221 41890 800939
rect 42014 792029 42074 802435
rect 42011 792028 42077 792029
rect 42011 791964 42012 792028
rect 42076 791964 42077 792028
rect 42011 791963 42077 791964
rect 42198 788765 42258 802707
rect 42195 788764 42261 788765
rect 42195 788700 42196 788764
rect 42260 788700 42261 788764
rect 42195 788699 42261 788700
rect 41827 788220 41893 788221
rect 41827 788156 41828 788220
rect 41892 788156 41893 788220
rect 41827 788155 41893 788156
rect 41643 788084 41709 788085
rect 41643 788020 41644 788084
rect 41708 788020 41709 788084
rect 41643 788019 41709 788020
rect 41459 786996 41525 786997
rect 41459 786932 41460 786996
rect 41524 786932 41525 786996
rect 41459 786931 41525 786932
rect 40171 773532 40237 773533
rect 40171 773468 40172 773532
rect 40236 773468 40237 773532
rect 40171 773467 40237 773468
rect 39987 771900 40053 771901
rect 39987 771836 39988 771900
rect 40052 771836 40053 771900
rect 39987 771835 40053 771836
rect 39987 771084 40053 771085
rect 39987 771020 39988 771084
rect 40052 771020 40053 771084
rect 39987 771019 40053 771020
rect 39990 728653 40050 771019
rect 40907 766188 40973 766189
rect 40907 766124 40908 766188
rect 40972 766124 40973 766188
rect 40907 766123 40973 766124
rect 40539 764964 40605 764965
rect 40539 764900 40540 764964
rect 40604 764900 40605 764964
rect 40539 764899 40605 764900
rect 40542 750413 40602 764899
rect 40723 764556 40789 764557
rect 40723 764492 40724 764556
rect 40788 764492 40789 764556
rect 40723 764491 40789 764492
rect 40726 754221 40786 764491
rect 40723 754220 40789 754221
rect 40723 754156 40724 754220
rect 40788 754156 40789 754220
rect 40723 754155 40789 754156
rect 40910 753133 40970 766123
rect 41643 758300 41709 758301
rect 41643 758236 41644 758300
rect 41708 758236 41709 758300
rect 41643 758235 41709 758236
rect 41459 757756 41525 757757
rect 41459 757692 41460 757756
rect 41524 757692 41525 757756
rect 41459 757691 41525 757692
rect 40907 753132 40973 753133
rect 40907 753068 40908 753132
rect 40972 753068 40973 753132
rect 40907 753067 40973 753068
rect 40539 750412 40605 750413
rect 40539 750348 40540 750412
rect 40604 750348 40605 750412
rect 40539 750347 40605 750348
rect 41462 742389 41522 757691
rect 41646 746605 41706 758235
rect 41827 757076 41893 757077
rect 41827 757012 41828 757076
rect 41892 757012 41893 757076
rect 41827 757011 41893 757012
rect 42379 757076 42445 757077
rect 42379 757012 42380 757076
rect 42444 757012 42445 757076
rect 42379 757011 42445 757012
rect 41830 754901 41890 757011
rect 41827 754900 41893 754901
rect 41827 754836 41828 754900
rect 41892 754836 41893 754900
rect 41827 754835 41893 754836
rect 42382 749325 42442 757011
rect 673870 752589 673930 872203
rect 675891 864788 675957 864789
rect 675891 864724 675892 864788
rect 675956 864724 675957 864788
rect 675891 864723 675957 864724
rect 675339 788084 675405 788085
rect 675339 788020 675340 788084
rect 675404 788020 675405 788084
rect 675339 788019 675405 788020
rect 675342 773941 675402 788019
rect 675707 786724 675773 786725
rect 675707 786660 675708 786724
rect 675772 786660 675773 786724
rect 675707 786659 675773 786660
rect 675523 784820 675589 784821
rect 675523 784756 675524 784820
rect 675588 784756 675589 784820
rect 675523 784755 675589 784756
rect 675339 773940 675405 773941
rect 675339 773876 675340 773940
rect 675404 773876 675405 773940
rect 675339 773875 675405 773876
rect 675526 773397 675586 784755
rect 675710 773397 675770 786659
rect 675894 774893 675954 864723
rect 675891 774892 675957 774893
rect 675891 774828 675892 774892
rect 675956 774828 675957 774892
rect 675891 774827 675957 774828
rect 675523 773396 675589 773397
rect 675523 773332 675524 773396
rect 675588 773332 675589 773396
rect 675523 773331 675589 773332
rect 675707 773396 675773 773397
rect 675707 773332 675708 773396
rect 675772 773332 675773 773396
rect 675707 773331 675773 773332
rect 676078 772717 676138 874107
rect 676630 772989 676690 876555
rect 676811 876484 676877 876485
rect 676811 876420 676812 876484
rect 676876 876420 676877 876484
rect 676811 876419 676877 876420
rect 676814 773125 676874 876419
rect 677179 872812 677245 872813
rect 677179 872748 677180 872812
rect 677244 872748 677245 872812
rect 677179 872747 677245 872748
rect 677182 866670 677242 872747
rect 677182 866610 677426 866670
rect 676995 784140 677061 784141
rect 676995 784076 676996 784140
rect 677060 784076 677061 784140
rect 676995 784075 677061 784076
rect 676811 773124 676877 773125
rect 676811 773060 676812 773124
rect 676876 773060 676877 773124
rect 676811 773059 676877 773060
rect 676627 772988 676693 772989
rect 676627 772924 676628 772988
rect 676692 772924 676693 772988
rect 676627 772923 676693 772924
rect 676075 772716 676141 772717
rect 676075 772652 676076 772716
rect 676140 772652 676141 772716
rect 676075 772651 676141 772652
rect 675155 766596 675221 766597
rect 675155 766532 675156 766596
rect 675220 766532 675221 766596
rect 675155 766531 675221 766532
rect 676075 766596 676141 766597
rect 676075 766532 676076 766596
rect 676140 766532 676141 766596
rect 676075 766531 676141 766532
rect 674971 765100 675037 765101
rect 674971 765036 674972 765100
rect 675036 765036 675037 765100
rect 674971 765035 675037 765036
rect 674787 759116 674853 759117
rect 674787 759052 674788 759116
rect 674852 759052 674853 759116
rect 674787 759051 674853 759052
rect 674790 757893 674850 759051
rect 674787 757892 674853 757893
rect 674787 757828 674788 757892
rect 674852 757828 674853 757892
rect 674787 757827 674853 757828
rect 673867 752588 673933 752589
rect 673867 752524 673868 752588
rect 673932 752524 673933 752588
rect 673867 752523 673933 752524
rect 42379 749324 42445 749325
rect 42379 749260 42380 749324
rect 42444 749260 42445 749324
rect 42379 749259 42445 749260
rect 41643 746604 41709 746605
rect 41643 746540 41644 746604
rect 41708 746540 41709 746604
rect 41643 746539 41709 746540
rect 41459 742388 41525 742389
rect 41459 742324 41460 742388
rect 41524 742324 41525 742388
rect 41459 742323 41525 742324
rect 40355 729468 40421 729469
rect 40355 729404 40356 729468
rect 40420 729404 40421 729468
rect 40355 729403 40421 729404
rect 39987 728652 40053 728653
rect 39987 728588 39988 728652
rect 40052 728588 40053 728652
rect 39987 728587 40053 728588
rect 40171 727836 40237 727837
rect 40171 727772 40172 727836
rect 40236 727772 40237 727836
rect 40171 727771 40237 727772
rect 40174 685541 40234 727771
rect 40358 687173 40418 729403
rect 674974 727293 675034 765035
rect 674971 727292 675037 727293
rect 674971 727228 674972 727292
rect 675036 727228 675037 727292
rect 674971 727227 675037 727228
rect 675158 726613 675218 766531
rect 675707 741708 675773 741709
rect 675707 741644 675708 741708
rect 675772 741644 675773 741708
rect 675707 741643 675773 741644
rect 675523 736132 675589 736133
rect 675523 736068 675524 736132
rect 675588 736068 675589 736132
rect 675523 736067 675589 736068
rect 675526 728381 675586 736067
rect 675710 728381 675770 741643
rect 675523 728380 675589 728381
rect 675523 728316 675524 728380
rect 675588 728316 675589 728380
rect 675523 728315 675589 728316
rect 675707 728380 675773 728381
rect 675707 728316 675708 728380
rect 675772 728316 675773 728380
rect 675707 728315 675773 728316
rect 675155 726612 675221 726613
rect 675155 726548 675156 726612
rect 675220 726548 675221 726612
rect 675155 726547 675221 726548
rect 41459 725388 41525 725389
rect 41459 725324 41460 725388
rect 41524 725324 41525 725388
rect 41459 725323 41525 725324
rect 40539 721308 40605 721309
rect 40539 721244 40540 721308
rect 40604 721244 40605 721308
rect 40539 721243 40605 721244
rect 40542 710837 40602 721243
rect 40539 710836 40605 710837
rect 40539 710772 40540 710836
rect 40604 710772 40605 710836
rect 40539 710771 40605 710772
rect 41462 702405 41522 725323
rect 676078 724437 676138 766531
rect 676627 734364 676693 734365
rect 676627 734300 676628 734364
rect 676692 734300 676693 734364
rect 676627 734299 676693 734300
rect 676075 724436 676141 724437
rect 676075 724372 676076 724436
rect 676140 724372 676141 724436
rect 676075 724371 676141 724372
rect 676630 723252 676690 734299
rect 676630 723182 676710 723252
rect 675891 721560 675957 721561
rect 675891 721496 675892 721560
rect 675956 721496 675957 721560
rect 675891 721495 675957 721496
rect 676075 721560 676141 721561
rect 676075 721496 676076 721560
rect 676140 721496 676141 721560
rect 676650 721528 676710 723182
rect 676075 721495 676141 721496
rect 41643 716140 41709 716141
rect 41643 716076 41644 716140
rect 41708 716076 41709 716140
rect 41643 716075 41709 716076
rect 41459 702404 41525 702405
rect 41459 702340 41460 702404
rect 41524 702340 41525 702404
rect 41459 702339 41525 702340
rect 41646 699413 41706 716075
rect 41827 715460 41893 715461
rect 41827 715396 41828 715460
rect 41892 715396 41893 715460
rect 41827 715395 41893 715396
rect 41830 703765 41890 715395
rect 42011 713828 42077 713829
rect 42011 713764 42012 713828
rect 42076 713764 42077 713828
rect 42011 713763 42077 713764
rect 42014 706757 42074 713763
rect 42195 713284 42261 713285
rect 42195 713220 42196 713284
rect 42260 713220 42261 713284
rect 42195 713219 42261 713220
rect 42198 708525 42258 713219
rect 42195 708524 42261 708525
rect 42195 708460 42196 708524
rect 42260 708460 42261 708524
rect 42195 708459 42261 708460
rect 42011 706756 42077 706757
rect 42011 706692 42012 706756
rect 42076 706692 42077 706756
rect 42011 706691 42077 706692
rect 41827 703764 41893 703765
rect 41827 703700 41828 703764
rect 41892 703700 41893 703764
rect 41827 703699 41893 703700
rect 41643 699412 41709 699413
rect 41643 699348 41644 699412
rect 41708 699348 41709 699412
rect 41643 699347 41709 699348
rect 675339 696964 675405 696965
rect 675339 696900 675340 696964
rect 675404 696900 675405 696964
rect 675339 696899 675405 696900
rect 40355 687172 40421 687173
rect 40355 687108 40356 687172
rect 40420 687108 40421 687172
rect 40355 687107 40421 687108
rect 40171 685540 40237 685541
rect 40171 685476 40172 685540
rect 40236 685476 40237 685540
rect 40171 685475 40237 685476
rect 39987 684724 40053 684725
rect 39987 684660 39988 684724
rect 40052 684660 40053 684724
rect 39987 684659 40053 684660
rect 30603 677788 30669 677789
rect 30603 677724 30604 677788
rect 30668 677724 30669 677788
rect 30603 677723 30669 677724
rect 30606 676565 30666 677723
rect 30603 676564 30669 676565
rect 30603 676500 30604 676564
rect 30668 676500 30669 676564
rect 30603 676499 30669 676500
rect 39990 642293 40050 684659
rect 675342 683365 675402 696899
rect 675523 694788 675589 694789
rect 675523 694724 675524 694788
rect 675588 694724 675589 694788
rect 675523 694723 675589 694724
rect 675526 683365 675586 694723
rect 675707 686220 675773 686221
rect 675707 686156 675708 686220
rect 675772 686156 675773 686220
rect 675707 686155 675773 686156
rect 675339 683364 675405 683365
rect 675339 683300 675340 683364
rect 675404 683300 675405 683364
rect 675339 683299 675405 683300
rect 675523 683364 675589 683365
rect 675523 683300 675524 683364
rect 675588 683300 675589 683364
rect 675523 683299 675589 683300
rect 675710 683229 675770 686155
rect 675707 683228 675773 683229
rect 675707 683164 675708 683228
rect 675772 683164 675773 683228
rect 675707 683163 675773 683164
rect 41459 682276 41525 682277
rect 41459 682212 41460 682276
rect 41524 682212 41525 682276
rect 41459 682211 41525 682212
rect 40539 679420 40605 679421
rect 40539 679356 40540 679420
rect 40604 679356 40605 679420
rect 40539 679355 40605 679356
rect 40542 664597 40602 679355
rect 40723 678196 40789 678197
rect 40723 678132 40724 678196
rect 40788 678132 40789 678196
rect 40723 678131 40789 678132
rect 40726 665413 40786 678131
rect 40723 665412 40789 665413
rect 40723 665348 40724 665412
rect 40788 665348 40789 665412
rect 40723 665347 40789 665348
rect 40539 664596 40605 664597
rect 40539 664532 40540 664596
rect 40604 664532 40605 664596
rect 40539 664531 40605 664532
rect 41462 661333 41522 682211
rect 675894 681869 675954 721495
rect 675891 681868 675957 681869
rect 675891 681804 675892 681868
rect 675956 681804 675957 681868
rect 675891 681803 675957 681804
rect 676078 678333 676138 721495
rect 676630 721462 676710 721528
rect 676443 694244 676509 694245
rect 676443 694180 676444 694244
rect 676508 694180 676509 694244
rect 676443 694179 676509 694180
rect 676446 683229 676506 694179
rect 676443 683228 676509 683229
rect 676443 683164 676444 683228
rect 676508 683164 676509 683228
rect 676443 683163 676509 683164
rect 676075 678332 676141 678333
rect 676075 678268 676076 678332
rect 676140 678268 676141 678332
rect 676075 678267 676141 678268
rect 676630 677964 676690 721462
rect 676998 713493 677058 784075
rect 677179 774892 677245 774893
rect 677179 774828 677180 774892
rect 677244 774828 677245 774892
rect 677179 774827 677245 774828
rect 677182 756805 677242 774827
rect 677179 756804 677245 756805
rect 677179 756740 677180 756804
rect 677244 756740 677245 756804
rect 677179 756739 677245 756740
rect 677366 753949 677426 866610
rect 677363 753948 677429 753949
rect 677363 753884 677364 753948
rect 677428 753884 677429 753948
rect 677363 753883 677429 753884
rect 677179 733004 677245 733005
rect 677179 732940 677180 733004
rect 677244 732940 677245 733004
rect 677179 732939 677245 732940
rect 676995 713492 677061 713493
rect 676995 713428 676996 713492
rect 677060 713428 677061 713492
rect 676995 713427 677061 713428
rect 676811 687444 676877 687445
rect 676811 687380 676812 687444
rect 676876 687380 676877 687444
rect 676811 687379 676877 687380
rect 676630 677892 676698 677964
rect 676638 676444 676698 677892
rect 675155 676428 675221 676429
rect 675155 676364 675156 676428
rect 675220 676364 675221 676428
rect 675155 676363 675221 676364
rect 675891 676428 675957 676429
rect 675891 676364 675892 676428
rect 675956 676364 675957 676428
rect 675891 676363 675957 676364
rect 676630 676376 676698 676444
rect 41643 671396 41709 671397
rect 41643 671332 41644 671396
rect 41708 671332 41709 671396
rect 41643 671331 41709 671332
rect 41459 661332 41525 661333
rect 41459 661268 41460 661332
rect 41524 661268 41525 661332
rect 41459 661267 41525 661268
rect 41646 658341 41706 671331
rect 42379 670988 42445 670989
rect 42379 670924 42380 670988
rect 42444 670924 42445 670988
rect 42379 670923 42445 670924
rect 41827 670716 41893 670717
rect 41827 670652 41828 670716
rect 41892 670652 41893 670716
rect 41827 670651 41893 670652
rect 42011 670716 42077 670717
rect 42011 670652 42012 670716
rect 42076 670652 42077 670716
rect 42011 670651 42077 670652
rect 41830 668541 41890 670651
rect 41827 668540 41893 668541
rect 41827 668476 41828 668540
rect 41892 668476 41893 668540
rect 41827 668475 41893 668476
rect 41827 668404 41893 668405
rect 41827 668340 41828 668404
rect 41892 668340 41893 668404
rect 41827 668339 41893 668340
rect 41830 660381 41890 668339
rect 42014 663373 42074 670651
rect 42195 670172 42261 670173
rect 42195 670108 42196 670172
rect 42260 670108 42261 670172
rect 42195 670107 42261 670108
rect 42011 663372 42077 663373
rect 42011 663308 42012 663372
rect 42076 663308 42077 663372
rect 42011 663307 42077 663308
rect 42198 660517 42258 670107
rect 42382 668405 42442 670923
rect 672947 669084 673013 669085
rect 672947 669020 672948 669084
rect 673012 669020 673013 669084
rect 672947 669019 673013 669020
rect 42379 668404 42445 668405
rect 42379 668340 42380 668404
rect 42444 668340 42445 668404
rect 42379 668339 42445 668340
rect 42195 660516 42261 660517
rect 42195 660452 42196 660516
rect 42260 660452 42261 660516
rect 42195 660451 42261 660452
rect 41827 660380 41893 660381
rect 41827 660316 41828 660380
rect 41892 660316 41893 660380
rect 41827 660315 41893 660316
rect 41643 658340 41709 658341
rect 41643 658276 41644 658340
rect 41708 658276 41709 658340
rect 41643 658275 41709 658276
rect 39987 642292 40053 642293
rect 39987 642228 39988 642292
rect 40052 642228 40053 642292
rect 39987 642227 40053 642228
rect 39987 641476 40053 641477
rect 39987 641412 39988 641476
rect 40052 641412 40053 641476
rect 39987 641411 40053 641412
rect 39990 599045 40050 641411
rect 41459 639436 41525 639437
rect 41459 639372 41460 639436
rect 41524 639372 41525 639436
rect 41459 639371 41525 639372
rect 40907 636580 40973 636581
rect 40907 636516 40908 636580
rect 40972 636516 40973 636580
rect 40907 636515 40973 636516
rect 40539 636172 40605 636173
rect 40539 636108 40540 636172
rect 40604 636108 40605 636172
rect 40539 636107 40605 636108
rect 40542 621485 40602 636107
rect 40723 634948 40789 634949
rect 40723 634884 40724 634948
rect 40788 634884 40789 634948
rect 40723 634883 40789 634884
rect 40726 623797 40786 634883
rect 40910 625293 40970 636515
rect 40907 625292 40973 625293
rect 40907 625228 40908 625292
rect 40972 625228 40973 625292
rect 40907 625227 40973 625228
rect 40723 623796 40789 623797
rect 40723 623732 40724 623796
rect 40788 623732 40789 623796
rect 40723 623731 40789 623732
rect 40539 621484 40605 621485
rect 40539 621420 40540 621484
rect 40604 621420 40605 621484
rect 40539 621419 40605 621420
rect 41462 614141 41522 639371
rect 41643 629916 41709 629917
rect 41643 629852 41644 629916
rect 41708 629852 41709 629916
rect 41643 629851 41709 629852
rect 41459 614140 41525 614141
rect 41459 614076 41460 614140
rect 41524 614076 41525 614140
rect 41459 614075 41525 614076
rect 41646 613461 41706 629851
rect 42195 629236 42261 629237
rect 42195 629172 42196 629236
rect 42260 629172 42261 629236
rect 42195 629171 42261 629172
rect 42011 629100 42077 629101
rect 42011 629036 42012 629100
rect 42076 629036 42077 629100
rect 42011 629035 42077 629036
rect 41827 628556 41893 628557
rect 41827 628492 41828 628556
rect 41892 628492 41893 628556
rect 41827 628491 41893 628492
rect 41830 616861 41890 628491
rect 42014 619037 42074 629035
rect 42011 619036 42077 619037
rect 42011 618972 42012 619036
rect 42076 618972 42077 619036
rect 42011 618971 42077 618972
rect 41827 616860 41893 616861
rect 41827 616796 41828 616860
rect 41892 616796 41893 616860
rect 41827 616795 41893 616796
rect 42198 616725 42258 629171
rect 42195 616724 42261 616725
rect 42195 616660 42196 616724
rect 42260 616660 42261 616724
rect 42195 616659 42261 616660
rect 41643 613460 41709 613461
rect 41643 613396 41644 613460
rect 41708 613396 41709 613460
rect 41643 613395 41709 613396
rect 39987 599044 40053 599045
rect 39987 598980 39988 599044
rect 40052 598980 40053 599044
rect 39987 598979 40053 598980
rect 39987 598228 40053 598229
rect 39987 598164 39988 598228
rect 40052 598164 40053 598228
rect 39987 598163 40053 598164
rect 39990 555933 40050 598163
rect 40539 592108 40605 592109
rect 40539 592044 40540 592108
rect 40604 592044 40605 592108
rect 40539 592043 40605 592044
rect 40542 577557 40602 592043
rect 40723 591700 40789 591701
rect 40723 591636 40724 591700
rect 40788 591636 40789 591700
rect 40723 591635 40789 591636
rect 40726 579053 40786 591635
rect 41459 587212 41525 587213
rect 41459 587148 41460 587212
rect 41524 587148 41525 587212
rect 41459 587147 41525 587148
rect 40907 585444 40973 585445
rect 40907 585380 40908 585444
rect 40972 585380 40973 585444
rect 40907 585379 40973 585380
rect 40910 581773 40970 585379
rect 40907 581772 40973 581773
rect 40907 581708 40908 581772
rect 40972 581708 40973 581772
rect 40907 581707 40973 581708
rect 40723 579052 40789 579053
rect 40723 578988 40724 579052
rect 40788 578988 40789 579052
rect 40723 578987 40789 578988
rect 40539 577556 40605 577557
rect 40539 577492 40540 577556
rect 40604 577492 40605 577556
rect 40539 577491 40605 577492
rect 41462 570485 41522 587147
rect 42379 585172 42445 585173
rect 42379 585108 42380 585172
rect 42444 585108 42445 585172
rect 42379 585107 42445 585108
rect 42011 584648 42077 584649
rect 42011 584584 42012 584648
rect 42076 584584 42077 584648
rect 42011 584583 42077 584584
rect 41643 584512 41709 584513
rect 41643 584448 41644 584512
rect 41708 584448 41709 584512
rect 41643 584447 41709 584448
rect 41646 580277 41706 584447
rect 41643 580276 41709 580277
rect 41643 580212 41644 580276
rect 41708 580212 41709 580276
rect 41643 580211 41709 580212
rect 42014 571573 42074 584583
rect 42382 574021 42442 585107
rect 42563 584220 42629 584221
rect 42563 584156 42564 584220
rect 42628 584156 42629 584220
rect 42563 584155 42629 584156
rect 42379 574020 42445 574021
rect 42379 573956 42380 574020
rect 42444 573956 42445 574020
rect 42379 573955 42445 573956
rect 42566 573885 42626 584155
rect 42563 573884 42629 573885
rect 42563 573820 42564 573884
rect 42628 573820 42629 573884
rect 42563 573819 42629 573820
rect 42011 571572 42077 571573
rect 42011 571508 42012 571572
rect 42076 571508 42077 571572
rect 42011 571507 42077 571508
rect 41459 570484 41525 570485
rect 41459 570420 41460 570484
rect 41524 570420 41525 570484
rect 41459 570419 41525 570420
rect 39987 555932 40053 555933
rect 39987 555868 39988 555932
rect 40052 555868 40053 555932
rect 39987 555867 40053 555868
rect 40723 550628 40789 550629
rect 40723 550564 40724 550628
rect 40788 550564 40789 550628
rect 40723 550563 40789 550564
rect 40539 549404 40605 549405
rect 40539 549340 40540 549404
rect 40604 549340 40605 549404
rect 40539 549339 40605 549340
rect 40542 531453 40602 549339
rect 40726 534173 40786 550563
rect 40907 548996 40973 548997
rect 40907 548932 40908 548996
rect 40972 548932 40973 548996
rect 40907 548931 40973 548932
rect 40910 534581 40970 548931
rect 41459 545188 41525 545189
rect 41459 545124 41460 545188
rect 41524 545124 41525 545188
rect 41459 545123 41525 545124
rect 40907 534580 40973 534581
rect 40907 534516 40908 534580
rect 40972 534516 40973 534580
rect 40907 534515 40973 534516
rect 40723 534172 40789 534173
rect 40723 534108 40724 534172
rect 40788 534108 40789 534172
rect 40723 534107 40789 534108
rect 40539 531452 40605 531453
rect 40539 531388 40540 531452
rect 40604 531388 40605 531452
rect 40539 531387 40605 531388
rect 41462 529957 41522 545123
rect 41643 543012 41709 543013
rect 41643 542948 41644 543012
rect 41708 542948 41709 543012
rect 41643 542947 41709 542948
rect 41459 529956 41525 529957
rect 41459 529892 41460 529956
rect 41524 529892 41525 529956
rect 41459 529891 41525 529892
rect 41646 529413 41706 542947
rect 41827 542876 41893 542877
rect 41827 542812 41828 542876
rect 41892 542812 41893 542876
rect 41827 542811 41893 542812
rect 41830 532677 41890 542811
rect 42011 542332 42077 542333
rect 42011 542268 42012 542332
rect 42076 542268 42077 542332
rect 42011 542267 42077 542268
rect 42014 535941 42074 542267
rect 42011 535940 42077 535941
rect 42011 535876 42012 535940
rect 42076 535876 42077 535940
rect 42011 535875 42077 535876
rect 41827 532676 41893 532677
rect 41827 532612 41828 532676
rect 41892 532612 41893 532676
rect 41827 532611 41893 532612
rect 41643 529412 41709 529413
rect 41643 529348 41644 529412
rect 41708 529348 41709 529412
rect 41643 529347 41709 529348
rect 672950 474877 673010 669019
rect 675158 637397 675218 676363
rect 675339 649908 675405 649909
rect 675339 649844 675340 649908
rect 675404 649844 675405 649908
rect 675339 649843 675405 649844
rect 675342 638757 675402 649843
rect 675523 645964 675589 645965
rect 675523 645900 675524 645964
rect 675588 645900 675589 645964
rect 675523 645899 675589 645900
rect 675339 638756 675405 638757
rect 675339 638692 675340 638756
rect 675404 638692 675405 638756
rect 675339 638691 675405 638692
rect 675526 638213 675586 645899
rect 675523 638212 675589 638213
rect 675523 638148 675524 638212
rect 675588 638148 675589 638212
rect 675523 638147 675589 638148
rect 675894 637533 675954 676363
rect 676630 662965 676690 676376
rect 676627 662964 676693 662965
rect 676627 662900 676628 662964
rect 676692 662900 676693 662964
rect 676627 662899 676693 662900
rect 676627 648684 676693 648685
rect 676627 648620 676628 648684
rect 676692 648620 676693 648684
rect 676627 648619 676693 648620
rect 676630 637941 676690 648619
rect 676627 637940 676693 637941
rect 676627 637876 676628 637940
rect 676692 637876 676693 637940
rect 676627 637875 676693 637876
rect 675891 637532 675957 637533
rect 675891 637468 675892 637532
rect 675956 637468 675957 637532
rect 675891 637467 675957 637468
rect 675155 637396 675221 637397
rect 675155 637332 675156 637396
rect 675220 637332 675221 637396
rect 675155 637331 675221 637332
rect 676075 631412 676141 631413
rect 676075 631348 676076 631412
rect 676140 631348 676141 631412
rect 676075 631347 676141 631348
rect 675339 606524 675405 606525
rect 675339 606460 675340 606524
rect 675404 606460 675405 606524
rect 675339 606459 675405 606460
rect 675342 592109 675402 606459
rect 675707 600948 675773 600949
rect 675707 600884 675708 600948
rect 675772 600884 675773 600948
rect 675707 600883 675773 600884
rect 675523 595372 675589 595373
rect 675523 595308 675524 595372
rect 675588 595308 675589 595372
rect 675523 595307 675589 595308
rect 675526 593061 675586 595307
rect 675710 593197 675770 600883
rect 675707 593196 675773 593197
rect 675707 593132 675708 593196
rect 675772 593132 675773 593196
rect 675707 593131 675773 593132
rect 675523 593060 675589 593061
rect 675523 592996 675524 593060
rect 675588 592996 675589 593060
rect 675523 592995 675589 592996
rect 675339 592108 675405 592109
rect 675339 592044 675340 592108
rect 675404 592044 675405 592108
rect 675339 592043 675405 592044
rect 676078 591429 676138 631347
rect 676814 618357 676874 687379
rect 676995 676428 677061 676429
rect 676995 676364 676996 676428
rect 677060 676364 677061 676428
rect 676995 676363 677061 676364
rect 676998 637941 677058 676363
rect 677182 663373 677242 732939
rect 677179 663372 677245 663373
rect 677179 663308 677180 663372
rect 677244 663308 677245 663372
rect 677179 663307 677245 663308
rect 677182 644950 677426 645010
rect 677182 644741 677242 644950
rect 677179 644740 677245 644741
rect 677179 644676 677180 644740
rect 677244 644676 677245 644740
rect 677179 644675 677245 644676
rect 677179 644604 677245 644605
rect 677179 644540 677180 644604
rect 677244 644540 677245 644604
rect 677179 644539 677245 644540
rect 676995 637940 677061 637941
rect 676995 637876 676996 637940
rect 677060 637876 677061 637940
rect 676995 637875 677061 637876
rect 676995 631412 677061 631413
rect 676995 631348 676996 631412
rect 677060 631348 677061 631412
rect 676995 631347 677061 631348
rect 676811 618356 676877 618357
rect 676811 618292 676812 618356
rect 676876 618292 676877 618356
rect 676811 618291 676877 618292
rect 676811 599044 676877 599045
rect 676811 598980 676812 599044
rect 676876 598980 676877 599044
rect 676811 598979 676877 598980
rect 676075 591428 676141 591429
rect 676075 591364 676076 591428
rect 676140 591364 676141 591428
rect 676075 591363 676141 591364
rect 675707 586260 675773 586261
rect 675707 586196 675708 586260
rect 675772 586196 675773 586260
rect 675707 586195 675773 586196
rect 676075 586260 676141 586261
rect 676075 586196 676076 586260
rect 676140 586196 676141 586260
rect 676075 586195 676141 586196
rect 675339 561236 675405 561237
rect 675339 561172 675340 561236
rect 675404 561172 675405 561236
rect 675339 561171 675405 561172
rect 675342 550357 675402 561171
rect 675523 559604 675589 559605
rect 675523 559540 675524 559604
rect 675588 559540 675589 559604
rect 675523 559539 675589 559540
rect 675526 554845 675586 559539
rect 675523 554844 675589 554845
rect 675523 554780 675524 554844
rect 675588 554780 675589 554844
rect 675523 554779 675589 554780
rect 675339 550356 675405 550357
rect 675339 550292 675340 550356
rect 675404 550292 675405 550356
rect 675339 550291 675405 550292
rect 675710 546821 675770 586195
rect 675891 584628 675957 584629
rect 675891 584564 675892 584628
rect 675956 584564 675957 584628
rect 675891 584563 675957 584564
rect 675707 546820 675773 546821
rect 675707 546756 675708 546820
rect 675772 546756 675773 546820
rect 675707 546755 675773 546756
rect 675894 546685 675954 584563
rect 675891 546684 675957 546685
rect 675891 546620 675892 546684
rect 675956 546620 675957 546684
rect 675891 546619 675957 546620
rect 676078 543013 676138 586195
rect 676627 562732 676693 562733
rect 676627 562668 676628 562732
rect 676692 562668 676693 562732
rect 676627 562667 676693 562668
rect 676630 546549 676690 562667
rect 676627 546548 676693 546549
rect 676627 546484 676628 546548
rect 676692 546484 676693 546548
rect 676627 546483 676693 546484
rect 676814 543693 676874 598979
rect 676998 592109 677058 631347
rect 676995 592108 677061 592109
rect 676995 592044 676996 592108
rect 677060 592044 677061 592108
rect 676995 592043 677061 592044
rect 677182 573205 677242 644539
rect 677179 573204 677245 573205
rect 677179 573140 677180 573204
rect 677244 573140 677245 573204
rect 677179 573139 677245 573140
rect 677366 572797 677426 644950
rect 677363 572796 677429 572797
rect 677363 572732 677364 572796
rect 677428 572732 677429 572796
rect 677363 572731 677429 572732
rect 677179 559060 677245 559061
rect 677179 558996 677180 559060
rect 677244 558996 677245 559060
rect 677179 558995 677245 558996
rect 677182 557550 677242 558995
rect 677182 557490 677426 557550
rect 677179 554028 677245 554029
rect 677179 553964 677180 554028
rect 677244 553964 677245 554028
rect 677179 553963 677245 553964
rect 676995 551988 677061 551989
rect 676995 551924 676996 551988
rect 677060 551924 677061 551988
rect 676995 551923 677061 551924
rect 676811 543692 676877 543693
rect 676811 543628 676812 543692
rect 676876 543628 676877 543692
rect 676811 543627 676877 543628
rect 676075 543012 676141 543013
rect 676075 542948 676076 543012
rect 676140 542948 676141 543012
rect 676075 542947 676141 542948
rect 676998 484530 677058 551923
rect 676078 484470 677058 484530
rect 676078 484125 676138 484470
rect 676075 484124 676141 484125
rect 676075 484060 676076 484124
rect 676140 484060 676141 484124
rect 676075 484059 676141 484060
rect 677182 483850 677242 553963
rect 677366 492421 677426 557490
rect 677363 492420 677429 492421
rect 677363 492356 677364 492420
rect 677428 492356 677429 492420
rect 677363 492355 677429 492356
rect 676078 483790 677242 483850
rect 676078 483717 676138 483790
rect 676075 483716 676141 483717
rect 676075 483652 676076 483716
rect 676140 483652 676141 483716
rect 676075 483651 676141 483652
rect 672947 474876 673013 474877
rect 672947 474812 672948 474876
rect 673012 474812 673013 474876
rect 672947 474811 673013 474812
rect 41827 426460 41893 426461
rect 41827 426396 41828 426460
rect 41892 426396 41893 426460
rect 41827 426395 41893 426396
rect 41830 426050 41890 426395
rect 40542 425990 41890 426050
rect 40054 420742 40120 420743
rect 40054 420678 40055 420742
rect 40119 420678 40120 420742
rect 40054 420677 40120 420678
rect 40058 419515 40118 420677
rect 40054 419514 40120 419515
rect 40054 419450 40055 419514
rect 40119 419450 40120 419514
rect 40054 419449 40120 419450
rect 40542 400077 40602 425990
rect 41827 425644 41893 425645
rect 41827 425580 41828 425644
rect 41892 425580 41893 425644
rect 41827 425579 41893 425580
rect 41830 425370 41890 425579
rect 40726 425310 41890 425370
rect 40539 400076 40605 400077
rect 40539 400012 40540 400076
rect 40604 400012 40605 400076
rect 40539 400011 40605 400012
rect 40726 398853 40786 425310
rect 42195 424828 42261 424829
rect 42195 424764 42196 424828
rect 42260 424764 42261 424828
rect 42195 424763 42261 424764
rect 41827 424012 41893 424013
rect 41827 424010 41828 424012
rect 40910 423950 41828 424010
rect 40910 399669 40970 423950
rect 41827 423948 41828 423950
rect 41892 423948 41893 424012
rect 41827 423947 41893 423948
rect 42011 423604 42077 423605
rect 42011 423540 42012 423604
rect 42076 423540 42077 423604
rect 42011 423539 42077 423540
rect 41827 422788 41893 422789
rect 41827 422724 41828 422788
rect 41892 422724 41893 422788
rect 41827 422723 41893 422724
rect 41830 422650 41890 422723
rect 41094 422590 41890 422650
rect 41094 409461 41154 422590
rect 42014 422310 42074 423539
rect 41830 422250 42074 422310
rect 41830 415309 41890 422250
rect 42198 418170 42258 424763
rect 42014 418110 42258 418170
rect 41827 415308 41893 415309
rect 41827 415244 41828 415308
rect 41892 415244 41893 415308
rect 41827 415243 41893 415244
rect 42014 415170 42074 418110
rect 41646 415110 42074 415170
rect 41459 414764 41525 414765
rect 41459 414700 41460 414764
rect 41524 414700 41525 414764
rect 41459 414699 41525 414700
rect 41091 409460 41157 409461
rect 41091 409396 41092 409460
rect 41156 409396 41157 409460
rect 41091 409395 41157 409396
rect 41462 401845 41522 414699
rect 41646 406333 41706 415110
rect 42011 415036 42077 415037
rect 42011 414972 42012 415036
rect 42076 414972 42077 415036
rect 42011 414971 42077 414972
rect 41827 414628 41893 414629
rect 41827 414564 41828 414628
rect 41892 414564 41893 414628
rect 41827 414563 41893 414564
rect 41830 411229 41890 414563
rect 41827 411228 41893 411229
rect 41827 411164 41828 411228
rect 41892 411164 41893 411228
rect 41827 411163 41893 411164
rect 41643 406332 41709 406333
rect 41643 406268 41644 406332
rect 41708 406268 41709 406332
rect 41643 406267 41709 406268
rect 42014 402525 42074 414971
rect 42011 402524 42077 402525
rect 42011 402460 42012 402524
rect 42076 402460 42077 402524
rect 42011 402459 42077 402460
rect 41459 401844 41525 401845
rect 41459 401780 41460 401844
rect 41524 401780 41525 401844
rect 41459 401779 41525 401780
rect 40907 399668 40973 399669
rect 40907 399604 40908 399668
rect 40972 399604 40973 399668
rect 40907 399603 40973 399604
rect 675891 399396 675957 399397
rect 675891 399332 675892 399396
rect 675956 399332 675957 399396
rect 675891 399331 675957 399332
rect 40723 398852 40789 398853
rect 40723 398788 40724 398852
rect 40788 398788 40789 398852
rect 40723 398787 40789 398788
rect 675523 388516 675589 388517
rect 675523 388452 675524 388516
rect 675588 388452 675589 388516
rect 675523 388451 675589 388452
rect 675339 387564 675405 387565
rect 675339 387500 675340 387564
rect 675404 387500 675405 387564
rect 675339 387499 675405 387500
rect 40723 383076 40789 383077
rect 40723 383012 40724 383076
rect 40788 383012 40789 383076
rect 40723 383011 40789 383012
rect 40539 382260 40605 382261
rect 40539 382196 40540 382260
rect 40604 382196 40605 382260
rect 40539 382195 40605 382196
rect 40542 355741 40602 382195
rect 40726 356965 40786 383011
rect 675342 382261 675402 387499
rect 675339 382260 675405 382261
rect 675339 382196 675340 382260
rect 675404 382196 675405 382260
rect 675339 382195 675405 382196
rect 41459 381852 41525 381853
rect 41459 381788 41460 381852
rect 41524 381788 41525 381852
rect 41459 381787 41525 381788
rect 40907 379812 40973 379813
rect 40907 379748 40908 379812
rect 40972 379748 40973 379812
rect 40907 379747 40973 379748
rect 40910 360229 40970 379747
rect 40907 360228 40973 360229
rect 40907 360164 40908 360228
rect 40972 360164 40973 360228
rect 40907 360163 40973 360164
rect 41462 358733 41522 381787
rect 675526 378725 675586 388451
rect 675707 387700 675773 387701
rect 675707 387636 675708 387700
rect 675772 387636 675773 387700
rect 675707 387635 675773 387636
rect 675523 378724 675589 378725
rect 675523 378660 675524 378724
rect 675588 378660 675589 378724
rect 675523 378659 675589 378660
rect 675710 375461 675770 387635
rect 675894 384981 675954 399331
rect 676259 398852 676325 398853
rect 676259 398788 676260 398852
rect 676324 398788 676325 398852
rect 676259 398787 676325 398788
rect 676075 395180 676141 395181
rect 676075 395116 676076 395180
rect 676140 395116 676141 395180
rect 676075 395115 676141 395116
rect 675891 384980 675957 384981
rect 675891 384916 675892 384980
rect 675956 384916 675957 384980
rect 675891 384915 675957 384916
rect 676078 377637 676138 395115
rect 676075 377636 676141 377637
rect 676075 377572 676076 377636
rect 676140 377572 676141 377636
rect 676075 377571 676141 377572
rect 675707 375460 675773 375461
rect 675707 375396 675708 375460
rect 675772 375396 675773 375460
rect 675707 375395 675773 375396
rect 676262 373693 676322 398787
rect 676443 397220 676509 397221
rect 676443 397156 676444 397220
rect 676508 397156 676509 397220
rect 676443 397155 676509 397156
rect 676259 373692 676325 373693
rect 676259 373628 676260 373692
rect 676324 373628 676325 373692
rect 676259 373627 676325 373628
rect 676446 372061 676506 397155
rect 676443 372060 676509 372061
rect 676443 371996 676444 372060
rect 676508 371996 676509 372060
rect 676443 371995 676509 371996
rect 42011 371924 42077 371925
rect 42011 371860 42012 371924
rect 42076 371860 42077 371924
rect 42011 371859 42077 371860
rect 41643 371380 41709 371381
rect 41643 371316 41644 371380
rect 41708 371316 41709 371380
rect 41643 371315 41709 371316
rect 41646 362949 41706 371315
rect 41827 370292 41893 370293
rect 41827 370228 41828 370292
rect 41892 370228 41893 370292
rect 41827 370227 41893 370228
rect 41830 366349 41890 370227
rect 41827 366348 41893 366349
rect 41827 366284 41828 366348
rect 41892 366284 41893 366348
rect 41827 366283 41893 366284
rect 42014 363765 42074 371859
rect 42011 363764 42077 363765
rect 42011 363700 42012 363764
rect 42076 363700 42077 363764
rect 42011 363699 42077 363700
rect 41643 362948 41709 362949
rect 41643 362884 41644 362948
rect 41708 362884 41709 362948
rect 41643 362883 41709 362884
rect 41459 358732 41525 358733
rect 41459 358668 41460 358732
rect 41524 358668 41525 358732
rect 41459 358667 41525 358668
rect 40723 356964 40789 356965
rect 40723 356900 40724 356964
rect 40788 356900 40789 356964
rect 40723 356899 40789 356900
rect 40539 355740 40605 355741
rect 40539 355676 40540 355740
rect 40604 355676 40605 355740
rect 40539 355675 40605 355676
rect 675523 354244 675589 354245
rect 675523 354180 675524 354244
rect 675588 354180 675589 354244
rect 675523 354179 675589 354180
rect 675339 353428 675405 353429
rect 675339 353364 675340 353428
rect 675404 353364 675405 353428
rect 675339 353363 675405 353364
rect 675342 345810 675402 353363
rect 675526 346490 675586 354179
rect 676078 353910 676506 353970
rect 676078 353701 676138 353910
rect 676075 353700 676141 353701
rect 676075 353636 676076 353700
rect 676140 353636 676141 353700
rect 676075 353635 676141 353636
rect 675891 353020 675957 353021
rect 675891 352956 675892 353020
rect 675956 352956 675957 353020
rect 675891 352955 675957 352956
rect 675894 350550 675954 352955
rect 676075 352068 676141 352069
rect 676075 352004 676076 352068
rect 676140 352004 676141 352068
rect 676075 352003 676141 352004
rect 676078 351930 676138 352003
rect 676078 351870 676322 351930
rect 675894 350490 676138 350550
rect 675526 346430 675954 346490
rect 675342 345750 675770 345810
rect 675523 343636 675589 343637
rect 675523 343572 675524 343636
rect 675588 343572 675589 343636
rect 675523 343571 675589 343572
rect 40723 339828 40789 339829
rect 40723 339764 40724 339828
rect 40788 339764 40789 339828
rect 40723 339763 40789 339764
rect 40539 339012 40605 339013
rect 40539 338948 40540 339012
rect 40604 338948 40605 339012
rect 40539 338947 40605 338948
rect 40542 312357 40602 338947
rect 40726 313853 40786 339763
rect 42011 338876 42077 338877
rect 42011 338812 42012 338876
rect 42076 338812 42077 338876
rect 42011 338811 42077 338812
rect 40907 337380 40973 337381
rect 40907 337316 40908 337380
rect 40972 337316 40973 337380
rect 40907 337315 40973 337316
rect 40723 313852 40789 313853
rect 40723 313788 40724 313852
rect 40788 313788 40789 313852
rect 40723 313787 40789 313788
rect 40910 313173 40970 337315
rect 41643 336972 41709 336973
rect 41643 336908 41644 336972
rect 41708 336908 41709 336972
rect 41643 336907 41709 336908
rect 41275 335748 41341 335749
rect 41275 335684 41276 335748
rect 41340 335684 41341 335748
rect 41275 335683 41341 335684
rect 41091 335340 41157 335341
rect 41091 335276 41092 335340
rect 41156 335276 41157 335340
rect 41091 335275 41157 335276
rect 41094 317389 41154 335275
rect 41278 321197 41338 335683
rect 41459 327860 41525 327861
rect 41459 327796 41460 327860
rect 41524 327796 41525 327860
rect 41459 327795 41525 327796
rect 41275 321196 41341 321197
rect 41275 321132 41276 321196
rect 41340 321132 41341 321196
rect 41275 321131 41341 321132
rect 41462 319973 41522 327795
rect 41459 319972 41525 319973
rect 41459 319908 41460 319972
rect 41524 319908 41525 319972
rect 41459 319907 41525 319908
rect 41091 317388 41157 317389
rect 41091 317324 41092 317388
rect 41156 317324 41157 317388
rect 41091 317323 41157 317324
rect 41646 315893 41706 336907
rect 41827 327724 41893 327725
rect 41827 327660 41828 327724
rect 41892 327660 41893 327724
rect 41827 327659 41893 327660
rect 41830 324869 41890 327659
rect 41827 324868 41893 324869
rect 41827 324804 41828 324868
rect 41892 324804 41893 324868
rect 41827 324803 41893 324804
rect 41643 315892 41709 315893
rect 41643 315828 41644 315892
rect 41708 315828 41709 315892
rect 41643 315827 41709 315828
rect 42014 315485 42074 338811
rect 675526 333573 675586 343571
rect 675710 340781 675770 345750
rect 675707 340780 675773 340781
rect 675707 340716 675708 340780
rect 675772 340716 675773 340780
rect 675707 340715 675773 340716
rect 675894 339421 675954 346430
rect 675891 339420 675957 339421
rect 675891 339356 675892 339420
rect 675956 339356 675957 339420
rect 675891 339355 675957 339356
rect 676078 337925 676138 350490
rect 676075 337924 676141 337925
rect 676075 337860 676076 337924
rect 676140 337860 676141 337924
rect 676075 337859 676141 337860
rect 675523 333572 675589 333573
rect 675523 333508 675524 333572
rect 675588 333508 675589 333572
rect 675523 333507 675589 333508
rect 676262 325549 676322 351870
rect 676446 325685 676506 353910
rect 676811 351150 676877 351151
rect 676811 351086 676812 351150
rect 676876 351086 676877 351150
rect 676811 351085 676877 351086
rect 676627 346628 676693 346629
rect 676627 346564 676628 346628
rect 676692 346564 676693 346628
rect 676627 346563 676693 346564
rect 676630 332621 676690 346563
rect 676814 335341 676874 351085
rect 677179 346492 677245 346493
rect 677179 346428 677180 346492
rect 677244 346428 677245 346492
rect 677179 346427 677245 346428
rect 677182 340890 677242 346427
rect 676998 340830 677242 340890
rect 676998 335885 677058 340830
rect 676995 335884 677061 335885
rect 676995 335820 676996 335884
rect 677060 335820 677061 335884
rect 676995 335819 677061 335820
rect 676811 335340 676877 335341
rect 676811 335276 676812 335340
rect 676876 335276 676877 335340
rect 676811 335275 676877 335276
rect 676627 332620 676693 332621
rect 676627 332556 676628 332620
rect 676692 332556 676693 332620
rect 676627 332555 676693 332556
rect 676443 325684 676509 325685
rect 676443 325620 676444 325684
rect 676508 325620 676509 325684
rect 676443 325619 676509 325620
rect 676259 325548 676325 325549
rect 676259 325484 676260 325548
rect 676324 325484 676325 325548
rect 676259 325483 676325 325484
rect 42011 315484 42077 315485
rect 42011 315420 42012 315484
rect 42076 315420 42077 315484
rect 42011 315419 42077 315420
rect 40907 313172 40973 313173
rect 40907 313108 40908 313172
rect 40972 313108 40973 313172
rect 40907 313107 40973 313108
rect 40539 312356 40605 312357
rect 40539 312292 40540 312356
rect 40604 312292 40605 312356
rect 40539 312291 40605 312292
rect 676443 308684 676509 308685
rect 676443 308620 676444 308684
rect 676508 308620 676509 308684
rect 676443 308619 676509 308620
rect 675891 308004 675957 308005
rect 675891 307940 675892 308004
rect 675956 307940 675957 308004
rect 675891 307939 675957 307940
rect 675894 306390 675954 307939
rect 676259 307052 676325 307053
rect 676259 306988 676260 307052
rect 676324 306988 676325 307052
rect 676259 306987 676325 306988
rect 675526 306330 675954 306390
rect 675339 297396 675405 297397
rect 675339 297332 675340 297396
rect 675404 297332 675405 297396
rect 675339 297331 675405 297332
rect 42747 296852 42813 296853
rect 42747 296788 42748 296852
rect 42812 296788 42813 296852
rect 42747 296787 42813 296788
rect 40542 296110 41890 296170
rect 40542 269109 40602 296110
rect 41830 296037 41890 296110
rect 41827 296036 41893 296037
rect 41827 295972 41828 296036
rect 41892 295972 41893 296036
rect 41827 295971 41893 295972
rect 42011 295628 42077 295629
rect 42011 295564 42012 295628
rect 42076 295564 42077 295628
rect 42011 295563 42077 295564
rect 41827 294404 41893 294405
rect 41827 294340 41828 294404
rect 41892 294340 41893 294404
rect 41827 294339 41893 294340
rect 41830 294130 41890 294339
rect 40726 294070 41890 294130
rect 40726 269789 40786 294070
rect 40910 293390 41890 293450
rect 40910 279853 40970 293390
rect 41830 293181 41890 293390
rect 41827 293180 41893 293181
rect 41827 293116 41828 293180
rect 41892 293116 41893 293180
rect 41827 293115 41893 293116
rect 41827 292772 41893 292773
rect 41827 292770 41828 292772
rect 41094 292710 41828 292770
rect 40907 279852 40973 279853
rect 40907 279788 40908 279852
rect 40972 279788 40973 279852
rect 40907 279787 40973 279788
rect 41094 278085 41154 292710
rect 41827 292708 41828 292710
rect 41892 292708 41893 292772
rect 41827 292707 41893 292708
rect 42014 292090 42074 295563
rect 42563 293996 42629 293997
rect 42563 293932 42564 293996
rect 42628 293932 42629 293996
rect 42563 293931 42629 293932
rect 41646 292030 42074 292090
rect 41459 284884 41525 284885
rect 41459 284820 41460 284884
rect 41524 284820 41525 284884
rect 41459 284819 41525 284820
rect 41462 281485 41522 284819
rect 41459 281484 41525 281485
rect 41459 281420 41460 281484
rect 41524 281420 41525 281484
rect 41459 281419 41525 281420
rect 41091 278084 41157 278085
rect 41091 278020 41092 278084
rect 41156 278020 41157 278084
rect 41091 278019 41157 278020
rect 41646 272237 41706 292030
rect 42566 290730 42626 293931
rect 41830 290670 42626 290730
rect 41830 273053 41890 290670
rect 42750 277410 42810 296787
rect 675342 292093 675402 297331
rect 675526 292637 675586 306330
rect 676075 305420 676141 305421
rect 676075 305356 676076 305420
rect 676140 305356 676141 305420
rect 676075 305355 676141 305356
rect 675707 299436 675773 299437
rect 675707 299372 675708 299436
rect 675772 299372 675773 299436
rect 675707 299371 675773 299372
rect 675710 294813 675770 299371
rect 675891 297940 675957 297941
rect 675891 297876 675892 297940
rect 675956 297876 675957 297940
rect 675891 297875 675957 297876
rect 675707 294812 675773 294813
rect 675707 294748 675708 294812
rect 675772 294748 675773 294812
rect 675707 294747 675773 294748
rect 675523 292636 675589 292637
rect 675523 292572 675524 292636
rect 675588 292572 675589 292636
rect 675894 292590 675954 297875
rect 675523 292571 675589 292572
rect 675710 292530 675954 292590
rect 675339 292092 675405 292093
rect 675339 292028 675340 292092
rect 675404 292028 675405 292092
rect 675339 292027 675405 292028
rect 675710 288421 675770 292530
rect 675707 288420 675773 288421
rect 675707 288356 675708 288420
rect 675772 288356 675773 288420
rect 675707 288355 675773 288356
rect 676078 285565 676138 305355
rect 676075 285564 676141 285565
rect 676075 285500 676076 285564
rect 676140 285500 676141 285564
rect 676075 285499 676141 285500
rect 676262 281485 676322 306987
rect 676446 283661 676506 308619
rect 676627 305012 676693 305013
rect 676627 304948 676628 305012
rect 676692 304948 676693 305012
rect 676627 304947 676693 304948
rect 676630 287333 676690 304947
rect 676627 287332 676693 287333
rect 676627 287268 676628 287332
rect 676692 287268 676693 287332
rect 676627 287267 676693 287268
rect 676443 283660 676509 283661
rect 676443 283596 676444 283660
rect 676508 283596 676509 283660
rect 676443 283595 676509 283596
rect 676259 281484 676325 281485
rect 676259 281420 676260 281484
rect 676324 281420 676325 281484
rect 676259 281419 676325 281420
rect 42014 277350 42810 277410
rect 41827 273052 41893 273053
rect 41827 272988 41828 273052
rect 41892 272988 41893 273052
rect 41827 272987 41893 272988
rect 41643 272236 41709 272237
rect 41643 272172 41644 272236
rect 41708 272172 41709 272236
rect 41643 272171 41709 272172
rect 42014 270469 42074 277350
rect 42011 270468 42077 270469
rect 42011 270404 42012 270468
rect 42076 270404 42077 270468
rect 42011 270403 42077 270404
rect 40723 269788 40789 269789
rect 40723 269724 40724 269788
rect 40788 269724 40789 269788
rect 40723 269723 40789 269724
rect 40539 269108 40605 269109
rect 40539 269044 40540 269108
rect 40604 269044 40605 269108
rect 40539 269043 40605 269044
rect 677179 260812 677245 260813
rect 677179 260748 677180 260812
rect 677244 260748 677245 260812
rect 677179 260747 677245 260748
rect 676995 260404 677061 260405
rect 676995 260340 676996 260404
rect 677060 260340 677061 260404
rect 676995 260339 677061 260340
rect 676811 259588 676877 259589
rect 676811 259524 676812 259588
rect 676876 259524 676877 259588
rect 676811 259523 676877 259524
rect 175043 253196 175109 253197
rect 175043 253132 175044 253196
rect 175108 253132 175109 253196
rect 175043 253131 175109 253132
rect 40539 250204 40605 250205
rect 40539 250140 40540 250204
rect 40604 250140 40605 250204
rect 40539 250139 40605 250140
rect 40542 232933 40602 250139
rect 40723 249796 40789 249797
rect 40723 249732 40724 249796
rect 40788 249732 40789 249796
rect 40723 249731 40789 249732
rect 40726 236741 40786 249731
rect 175046 241637 175106 253131
rect 675155 251564 675221 251565
rect 675155 251500 675156 251564
rect 675220 251500 675221 251564
rect 675155 251499 675221 251500
rect 675158 249661 675218 251499
rect 675155 249660 675221 249661
rect 675155 249596 675156 249660
rect 675220 249596 675221 249660
rect 675155 249595 675221 249596
rect 675707 245716 675773 245717
rect 675707 245652 675708 245716
rect 675772 245652 675773 245716
rect 675707 245651 675773 245652
rect 175043 241636 175109 241637
rect 175043 241572 175044 241636
rect 175108 241572 175109 241636
rect 175043 241571 175109 241572
rect 42011 238100 42077 238101
rect 42011 238036 42012 238100
rect 42076 238036 42077 238100
rect 42011 238035 42077 238036
rect 40723 236740 40789 236741
rect 40723 236676 40724 236740
rect 40788 236676 40789 236740
rect 40723 236675 40789 236676
rect 40539 232932 40605 232933
rect 40539 232868 40540 232932
rect 40604 232868 40605 232932
rect 40539 232867 40605 232868
rect 42014 227357 42074 238035
rect 42195 237420 42261 237421
rect 42195 237356 42196 237420
rect 42260 237356 42261 237420
rect 42195 237355 42261 237356
rect 42198 228989 42258 237355
rect 675710 236877 675770 245651
rect 676814 245445 676874 259523
rect 676811 245444 676877 245445
rect 676811 245380 676812 245444
rect 676876 245380 676877 245444
rect 676811 245379 676877 245380
rect 676998 238645 677058 260339
rect 677182 246669 677242 260747
rect 677179 246668 677245 246669
rect 677179 246604 677180 246668
rect 677244 246604 677245 246668
rect 677179 246603 677245 246604
rect 676995 238644 677061 238645
rect 676995 238580 676996 238644
rect 677060 238580 677061 238644
rect 676995 238579 677061 238580
rect 675707 236876 675773 236877
rect 675707 236812 675708 236876
rect 675772 236812 675773 236876
rect 675707 236811 675773 236812
rect 647371 231164 647437 231165
rect 647371 231100 647372 231164
rect 647436 231100 647437 231164
rect 647371 231099 647437 231100
rect 646451 229668 646517 229669
rect 646451 229604 646452 229668
rect 646516 229604 646517 229668
rect 646451 229603 646517 229604
rect 42195 228988 42261 228989
rect 42195 228924 42196 228988
rect 42260 228924 42261 228988
rect 42195 228923 42261 228924
rect 42011 227356 42077 227357
rect 42011 227292 42012 227356
rect 42076 227292 42077 227356
rect 42011 227291 42077 227292
rect 646454 213077 646514 229603
rect 647374 213077 647434 231099
rect 675891 218652 675957 218653
rect 675891 218588 675892 218652
rect 675956 218588 675957 218652
rect 675891 218587 675957 218588
rect 675707 218244 675773 218245
rect 675707 218180 675708 218244
rect 675772 218180 675773 218244
rect 675707 218179 675773 218180
rect 675523 217836 675589 217837
rect 675523 217772 675524 217836
rect 675588 217772 675589 217836
rect 675523 217771 675589 217772
rect 646451 213076 646517 213077
rect 646451 213012 646452 213076
rect 646516 213012 646517 213076
rect 646451 213011 646517 213012
rect 647371 213076 647437 213077
rect 647371 213012 647372 213076
rect 647436 213012 647437 213076
rect 647371 213011 647437 213012
rect 41643 209812 41709 209813
rect 41643 209748 41644 209812
rect 41708 209748 41709 209812
rect 41643 209747 41709 209748
rect 40539 209404 40605 209405
rect 40539 209340 40540 209404
rect 40604 209340 40605 209404
rect 40539 209339 40605 209340
rect 40542 183021 40602 209339
rect 41459 208588 41525 208589
rect 41459 208524 41460 208588
rect 41524 208524 41525 208588
rect 41459 208523 41525 208524
rect 40723 206956 40789 206957
rect 40723 206892 40724 206956
rect 40788 206892 40789 206956
rect 40723 206891 40789 206892
rect 40726 195397 40786 206891
rect 40723 195396 40789 195397
rect 40723 195332 40724 195396
rect 40788 195332 40789 195396
rect 40723 195331 40789 195332
rect 41462 190229 41522 208523
rect 41646 195261 41706 209747
rect 675339 207228 675405 207229
rect 675339 207164 675340 207228
rect 675404 207164 675405 207228
rect 675339 207163 675405 207164
rect 675342 200130 675402 207163
rect 675526 202741 675586 217771
rect 675710 209949 675770 218179
rect 675894 214570 675954 218587
rect 676627 215558 676693 215559
rect 676627 215494 676628 215558
rect 676692 215494 676693 215558
rect 676627 215493 676693 215494
rect 675894 214510 676322 214570
rect 676075 214028 676141 214029
rect 676075 213964 676076 214028
rect 676140 213964 676141 214028
rect 676075 213963 676141 213964
rect 675707 209948 675773 209949
rect 675707 209884 675708 209948
rect 675772 209884 675773 209948
rect 675707 209883 675773 209884
rect 676078 209810 676138 213963
rect 675710 209750 676138 209810
rect 675710 204237 675770 209750
rect 675891 209676 675957 209677
rect 675891 209612 675892 209676
rect 675956 209612 675957 209676
rect 675891 209611 675957 209612
rect 675894 205597 675954 209611
rect 676075 208316 676141 208317
rect 676075 208252 676076 208316
rect 676140 208252 676141 208316
rect 676075 208251 676141 208252
rect 675891 205596 675957 205597
rect 675891 205532 675892 205596
rect 675956 205532 675957 205596
rect 675891 205531 675957 205532
rect 676078 205053 676138 208251
rect 676075 205052 676141 205053
rect 676075 204988 676076 205052
rect 676140 204988 676141 205052
rect 676075 204987 676141 204988
rect 675707 204236 675773 204237
rect 675707 204172 675708 204236
rect 675772 204172 675773 204236
rect 675707 204171 675773 204172
rect 675523 202740 675589 202741
rect 675523 202676 675524 202740
rect 675588 202676 675589 202740
rect 675523 202675 675589 202676
rect 675342 200070 676138 200130
rect 41827 199340 41893 199341
rect 41827 199276 41828 199340
rect 41892 199276 41893 199340
rect 41827 199275 41893 199276
rect 41643 195260 41709 195261
rect 41643 195196 41644 195260
rect 41708 195196 41709 195260
rect 41643 195195 41709 195196
rect 41459 190228 41525 190229
rect 41459 190164 41460 190228
rect 41524 190164 41525 190228
rect 41459 190163 41525 190164
rect 41830 184245 41890 199275
rect 676078 198389 676138 200070
rect 676075 198388 676141 198389
rect 676075 198324 676076 198388
rect 676140 198324 676141 198388
rect 676075 198323 676141 198324
rect 42195 195396 42261 195397
rect 42195 195332 42196 195396
rect 42260 195332 42261 195396
rect 42195 195331 42261 195332
rect 42198 187373 42258 195331
rect 676262 190229 676322 214510
rect 676443 211308 676509 211309
rect 676443 211244 676444 211308
rect 676508 211244 676509 211308
rect 676443 211243 676509 211244
rect 676446 190365 676506 211243
rect 676630 195397 676690 215493
rect 676995 214334 677061 214335
rect 676995 214270 676996 214334
rect 677060 214270 677061 214334
rect 676995 214269 677061 214270
rect 676811 211444 676877 211445
rect 676811 211380 676812 211444
rect 676876 211380 676877 211444
rect 676811 211379 676877 211380
rect 676814 201381 676874 211379
rect 676998 202877 677058 214269
rect 676995 202876 677061 202877
rect 676995 202812 676996 202876
rect 677060 202812 677061 202876
rect 676995 202811 677061 202812
rect 676811 201380 676877 201381
rect 676811 201316 676812 201380
rect 676876 201316 676877 201380
rect 676811 201315 676877 201316
rect 676627 195396 676693 195397
rect 676627 195332 676628 195396
rect 676692 195332 676693 195396
rect 676627 195331 676693 195332
rect 676443 190364 676509 190365
rect 676443 190300 676444 190364
rect 676508 190300 676509 190364
rect 676443 190299 676509 190300
rect 676259 190228 676325 190229
rect 676259 190164 676260 190228
rect 676324 190164 676325 190228
rect 676259 190163 676325 190164
rect 42195 187372 42261 187373
rect 42195 187308 42196 187372
rect 42260 187308 42261 187372
rect 42195 187307 42261 187308
rect 41827 184244 41893 184245
rect 41827 184180 41828 184244
rect 41892 184180 41893 184244
rect 41827 184179 41893 184180
rect 40539 183020 40605 183021
rect 40539 182956 40540 183020
rect 40604 182956 40605 183020
rect 40539 182955 40605 182956
rect 675339 174044 675405 174045
rect 675339 173980 675340 174044
rect 675404 173980 675405 174044
rect 675339 173979 675405 173980
rect 675342 159493 675402 173979
rect 676078 173710 676322 173770
rect 676078 173501 676138 173710
rect 676075 173500 676141 173501
rect 676075 173436 676076 173500
rect 676140 173436 676141 173500
rect 676075 173435 676141 173436
rect 676262 173090 676322 173710
rect 676262 173030 676506 173090
rect 676075 171868 676141 171869
rect 676075 171804 676076 171868
rect 676140 171804 676141 171868
rect 676075 171803 676141 171804
rect 676078 171730 676138 171803
rect 676078 171670 676322 171730
rect 675891 170780 675957 170781
rect 675891 170716 675892 170780
rect 675956 170716 675957 170780
rect 675891 170715 675957 170716
rect 675707 169692 675773 169693
rect 675707 169628 675708 169692
rect 675772 169628 675773 169692
rect 675707 169627 675773 169628
rect 675523 162620 675589 162621
rect 675523 162556 675524 162620
rect 675588 162556 675589 162620
rect 675523 162555 675589 162556
rect 675339 159492 675405 159493
rect 675339 159428 675340 159492
rect 675404 159428 675405 159492
rect 675339 159427 675405 159428
rect 675526 157045 675586 162555
rect 675710 157453 675770 169627
rect 675707 157452 675773 157453
rect 675707 157388 675708 157452
rect 675772 157388 675773 157452
rect 675707 157387 675773 157388
rect 675523 157044 675589 157045
rect 675523 156980 675524 157044
rect 675588 156980 675589 157044
rect 675523 156979 675589 156980
rect 675894 156365 675954 170715
rect 676075 162756 676141 162757
rect 676075 162692 676076 162756
rect 676140 162692 676141 162756
rect 676075 162691 676141 162692
rect 675891 156364 675957 156365
rect 675891 156300 675892 156364
rect 675956 156300 675957 156364
rect 675891 156299 675957 156300
rect 676078 153101 676138 162691
rect 676075 153100 676141 153101
rect 676075 153036 676076 153100
rect 676140 153036 676141 153100
rect 676075 153035 676141 153036
rect 676262 146301 676322 171670
rect 676446 148477 676506 173030
rect 676627 166428 676693 166429
rect 676627 166364 676628 166428
rect 676692 166364 676693 166428
rect 676627 166363 676693 166364
rect 676811 166428 676877 166429
rect 676811 166364 676812 166428
rect 676876 166364 676877 166428
rect 676811 166363 676877 166364
rect 676630 151605 676690 166363
rect 676814 160037 676874 166363
rect 676811 160036 676877 160037
rect 676811 159972 676812 160036
rect 676876 159972 676877 160036
rect 676811 159971 676877 159972
rect 676627 151604 676693 151605
rect 676627 151540 676628 151604
rect 676692 151540 676693 151604
rect 676627 151539 676693 151540
rect 676443 148476 676509 148477
rect 676443 148412 676444 148476
rect 676508 148412 676509 148476
rect 676443 148411 676509 148412
rect 676259 146300 676325 146301
rect 676259 146236 676260 146300
rect 676324 146236 676325 146300
rect 676259 146235 676325 146236
rect 675339 128892 675405 128893
rect 675339 128828 675340 128892
rect 675404 128828 675405 128892
rect 675339 128827 675405 128828
rect 675342 114205 675402 128827
rect 676259 126580 676325 126581
rect 676259 126516 676260 126580
rect 676324 126516 676325 126580
rect 676259 126515 676325 126516
rect 675707 124948 675773 124949
rect 675707 124884 675708 124948
rect 675772 124884 675773 124948
rect 675707 124883 675773 124884
rect 675523 117196 675589 117197
rect 675523 117132 675524 117196
rect 675588 117132 675589 117196
rect 675523 117131 675589 117132
rect 675339 114204 675405 114205
rect 675339 114140 675340 114204
rect 675404 114140 675405 114204
rect 675339 114139 675405 114140
rect 675526 111757 675586 117131
rect 675710 112573 675770 124883
rect 676075 118012 676141 118013
rect 676075 117948 676076 118012
rect 676140 117948 676141 118012
rect 676075 117947 676141 117948
rect 675891 117332 675957 117333
rect 675891 117268 675892 117332
rect 675956 117268 675957 117332
rect 675891 117267 675957 117268
rect 675707 112572 675773 112573
rect 675707 112508 675708 112572
rect 675772 112508 675773 112572
rect 675707 112507 675773 112508
rect 675523 111756 675589 111757
rect 675523 111692 675524 111756
rect 675588 111692 675589 111756
rect 675523 111691 675589 111692
rect 675894 104821 675954 117267
rect 676078 108221 676138 117947
rect 676075 108220 676141 108221
rect 676075 108156 676076 108220
rect 676140 108156 676141 108220
rect 676075 108155 676141 108156
rect 675891 104820 675957 104821
rect 675891 104756 675892 104820
rect 675956 104756 675957 104820
rect 675891 104755 675957 104756
rect 676262 101421 676322 126515
rect 676443 124540 676509 124541
rect 676443 124476 676444 124540
rect 676508 124476 676509 124540
rect 676443 124475 676509 124476
rect 676446 109037 676506 124475
rect 676811 121684 676877 121685
rect 676811 121620 676812 121684
rect 676876 121620 676877 121684
rect 676811 121619 676877 121620
rect 676443 109036 676509 109037
rect 676443 108972 676444 109036
rect 676508 108972 676509 109036
rect 676443 108971 676509 108972
rect 676814 103189 676874 121619
rect 676811 103188 676877 103189
rect 676811 103124 676812 103188
rect 676876 103124 676877 103188
rect 676811 103123 676877 103124
rect 676259 101420 676325 101421
rect 676259 101356 676260 101420
rect 676324 101356 676325 101420
rect 676259 101355 676325 101356
rect 639827 96524 639893 96525
rect 639827 96460 639828 96524
rect 639892 96460 639893 96524
rect 639827 96459 639893 96460
rect 634675 95844 634741 95845
rect 634675 95780 634676 95844
rect 634740 95780 634741 95844
rect 634675 95779 634741 95780
rect 634678 77757 634738 95779
rect 639830 77757 639890 96459
rect 634675 77756 634741 77757
rect 634675 77692 634676 77756
rect 634740 77692 634741 77756
rect 634675 77691 634741 77692
rect 639827 77756 639893 77757
rect 639827 77692 639828 77756
rect 639892 77692 639893 77756
rect 639827 77691 639893 77692
rect 638907 75172 638973 75173
rect 638907 75108 638908 75172
rect 638972 75108 638973 75172
rect 638907 75107 638973 75108
rect 638910 52461 638970 75107
rect 638907 52460 638973 52461
rect 638907 52396 638908 52460
rect 638972 52396 638973 52460
rect 638907 52395 638973 52396
rect 520227 50556 520293 50557
rect 520227 50492 520228 50556
rect 520292 50492 520293 50556
rect 520227 50491 520293 50492
rect 514707 50284 514773 50285
rect 514707 50220 514708 50284
rect 514772 50220 514773 50284
rect 514707 50219 514773 50220
rect 187555 47564 187621 47565
rect 187555 47500 187556 47564
rect 187620 47500 187621 47564
rect 187555 47499 187621 47500
rect 141923 44028 141989 44029
rect 141923 43964 141924 44028
rect 141988 43964 141989 44028
rect 141923 43963 141989 43964
rect 141926 40357 141986 43963
rect 187558 42125 187618 47499
rect 471651 46612 471717 46613
rect 471651 46548 471652 46612
rect 471716 46548 471717 46612
rect 471651 46547 471717 46548
rect 460611 46340 460677 46341
rect 460611 46276 460612 46340
rect 460676 46276 460677 46340
rect 460611 46275 460677 46276
rect 365115 45116 365181 45117
rect 365115 45052 365116 45116
rect 365180 45052 365181 45116
rect 365115 45051 365181 45052
rect 361987 44980 362053 44981
rect 361987 44916 361988 44980
rect 362052 44916 362053 44980
rect 361987 44915 362053 44916
rect 310099 44844 310165 44845
rect 310099 44780 310100 44844
rect 310164 44780 310165 44844
rect 310099 44779 310165 44780
rect 310102 42397 310162 44779
rect 310099 42396 310165 42397
rect 310099 42332 310100 42396
rect 310164 42332 310165 42396
rect 310099 42331 310165 42332
rect 361990 42125 362050 44915
rect 365118 42125 365178 45051
rect 460614 42125 460674 46275
rect 471654 42125 471714 46547
rect 514710 42125 514770 50219
rect 518571 46748 518637 46749
rect 518571 46684 518572 46748
rect 518636 46684 518637 46748
rect 518571 46683 518637 46684
rect 518574 42397 518634 46683
rect 518571 42396 518637 42397
rect 518571 42332 518572 42396
rect 518636 42332 518637 42396
rect 518571 42331 518637 42332
rect 520230 42125 520290 50491
rect 521699 50420 521765 50421
rect 521699 50356 521700 50420
rect 521764 50356 521765 50420
rect 521699 50355 521765 50356
rect 521702 42125 521762 50355
rect 529795 50284 529861 50285
rect 529795 50220 529796 50284
rect 529860 50220 529861 50284
rect 529795 50219 529861 50220
rect 529798 42125 529858 50219
rect 187555 42124 187621 42125
rect 187555 42060 187556 42124
rect 187620 42060 187621 42124
rect 187555 42059 187621 42060
rect 361987 42124 362053 42125
rect 361987 42060 361988 42124
rect 362052 42060 362053 42124
rect 361987 42059 362053 42060
rect 365115 42124 365181 42125
rect 365115 42060 365116 42124
rect 365180 42060 365181 42124
rect 365115 42059 365181 42060
rect 460611 42124 460677 42125
rect 460611 42060 460612 42124
rect 460676 42060 460677 42124
rect 460611 42059 460677 42060
rect 471651 42124 471717 42125
rect 471651 42060 471652 42124
rect 471716 42060 471717 42124
rect 471651 42059 471717 42060
rect 514707 42124 514773 42125
rect 514707 42060 514708 42124
rect 514772 42060 514773 42124
rect 514707 42059 514773 42060
rect 520227 42124 520293 42125
rect 520227 42060 520228 42124
rect 520292 42060 520293 42124
rect 520227 42059 520293 42060
rect 521699 42124 521765 42125
rect 521699 42060 521700 42124
rect 521764 42060 521765 42124
rect 521699 42059 521765 42060
rect 529795 42124 529861 42125
rect 529795 42060 529796 42124
rect 529860 42060 529861 42124
rect 529795 42059 529861 42060
rect 141923 40356 141989 40357
rect 141923 40292 141924 40356
rect 141988 40292 141989 40356
rect 141923 40291 141989 40292
<< via4 >>
rect 240278 997102 240514 997338
rect 246350 997324 246436 997338
rect 246436 997324 246500 997338
rect 246500 997324 246586 997338
rect 246350 997102 246586 997324
rect 485550 997102 485786 997338
rect 505054 997102 505290 997338
rect 536518 997102 536754 997338
rect 554550 997102 554786 997338
<< metal5 >>
rect 78440 1018512 90960 1031002
rect 129840 1018512 142360 1031002
rect 181240 1018512 193760 1031002
rect 232640 1018512 245160 1031002
rect 284240 1018512 296760 1031002
rect 334810 1018624 346978 1030789
rect 386040 1018512 398560 1031002
rect 475040 1018512 487560 1031002
rect 526440 1018512 538960 1031002
rect 577010 1018624 589178 1030789
rect 628240 1018512 640760 1031002
rect 240236 997338 246628 997380
rect 240236 997102 240278 997338
rect 240514 997102 246350 997338
rect 246586 997102 246628 997338
rect 240236 997060 246628 997102
rect 485508 997338 505332 997380
rect 485508 997102 485550 997338
rect 485786 997102 505054 997338
rect 505290 997102 505332 997338
rect 485508 997060 505332 997102
rect 536476 997338 554828 997380
rect 536476 997102 536518 997338
rect 536754 997102 554550 997338
rect 554786 997102 554828 997338
rect 536476 997060 554828 997102
rect 6598 956440 19088 968960
rect 698512 952840 711002 965360
rect 6167 914054 19620 924934
rect 697980 909666 711433 920546
rect 6811 871210 18976 883378
rect 698512 863640 711002 876160
rect 6811 829010 18976 841178
rect 698624 819822 710789 831990
rect 6598 786640 19088 799160
rect 698512 774440 711002 786960
rect 6598 743440 19088 755960
rect 698512 729440 711002 741960
rect 6598 700240 19088 712760
rect 698512 684440 711002 696960
rect 6598 657040 19088 669560
rect 698512 639240 711002 651760
rect 6598 613840 19088 626360
rect 698512 594240 711002 606760
rect 6598 570640 19088 583160
rect 698512 549040 711002 561560
rect 6598 527440 19088 539960
rect 698624 505222 710789 517390
rect 6811 484410 18976 496578
rect 697980 461866 711433 472746
rect 6167 442854 19620 453734
rect 698624 417022 710789 429190
rect 6598 399840 19088 412360
rect 698512 371840 711002 384360
rect 6598 356640 19088 369160
rect 698512 326640 711002 339160
rect 6598 313440 19088 325960
rect 6598 270240 19088 282760
rect 698512 281640 711002 294160
rect 6598 227040 19088 239560
rect 698512 236640 711002 249160
rect 6598 183840 19088 196360
rect 698512 191440 711002 203960
rect 698512 146440 711002 158960
rect 6811 111610 18976 123778
rect 698512 101240 711002 113760
rect 6167 70054 19620 80934
rect 80222 6811 92390 18976
rect 136713 7143 144150 18309
rect 187640 6598 200160 19088
rect 243266 6167 254146 19620
rect 296240 6598 308760 19088
rect 351040 6598 363560 19088
rect 405840 6598 418360 19088
rect 460640 6598 473160 19088
rect 515440 6598 527960 19088
rect 570422 6811 582590 18976
rect 624222 6811 636390 18976
use caravel_logo  caravel_logo_0
timestamp 1638586901
transform 1 0 269006 0 1 5020
box -2520 0 15000 15560
use caravel_motto  caravel_motto_0
timestamp 1637698310
transform 1 0 -52778 0 1 -5036
box 373080 14838 395618 19242
use caravel_power_routing  caravel_power_routing_0
timestamp 1650914956
transform 1 0 0 0 1 0
box 0 0 717600 1037600
use caravel_clocking  clocking
timestamp 1638876627
transform 1 0 626764 0 1 63284
box -38 -48 20000 12000
use copyright_block  copyright_block_0
timestamp 1649268499
transform 1 0 149554 0 1 16026
box -262 -10348 35048 2764
use gpio_control_block  gpio_control_bidir_1\[0\]
timestamp 1650900217
transform -1 0 710203 0 1 121000
box 882 416 34000 13000
use gpio_control_block  gpio_control_bidir_1\[1\]
timestamp 1650900217
transform -1 0 710203 0 1 166200
box 882 416 34000 13000
use gpio_control_block  gpio_control_bidir_2\[0\]
timestamp 1650900217
transform 1 0 7631 0 1 289000
box 882 416 34000 13000
use gpio_control_block  gpio_control_bidir_2\[1\]
timestamp 1650900217
transform 1 0 7631 0 1 245800
box 882 416 34000 13000
use gpio_control_block  gpio_control_bidir_2\[2\]
timestamp 1650900217
transform 1 0 7631 0 1 202600
box 882 416 34000 13000
use gpio_control_block  gpio_control_in_1\[0\]
timestamp 1650900217
transform -1 0 710203 0 1 523800
box 882 416 34000 13000
use gpio_control_block  gpio_control_in_1\[1\]
timestamp 1650900217
transform -1 0 710203 0 1 568800
box 882 416 34000 13000
use gpio_control_block  gpio_control_in_1\[2\]
timestamp 1650900217
transform -1 0 710203 0 1 614000
box 882 416 34000 13000
use gpio_control_block  gpio_control_in_1\[3\]
timestamp 1650900217
transform -1 0 710203 0 1 659000
box 882 416 34000 13000
use gpio_control_block  gpio_control_in_1\[4\]
timestamp 1650900217
transform -1 0 710203 0 1 704200
box 882 416 34000 13000
use gpio_control_block  gpio_control_in_1\[5\]
timestamp 1650900217
transform -1 0 710203 0 1 749200
box 882 416 34000 13000
use gpio_control_block  gpio_control_in_1\[6\]
timestamp 1650900217
transform -1 0 710203 0 1 927600
box 882 416 34000 13000
use gpio_control_block  gpio_control_in_1\[7\]
timestamp 1650900217
transform 0 1 549200 -1 0 1030077
box 882 416 34000 13000
use gpio_control_block  gpio_control_in_1\[8\]
timestamp 1650900217
transform 0 1 497800 -1 0 1030077
box 882 416 34000 13000
use gpio_control_block  gpio_control_in_1\[9\]
timestamp 1650900217
transform 0 1 420800 -1 0 1030077
box 882 416 34000 13000
use gpio_control_block  gpio_control_in_1\[10\]
timestamp 1650900217
transform 0 1 353400 -1 0 1030077
box 882 416 34000 13000
use gpio_control_block  gpio_control_in_1a\[0\]
timestamp 1650900217
transform -1 0 710203 0 1 211200
box 882 416 34000 13000
use gpio_control_block  gpio_control_in_1a\[1\]
timestamp 1650900217
transform -1 0 710203 0 1 256400
box 882 416 34000 13000
use gpio_control_block  gpio_control_in_1a\[2\]
timestamp 1650900217
transform -1 0 710203 0 1 301400
box 882 416 34000 13000
use gpio_control_block  gpio_control_in_1a\[3\]
timestamp 1650900217
transform -1 0 710203 0 1 346400
box 882 416 34000 13000
use gpio_control_block  gpio_control_in_1a\[4\]
timestamp 1650900217
transform -1 0 710203 0 1 391600
box 882 416 34000 13000
use gpio_control_block  gpio_control_in_1a\[5\]
timestamp 1650900217
transform -1 0 710203 0 1 479800
box 882 416 34000 13000
use gpio_control_block  gpio_control_in_2\[0\]
timestamp 1650900217
transform 0 1 303000 -1 0 1030077
box 882 416 34000 13000
use gpio_control_block  gpio_control_in_2\[1\]
timestamp 1650900217
transform 0 1 251400 -1 0 1030077
box 882 416 34000 13000
use gpio_control_block  gpio_control_in_2\[2\]
timestamp 1650900217
transform 0 1 200000 -1 0 1030077
box 882 416 34000 13000
use gpio_control_block  gpio_control_in_2\[3\]
timestamp 1650900217
transform 0 1 148600 -1 0 1030077
box 882 416 34000 13000
use gpio_control_block  gpio_control_in_2\[4\]
timestamp 1650900217
transform 0 1 97200 -1 0 1030077
box 882 416 34000 13000
use gpio_control_block  gpio_control_in_2\[5\]
timestamp 1650900217
transform 1 0 7631 0 1 931200
box 882 416 34000 13000
use gpio_control_block  gpio_control_in_2\[6\]
timestamp 1650900217
transform 1 0 7631 0 1 805400
box 882 416 34000 13000
use gpio_control_block  gpio_control_in_2\[7\]
timestamp 1650900217
transform 1 0 7631 0 1 762200
box 882 416 34000 13000
use gpio_control_block  gpio_control_in_2\[8\]
timestamp 1650900217
transform 1 0 7631 0 1 719000
box 882 416 34000 13000
use gpio_control_block  gpio_control_in_2\[9\]
timestamp 1650900217
transform 1 0 7631 0 1 675800
box 882 416 34000 13000
use gpio_control_block  gpio_control_in_2\[10\]
timestamp 1650900217
transform 1 0 7631 0 1 632600
box 882 416 34000 13000
use gpio_control_block  gpio_control_in_2\[11\]
timestamp 1650900217
transform 1 0 7631 0 1 589400
box 882 416 34000 13000
use gpio_control_block  gpio_control_in_2\[12\]
timestamp 1650900217
transform 1 0 7631 0 1 546200
box 882 416 34000 13000
use gpio_control_block  gpio_control_in_2\[13\]
timestamp 1650900217
transform 1 0 7631 0 1 418600
box 882 416 34000 13000
use gpio_control_block  gpio_control_in_2\[14\]
timestamp 1650900217
transform 1 0 7631 0 1 375400
box 882 416 34000 13000
use gpio_control_block  gpio_control_in_2\[15\]
timestamp 1650900217
transform 1 0 7631 0 1 332200
box 882 416 34000 13000
use gpio_defaults_block  gpio_defaults_block_0\[0\]
timestamp 1638587925
transform -1 0 709467 0 1 134000
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_0\[1\]
timestamp 1638587925
transform -1 0 709467 0 1 179200
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_2\[0\]
timestamp 1638587925
transform -1 0 709467 0 1 224200
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_2\[1\]
timestamp 1638587925
transform -1 0 709467 0 1 269400
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_2\[2\]
timestamp 1638587925
transform -1 0 709467 0 1 314400
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_5
timestamp 1638587925
transform -1 0 709467 0 1 359400
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_6
timestamp 1638587925
transform -1 0 709467 0 1 404600
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_7
timestamp 1638587925
transform -1 0 709467 0 1 492800
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_8
timestamp 1638587925
transform -1 0 709467 0 1 536800
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_9
timestamp 1638587925
transform -1 0 709467 0 1 581800
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_10
timestamp 1638587925
transform -1 0 709467 0 1 627000
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_11
timestamp 1638587925
transform -1 0 709467 0 1 672000
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_12
timestamp 1638587925
transform -1 0 709467 0 1 717200
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_13
timestamp 1638587925
transform -1 0 709467 0 1 762200
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_14
timestamp 1638587925
transform -1 0 709467 0 1 940600
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_15
timestamp 1638587925
transform 0 1 562194 -1 0 1029341
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_16
timestamp 1638587925
transform 0 1 510794 -1 0 1029341
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_17
timestamp 1638587925
transform 0 1 433794 -1 0 1029341
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_18
timestamp 1638587925
transform 0 1 366394 -1 0 1029341
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_19
timestamp 1638587925
transform 0 1 315994 -1 0 1029341
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_20
timestamp 1638587925
transform 0 1 264394 -1 0 1029341
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_21
timestamp 1638587925
transform 0 1 212994 -1 0 1029341
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_22
timestamp 1638587925
transform 0 1 161594 -1 0 1029341
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_23
timestamp 1638587925
transform 0 1 110194 -1 0 1029341
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_24
timestamp 1638587925
transform 1 0 8367 0 1 944200
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_25
timestamp 1638587925
transform 1 0 8367 0 1 818400
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_26
timestamp 1638587925
transform 1 0 8367 0 1 775200
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_27
timestamp 1638587925
transform 1 0 8367 0 1 732000
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_28
timestamp 1638587925
transform 1 0 8367 0 1 688800
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_29
timestamp 1638587925
transform 1 0 8367 0 1 645600
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_30
timestamp 1638587925
transform 1 0 8367 0 1 602400
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_31
timestamp 1638587925
transform 1 0 8367 0 1 559200
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_32
timestamp 1638587925
transform 1 0 8367 0 1 431600
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_33
timestamp 1638587925
transform 1 0 8367 0 1 388400
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_34
timestamp 1638587925
transform 1 0 8367 0 1 345200
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_35
timestamp 1638587925
transform 1 0 8367 0 1 302000
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_36
timestamp 1638587925
transform 1 0 8367 0 1 258800
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_37
timestamp 1638587925
transform 1 0 8367 0 1 215600
box -38 0 6018 2224
use housekeeping  housekeeping
timestamp 1638464048
transform 1 0 606434 0 1 100002
box 0 0 60046 110190
use mgmt_protect  mgmt_buffers
timestamp 1649962643
transform 1 0 192180 0 1 232036
box -400 -400 220400 32400
use user_project_wrapper  mprj
timestamp 1637147503
transform 1 0 65308 0 1 278718
box -8726 -7654 592650 711590
use open_source  open_source_0 hexdigits
timestamp 1638586442
transform 1 0 206830 0 1 2016
box 752 5164 29030 16242
use chip_io  padframe
timestamp 1638030917
transform 1 0 0 0 1 0
box 0 0 717600 1037600
use digital_pll  pll
timestamp 1638875307
transform 1 0 628146 0 1 80944
box 0 0 15000 15000
use simple_por  por
timestamp 1650914729
transform 1 0 650146 0 -1 55282
box -52 -62 11344 8684
use xres_buf  rstb_level
timestamp 1649268499
transform -1 0 145710 0 -1 50488
box 374 -400 3540 3800
use mgmt_core_wrapper  soc
timestamp 1638280046
transform 1 0 52034 0 1 53002
box 382 -400 524400 164400
use spare_logic_block  spare_logic\[0\]
timestamp 1638030917
transform 1 0 88632 0 1 232528
box 0 0 9000 9000
use spare_logic_block  spare_logic\[1\]
timestamp 1638030917
transform 1 0 168632 0 1 232528
box 0 0 9000 9000
use spare_logic_block  spare_logic\[2\]
timestamp 1638030917
transform 1 0 640874 0 1 220592
box 0 0 9000 9000
use spare_logic_block  spare_logic\[3\]
timestamp 1638030917
transform 1 0 428632 0 1 232528
box 0 0 9000 9000
use user_id_textblock  user_id_textblock_0
timestamp 1608324878
transform 1 0 96286 0 1 6596
box -656 1508 33720 10344
use user_id_programming  user_id_value
timestamp 1650371074
transform 1 0 656624 0 1 88126
box 0 0 7109 7077
<< labels >>
flabel metal5 s 187640 6598 200160 19088 0 FreeSans 25000 0 0 0 clock
port 0 nsew signal input
flabel metal5 s 351040 6598 363560 19088 0 FreeSans 25000 0 0 0 flash_clk
port 1 nsew signal tristate
flabel metal5 s 296240 6598 308760 19088 0 FreeSans 25000 0 0 0 flash_csb
port 2 nsew signal tristate
flabel metal5 s 405840 6598 418360 19088 0 FreeSans 25000 0 0 0 flash_io0
port 3 nsew signal tristate
flabel metal5 s 460640 6598 473160 19088 0 FreeSans 25000 0 0 0 flash_io1
port 4 nsew signal tristate
flabel metal5 s 515440 6598 527960 19088 0 FreeSans 25000 0 0 0 gpio
port 5 nsew signal bidirectional
flabel metal5 s 698512 101240 711002 113760 0 FreeSans 25000 0 0 0 mprj_io[0]
port 6 nsew signal bidirectional
flabel metal5 s 698512 684440 711002 696960 0 FreeSans 25000 0 0 0 mprj_io[10]
port 7 nsew signal bidirectional
flabel metal5 s 698512 729440 711002 741960 0 FreeSans 25000 0 0 0 mprj_io[11]
port 8 nsew signal bidirectional
flabel metal5 s 698512 774440 711002 786960 0 FreeSans 25000 0 0 0 mprj_io[12]
port 9 nsew signal bidirectional
flabel metal5 s 698512 863640 711002 876160 0 FreeSans 25000 0 0 0 mprj_io[13]
port 10 nsew signal bidirectional
flabel metal5 s 698512 952840 711002 965360 0 FreeSans 25000 0 0 0 mprj_io[14]
port 11 nsew signal bidirectional
flabel metal5 s 628240 1018512 640760 1031002 0 FreeSans 25000 0 0 0 mprj_io[15]
port 12 nsew signal bidirectional
flabel metal5 s 526440 1018512 538960 1031002 0 FreeSans 25000 0 0 0 mprj_io[16]
port 13 nsew signal bidirectional
flabel metal5 s 475040 1018512 487560 1031002 0 FreeSans 25000 0 0 0 mprj_io[17]
port 14 nsew signal bidirectional
flabel metal5 s 386040 1018512 398560 1031002 0 FreeSans 25000 0 0 0 mprj_io[18]
port 15 nsew signal bidirectional
flabel metal5 s 284240 1018512 296760 1031002 0 FreeSans 25000 0 0 0 mprj_io[19]
port 16 nsew signal bidirectional
flabel metal5 s 698512 146440 711002 158960 0 FreeSans 25000 0 0 0 mprj_io[1]
port 17 nsew signal bidirectional
flabel metal5 s 232640 1018512 245160 1031002 0 FreeSans 25000 0 0 0 mprj_io[20]
port 18 nsew signal bidirectional
flabel metal5 s 181240 1018512 193760 1031002 0 FreeSans 25000 0 0 0 mprj_io[21]
port 19 nsew signal bidirectional
flabel metal5 s 129840 1018512 142360 1031002 0 FreeSans 25000 0 0 0 mprj_io[22]
port 20 nsew signal bidirectional
flabel metal5 s 78440 1018512 90960 1031002 0 FreeSans 25000 0 0 0 mprj_io[23]
port 21 nsew signal bidirectional
flabel metal5 s 6598 956440 19088 968960 0 FreeSans 25000 0 0 0 mprj_io[24]
port 22 nsew signal bidirectional
flabel metal5 s 6598 786640 19088 799160 0 FreeSans 25000 0 0 0 mprj_io[25]
port 23 nsew signal bidirectional
flabel metal5 s 6598 743440 19088 755960 0 FreeSans 25000 0 0 0 mprj_io[26]
port 24 nsew signal bidirectional
flabel metal5 s 6598 700240 19088 712760 0 FreeSans 25000 0 0 0 mprj_io[27]
port 25 nsew signal bidirectional
flabel metal5 s 6598 657040 19088 669560 0 FreeSans 25000 0 0 0 mprj_io[28]
port 26 nsew signal bidirectional
flabel metal5 s 6598 613840 19088 626360 0 FreeSans 25000 0 0 0 mprj_io[29]
port 27 nsew signal bidirectional
flabel metal5 s 698512 191440 711002 203960 0 FreeSans 25000 0 0 0 mprj_io[2]
port 28 nsew signal bidirectional
flabel metal5 s 6598 570640 19088 583160 0 FreeSans 25000 0 0 0 mprj_io[30]
port 29 nsew signal bidirectional
flabel metal5 s 6598 527440 19088 539960 0 FreeSans 25000 0 0 0 mprj_io[31]
port 30 nsew signal bidirectional
flabel metal5 s 6598 399840 19088 412360 0 FreeSans 25000 0 0 0 mprj_io[32]
port 31 nsew signal bidirectional
flabel metal5 s 6598 356640 19088 369160 0 FreeSans 25000 0 0 0 mprj_io[33]
port 32 nsew signal bidirectional
flabel metal5 s 6598 313440 19088 325960 0 FreeSans 25000 0 0 0 mprj_io[34]
port 33 nsew signal bidirectional
flabel metal5 s 6598 270240 19088 282760 0 FreeSans 25000 0 0 0 mprj_io[35]
port 34 nsew signal bidirectional
flabel metal5 s 6598 227040 19088 239560 0 FreeSans 25000 0 0 0 mprj_io[36]
port 35 nsew signal bidirectional
flabel metal5 s 6598 183840 19088 196360 0 FreeSans 25000 0 0 0 mprj_io[37]
port 36 nsew signal bidirectional
flabel metal5 s 698512 236640 711002 249160 0 FreeSans 25000 0 0 0 mprj_io[3]
port 37 nsew signal bidirectional
flabel metal5 s 698512 281640 711002 294160 0 FreeSans 25000 0 0 0 mprj_io[4]
port 38 nsew signal bidirectional
flabel metal5 s 698512 326640 711002 339160 0 FreeSans 25000 0 0 0 mprj_io[5]
port 39 nsew signal bidirectional
flabel metal5 s 698512 371840 711002 384360 0 FreeSans 25000 0 0 0 mprj_io[6]
port 40 nsew signal bidirectional
flabel metal5 s 698512 549040 711002 561560 0 FreeSans 25000 0 0 0 mprj_io[7]
port 41 nsew signal bidirectional
flabel metal5 s 698512 594240 711002 606760 0 FreeSans 25000 0 0 0 mprj_io[8]
port 42 nsew signal bidirectional
flabel metal5 s 698512 639240 711002 651760 0 FreeSans 25000 0 0 0 mprj_io[9]
port 43 nsew signal bidirectional
flabel metal5 s 136713 7143 144150 18309 0 FreeSans 25000 0 0 0 resetb
port 44 nsew signal input
flabel metal5 s 6167 70054 19620 80934 0 FreeSans 25000 0 0 0 vccd
port 45 nsew signal bidirectional
flabel metal5 s 697980 909666 711433 920546 0 FreeSans 25000 0 0 0 vccd1
port 46 nsew signal bidirectional
flabel metal5 s 6167 914054 19620 924934 0 FreeSans 25000 0 0 0 vccd2
port 47 nsew signal bidirectional
flabel metal5 s 624222 6811 636390 18976 0 FreeSans 25000 0 0 0 vdda
port 48 nsew signal bidirectional
flabel metal5 s 698624 819822 710789 831990 0 FreeSans 25000 0 0 0 vdda1
port 49 nsew signal bidirectional
flabel metal5 s 698624 505222 710789 517390 0 FreeSans 25000 0 0 0 vdda1_2
port 50 nsew signal bidirectional
flabel metal5 s 6811 484410 18976 496578 0 FreeSans 25000 0 0 0 vdda2
port 51 nsew signal bidirectional
flabel metal5 s 6811 111610 18976 123778 0 FreeSans 25000 0 0 0 vddio
port 52 nsew signal bidirectional
flabel metal5 s 6811 871210 18976 883378 0 FreeSans 25000 0 0 0 vddio_2
port 53 nsew signal bidirectional
flabel metal5 s 80222 6811 92390 18976 0 FreeSans 25000 0 0 0 vssa
port 54 nsew signal bidirectional
flabel metal5 s 577010 1018624 589178 1030789 0 FreeSans 25000 0 0 0 vssa1
port 55 nsew signal bidirectional
flabel metal5 s 698624 417022 710789 429190 0 FreeSans 25000 0 0 0 vssa1_2
port 56 nsew signal bidirectional
flabel metal5 s 6811 829010 18976 841178 0 FreeSans 25000 0 0 0 vssa2
port 57 nsew signal bidirectional
flabel metal5 s 243266 6167 254146 19620 0 FreeSans 25000 0 0 0 vssd
port 58 nsew signal bidirectional
flabel metal5 s 697980 461866 711433 472746 0 FreeSans 25000 0 0 0 vssd1
port 59 nsew signal bidirectional
flabel metal5 s 6167 442854 19620 453734 0 FreeSans 25000 0 0 0 vssd2
port 60 nsew signal bidirectional
flabel metal5 s 570422 6811 582590 18976 0 FreeSans 25000 0 0 0 vssio
port 61 nsew signal bidirectional
flabel metal5 s 334810 1018624 346978 1030789 0 FreeSans 25000 0 0 0 vssio_2
port 62 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 0 0 717600 1037600
<< end >>
