magic
tech sky130A
magscale 36 1
timestamp 1598763267
<< metal5 >>
rect 0 100 35 105
rect 0 95 40 100
rect 0 85 45 95
rect 0 60 15 85
rect 30 60 45 85
rect 0 45 45 60
rect 0 20 15 45
rect 30 20 45 45
rect 0 10 45 20
rect 0 5 40 10
rect 0 0 35 5
<< properties >>
string FIXED_BBOX 0 -30 60 105
<< end >>
