VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO caravan_signal_routing
  CLASS BLOCK ;
  FOREIGN caravan_signal_routing ;
  ORIGIN 0.000 0.000 ;
  SIZE 1.000 BY 1.000 ;
  OBS
      LAYER met3 ;
        POLYGON 199.220 4710.300 199.220 4707.090 196.010 4707.090 ;
        RECT 199.220 4709.800 224.220 4778.310 ;
        RECT 199.220 4707.090 221.010 4709.800 ;
        RECT 196.010 4703.090 221.010 4707.090 ;
        POLYGON 221.010 4709.800 224.220 4709.800 221.010 4706.590 ;
        RECT 456.220 4707.090 481.220 4778.360 ;
        RECT 456.010 4706.410 481.220 4707.090 ;
        RECT 713.220 4707.090 738.220 4778.180 ;
        RECT 893.500 4756.600 964.895 4778.180 ;
        POLYGON 893.500 4756.600 943.010 4756.600 943.010 4707.090 ;
        RECT 943.010 4707.090 964.895 4756.600 ;
        RECT 966.395 4710.205 977.395 4778.180 ;
        POLYGON 966.395 4710.205 969.510 4710.205 969.510 4707.090 ;
        RECT 969.510 4707.090 977.395 4710.205 ;
        RECT 978.390 4710.710 989.390 4778.180 ;
        POLYGON 978.390 4710.710 980.260 4710.710 980.260 4708.840 ;
        RECT 980.260 4708.840 989.390 4710.710 ;
        RECT 990.890 4750.080 1062.500 4778.180 ;
        RECT 990.890 4710.710 1019.510 4750.080 ;
        POLYGON 990.890 4710.710 992.760 4710.710 992.760 4708.840 ;
        RECT 992.760 4708.840 1019.510 4710.710 ;
        POLYGON 977.395 4708.840 979.145 4707.090 977.395 4707.090 ;
        POLYGON 980.260 4708.840 982.010 4708.840 982.010 4707.090 ;
        RECT 982.010 4707.090 989.390 4708.840 ;
        POLYGON 989.390 4708.840 991.140 4707.090 989.390 4707.090 ;
        POLYGON 992.760 4708.840 994.510 4708.840 994.510 4707.090 ;
        RECT 713.220 4706.760 741.010 4707.090 ;
        RECT 456.010 4703.090 481.010 4706.410 ;
        RECT 716.010 4703.090 741.010 4706.760 ;
        RECT 943.010 4703.090 968.010 4707.090 ;
        RECT 969.510 4703.090 980.510 4707.090 ;
        RECT 982.010 4703.090 993.010 4707.090 ;
        RECT 994.510 4703.090 1019.510 4708.840 ;
        POLYGON 1019.510 4750.080 1062.500 4750.080 1019.510 4707.090 ;
        RECT 1156.500 4752.100 1227.895 4778.270 ;
        POLYGON 1156.500 4752.100 1201.510 4752.100 1201.510 4707.090 ;
        RECT 1201.510 4708.475 1227.895 4752.100 ;
        RECT 1201.510 4703.090 1226.510 4708.475 ;
        POLYGON 1226.510 4708.475 1227.895 4708.475 1226.510 4707.090 ;
        RECT 1229.395 4708.475 1240.395 4778.270 ;
        POLYGON 1229.395 4708.090 1229.395 4707.090 1228.395 4707.090 ;
        RECT 1229.395 4707.090 1239.010 4708.475 ;
        POLYGON 1239.010 4708.475 1240.395 4708.475 1239.010 4707.090 ;
        RECT 1241.390 4707.970 1252.390 4778.270 ;
        POLYGON 1241.390 4707.970 1241.390 4707.090 1240.510 4707.090 ;
        RECT 1241.390 4707.090 1251.510 4707.970 ;
        POLYGON 1251.510 4707.970 1252.390 4707.970 1251.510 4707.090 ;
        RECT 1253.890 4754.580 1325.500 4778.270 ;
        RECT 1253.890 4707.090 1278.010 4754.580 ;
        POLYGON 1278.010 4754.580 1325.500 4754.580 1278.010 4707.090 ;
        RECT 1665.500 4751.600 1736.895 4778.110 ;
        POLYGON 1665.500 4751.600 1710.010 4751.600 1710.010 4707.090 ;
        RECT 1710.010 4708.975 1736.895 4751.600 ;
        RECT 1228.010 4703.090 1239.010 4707.090 ;
        RECT 1240.510 4703.090 1251.510 4707.090 ;
        RECT 1253.010 4703.090 1278.010 4707.090 ;
        RECT 1710.010 4703.090 1735.010 4708.975 ;
        POLYGON 1735.010 4708.975 1736.895 4708.975 1735.010 4707.090 ;
        RECT 1738.395 4708.975 1749.395 4778.110 ;
        POLYGON 1738.395 4708.490 1738.395 4707.090 1736.995 4707.090 ;
        RECT 1738.395 4708.470 1748.890 4708.975 ;
        POLYGON 1748.890 4708.975 1749.395 4708.975 1748.890 4708.470 ;
        RECT 1750.390 4708.470 1761.390 4778.110 ;
        RECT 1738.395 4707.090 1747.510 4708.470 ;
        POLYGON 1747.510 4708.470 1748.890 4708.470 1747.510 4707.090 ;
        POLYGON 1750.390 4708.470 1750.390 4707.090 1749.010 4707.090 ;
        RECT 1750.390 4707.090 1760.010 4708.470 ;
        POLYGON 1760.010 4708.470 1761.390 4708.470 1760.010 4707.090 ;
        RECT 1762.890 4755.080 1834.500 4778.110 ;
        RECT 1762.890 4707.090 1786.510 4755.080 ;
        POLYGON 1786.510 4755.080 1834.500 4755.080 1786.510 4707.090 ;
        RECT 2182.220 4707.090 2207.220 4778.020 ;
        RECT 1736.510 4703.090 1747.510 4707.090 ;
        RECT 1749.010 4703.090 1760.010 4707.090 ;
        RECT 1761.510 4703.090 1786.510 4707.090 ;
        RECT 2182.010 4706.420 2207.220 4707.090 ;
        RECT 2439.220 4709.820 2464.220 4778.460 ;
        POLYGON 2439.220 4709.820 2442.010 4709.820 2442.010 4707.030 ;
        RECT 2442.010 4707.090 2464.220 4709.820 ;
        POLYGON 2464.220 4709.880 2467.010 4707.090 2464.220 4707.090 ;
        RECT 2182.010 4703.090 2207.010 4706.420 ;
        RECT 2442.010 4703.090 2467.010 4707.090 ;
        RECT 2667.000 4707.890 2690.895 4777.960 ;
        POLYGON 2667.000 4707.890 2668.010 4707.890 2668.010 4706.880 ;
        RECT 2668.010 4707.090 2690.895 4707.890 ;
        POLYGON 2690.895 4708.205 2692.010 4707.090 2690.895 4707.090 ;
        RECT 2668.010 4703.090 2692.010 4707.090 ;
        RECT 2716.890 4708.000 2740.790 4777.960 ;
        POLYGON 2716.890 4708.000 2718.010 4708.000 2718.010 4706.880 ;
        RECT 2718.010 4707.090 2740.790 4708.000 ;
        POLYGON 2740.790 4708.310 2742.010 4707.090 2740.790 4707.090 ;
        RECT 2948.220 4707.090 2973.220 4778.730 ;
        RECT 2718.010 4703.090 2742.010 4707.090 ;
        RECT 2948.010 4706.370 2973.220 4707.090 ;
        RECT 2948.010 4703.090 2973.010 4706.370 ;
        RECT -12.680 4609.300 105.820 4615.220 ;
        POLYGON 105.820 4615.220 111.740 4609.300 105.820 4609.300 ;
        RECT -12.680 4590.220 115.040 4609.300 ;
        POLYGON 105.125 4590.220 111.040 4590.220 111.040 4584.305 ;
        RECT 111.040 4584.300 115.040 4590.220 ;
        RECT 3035.040 4597.780 3039.040 4598.010 ;
        RECT 3035.040 4573.010 3177.530 4597.780 ;
        RECT 3038.580 4572.780 3177.530 4573.010 ;
        RECT 111.040 4424.200 115.040 4426.300 ;
        RECT -6.220 4402.300 115.040 4424.200 ;
        RECT -6.220 4400.255 111.260 4402.300 ;
        RECT 3035.040 4402.010 3039.040 4406.010 ;
        POLYGON 3039.040 4406.010 3043.040 4402.010 3039.040 4402.010 ;
        RECT 3035.040 4382.010 3170.900 4402.010 ;
        POLYGON 3038.130 4382.010 3042.140 4382.010 3042.140 4378.000 ;
        RECT 3042.140 4378.000 3170.900 4382.010 ;
        RECT 111.040 4374.000 115.040 4376.305 ;
        RECT -6.220 4352.300 115.040 4374.000 ;
        RECT -6.220 4350.000 111.300 4352.300 ;
        RECT 3035.040 4351.745 3039.040 4356.010 ;
        POLYGON 3039.040 4356.010 3043.305 4351.745 3039.040 4351.745 ;
        RECT 3035.040 4332.010 3170.900 4351.745 ;
        POLYGON 3038.170 4332.010 3042.380 4332.010 3042.380 4327.800 ;
        RECT 3042.380 4327.800 3170.900 4332.010 ;
        POLYGON 111.040 4004.300 111.040 4001.790 108.530 4001.790 ;
        RECT 111.040 4001.790 115.040 4004.300 ;
        RECT -12.000 3980.300 115.040 4001.790 ;
        RECT -12.000 3977.890 109.260 3980.300 ;
        POLYGON 109.260 3980.300 111.670 3980.300 109.260 3977.890 ;
        RECT 3035.040 3956.005 3039.040 3959.900 ;
        POLYGON 111.040 3954.300 111.040 3951.895 108.635 3951.895 ;
        RECT 111.040 3951.895 115.040 3954.300 ;
        RECT -12.000 3930.300 115.040 3951.895 ;
        RECT 3035.040 3935.900 3176.660 3956.005 ;
        RECT 3037.790 3932.105 3176.660 3935.900 ;
        RECT 37.960 3930.295 111.670 3930.300 ;
        RECT -12.000 3927.995 109.370 3930.295 ;
        POLYGON 109.370 3930.295 111.670 3930.295 109.370 3927.995 ;
        RECT 3035.040 3906.110 3039.040 3909.900 ;
        RECT 3035.040 3885.900 3176.660 3906.110 ;
        RECT 3037.790 3882.210 3176.660 3885.900 ;
        RECT 3035.040 2383.005 3039.040 2383.240 ;
        RECT 3035.040 2359.240 3176.660 2383.005 ;
        RECT 3038.790 2359.105 3124.080 2359.240 ;
        RECT 3035.040 2333.110 3039.040 2333.240 ;
        RECT 3035.040 2309.240 3176.660 2333.110 ;
        RECT 3038.830 2309.210 3124.120 2309.240 ;
        POLYGON 111.040 2281.530 111.040 2278.790 108.300 2278.790 ;
        RECT 111.040 2278.790 115.040 2281.530 ;
        RECT -12.000 2257.530 115.040 2278.790 ;
        RECT -12.000 2254.890 108.560 2257.530 ;
        POLYGON 108.560 2257.530 111.200 2257.530 108.560 2254.890 ;
        POLYGON 111.040 2231.525 111.040 2228.895 108.410 2228.895 ;
        RECT 111.040 2228.895 115.040 2231.530 ;
        RECT -12.000 2207.530 115.040 2228.895 ;
        RECT -12.000 2204.995 108.705 2207.530 ;
        POLYGON 108.705 2207.530 111.240 2207.530 108.705 2204.995 ;
        RECT 3035.040 2163.000 3039.040 2164.240 ;
        RECT 3035.040 2140.240 3169.390 2163.000 ;
        RECT 3038.710 2139.000 3169.390 2140.240 ;
        RECT 3035.040 2112.745 3039.040 2114.240 ;
        RECT 3035.040 2090.240 3169.390 2112.745 ;
        RECT 3038.710 2088.800 3169.390 2090.240 ;
        POLYGON 111.040 2071.530 111.040 2068.200 107.710 2068.200 ;
        RECT 111.040 2068.200 115.040 2071.530 ;
        RECT -4.500 2047.530 115.040 2068.200 ;
        RECT -4.500 2044.255 108.135 2047.530 ;
        POLYGON 108.135 2047.530 111.410 2047.530 108.135 2044.255 ;
        POLYGON 111.040 2021.530 111.040 2018.000 107.510 2018.000 ;
        RECT 111.040 2018.000 115.040 2021.530 ;
        RECT -4.500 1997.530 115.040 2018.000 ;
        RECT -4.500 1994.000 107.790 1997.530 ;
        POLYGON 107.790 1997.530 111.320 1997.530 107.790 1994.000 ;
        RECT 3038.840 1941.240 3176.880 1942.005 ;
        RECT 3035.040 1918.105 3176.880 1941.240 ;
        RECT 3035.040 1917.310 3173.620 1918.105 ;
        RECT 3035.040 1917.240 3039.040 1917.310 ;
        RECT 3038.790 1891.240 3176.880 1892.110 ;
        RECT 3035.040 1868.210 3176.880 1891.240 ;
        RECT 3035.040 1867.240 3039.040 1868.210 ;
      LAYER via3 ;
        RECT 895.635 4758.740 962.755 4767.460 ;
        RECT 993.025 4758.740 1060.145 4767.460 ;
        RECT 1158.635 4758.740 1225.755 4767.460 ;
        RECT 1256.025 4758.740 1323.145 4767.460 ;
        RECT 1667.635 4758.740 1734.755 4767.460 ;
        RECT 1765.025 4758.740 1832.145 4767.460 ;
        RECT 2667.925 4711.955 2689.845 4723.475 ;
        RECT 2717.925 4711.955 2739.845 4723.475 ;
        RECT 91.780 3979.040 103.300 4000.960 ;
        RECT 91.780 3929.040 103.300 3950.960 ;
        RECT 3068.125 3933.255 3079.645 3955.175 ;
        RECT 3068.125 3883.255 3079.645 3905.175 ;
        RECT 3068.125 2360.255 3079.645 2382.175 ;
        RECT 3068.125 2310.255 3079.645 2332.175 ;
        RECT 67.780 2256.040 79.300 2277.960 ;
        RECT 67.780 2206.040 79.300 2227.960 ;
        RECT 3044.125 1919.255 3055.645 1941.175 ;
        RECT 3044.125 1869.255 3055.645 1891.175 ;
      LAYER met4 ;
        RECT 893.500 4756.600 964.895 4769.600 ;
        POLYGON 893.500 4756.600 943.010 4756.600 943.010 4707.090 ;
        RECT 943.010 4707.090 964.895 4756.600 ;
        RECT 990.890 4758.600 1062.285 4769.600 ;
        RECT 990.890 4750.080 1062.500 4758.600 ;
        RECT 990.890 4710.710 1019.510 4750.080 ;
        POLYGON 990.890 4710.710 994.510 4710.710 994.510 4707.090 ;
        RECT 943.010 4703.090 968.010 4707.090 ;
        RECT 994.510 4703.090 1019.510 4710.710 ;
        POLYGON 1019.510 4750.080 1062.500 4750.080 1019.510 4707.090 ;
        RECT 1156.500 4752.100 1227.895 4769.600 ;
        POLYGON 1156.500 4752.100 1201.510 4752.100 1201.510 4707.090 ;
        RECT 1201.510 4708.475 1227.895 4752.100 ;
        RECT 1201.510 4703.090 1226.510 4708.475 ;
        POLYGON 1226.510 4708.475 1227.895 4708.475 1226.510 4707.090 ;
        RECT 1253.890 4758.600 1325.285 4769.600 ;
        RECT 1253.890 4754.580 1325.500 4758.600 ;
        RECT 1253.890 4707.090 1278.010 4754.580 ;
        POLYGON 1278.010 4754.580 1325.500 4754.580 1278.010 4707.090 ;
        RECT 1665.500 4751.600 1736.895 4769.600 ;
        POLYGON 1665.500 4751.600 1710.010 4751.600 1710.010 4707.090 ;
        RECT 1710.010 4708.975 1736.895 4751.600 ;
        RECT 1253.010 4703.090 1278.010 4707.090 ;
        RECT 1710.010 4703.090 1735.010 4708.975 ;
        POLYGON 1735.010 4708.975 1736.895 4708.975 1735.010 4707.090 ;
        RECT 1762.890 4758.600 1834.285 4769.600 ;
        RECT 1762.890 4755.080 1834.500 4758.600 ;
        RECT 1762.890 4707.090 1786.510 4755.080 ;
        POLYGON 1786.510 4755.080 1834.500 4755.080 1786.510 4707.090 ;
        RECT 2667.005 4711.410 2690.895 4724.420 ;
        RECT 2716.890 4711.410 2740.790 4724.405 ;
        RECT 1761.510 4703.090 1786.510 4707.090 ;
        RECT 90.955 3977.890 103.955 4001.790 ;
        RECT 90.955 3927.995 103.955 3951.895 ;
        RECT 3067.300 3932.105 3080.300 3956.005 ;
        RECT 3067.300 3882.210 3080.300 3906.110 ;
        RECT 3067.300 2359.105 3080.300 2383.005 ;
        RECT 3067.300 2309.210 3080.300 2333.110 ;
        RECT 66.955 2254.890 79.955 2278.790 ;
        RECT 66.955 2204.995 79.955 2228.895 ;
        RECT 3043.300 1917.310 3056.300 1942.005 ;
        RECT 3043.300 1868.210 3056.300 1892.110 ;
        RECT 66.950 1144.180 79.950 1218.290 ;
        RECT 3043.300 1132.580 3056.300 1218.290 ;
        RECT 3067.300 1120.980 3080.300 1218.290 ;
      LAYER met5 ;
        RECT 893.500 4756.600 964.895 4769.600 ;
        POLYGON 893.500 4756.600 943.010 4756.600 943.010 4707.090 ;
        RECT 943.010 4707.090 964.895 4756.600 ;
        RECT 990.890 4758.600 1062.285 4769.600 ;
        RECT 990.890 4750.080 1062.500 4758.600 ;
        RECT 990.890 4710.710 1019.510 4750.080 ;
        POLYGON 990.890 4710.710 994.510 4710.710 994.510 4707.090 ;
        RECT 943.010 4703.090 968.010 4707.090 ;
        RECT 994.510 4703.090 1019.510 4710.710 ;
        POLYGON 1019.510 4750.080 1062.500 4750.080 1019.510 4707.090 ;
        RECT 1156.500 4752.100 1227.895 4769.600 ;
        POLYGON 1156.500 4752.100 1201.510 4752.100 1201.510 4707.090 ;
        RECT 1201.510 4708.475 1227.895 4752.100 ;
        RECT 1201.510 4703.090 1226.510 4708.475 ;
        POLYGON 1226.510 4708.475 1227.895 4708.475 1226.510 4707.090 ;
        RECT 1253.890 4758.600 1325.285 4769.600 ;
        RECT 1253.890 4754.580 1325.500 4758.600 ;
        RECT 1253.890 4707.090 1278.010 4754.580 ;
        POLYGON 1278.010 4754.580 1325.500 4754.580 1278.010 4707.090 ;
        RECT 1665.500 4751.600 1736.895 4769.600 ;
        POLYGON 1665.500 4751.600 1710.010 4751.600 1710.010 4707.090 ;
        RECT 1710.010 4708.975 1736.895 4751.600 ;
        RECT 1253.010 4703.090 1278.010 4707.090 ;
        RECT 1710.010 4703.090 1735.010 4708.975 ;
        POLYGON 1735.010 4708.975 1736.895 4708.975 1735.010 4707.090 ;
        RECT 1762.890 4758.600 1834.285 4769.600 ;
        RECT 1762.890 4755.080 1834.500 4758.600 ;
        RECT 1762.890 4707.090 1786.510 4755.080 ;
        POLYGON 1786.510 4755.080 1834.500 4755.080 1786.510 4707.090 ;
        RECT 2667.000 4711.410 3056.300 4724.410 ;
        RECT 1761.510 4703.090 1786.510 4707.090 ;
        RECT 66.955 1195.000 79.955 2278.790 ;
        RECT 3043.300 1195.000 3056.300 4711.410 ;
        RECT 3067.300 1195.000 3080.300 3956.005 ;
  END
END caravan_signal_routing
END LIBRARY

