magic
tech sky130A
magscale 1 2
timestamp 1666101174
<< viali >>
rect 3893 13481 3927 13515
rect 7849 13413 7883 13447
rect 13737 13413 13771 13447
rect 14749 13345 14783 13379
rect 16221 13345 16255 13379
rect 18061 13345 18095 13379
rect 2881 13277 2915 13311
rect 3525 13277 3559 13311
rect 4813 13277 4847 13311
rect 6469 13277 6503 13311
rect 6745 13277 6779 13311
rect 8033 13277 8067 13311
rect 9137 13277 9171 13311
rect 10149 13277 10183 13311
rect 11805 13277 11839 13311
rect 12449 13277 12483 13311
rect 13277 13277 13311 13311
rect 14197 13277 14231 13311
rect 15209 13277 15243 13311
rect 15669 13277 15703 13311
rect 16129 13277 16163 13311
rect 16773 13277 16807 13311
rect 3433 13209 3467 13243
rect 4261 13209 4295 13243
rect 4353 13209 4387 13243
rect 5549 13209 5583 13243
rect 6929 13209 6963 13243
rect 7481 13209 7515 13243
rect 8677 13209 8711 13243
rect 9597 13209 9631 13243
rect 9689 13209 9723 13243
rect 10977 13209 11011 13243
rect 12265 13209 12299 13243
rect 12725 13209 12759 13243
rect 13829 13209 13863 13243
rect 14657 13209 14691 13243
rect 17233 13209 17267 13243
rect 17325 13209 17359 13243
rect 17601 13209 17635 13243
rect 2237 13141 2271 13175
rect 2329 13141 2363 13175
rect 2697 13141 2731 13175
rect 5181 13141 5215 13175
rect 5641 13141 5675 13175
rect 6101 13141 6135 13175
rect 6561 13141 6595 13175
rect 7389 13141 7423 13175
rect 8585 13141 8619 13175
rect 9965 13141 9999 13175
rect 10609 13141 10643 13175
rect 10701 13141 10735 13175
rect 11621 13141 11655 13175
rect 12633 13141 12667 13175
rect 15025 13141 15059 13175
rect 15761 13141 15795 13175
rect 17785 13141 17819 13175
rect 14381 12937 14415 12971
rect 2329 12869 2363 12903
rect 4997 12869 5031 12903
rect 7205 12869 7239 12903
rect 9965 12869 9999 12903
rect 10701 12869 10735 12903
rect 11805 12869 11839 12903
rect 13829 12869 13863 12903
rect 14473 12869 14507 12903
rect 17969 12869 18003 12903
rect 1685 12801 1719 12835
rect 2605 12801 2639 12835
rect 3617 12801 3651 12835
rect 4537 12801 4571 12835
rect 4813 12801 4847 12835
rect 5733 12801 5767 12835
rect 6101 12801 6135 12835
rect 7481 12801 7515 12835
rect 8401 12801 8435 12835
rect 9321 12801 9355 12835
rect 10241 12801 10275 12835
rect 10793 12801 10827 12835
rect 11621 12801 11655 12835
rect 12541 12801 12575 12835
rect 13093 12801 13127 12835
rect 14013 12801 14047 12835
rect 14841 12801 14875 12835
rect 15761 12801 15795 12835
rect 17049 12801 17083 12835
rect 17785 12801 17819 12835
rect 18429 12801 18463 12835
rect 6653 12733 6687 12767
rect 11253 12733 11287 12767
rect 3249 12665 3283 12699
rect 7113 12665 7147 12699
rect 8953 12665 8987 12699
rect 16129 12665 16163 12699
rect 18245 12597 18279 12631
rect 3433 12393 3467 12427
rect 4353 12393 4387 12427
rect 9229 12393 9263 12427
rect 11621 12393 11655 12427
rect 13001 12393 13035 12427
rect 17141 12393 17175 12427
rect 2237 12325 2271 12359
rect 3157 12325 3191 12359
rect 4905 12325 4939 12359
rect 7573 12325 7607 12359
rect 10241 12325 10275 12359
rect 15485 12325 15519 12359
rect 17969 12325 18003 12359
rect 1777 12257 1811 12291
rect 2329 12257 2363 12291
rect 4813 12257 4847 12291
rect 8125 12257 8159 12291
rect 8677 12257 8711 12291
rect 9781 12257 9815 12291
rect 17509 12257 17543 12291
rect 18061 12257 18095 12291
rect 3893 12189 3927 12223
rect 4169 12189 4203 12223
rect 5365 12189 5399 12223
rect 6009 12189 6043 12223
rect 6285 12189 6319 12223
rect 7757 12189 7791 12223
rect 9459 12189 9493 12223
rect 10420 12189 10454 12223
rect 10609 12189 10643 12223
rect 10793 12189 10827 12223
rect 11069 12189 11103 12223
rect 11253 12189 11287 12223
rect 11489 12189 11523 12223
rect 12449 12189 12483 12223
rect 12725 12189 12759 12223
rect 12869 12189 12903 12223
rect 13461 12189 13495 12223
rect 13645 12189 13679 12223
rect 14197 12189 14231 12223
rect 15393 12189 15427 12223
rect 16221 12189 16255 12223
rect 16957 12189 16991 12223
rect 18337 12189 18371 12223
rect 2973 12121 3007 12155
rect 8585 12121 8619 12155
rect 9229 12121 9263 12155
rect 10517 12121 10551 12155
rect 11342 12121 11376 12155
rect 12633 12121 12667 12155
rect 16681 12121 16715 12155
rect 3985 12053 4019 12087
rect 5825 12053 5859 12087
rect 9597 12053 9631 12087
rect 9689 12053 9723 12087
rect 11989 12053 12023 12087
rect 13645 12053 13679 12087
rect 16313 12053 16347 12087
rect 16773 12053 16807 12087
rect 2973 11849 3007 11883
rect 5641 11849 5675 11883
rect 6929 11849 6963 11883
rect 9137 11849 9171 11883
rect 9505 11849 9539 11883
rect 9781 11849 9815 11883
rect 10885 11849 10919 11883
rect 13277 11849 13311 11883
rect 15393 11849 15427 11883
rect 2329 11781 2363 11815
rect 3433 11781 3467 11815
rect 5273 11781 5307 11815
rect 6009 11781 6043 11815
rect 6561 11781 6595 11815
rect 7757 11781 7791 11815
rect 8585 11781 8619 11815
rect 11897 11781 11931 11815
rect 13093 11781 13127 11815
rect 13921 11781 13955 11815
rect 14289 11781 14323 11815
rect 15025 11781 15059 11815
rect 3065 11713 3099 11747
rect 3525 11713 3559 11747
rect 3709 11713 3743 11747
rect 4813 11713 4847 11747
rect 5089 11713 5123 11747
rect 5549 11713 5583 11747
rect 5825 11713 5859 11747
rect 7113 11713 7147 11747
rect 7389 11713 7423 11747
rect 8309 11713 8343 11747
rect 8493 11713 8527 11747
rect 10057 11713 10091 11747
rect 10241 11713 10275 11747
rect 10701 11713 10735 11747
rect 11621 11713 11655 11747
rect 11805 11713 11839 11747
rect 11994 11713 12028 11747
rect 12541 11713 12575 11747
rect 13553 11713 13587 11747
rect 14105 11713 14139 11747
rect 14381 11713 14415 11747
rect 15281 11713 15315 11747
rect 16221 11713 16255 11747
rect 16865 11713 16899 11747
rect 17785 11713 17819 11747
rect 1777 11645 1811 11679
rect 3893 11645 3927 11679
rect 4261 11645 4295 11679
rect 8125 11645 8159 11679
rect 9689 11645 9723 11679
rect 9965 11645 9999 11679
rect 10517 11645 10551 11679
rect 15485 11645 15519 11679
rect 15577 11645 15611 11679
rect 2237 11577 2271 11611
rect 4721 11577 4755 11611
rect 7297 11577 7331 11611
rect 12173 11577 12207 11611
rect 14841 11577 14875 11611
rect 15853 11577 15887 11611
rect 18153 11577 18187 11611
rect 12633 11509 12667 11543
rect 13277 11509 13311 11543
rect 16405 11509 16439 11543
rect 3433 11305 3467 11339
rect 7113 11305 7147 11339
rect 13737 11305 13771 11339
rect 15301 11305 15335 11339
rect 2789 11237 2823 11271
rect 5181 11237 5215 11271
rect 8677 11237 8711 11271
rect 10057 11237 10091 11271
rect 10609 11237 10643 11271
rect 14933 11237 14967 11271
rect 17969 11237 18003 11271
rect 7573 11169 7607 11203
rect 7665 11169 7699 11203
rect 11069 11169 11103 11203
rect 11529 11169 11563 11203
rect 12541 11169 12575 11203
rect 13277 11169 13311 11203
rect 14565 11169 14599 11203
rect 17141 11169 17175 11203
rect 17693 11169 17727 11203
rect 1501 11101 1535 11135
rect 2973 11101 3007 11135
rect 3893 11101 3927 11135
rect 5365 11101 5399 11135
rect 5917 11101 5951 11135
rect 6653 11101 6687 11135
rect 7369 11101 7403 11135
rect 8033 11101 8067 11135
rect 8217 11101 8251 11135
rect 8322 11079 8356 11113
rect 8435 11101 8469 11135
rect 9287 11101 9321 11135
rect 9413 11101 9447 11135
rect 9504 11101 9538 11135
rect 9689 11101 9723 11135
rect 10425 11101 10459 11135
rect 10609 11101 10643 11135
rect 10977 11101 11011 11135
rect 11253 11101 11287 11135
rect 11345 11101 11379 11135
rect 11897 11101 11931 11135
rect 12081 11101 12115 11135
rect 12173 11101 12207 11135
rect 12299 11101 12333 11135
rect 13185 11101 13219 11135
rect 13461 11101 13495 11135
rect 13553 11101 13587 11135
rect 14197 11101 14231 11135
rect 14362 11101 14396 11135
rect 14473 11101 14507 11135
rect 14749 11101 14783 11135
rect 15209 11101 15243 11135
rect 15393 11101 15427 11135
rect 15945 11101 15979 11135
rect 16681 11101 16715 11135
rect 17233 11101 17267 11135
rect 18153 11101 18187 11135
rect 5733 11033 5767 11067
rect 7113 11033 7147 11067
rect 9045 11033 9079 11067
rect 16865 11033 16899 11067
rect 7481 10965 7515 10999
rect 12817 10965 12851 10999
rect 8493 10761 8527 10795
rect 15209 10761 15243 10795
rect 15301 10761 15335 10795
rect 16405 10761 16439 10795
rect 1869 10693 1903 10727
rect 2329 10693 2363 10727
rect 2605 10693 2639 10727
rect 4905 10693 4939 10727
rect 5089 10693 5123 10727
rect 5549 10693 5583 10727
rect 6745 10693 6779 10727
rect 10793 10693 10827 10727
rect 12541 10693 12575 10727
rect 13461 10693 13495 10727
rect 14289 10693 14323 10727
rect 14473 10693 14507 10727
rect 15853 10693 15887 10727
rect 17509 10693 17543 10727
rect 18245 10693 18279 10727
rect 2053 10625 2087 10659
rect 2237 10625 2271 10659
rect 3709 10625 3743 10659
rect 4077 10625 4111 10659
rect 5641 10625 5675 10659
rect 6101 10625 6135 10659
rect 7297 10625 7331 10659
rect 7481 10625 7515 10659
rect 7573 10625 7607 10659
rect 8033 10625 8067 10659
rect 8325 10625 8359 10659
rect 8953 10625 8987 10659
rect 9137 10625 9171 10659
rect 9321 10625 9355 10659
rect 10517 10625 10551 10659
rect 10701 10625 10735 10659
rect 10937 10625 10971 10659
rect 11989 10625 12023 10659
rect 12173 10625 12207 10659
rect 12633 10625 12667 10659
rect 12817 10625 12851 10659
rect 13277 10625 13311 10659
rect 14749 10625 14783 10659
rect 15117 10625 15151 10659
rect 15439 10625 15473 10659
rect 15669 10625 15703 10659
rect 16313 10625 16347 10659
rect 18337 10625 18371 10659
rect 3985 10557 4019 10591
rect 4537 10557 4571 10591
rect 10149 10557 10183 10591
rect 13553 10557 13587 10591
rect 16957 10557 16991 10591
rect 17785 10557 17819 10591
rect 8125 10489 8159 10523
rect 9781 10489 9815 10523
rect 11069 10489 11103 10523
rect 12173 10489 12207 10523
rect 17417 10489 17451 10523
rect 3157 10421 3191 10455
rect 3617 10421 3651 10455
rect 7113 10421 7147 10455
rect 9689 10421 9723 10455
rect 14473 10421 14507 10455
rect 5089 10217 5123 10251
rect 11897 10217 11931 10251
rect 12081 10217 12115 10251
rect 14289 10217 14323 10251
rect 18061 10217 18095 10251
rect 3433 10149 3467 10183
rect 7205 10149 7239 10183
rect 3525 10081 3559 10115
rect 6469 10081 6503 10115
rect 7941 10081 7975 10115
rect 8401 10081 8435 10115
rect 10057 10081 10091 10115
rect 15393 10081 15427 10115
rect 2421 10013 2455 10047
rect 2605 10013 2639 10047
rect 2973 10013 3007 10047
rect 4077 10013 4111 10047
rect 4813 10013 4847 10047
rect 5273 10013 5307 10047
rect 5825 10013 5859 10047
rect 6101 10013 6135 10047
rect 6377 10013 6411 10047
rect 7021 10013 7055 10047
rect 8107 10013 8141 10047
rect 8217 10013 8251 10047
rect 8493 10013 8527 10047
rect 9229 10013 9263 10047
rect 9413 10013 9447 10047
rect 9873 10013 9907 10047
rect 10701 10013 10735 10047
rect 10885 10013 10919 10047
rect 11161 10013 11195 10047
rect 11345 10013 11379 10047
rect 11437 10013 11471 10047
rect 12725 10013 12759 10047
rect 13093 10013 13127 10047
rect 13277 10013 13311 10047
rect 13461 10013 13495 10047
rect 14473 10013 14507 10047
rect 14565 10013 14599 10047
rect 14749 10013 14783 10047
rect 14841 10013 14875 10047
rect 15117 10013 15151 10047
rect 15301 10013 15335 10047
rect 15669 10013 15703 10047
rect 16037 10013 16071 10047
rect 16773 10013 16807 10047
rect 17693 10013 17727 10047
rect 18153 10013 18187 10047
rect 2145 9945 2179 9979
rect 3893 9945 3927 9979
rect 6745 9945 6779 9979
rect 9045 9945 9079 9979
rect 10149 9945 10183 9979
rect 10241 9945 10275 9979
rect 12265 9945 12299 9979
rect 17417 9945 17451 9979
rect 1777 9877 1811 9911
rect 2237 9877 2271 9911
rect 5641 9877 5675 9911
rect 6837 9877 6871 9911
rect 10609 9877 10643 9911
rect 12081 9877 12115 9911
rect 12633 9877 12667 9911
rect 13829 9877 13863 9911
rect 16221 9877 16255 9911
rect 11161 9673 11195 9707
rect 9137 9605 9171 9639
rect 10158 9605 10192 9639
rect 15301 9605 15335 9639
rect 16405 9605 16439 9639
rect 16865 9605 16899 9639
rect 17233 9605 17267 9639
rect 2237 9537 2271 9571
rect 2789 9537 2823 9571
rect 4261 9537 4295 9571
rect 5089 9537 5123 9571
rect 5641 9537 5675 9571
rect 6101 9537 6135 9571
rect 6469 9537 6503 9571
rect 7113 9537 7147 9571
rect 7297 9537 7331 9571
rect 7389 9537 7423 9571
rect 8033 9537 8067 9571
rect 8309 9537 8343 9571
rect 8493 9537 8527 9571
rect 9321 9537 9355 9571
rect 9505 9537 9539 9571
rect 9781 9537 9815 9571
rect 10425 9537 10459 9571
rect 10793 9537 10827 9571
rect 10977 9537 11011 9571
rect 11713 9537 11747 9571
rect 11989 9537 12023 9571
rect 12449 9537 12483 9571
rect 13001 9537 13035 9571
rect 13185 9537 13219 9571
rect 13645 9537 13679 9571
rect 14289 9537 14323 9571
rect 14381 9537 14415 9571
rect 14565 9537 14599 9571
rect 15209 9537 15243 9571
rect 15393 9537 15427 9571
rect 15669 9537 15703 9571
rect 17049 9537 17083 9571
rect 17325 9537 17359 9571
rect 6009 9469 6043 9503
rect 7941 9469 7975 9503
rect 11621 9469 11655 9503
rect 12265 9469 12299 9503
rect 13369 9469 13403 9503
rect 17601 9469 17635 9503
rect 18153 9469 18187 9503
rect 4077 9401 4111 9435
rect 7205 9401 7239 9435
rect 12633 9401 12667 9435
rect 14473 9401 14507 9435
rect 16313 9401 16347 9435
rect 18061 9401 18095 9435
rect 2053 9333 2087 9367
rect 4905 9333 4939 9367
rect 6653 9333 6687 9367
rect 7573 9333 7607 9367
rect 8769 9333 8803 9367
rect 10149 9333 10183 9367
rect 13737 9333 13771 9367
rect 3525 9129 3559 9163
rect 10517 9129 10551 9163
rect 11713 9129 11747 9163
rect 5089 9061 5123 9095
rect 9597 9061 9631 9095
rect 12173 9061 12207 9095
rect 14381 9061 14415 9095
rect 14749 9061 14783 9095
rect 15669 9061 15703 9095
rect 18153 9061 18187 9095
rect 3985 8993 4019 9027
rect 5733 8993 5767 9027
rect 6193 8993 6227 9027
rect 7113 8993 7147 9027
rect 2053 8925 2087 8959
rect 4905 8925 4939 8959
rect 6009 8925 6043 8959
rect 6837 8925 6871 8959
rect 7205 8925 7239 8959
rect 7481 8925 7515 8959
rect 7757 8925 7791 8959
rect 8033 8925 8067 8959
rect 8493 8925 8527 8959
rect 9413 8925 9447 8959
rect 9597 8925 9631 8959
rect 10701 8925 10735 8959
rect 10792 8925 10826 8959
rect 10948 8925 10982 8959
rect 11081 8925 11115 8959
rect 11805 8925 11839 8959
rect 12173 8925 12207 8959
rect 12357 8925 12391 8959
rect 13093 8925 13127 8959
rect 13185 8925 13219 8959
rect 13277 8925 13311 8959
rect 13369 8925 13403 8959
rect 14289 8925 14323 8959
rect 14473 8925 14507 8959
rect 14565 8925 14599 8959
rect 15117 8925 15151 8959
rect 15537 8925 15571 8959
rect 16037 8925 16071 8959
rect 16681 8925 16715 8959
rect 17693 8925 17727 8959
rect 1501 8857 1535 8891
rect 4445 8857 4479 8891
rect 4537 8857 4571 8891
rect 5641 8857 5675 8891
rect 9965 8857 9999 8891
rect 15301 8857 15335 8891
rect 15393 8857 15427 8891
rect 6653 8789 6687 8823
rect 7849 8789 7883 8823
rect 8585 8789 8619 8823
rect 13553 8789 13587 8823
rect 6653 8585 6687 8619
rect 7757 8585 7791 8619
rect 12817 8585 12851 8619
rect 4169 8517 4203 8551
rect 4445 8517 4479 8551
rect 5733 8517 5767 8551
rect 10885 8517 10919 8551
rect 14381 8517 14415 8551
rect 15393 8517 15427 8551
rect 15485 8517 15519 8551
rect 17969 8517 18003 8551
rect 2605 8449 2639 8483
rect 4077 8449 4111 8483
rect 4629 8449 4663 8483
rect 5365 8449 5399 8483
rect 5825 8449 5859 8483
rect 6009 8449 6043 8483
rect 6469 8449 6503 8483
rect 7113 8449 7147 8483
rect 7297 8449 7331 8483
rect 8309 8449 8343 8483
rect 8493 8449 8527 8483
rect 9045 8449 9079 8483
rect 9321 8449 9355 8483
rect 9597 8449 9631 8483
rect 9781 8449 9815 8483
rect 10057 8449 10091 8483
rect 10333 8449 10367 8483
rect 10425 8449 10459 8483
rect 11161 8449 11195 8483
rect 11897 8449 11931 8483
rect 12357 8449 12391 8483
rect 13368 8471 13402 8505
rect 13460 8439 13494 8473
rect 13553 8449 13587 8483
rect 13737 8449 13771 8483
rect 14105 8449 14139 8483
rect 14197 8449 14231 8483
rect 14933 8449 14967 8483
rect 15209 8449 15243 8483
rect 15629 8449 15663 8483
rect 16313 8449 16347 8483
rect 7481 8381 7515 8415
rect 8125 8381 8159 8415
rect 16768 8381 16802 8415
rect 17325 8381 17359 8415
rect 11713 8313 11747 8347
rect 13093 8313 13127 8347
rect 14749 8313 14783 8347
rect 15761 8313 15795 8347
rect 17233 8313 17267 8347
rect 18429 8313 18463 8347
rect 1869 8245 1903 8279
rect 9229 8245 9263 8279
rect 12265 8245 12299 8279
rect 16221 8245 16255 8279
rect 17877 8245 17911 8279
rect 5457 8041 5491 8075
rect 5917 8041 5951 8075
rect 10057 8041 10091 8075
rect 10609 8041 10643 8075
rect 11621 8041 11655 8075
rect 13829 8041 13863 8075
rect 4629 7973 4663 8007
rect 11805 7973 11839 8007
rect 14197 7973 14231 8007
rect 16497 7973 16531 8007
rect 18153 7973 18187 8007
rect 6377 7905 6411 7939
rect 7297 7905 7331 7939
rect 8125 7905 8159 7939
rect 9505 7905 9539 7939
rect 14749 7905 14783 7939
rect 16037 7905 16071 7939
rect 1501 7837 1535 7871
rect 4537 7837 4571 7871
rect 5089 7837 5123 7871
rect 5365 7837 5399 7871
rect 6653 7837 6687 7871
rect 7849 7837 7883 7871
rect 9045 7837 9079 7871
rect 9321 7837 9355 7871
rect 9873 7837 9907 7871
rect 10885 7837 10919 7871
rect 11253 7837 11287 7871
rect 12725 7837 12759 7871
rect 13001 7837 13035 7871
rect 14841 7837 14875 7871
rect 16865 7837 16899 7871
rect 17877 7837 17911 7871
rect 3065 7769 3099 7803
rect 10425 7769 10459 7803
rect 11630 7769 11664 7803
rect 16589 7769 16623 7803
rect 4261 7701 4295 7735
rect 8677 7701 8711 7735
rect 9137 7701 9171 7735
rect 10609 7701 10643 7735
rect 12173 7701 12207 7735
rect 15669 7701 15703 7735
rect 2329 7497 2363 7531
rect 4353 7497 4387 7531
rect 5549 7497 5583 7531
rect 6009 7497 6043 7531
rect 7389 7497 7423 7531
rect 7849 7497 7883 7531
rect 7941 7497 7975 7531
rect 11805 7497 11839 7531
rect 15577 7497 15611 7531
rect 16313 7497 16347 7531
rect 17969 7497 18003 7531
rect 8309 7429 8343 7463
rect 13093 7429 13127 7463
rect 16405 7429 16439 7463
rect 17417 7429 17451 7463
rect 17693 7429 17727 7463
rect 1593 7361 1627 7395
rect 1869 7361 1903 7395
rect 2053 7361 2087 7395
rect 3157 7361 3191 7395
rect 3525 7361 3559 7395
rect 3801 7361 3835 7395
rect 4445 7361 4479 7395
rect 4813 7361 4847 7395
rect 5089 7361 5123 7395
rect 6745 7361 6779 7395
rect 7205 7361 7239 7395
rect 7757 7361 7791 7395
rect 8053 7361 8087 7395
rect 8953 7361 8987 7395
rect 9137 7361 9171 7395
rect 9781 7361 9815 7395
rect 10425 7361 10459 7395
rect 10517 7361 10551 7395
rect 11713 7361 11747 7395
rect 11943 7361 11977 7395
rect 12173 7361 12207 7395
rect 12357 7361 12391 7395
rect 13921 7361 13955 7395
rect 14657 7361 14691 7395
rect 15025 7361 15059 7395
rect 15761 7361 15795 7395
rect 16773 7361 16807 7395
rect 18153 7361 18187 7395
rect 2421 7293 2455 7327
rect 2789 7293 2823 7327
rect 3433 7293 3467 7327
rect 5181 7293 5215 7327
rect 9597 7293 9631 7327
rect 11621 7293 11655 7327
rect 13001 7293 13035 7327
rect 13185 7293 13219 7327
rect 14841 7293 14875 7327
rect 9229 7225 9263 7259
rect 13553 7225 13587 7259
rect 15025 7225 15059 7259
rect 6561 7157 6595 7191
rect 8493 7157 8527 7191
rect 9965 7157 9999 7191
rect 10701 7157 10735 7191
rect 14105 7157 14139 7191
rect 3157 6953 3191 6987
rect 2145 6885 2179 6919
rect 13461 6885 13495 6919
rect 2513 6817 2547 6851
rect 7481 6817 7515 6851
rect 10609 6817 10643 6851
rect 15209 6817 15243 6851
rect 18061 6817 18095 6851
rect 1961 6749 1995 6783
rect 2237 6749 2271 6783
rect 3341 6749 3375 6783
rect 3525 6749 3559 6783
rect 4813 6749 4847 6783
rect 5273 6749 5307 6783
rect 5825 6749 5859 6783
rect 6837 6749 6871 6783
rect 10057 6749 10091 6783
rect 10839 6749 10873 6783
rect 10977 6749 11011 6783
rect 11529 6749 11563 6783
rect 11897 6749 11931 6783
rect 13031 6749 13065 6783
rect 13553 6749 13587 6783
rect 14289 6749 14323 6783
rect 14657 6749 14691 6783
rect 15577 6749 15611 6783
rect 15761 6749 15795 6783
rect 16405 6749 16439 6783
rect 17141 6749 17175 6783
rect 17601 6749 17635 6783
rect 4445 6681 4479 6715
rect 8309 6681 8343 6715
rect 9045 6681 9079 6715
rect 17325 6681 17359 6715
rect 18153 6681 18187 6715
rect 1593 6613 1627 6647
rect 2421 6613 2455 6647
rect 2697 6613 2731 6647
rect 4077 6613 4111 6647
rect 10977 6613 11011 6647
rect 12541 6613 12575 6647
rect 12909 6613 12943 6647
rect 13093 6613 13127 6647
rect 15945 6613 15979 6647
rect 4353 6409 4387 6443
rect 8493 6409 8527 6443
rect 9137 6409 9171 6443
rect 12173 6409 12207 6443
rect 15761 6409 15795 6443
rect 3985 6341 4019 6375
rect 10885 6341 10919 6375
rect 12265 6341 12299 6375
rect 16037 6341 16071 6375
rect 16221 6341 16255 6375
rect 1961 6273 1995 6307
rect 2513 6273 2547 6307
rect 2605 6273 2639 6307
rect 2789 6273 2823 6307
rect 3341 6273 3375 6307
rect 3525 6273 3559 6307
rect 3617 6273 3651 6307
rect 3710 6273 3744 6307
rect 4261 6273 4295 6307
rect 4445 6273 4479 6307
rect 5147 6273 5181 6307
rect 5273 6273 5307 6307
rect 5365 6273 5399 6307
rect 5549 6273 5583 6307
rect 5825 6273 5859 6307
rect 6653 6273 6687 6307
rect 6837 6273 6871 6307
rect 7665 6273 7699 6307
rect 8585 6273 8619 6307
rect 9045 6273 9079 6307
rect 9965 6273 9999 6307
rect 10517 6273 10551 6307
rect 10701 6273 10735 6307
rect 13185 6273 13219 6307
rect 14197 6273 14231 6307
rect 14289 6273 14323 6307
rect 15025 6273 15059 6307
rect 15117 6273 15151 6307
rect 16405 6273 16439 6307
rect 16865 6273 16899 6307
rect 18061 6273 18095 6307
rect 2693 6205 2727 6239
rect 6469 6205 6503 6239
rect 8493 6205 8527 6239
rect 9137 6205 9171 6239
rect 12173 6205 12207 6239
rect 13277 6205 13311 6239
rect 13461 6205 13495 6239
rect 14013 6205 14047 6239
rect 14749 6205 14783 6239
rect 14841 6205 14875 6239
rect 4905 6137 4939 6171
rect 8033 6137 8067 6171
rect 9597 6137 9631 6171
rect 18153 6137 18187 6171
rect 1593 6069 1627 6103
rect 2053 6069 2087 6103
rect 2973 6069 3007 6103
rect 5917 6069 5951 6103
rect 7481 6069 7515 6103
rect 10149 6069 10183 6103
rect 11713 6069 11747 6103
rect 13645 6069 13679 6103
rect 15301 6069 15335 6103
rect 2145 5865 2179 5899
rect 3157 5865 3191 5899
rect 4077 5865 4111 5899
rect 4261 5865 4295 5899
rect 13369 5865 13403 5899
rect 18061 5865 18095 5899
rect 4721 5797 4755 5831
rect 7205 5797 7239 5831
rect 17509 5797 17543 5831
rect 18337 5797 18371 5831
rect 2973 5729 3007 5763
rect 5641 5729 5675 5763
rect 8125 5729 8159 5763
rect 10057 5729 10091 5763
rect 15209 5729 15243 5763
rect 17049 5729 17083 5763
rect 2053 5661 2087 5695
rect 2237 5661 2271 5695
rect 2513 5661 2547 5695
rect 2697 5661 2731 5695
rect 2789 5661 2823 5695
rect 2881 5661 2915 5695
rect 5549 5661 5583 5695
rect 6009 5661 6043 5695
rect 6377 5661 6411 5695
rect 7481 5661 7515 5695
rect 8309 5661 8343 5695
rect 8493 5661 8527 5695
rect 9689 5661 9723 5695
rect 9965 5661 9999 5695
rect 11529 5661 11563 5695
rect 13185 5661 13219 5695
rect 14197 5661 14231 5695
rect 14381 5661 14415 5695
rect 14933 5661 14967 5695
rect 17877 5661 17911 5695
rect 4261 5593 4295 5627
rect 4445 5593 4479 5627
rect 4905 5593 4939 5627
rect 5273 5593 5307 5627
rect 7757 5593 7791 5627
rect 17601 5593 17635 5627
rect 1593 5525 1627 5559
rect 4997 5525 5031 5559
rect 5089 5525 5123 5559
rect 6561 5525 6595 5559
rect 7665 5525 7699 5559
rect 11345 5525 11379 5559
rect 14473 5525 14507 5559
rect 16681 5525 16715 5559
rect 3525 5321 3559 5355
rect 4077 5321 4111 5355
rect 4537 5321 4571 5355
rect 5365 5321 5399 5355
rect 8769 5321 8803 5355
rect 10885 5321 10919 5355
rect 13369 5321 13403 5355
rect 15485 5321 15519 5355
rect 15853 5321 15887 5355
rect 16405 5321 16439 5355
rect 16773 5321 16807 5355
rect 17325 5321 17359 5355
rect 7297 5253 7331 5287
rect 9413 5253 9447 5287
rect 11897 5253 11931 5287
rect 14013 5253 14047 5287
rect 17509 5253 17543 5287
rect 2513 5185 2547 5219
rect 2881 5185 2915 5219
rect 3157 5185 3191 5219
rect 3985 5185 4019 5219
rect 4169 5185 4203 5219
rect 4445 5185 4479 5219
rect 4813 5185 4847 5219
rect 5549 5185 5583 5219
rect 6745 5185 6779 5219
rect 13737 5185 13771 5219
rect 4997 5117 5031 5151
rect 5733 5117 5767 5151
rect 7021 5117 7055 5151
rect 9137 5117 9171 5151
rect 11621 5117 11655 5151
rect 17969 5117 18003 5151
rect 2513 4981 2547 5015
rect 6009 4981 6043 5015
rect 6561 4981 6595 5015
rect 2513 4777 2547 4811
rect 2973 4777 3007 4811
rect 7941 4777 7975 4811
rect 11253 4777 11287 4811
rect 14381 4777 14415 4811
rect 16497 4777 16531 4811
rect 10149 4709 10183 4743
rect 13737 4709 13771 4743
rect 1685 4641 1719 4675
rect 5273 4641 5307 4675
rect 6469 4641 6503 4675
rect 9229 4641 9263 4675
rect 13001 4641 13035 4675
rect 14749 4641 14783 4675
rect 17693 4641 17727 4675
rect 1869 4573 1903 4607
rect 2605 4573 2639 4607
rect 3525 4573 3559 4607
rect 4261 4573 4295 4607
rect 4445 4573 4479 4607
rect 4905 4573 4939 4607
rect 5089 4573 5123 4607
rect 5641 4573 5675 4607
rect 5917 4573 5951 4607
rect 6193 4573 6227 4607
rect 8401 4573 8435 4607
rect 8677 4573 8711 4607
rect 9321 4573 9355 4607
rect 9597 4573 9631 4607
rect 9965 4573 9999 4607
rect 10057 4573 10091 4607
rect 13553 4573 13587 4607
rect 13737 4573 13771 4607
rect 14197 4573 14231 4607
rect 17141 4573 17175 4607
rect 17233 4573 17267 4607
rect 17601 4573 17635 4607
rect 18061 4573 18095 4607
rect 4629 4505 4663 4539
rect 8309 4505 8343 4539
rect 12725 4505 12759 4539
rect 15025 4505 15059 4539
rect 16957 4505 16991 4539
rect 2053 4437 2087 4471
rect 3341 4437 3375 4471
rect 3985 4437 4019 4471
rect 5641 4437 5675 4471
rect 4169 4233 4203 4267
rect 5089 4233 5123 4267
rect 11989 4233 12023 4267
rect 12633 4233 12667 4267
rect 14197 4233 14231 4267
rect 16865 4233 16899 4267
rect 1685 4165 1719 4199
rect 2145 4165 2179 4199
rect 17969 4165 18003 4199
rect 1869 4097 1903 4131
rect 2053 4097 2087 4131
rect 2421 4097 2455 4131
rect 5641 4097 5675 4131
rect 5825 4097 5859 4131
rect 8585 4097 8619 4131
rect 9137 4097 9171 4131
rect 9873 4097 9907 4131
rect 10057 4097 10091 4131
rect 10609 4097 10643 4131
rect 11805 4097 11839 4131
rect 12081 4097 12115 4131
rect 12449 4097 12483 4131
rect 12633 4097 12667 4131
rect 13185 4097 13219 4131
rect 13369 4097 13403 4131
rect 14013 4097 14047 4131
rect 14197 4097 14231 4131
rect 17049 4097 17083 4131
rect 17693 4097 17727 4131
rect 18061 4097 18095 4131
rect 18245 4097 18279 4131
rect 2697 4029 2731 4063
rect 4997 4029 5031 4063
rect 5181 4029 5215 4063
rect 5549 4029 5583 4063
rect 6469 4029 6503 4063
rect 6745 4029 6779 4063
rect 9689 4029 9723 4063
rect 10793 4029 10827 4063
rect 13001 4029 13035 4063
rect 14565 4029 14599 4063
rect 14841 4029 14875 4063
rect 17325 4029 17359 4063
rect 4629 3961 4663 3995
rect 9321 3961 9355 3995
rect 8217 3893 8251 3927
rect 8769 3893 8803 3927
rect 10425 3893 10459 3927
rect 16313 3893 16347 3927
rect 17693 3893 17727 3927
rect 2789 3689 2823 3723
rect 6285 3689 6319 3723
rect 13369 3689 13403 3723
rect 16865 3689 16899 3723
rect 18337 3689 18371 3723
rect 6745 3621 6779 3655
rect 2145 3553 2179 3587
rect 2421 3553 2455 3587
rect 3893 3553 3927 3587
rect 5733 3553 5767 3587
rect 7481 3553 7515 3587
rect 11621 3553 11655 3587
rect 15393 3553 15427 3587
rect 17877 3553 17911 3587
rect 1685 3485 1719 3519
rect 3341 3485 3375 3519
rect 4629 3485 4663 3519
rect 4905 3485 4939 3519
rect 6653 3485 6687 3519
rect 7113 3485 7147 3519
rect 7665 3485 7699 3519
rect 7849 3485 7883 3519
rect 8493 3485 8527 3519
rect 8677 3485 8711 3519
rect 9045 3485 9079 3519
rect 9137 3485 9171 3519
rect 9321 3485 9355 3519
rect 9965 3485 9999 3519
rect 10241 3485 10275 3519
rect 10701 3485 10735 3519
rect 10885 3485 10919 3519
rect 10977 3485 11011 3519
rect 11086 3485 11120 3519
rect 14197 3485 14231 3519
rect 14381 3485 14415 3519
rect 15117 3485 15151 3519
rect 17969 3485 18003 3519
rect 2605 3417 2639 3451
rect 5273 3417 5307 3451
rect 6009 3417 6043 3451
rect 10149 3417 10183 3451
rect 11345 3417 11379 3451
rect 11897 3417 11931 3451
rect 1777 3349 1811 3383
rect 2513 3349 2547 3383
rect 3249 3349 3283 3383
rect 5825 3349 5859 3383
rect 8585 3349 8619 3383
rect 9505 3349 9539 3383
rect 14289 3349 14323 3383
rect 17399 3349 17433 3383
rect 17877 3349 17911 3383
rect 2697 3145 2731 3179
rect 4353 3145 4387 3179
rect 4813 3145 4847 3179
rect 5825 3145 5859 3179
rect 7481 3145 7515 3179
rect 8033 3145 8067 3179
rect 16313 3145 16347 3179
rect 17877 3145 17911 3179
rect 17969 3145 18003 3179
rect 2053 3077 2087 3111
rect 9505 3077 9539 3111
rect 14289 3077 14323 3111
rect 17509 3077 17543 3111
rect 1777 3009 1811 3043
rect 2237 3009 2271 3043
rect 2973 3009 3007 3043
rect 3801 3009 3835 3043
rect 3985 3009 4019 3043
rect 4997 3009 5031 3043
rect 5089 3009 5123 3043
rect 5273 3009 5307 3043
rect 5365 3009 5399 3043
rect 5825 3009 5859 3043
rect 6101 3009 6135 3043
rect 6745 3009 6779 3043
rect 7665 3009 7699 3043
rect 9781 3009 9815 3043
rect 10793 3009 10827 3043
rect 11621 3009 11655 3043
rect 11805 3009 11839 3043
rect 12449 3009 12483 3043
rect 12725 3009 12759 3043
rect 13369 3009 13403 3043
rect 13645 3009 13679 3043
rect 13921 3009 13955 3043
rect 14105 3009 14139 3043
rect 17233 3009 17267 3043
rect 6561 2941 6595 2975
rect 6929 2941 6963 2975
rect 10609 2941 10643 2975
rect 11161 2941 11195 2975
rect 14565 2941 14599 2975
rect 14841 2941 14875 2975
rect 17785 2941 17819 2975
rect 18245 2941 18279 2975
rect 11069 2873 11103 2907
rect 12449 2873 12483 2907
rect 13369 2873 13403 2907
rect 11989 2805 12023 2839
rect 17049 2805 17083 2839
rect 2513 2601 2547 2635
rect 7941 2601 7975 2635
rect 10241 2601 10275 2635
rect 11253 2601 11287 2635
rect 13737 2601 13771 2635
rect 14381 2601 14415 2635
rect 3249 2533 3283 2567
rect 4445 2533 4479 2567
rect 17601 2533 17635 2567
rect 4537 2465 4571 2499
rect 5733 2465 5767 2499
rect 7481 2465 7515 2499
rect 10793 2465 10827 2499
rect 11989 2465 12023 2499
rect 15117 2465 15151 2499
rect 15393 2465 15427 2499
rect 1869 2397 1903 2431
rect 2329 2397 2363 2431
rect 2697 2397 2731 2431
rect 2789 2397 2823 2431
rect 3249 2397 3283 2431
rect 3525 2397 3559 2431
rect 3985 2397 4019 2431
rect 4169 2397 4203 2431
rect 5089 2397 5123 2431
rect 5273 2397 5307 2431
rect 5457 2397 5491 2431
rect 8125 2397 8159 2431
rect 8217 2397 8251 2431
rect 9137 2397 9171 2431
rect 9321 2397 9355 2431
rect 10517 2397 10551 2431
rect 10977 2397 11011 2431
rect 14197 2397 14231 2431
rect 6009 2329 6043 2363
rect 10057 2329 10091 2363
rect 11345 2329 11379 2363
rect 12265 2329 12299 2363
rect 17877 2329 17911 2363
rect 18061 2329 18095 2363
rect 18153 2329 18187 2363
rect 1685 2261 1719 2295
rect 9229 2261 9263 2295
rect 10241 2261 10275 2295
rect 14841 2261 14875 2295
rect 16865 2261 16899 2295
rect 5089 2057 5123 2091
rect 6009 2057 6043 2091
rect 6561 2057 6595 2091
rect 8401 2057 8435 2091
rect 18153 2057 18187 2091
rect 1685 1989 1719 2023
rect 2421 1989 2455 2023
rect 3617 1989 3651 2023
rect 1869 1921 1903 1955
rect 1961 1921 1995 1955
rect 2329 1921 2363 1955
rect 2697 1921 2731 1955
rect 3341 1921 3375 1955
rect 5825 1921 5859 1955
rect 6009 1921 6043 1955
rect 6469 1921 6503 1955
rect 10149 1921 10183 1955
rect 10517 1921 10551 1955
rect 11069 1921 11103 1955
rect 13461 1921 13495 1955
rect 15577 1921 15611 1955
rect 15945 1921 15979 1955
rect 16129 1921 16163 1955
rect 17141 1921 17175 1955
rect 17325 1921 17359 1955
rect 2881 1853 2915 1887
rect 6929 1853 6963 1887
rect 7757 1853 7791 1887
rect 9873 1853 9907 1887
rect 11161 1853 11195 1887
rect 13185 1853 13219 1887
rect 15301 1853 15335 1887
rect 10793 1785 10827 1819
rect 15945 1785 15979 1819
rect 11713 1717 11747 1751
rect 13829 1717 13863 1751
rect 3985 1513 4019 1547
rect 5917 1513 5951 1547
rect 12173 1513 12207 1547
rect 1501 1377 1535 1411
rect 4445 1377 4479 1411
rect 7481 1377 7515 1411
rect 9413 1377 9447 1411
rect 10333 1377 10367 1411
rect 11161 1377 11195 1411
rect 14565 1377 14599 1411
rect 14841 1377 14875 1411
rect 3249 1309 3283 1343
rect 5181 1309 5215 1343
rect 5365 1309 5399 1343
rect 5549 1309 5583 1343
rect 6101 1309 6135 1343
rect 7003 1309 7037 1343
rect 8401 1309 8435 1343
rect 9045 1309 9079 1343
rect 9229 1309 9263 1343
rect 9597 1309 9631 1343
rect 10517 1309 10551 1343
rect 11989 1309 12023 1343
rect 16773 1309 16807 1343
rect 16957 1309 16991 1343
rect 17601 1309 17635 1343
rect 18153 1309 18187 1343
rect 4537 1241 4571 1275
rect 7481 1241 7515 1275
rect 7573 1241 7607 1275
rect 4445 1173 4479 1207
rect 6469 1173 6503 1207
rect 8585 1173 8619 1207
rect 16313 1173 16347 1207
rect 16865 1173 16899 1207
rect 17785 1173 17819 1207
rect 18337 1173 18371 1207
<< metal1 >>
rect 12710 13676 12716 13728
rect 12768 13716 12774 13728
rect 17310 13716 17316 13728
rect 12768 13688 17316 13716
rect 12768 13676 12774 13688
rect 17310 13676 17316 13688
rect 17368 13676 17374 13728
rect 1104 13626 18860 13648
rect 1104 13574 4214 13626
rect 4266 13574 4278 13626
rect 4330 13574 4342 13626
rect 4394 13574 4406 13626
rect 4458 13574 4470 13626
rect 4522 13574 12214 13626
rect 12266 13574 12278 13626
rect 12330 13574 12342 13626
rect 12394 13574 12406 13626
rect 12458 13574 12470 13626
rect 12522 13574 18860 13626
rect 1104 13552 18860 13574
rect 1302 13472 1308 13524
rect 1360 13512 1366 13524
rect 3881 13515 3939 13521
rect 3881 13512 3893 13515
rect 1360 13484 3893 13512
rect 1360 13472 1366 13484
rect 3881 13481 3893 13484
rect 3927 13481 3939 13515
rect 3881 13475 3939 13481
rect 3896 13376 3924 13475
rect 7098 13472 7104 13524
rect 7156 13512 7162 13524
rect 8478 13512 8484 13524
rect 7156 13484 8484 13512
rect 7156 13472 7162 13484
rect 8478 13472 8484 13484
rect 8536 13472 8542 13524
rect 5534 13404 5540 13456
rect 5592 13444 5598 13456
rect 7837 13447 7895 13453
rect 7837 13444 7849 13447
rect 5592 13416 7849 13444
rect 5592 13404 5598 13416
rect 7837 13413 7849 13416
rect 7883 13413 7895 13447
rect 7837 13407 7895 13413
rect 13725 13447 13783 13453
rect 13725 13413 13737 13447
rect 13771 13444 13783 13447
rect 13814 13444 13820 13456
rect 13771 13416 13820 13444
rect 13771 13413 13783 13416
rect 13725 13407 13783 13413
rect 13814 13404 13820 13416
rect 13872 13444 13878 13456
rect 13872 13416 16344 13444
rect 13872 13404 13878 13416
rect 3896 13348 6500 13376
rect 2869 13311 2927 13317
rect 2869 13277 2881 13311
rect 2915 13308 2927 13311
rect 2958 13308 2964 13320
rect 2915 13280 2964 13308
rect 2915 13277 2927 13280
rect 2869 13271 2927 13277
rect 2958 13268 2964 13280
rect 3016 13268 3022 13320
rect 3513 13311 3571 13317
rect 3513 13277 3525 13311
rect 3559 13308 3571 13311
rect 4430 13308 4436 13320
rect 3559 13280 4436 13308
rect 3559 13277 3571 13280
rect 3513 13271 3571 13277
rect 4430 13268 4436 13280
rect 4488 13268 4494 13320
rect 4522 13268 4528 13320
rect 4580 13308 4586 13320
rect 6472 13317 6500 13348
rect 6546 13336 6552 13388
rect 6604 13376 6610 13388
rect 6604 13348 8064 13376
rect 6604 13336 6610 13348
rect 4801 13311 4859 13317
rect 4801 13308 4813 13311
rect 4580 13280 4813 13308
rect 4580 13268 4586 13280
rect 4801 13277 4813 13280
rect 4847 13277 4859 13311
rect 4801 13271 4859 13277
rect 6457 13311 6515 13317
rect 6457 13277 6469 13311
rect 6503 13277 6515 13311
rect 6457 13271 6515 13277
rect 6733 13311 6791 13317
rect 6733 13277 6745 13311
rect 6779 13308 6791 13311
rect 7006 13308 7012 13320
rect 6779 13280 7012 13308
rect 6779 13277 6791 13280
rect 6733 13271 6791 13277
rect 7006 13268 7012 13280
rect 7064 13268 7070 13320
rect 8036 13317 8064 13348
rect 8938 13336 8944 13388
rect 8996 13376 9002 13388
rect 14737 13379 14795 13385
rect 8996 13348 14320 13376
rect 8996 13336 9002 13348
rect 8021 13311 8079 13317
rect 8021 13277 8033 13311
rect 8067 13277 8079 13311
rect 8021 13271 8079 13277
rect 9125 13311 9183 13317
rect 9125 13277 9137 13311
rect 9171 13308 9183 13311
rect 9306 13308 9312 13320
rect 9171 13280 9312 13308
rect 9171 13277 9183 13280
rect 9125 13271 9183 13277
rect 9306 13268 9312 13280
rect 9364 13268 9370 13320
rect 10134 13308 10140 13320
rect 10095 13280 10140 13308
rect 10134 13268 10140 13280
rect 10192 13268 10198 13320
rect 11606 13268 11612 13320
rect 11664 13308 11670 13320
rect 11793 13311 11851 13317
rect 11793 13308 11805 13311
rect 11664 13280 11805 13308
rect 11664 13268 11670 13280
rect 11793 13277 11805 13280
rect 11839 13277 11851 13311
rect 11793 13271 11851 13277
rect 12437 13311 12495 13317
rect 12437 13277 12449 13311
rect 12483 13308 12495 13311
rect 12618 13308 12624 13320
rect 12483 13280 12624 13308
rect 12483 13277 12495 13280
rect 12437 13271 12495 13277
rect 12618 13268 12624 13280
rect 12676 13268 12682 13320
rect 13078 13268 13084 13320
rect 13136 13308 13142 13320
rect 13265 13311 13323 13317
rect 13265 13308 13277 13311
rect 13136 13280 13277 13308
rect 13136 13268 13142 13280
rect 13265 13277 13277 13280
rect 13311 13277 13323 13311
rect 14182 13308 14188 13320
rect 14143 13280 14188 13308
rect 13265 13271 13323 13277
rect 14182 13268 14188 13280
rect 14240 13268 14246 13320
rect 14292 13308 14320 13348
rect 14737 13345 14749 13379
rect 14783 13376 14795 13379
rect 16209 13379 16267 13385
rect 16209 13376 16221 13379
rect 14783 13348 16221 13376
rect 14783 13345 14795 13348
rect 14737 13339 14795 13345
rect 16209 13345 16221 13348
rect 16255 13345 16267 13379
rect 16209 13339 16267 13345
rect 15197 13311 15255 13317
rect 14292 13280 15148 13308
rect 3421 13243 3479 13249
rect 3421 13209 3433 13243
rect 3467 13240 3479 13243
rect 4249 13243 4307 13249
rect 4249 13240 4261 13243
rect 3467 13212 4261 13240
rect 3467 13209 3479 13212
rect 3421 13203 3479 13209
rect 4249 13209 4261 13212
rect 4295 13209 4307 13243
rect 4249 13203 4307 13209
rect 4338 13200 4344 13252
rect 4396 13240 4402 13252
rect 5537 13243 5595 13249
rect 5537 13240 5549 13243
rect 4396 13212 5549 13240
rect 4396 13200 4402 13212
rect 5537 13209 5549 13212
rect 5583 13209 5595 13243
rect 5537 13203 5595 13209
rect 5994 13200 6000 13252
rect 6052 13240 6058 13252
rect 6917 13243 6975 13249
rect 6052 13212 6684 13240
rect 6052 13200 6058 13212
rect 2222 13172 2228 13184
rect 2183 13144 2228 13172
rect 2222 13132 2228 13144
rect 2280 13132 2286 13184
rect 2314 13132 2320 13184
rect 2372 13172 2378 13184
rect 2682 13172 2688 13184
rect 2372 13144 2417 13172
rect 2643 13144 2688 13172
rect 2372 13132 2378 13144
rect 2682 13132 2688 13144
rect 2740 13132 2746 13184
rect 5166 13172 5172 13184
rect 5127 13144 5172 13172
rect 5166 13132 5172 13144
rect 5224 13132 5230 13184
rect 5626 13172 5632 13184
rect 5587 13144 5632 13172
rect 5626 13132 5632 13144
rect 5684 13132 5690 13184
rect 6086 13172 6092 13184
rect 6047 13144 6092 13172
rect 6086 13132 6092 13144
rect 6144 13132 6150 13184
rect 6178 13132 6184 13184
rect 6236 13172 6242 13184
rect 6549 13175 6607 13181
rect 6549 13172 6561 13175
rect 6236 13144 6561 13172
rect 6236 13132 6242 13144
rect 6549 13141 6561 13144
rect 6595 13141 6607 13175
rect 6656 13172 6684 13212
rect 6917 13209 6929 13243
rect 6963 13240 6975 13243
rect 7282 13240 7288 13252
rect 6963 13212 7288 13240
rect 6963 13209 6975 13212
rect 6917 13203 6975 13209
rect 7282 13200 7288 13212
rect 7340 13200 7346 13252
rect 7469 13243 7527 13249
rect 7469 13209 7481 13243
rect 7515 13240 7527 13243
rect 7558 13240 7564 13252
rect 7515 13212 7564 13240
rect 7515 13209 7527 13212
rect 7469 13203 7527 13209
rect 7558 13200 7564 13212
rect 7616 13200 7622 13252
rect 8665 13243 8723 13249
rect 8665 13209 8677 13243
rect 8711 13240 8723 13243
rect 9582 13240 9588 13252
rect 8711 13212 9588 13240
rect 8711 13209 8723 13212
rect 8665 13203 8723 13209
rect 9582 13200 9588 13212
rect 9640 13200 9646 13252
rect 9677 13243 9735 13249
rect 9677 13209 9689 13243
rect 9723 13209 9735 13243
rect 9677 13203 9735 13209
rect 7377 13175 7435 13181
rect 7377 13172 7389 13175
rect 6656 13144 7389 13172
rect 6549 13135 6607 13141
rect 7377 13141 7389 13144
rect 7423 13141 7435 13175
rect 8570 13172 8576 13184
rect 8531 13144 8576 13172
rect 7377 13135 7435 13141
rect 8570 13132 8576 13144
rect 8628 13132 8634 13184
rect 9692 13172 9720 13203
rect 9766 13200 9772 13252
rect 9824 13240 9830 13252
rect 10965 13243 11023 13249
rect 10965 13240 10977 13243
rect 9824 13212 10977 13240
rect 9824 13200 9830 13212
rect 10965 13209 10977 13212
rect 11011 13209 11023 13243
rect 10965 13203 11023 13209
rect 11330 13200 11336 13252
rect 11388 13240 11394 13252
rect 12250 13240 12256 13252
rect 11388 13212 12020 13240
rect 12211 13212 12256 13240
rect 11388 13200 11394 13212
rect 9953 13175 10011 13181
rect 9953 13172 9965 13175
rect 9692 13144 9965 13172
rect 9953 13141 9965 13144
rect 9999 13141 10011 13175
rect 10594 13172 10600 13184
rect 10555 13144 10600 13172
rect 9953 13135 10011 13141
rect 10594 13132 10600 13144
rect 10652 13132 10658 13184
rect 10689 13175 10747 13181
rect 10689 13141 10701 13175
rect 10735 13172 10747 13175
rect 10778 13172 10784 13184
rect 10735 13144 10784 13172
rect 10735 13141 10747 13144
rect 10689 13135 10747 13141
rect 10778 13132 10784 13144
rect 10836 13132 10842 13184
rect 11054 13132 11060 13184
rect 11112 13172 11118 13184
rect 11609 13175 11667 13181
rect 11609 13172 11621 13175
rect 11112 13144 11621 13172
rect 11112 13132 11118 13144
rect 11609 13141 11621 13144
rect 11655 13141 11667 13175
rect 11992 13172 12020 13212
rect 12250 13200 12256 13212
rect 12308 13200 12314 13252
rect 12710 13240 12716 13252
rect 12671 13212 12716 13240
rect 12710 13200 12716 13212
rect 12768 13200 12774 13252
rect 13817 13243 13875 13249
rect 13817 13209 13829 13243
rect 13863 13209 13875 13243
rect 14642 13240 14648 13252
rect 14603 13212 14648 13240
rect 13817 13203 13875 13209
rect 12621 13175 12679 13181
rect 12621 13172 12633 13175
rect 11992 13144 12633 13172
rect 11609 13135 11667 13141
rect 12621 13141 12633 13144
rect 12667 13172 12679 13175
rect 13722 13172 13728 13184
rect 12667 13144 13728 13172
rect 12667 13141 12679 13144
rect 12621 13135 12679 13141
rect 13722 13132 13728 13144
rect 13780 13132 13786 13184
rect 13832 13172 13860 13203
rect 14642 13200 14648 13212
rect 14700 13200 14706 13252
rect 15013 13175 15071 13181
rect 15013 13172 15025 13175
rect 13832 13144 15025 13172
rect 15013 13141 15025 13144
rect 15059 13141 15071 13175
rect 15120 13172 15148 13280
rect 15197 13277 15209 13311
rect 15243 13304 15255 13311
rect 15378 13308 15384 13320
rect 15304 13304 15384 13308
rect 15243 13280 15384 13304
rect 15243 13277 15332 13280
rect 15197 13276 15332 13277
rect 15197 13271 15255 13276
rect 15378 13268 15384 13280
rect 15436 13268 15442 13320
rect 15657 13311 15715 13317
rect 15657 13277 15669 13311
rect 15703 13277 15715 13311
rect 15657 13271 15715 13277
rect 16117 13311 16175 13317
rect 16117 13277 16129 13311
rect 16163 13308 16175 13311
rect 16316 13308 16344 13416
rect 17218 13336 17224 13388
rect 17276 13376 17282 13388
rect 18049 13379 18107 13385
rect 18049 13376 18061 13379
rect 17276 13348 18061 13376
rect 17276 13336 17282 13348
rect 18049 13345 18061 13348
rect 18095 13345 18107 13379
rect 18049 13339 18107 13345
rect 16758 13308 16764 13320
rect 16163 13280 16344 13308
rect 16719 13280 16764 13308
rect 16163 13277 16175 13280
rect 16117 13271 16175 13277
rect 15672 13240 15700 13271
rect 16758 13268 16764 13280
rect 16816 13268 16822 13320
rect 15488 13212 15700 13240
rect 15488 13172 15516 13212
rect 16022 13200 16028 13252
rect 16080 13240 16086 13252
rect 17221 13243 17279 13249
rect 17221 13240 17233 13243
rect 16080 13212 17233 13240
rect 16080 13200 16086 13212
rect 17221 13209 17233 13212
rect 17267 13209 17279 13243
rect 17221 13203 17279 13209
rect 17313 13243 17371 13249
rect 17313 13209 17325 13243
rect 17359 13240 17371 13243
rect 17589 13243 17647 13249
rect 17589 13240 17601 13243
rect 17359 13212 17601 13240
rect 17359 13209 17371 13212
rect 17313 13203 17371 13209
rect 17589 13209 17601 13212
rect 17635 13209 17647 13243
rect 17589 13203 17647 13209
rect 15746 13172 15752 13184
rect 15120 13144 15516 13172
rect 15707 13144 15752 13172
rect 15013 13135 15071 13141
rect 15746 13132 15752 13144
rect 15804 13132 15810 13184
rect 17770 13172 17776 13184
rect 17731 13144 17776 13172
rect 17770 13132 17776 13144
rect 17828 13132 17834 13184
rect 1104 13082 18860 13104
rect 1104 13030 8214 13082
rect 8266 13030 8278 13082
rect 8330 13030 8342 13082
rect 8394 13030 8406 13082
rect 8458 13030 8470 13082
rect 8522 13030 16214 13082
rect 16266 13030 16278 13082
rect 16330 13030 16342 13082
rect 16394 13030 16406 13082
rect 16458 13030 16470 13082
rect 16522 13030 18860 13082
rect 1104 13008 18860 13030
rect 6086 12928 6092 12980
rect 6144 12968 6150 12980
rect 6914 12968 6920 12980
rect 6144 12940 6920 12968
rect 6144 12928 6150 12940
rect 6914 12928 6920 12940
rect 6972 12928 6978 12980
rect 10594 12968 10600 12980
rect 7208 12940 10600 12968
rect 2222 12860 2228 12912
rect 2280 12900 2286 12912
rect 2317 12903 2375 12909
rect 2317 12900 2329 12903
rect 2280 12872 2329 12900
rect 2280 12860 2286 12872
rect 2317 12869 2329 12872
rect 2363 12869 2375 12903
rect 2317 12863 2375 12869
rect 4430 12860 4436 12912
rect 4488 12900 4494 12912
rect 4890 12900 4896 12912
rect 4488 12872 4896 12900
rect 4488 12860 4494 12872
rect 4890 12860 4896 12872
rect 4948 12900 4954 12912
rect 4985 12903 5043 12909
rect 4985 12900 4997 12903
rect 4948 12872 4997 12900
rect 4948 12860 4954 12872
rect 4985 12869 4997 12872
rect 5031 12869 5043 12903
rect 4985 12863 5043 12869
rect 5626 12860 5632 12912
rect 5684 12900 5690 12912
rect 7208 12909 7236 12940
rect 10594 12928 10600 12940
rect 10652 12928 10658 12980
rect 11606 12928 11612 12980
rect 11664 12968 11670 12980
rect 14369 12971 14427 12977
rect 14369 12968 14381 12971
rect 11664 12940 14381 12968
rect 11664 12928 11670 12940
rect 14369 12937 14381 12940
rect 14415 12937 14427 12971
rect 16758 12968 16764 12980
rect 14369 12931 14427 12937
rect 15580 12940 16764 12968
rect 7193 12903 7251 12909
rect 5684 12872 7144 12900
rect 5684 12860 5690 12872
rect 1673 12835 1731 12841
rect 1673 12801 1685 12835
rect 1719 12801 1731 12835
rect 1673 12795 1731 12801
rect 2593 12835 2651 12841
rect 2593 12801 2605 12835
rect 2639 12832 2651 12835
rect 2958 12832 2964 12844
rect 2639 12804 2964 12832
rect 2639 12801 2651 12804
rect 2593 12795 2651 12801
rect 1688 12628 1716 12795
rect 2958 12792 2964 12804
rect 3016 12792 3022 12844
rect 3605 12835 3663 12841
rect 3605 12801 3617 12835
rect 3651 12801 3663 12835
rect 4522 12832 4528 12844
rect 4483 12804 4528 12832
rect 3605 12795 3663 12801
rect 3142 12724 3148 12776
rect 3200 12764 3206 12776
rect 3620 12764 3648 12795
rect 4522 12792 4528 12804
rect 4580 12792 4586 12844
rect 4801 12835 4859 12841
rect 4801 12801 4813 12835
rect 4847 12801 4859 12835
rect 4801 12795 4859 12801
rect 5721 12835 5779 12841
rect 5721 12801 5733 12835
rect 5767 12832 5779 12835
rect 5902 12832 5908 12844
rect 5767 12804 5908 12832
rect 5767 12801 5779 12804
rect 5721 12795 5779 12801
rect 4816 12764 4844 12795
rect 5902 12792 5908 12804
rect 5960 12792 5966 12844
rect 6089 12835 6147 12841
rect 6089 12801 6101 12835
rect 6135 12832 6147 12835
rect 6822 12832 6828 12844
rect 6135 12804 6828 12832
rect 6135 12801 6147 12804
rect 6089 12795 6147 12801
rect 6822 12792 6828 12804
rect 6880 12792 6886 12844
rect 7116 12832 7144 12872
rect 7193 12869 7205 12903
rect 7239 12869 7251 12903
rect 7193 12863 7251 12869
rect 7300 12872 9444 12900
rect 7116 12822 7236 12832
rect 7300 12822 7328 12872
rect 7116 12804 7328 12822
rect 7208 12794 7328 12804
rect 7374 12792 7380 12844
rect 7432 12832 7438 12844
rect 8404 12841 8432 12872
rect 7469 12835 7527 12841
rect 7469 12832 7481 12835
rect 7432 12804 7481 12832
rect 7432 12792 7438 12804
rect 7469 12801 7481 12804
rect 7515 12801 7527 12835
rect 7469 12795 7527 12801
rect 8389 12835 8447 12841
rect 8389 12801 8401 12835
rect 8435 12801 8447 12835
rect 9306 12832 9312 12844
rect 9267 12804 9312 12832
rect 8389 12795 8447 12801
rect 9306 12792 9312 12804
rect 9364 12792 9370 12844
rect 9416 12832 9444 12872
rect 9582 12860 9588 12912
rect 9640 12900 9646 12912
rect 9953 12903 10011 12909
rect 9953 12900 9965 12903
rect 9640 12872 9965 12900
rect 9640 12860 9646 12872
rect 9953 12869 9965 12872
rect 9999 12869 10011 12903
rect 9953 12863 10011 12869
rect 10689 12903 10747 12909
rect 10689 12869 10701 12903
rect 10735 12900 10747 12903
rect 11054 12900 11060 12912
rect 10735 12872 11060 12900
rect 10735 12869 10747 12872
rect 10689 12863 10747 12869
rect 11054 12860 11060 12872
rect 11112 12860 11118 12912
rect 11793 12903 11851 12909
rect 11793 12900 11805 12903
rect 11164 12872 11805 12900
rect 10134 12832 10140 12844
rect 9416 12804 10140 12832
rect 10134 12792 10140 12804
rect 10192 12832 10198 12844
rect 10229 12835 10287 12841
rect 10229 12832 10241 12835
rect 10192 12804 10241 12832
rect 10192 12792 10198 12804
rect 10229 12801 10241 12804
rect 10275 12801 10287 12835
rect 10778 12832 10784 12844
rect 10739 12804 10784 12832
rect 10229 12795 10287 12801
rect 10778 12792 10784 12804
rect 10836 12832 10842 12844
rect 11164 12832 11192 12872
rect 11793 12869 11805 12872
rect 11839 12869 11851 12903
rect 13814 12900 13820 12912
rect 11793 12863 11851 12869
rect 12544 12872 13216 12900
rect 13775 12872 13820 12900
rect 11606 12832 11612 12844
rect 10836 12804 11192 12832
rect 11567 12804 11612 12832
rect 10836 12792 10842 12804
rect 11606 12792 11612 12804
rect 11664 12792 11670 12844
rect 12544 12841 12572 12872
rect 12529 12835 12587 12841
rect 12529 12832 12541 12835
rect 11992 12804 12541 12832
rect 3200 12736 4844 12764
rect 3200 12724 3206 12736
rect 3237 12699 3295 12705
rect 3237 12665 3249 12699
rect 3283 12696 3295 12699
rect 4338 12696 4344 12708
rect 3283 12668 4344 12696
rect 3283 12665 3295 12668
rect 3237 12659 3295 12665
rect 4338 12656 4344 12668
rect 4396 12656 4402 12708
rect 4816 12696 4844 12736
rect 6270 12724 6276 12776
rect 6328 12764 6334 12776
rect 6641 12767 6699 12773
rect 6641 12764 6653 12767
rect 6328 12736 6653 12764
rect 6328 12724 6334 12736
rect 6641 12733 6653 12736
rect 6687 12733 6699 12767
rect 6641 12727 6699 12733
rect 6914 12724 6920 12776
rect 6972 12764 6978 12776
rect 11241 12767 11299 12773
rect 6972 12736 11192 12764
rect 6972 12724 6978 12736
rect 6546 12696 6552 12708
rect 4816 12668 6552 12696
rect 6546 12656 6552 12668
rect 6604 12656 6610 12708
rect 7101 12699 7159 12705
rect 7101 12665 7113 12699
rect 7147 12696 7159 12699
rect 7558 12696 7564 12708
rect 7147 12668 7564 12696
rect 7147 12665 7159 12668
rect 7101 12659 7159 12665
rect 7558 12656 7564 12668
rect 7616 12656 7622 12708
rect 8938 12696 8944 12708
rect 8899 12668 8944 12696
rect 8938 12656 8944 12668
rect 8996 12656 9002 12708
rect 11164 12696 11192 12736
rect 11241 12733 11253 12767
rect 11287 12764 11299 12767
rect 11992 12764 12020 12804
rect 12529 12801 12541 12804
rect 12575 12801 12587 12835
rect 13078 12832 13084 12844
rect 13039 12804 13084 12832
rect 12529 12795 12587 12801
rect 13078 12792 13084 12804
rect 13136 12792 13142 12844
rect 13188 12832 13216 12872
rect 13814 12860 13820 12872
rect 13872 12860 13878 12912
rect 14461 12903 14519 12909
rect 14461 12869 14473 12903
rect 14507 12900 14519 12903
rect 14642 12900 14648 12912
rect 14507 12872 14648 12900
rect 14507 12869 14519 12872
rect 14461 12863 14519 12869
rect 14642 12860 14648 12872
rect 14700 12900 14706 12912
rect 15470 12900 15476 12912
rect 14700 12872 15476 12900
rect 14700 12860 14706 12872
rect 15470 12860 15476 12872
rect 15528 12860 15534 12912
rect 13906 12832 13912 12844
rect 13188 12804 13912 12832
rect 13906 12792 13912 12804
rect 13964 12792 13970 12844
rect 13998 12792 14004 12844
rect 14056 12832 14062 12844
rect 14829 12835 14887 12841
rect 14056 12804 14101 12832
rect 14056 12792 14062 12804
rect 14829 12801 14841 12835
rect 14875 12832 14887 12835
rect 15580 12832 15608 12940
rect 16758 12928 16764 12940
rect 16816 12928 16822 12980
rect 17957 12903 18015 12909
rect 17957 12900 17969 12903
rect 16546 12872 17969 12900
rect 15746 12832 15752 12844
rect 14875 12804 15608 12832
rect 15707 12804 15752 12832
rect 14875 12801 14887 12804
rect 14829 12795 14887 12801
rect 11287 12736 12020 12764
rect 11287 12733 11299 12736
rect 11241 12727 11299 12733
rect 12066 12724 12072 12776
rect 12124 12764 12130 12776
rect 14844 12764 14872 12795
rect 15746 12792 15752 12804
rect 15804 12832 15810 12844
rect 16546 12832 16574 12872
rect 17957 12869 17969 12872
rect 18003 12900 18015 12903
rect 18003 12872 18460 12900
rect 18003 12869 18015 12872
rect 17957 12863 18015 12869
rect 17034 12832 17040 12844
rect 15804 12804 16574 12832
rect 16995 12804 17040 12832
rect 15804 12792 15810 12804
rect 17034 12792 17040 12804
rect 17092 12792 17098 12844
rect 17770 12832 17776 12844
rect 17731 12804 17776 12832
rect 17770 12792 17776 12804
rect 17828 12792 17834 12844
rect 18432 12841 18460 12872
rect 18417 12835 18475 12841
rect 18417 12801 18429 12835
rect 18463 12801 18475 12835
rect 18417 12795 18475 12801
rect 12124 12736 14872 12764
rect 12124 12724 12130 12736
rect 12710 12696 12716 12708
rect 11164 12668 12716 12696
rect 12710 12656 12716 12668
rect 12768 12656 12774 12708
rect 16022 12656 16028 12708
rect 16080 12696 16086 12708
rect 16117 12699 16175 12705
rect 16117 12696 16129 12699
rect 16080 12668 16129 12696
rect 16080 12656 16086 12668
rect 16117 12665 16129 12668
rect 16163 12665 16175 12699
rect 16117 12659 16175 12665
rect 1762 12628 1768 12640
rect 1675 12600 1768 12628
rect 1762 12588 1768 12600
rect 1820 12628 1826 12640
rect 12250 12628 12256 12640
rect 1820 12600 12256 12628
rect 1820 12588 1826 12600
rect 12250 12588 12256 12600
rect 12308 12588 12314 12640
rect 13998 12588 14004 12640
rect 14056 12628 14062 12640
rect 15378 12628 15384 12640
rect 14056 12600 15384 12628
rect 14056 12588 14062 12600
rect 15378 12588 15384 12600
rect 15436 12588 15442 12640
rect 18230 12628 18236 12640
rect 18191 12600 18236 12628
rect 18230 12588 18236 12600
rect 18288 12588 18294 12640
rect 1104 12538 18860 12560
rect 1104 12486 4214 12538
rect 4266 12486 4278 12538
rect 4330 12486 4342 12538
rect 4394 12486 4406 12538
rect 4458 12486 4470 12538
rect 4522 12486 12214 12538
rect 12266 12486 12278 12538
rect 12330 12486 12342 12538
rect 12394 12486 12406 12538
rect 12458 12486 12470 12538
rect 12522 12486 18860 12538
rect 1104 12464 18860 12486
rect 3418 12424 3424 12436
rect 3379 12396 3424 12424
rect 3418 12384 3424 12396
rect 3476 12384 3482 12436
rect 4341 12427 4399 12433
rect 4341 12393 4353 12427
rect 4387 12424 4399 12427
rect 4614 12424 4620 12436
rect 4387 12396 4620 12424
rect 4387 12393 4399 12396
rect 4341 12387 4399 12393
rect 4614 12384 4620 12396
rect 4672 12384 4678 12436
rect 7208 12396 7696 12424
rect 2222 12356 2228 12368
rect 2183 12328 2228 12356
rect 2222 12316 2228 12328
rect 2280 12316 2286 12368
rect 3142 12356 3148 12368
rect 3103 12328 3148 12356
rect 3142 12316 3148 12328
rect 3200 12316 3206 12368
rect 4890 12356 4896 12368
rect 4851 12328 4896 12356
rect 4890 12316 4896 12328
rect 4948 12316 4954 12368
rect 1762 12288 1768 12300
rect 1723 12260 1768 12288
rect 1762 12248 1768 12260
rect 1820 12248 1826 12300
rect 2317 12291 2375 12297
rect 2317 12257 2329 12291
rect 2363 12288 2375 12291
rect 2682 12288 2688 12300
rect 2363 12260 2688 12288
rect 2363 12257 2375 12260
rect 2317 12251 2375 12257
rect 2682 12248 2688 12260
rect 2740 12248 2746 12300
rect 4801 12291 4859 12297
rect 4801 12257 4813 12291
rect 4847 12288 4859 12291
rect 5534 12288 5540 12300
rect 4847 12260 5540 12288
rect 4847 12257 4859 12260
rect 4801 12251 4859 12257
rect 5534 12248 5540 12260
rect 5592 12248 5598 12300
rect 5902 12288 5908 12300
rect 5815 12260 5908 12288
rect 3418 12180 3424 12232
rect 3476 12220 3482 12232
rect 3881 12223 3939 12229
rect 3881 12220 3893 12223
rect 3476 12192 3893 12220
rect 3476 12180 3482 12192
rect 3881 12189 3893 12192
rect 3927 12189 3939 12223
rect 3881 12183 3939 12189
rect 4157 12223 4215 12229
rect 4157 12189 4169 12223
rect 4203 12189 4215 12223
rect 4157 12183 4215 12189
rect 5353 12223 5411 12229
rect 5353 12189 5365 12223
rect 5399 12220 5411 12223
rect 5828 12220 5856 12260
rect 5902 12248 5908 12260
rect 5960 12288 5966 12300
rect 7208 12288 7236 12396
rect 7558 12356 7564 12368
rect 7519 12328 7564 12356
rect 7558 12316 7564 12328
rect 7616 12316 7622 12368
rect 7668 12356 7696 12396
rect 7742 12384 7748 12436
rect 7800 12424 7806 12436
rect 9122 12424 9128 12436
rect 7800 12396 9128 12424
rect 7800 12384 7806 12396
rect 9122 12384 9128 12396
rect 9180 12384 9186 12436
rect 9217 12427 9275 12433
rect 9217 12393 9229 12427
rect 9263 12424 9275 12427
rect 9306 12424 9312 12436
rect 9263 12396 9312 12424
rect 9263 12393 9275 12396
rect 9217 12387 9275 12393
rect 9306 12384 9312 12396
rect 9364 12384 9370 12436
rect 9490 12384 9496 12436
rect 9548 12424 9554 12436
rect 11330 12424 11336 12436
rect 9548 12396 11336 12424
rect 9548 12384 9554 12396
rect 11330 12384 11336 12396
rect 11388 12384 11394 12436
rect 11609 12427 11667 12433
rect 11609 12393 11621 12427
rect 11655 12424 11667 12427
rect 12066 12424 12072 12436
rect 11655 12396 12072 12424
rect 11655 12393 11667 12396
rect 11609 12387 11667 12393
rect 12066 12384 12072 12396
rect 12124 12384 12130 12436
rect 12802 12424 12808 12436
rect 12636 12396 12808 12424
rect 10229 12359 10287 12365
rect 10229 12356 10241 12359
rect 7668 12328 10241 12356
rect 10229 12325 10241 12328
rect 10275 12325 10287 12359
rect 11790 12356 11796 12368
rect 10229 12319 10287 12325
rect 10336 12328 11796 12356
rect 5960 12260 7236 12288
rect 5960 12248 5966 12260
rect 7374 12248 7380 12300
rect 7432 12288 7438 12300
rect 8113 12291 8171 12297
rect 8113 12288 8125 12291
rect 7432 12260 8125 12288
rect 7432 12248 7438 12260
rect 8113 12257 8125 12260
rect 8159 12257 8171 12291
rect 8113 12251 8171 12257
rect 8570 12248 8576 12300
rect 8628 12288 8634 12300
rect 8665 12291 8723 12297
rect 8665 12288 8677 12291
rect 8628 12260 8677 12288
rect 8628 12248 8634 12260
rect 8665 12257 8677 12260
rect 8711 12257 8723 12291
rect 8665 12251 8723 12257
rect 9122 12248 9128 12300
rect 9180 12288 9186 12300
rect 9769 12291 9827 12297
rect 9769 12288 9781 12291
rect 9180 12260 9781 12288
rect 9180 12248 9186 12260
rect 9769 12257 9781 12260
rect 9815 12257 9827 12291
rect 10336 12288 10364 12328
rect 11790 12316 11796 12328
rect 11848 12316 11854 12368
rect 11882 12316 11888 12368
rect 11940 12356 11946 12368
rect 12636 12356 12664 12396
rect 12802 12384 12808 12396
rect 12860 12384 12866 12436
rect 12989 12427 13047 12433
rect 12989 12393 13001 12427
rect 13035 12424 13047 12427
rect 13078 12424 13084 12436
rect 13035 12396 13084 12424
rect 13035 12393 13047 12396
rect 12989 12387 13047 12393
rect 13078 12384 13084 12396
rect 13136 12384 13142 12436
rect 13722 12384 13728 12436
rect 13780 12424 13786 12436
rect 14274 12424 14280 12436
rect 13780 12396 14280 12424
rect 13780 12384 13786 12396
rect 14274 12384 14280 12396
rect 14332 12384 14338 12436
rect 17034 12384 17040 12436
rect 17092 12424 17098 12436
rect 17129 12427 17187 12433
rect 17129 12424 17141 12427
rect 17092 12396 17141 12424
rect 17092 12384 17098 12396
rect 17129 12393 17141 12396
rect 17175 12393 17187 12427
rect 17129 12387 17187 12393
rect 11940 12328 12664 12356
rect 11940 12316 11946 12328
rect 12710 12316 12716 12368
rect 12768 12356 12774 12368
rect 12768 12328 12848 12356
rect 12768 12316 12774 12328
rect 9769 12251 9827 12257
rect 10244 12260 10364 12288
rect 5994 12220 6000 12232
rect 5399 12192 5856 12220
rect 5955 12192 6000 12220
rect 5399 12189 5411 12192
rect 5353 12183 5411 12189
rect 2222 12112 2228 12164
rect 2280 12152 2286 12164
rect 2961 12155 3019 12161
rect 2961 12152 2973 12155
rect 2280 12124 2973 12152
rect 2280 12112 2286 12124
rect 2961 12121 2973 12124
rect 3007 12121 3019 12155
rect 4172 12152 4200 12183
rect 5994 12180 6000 12192
rect 6052 12180 6058 12232
rect 6270 12220 6276 12232
rect 6231 12192 6276 12220
rect 6270 12180 6276 12192
rect 6328 12180 6334 12232
rect 7745 12223 7803 12229
rect 7745 12189 7757 12223
rect 7791 12220 7803 12223
rect 7791 12192 9352 12220
rect 7791 12189 7803 12192
rect 7745 12183 7803 12189
rect 8478 12152 8484 12164
rect 4172 12124 8484 12152
rect 2961 12115 3019 12121
rect 8478 12112 8484 12124
rect 8536 12112 8542 12164
rect 8573 12155 8631 12161
rect 8573 12121 8585 12155
rect 8619 12152 8631 12155
rect 8938 12152 8944 12164
rect 8619 12124 8944 12152
rect 8619 12121 8631 12124
rect 8573 12115 8631 12121
rect 8938 12112 8944 12124
rect 8996 12112 9002 12164
rect 9214 12152 9220 12164
rect 9175 12124 9220 12152
rect 9214 12112 9220 12124
rect 9272 12112 9278 12164
rect 9324 12152 9352 12192
rect 9398 12180 9404 12232
rect 9456 12229 9462 12232
rect 9456 12223 9505 12229
rect 9456 12189 9459 12223
rect 9493 12220 9505 12223
rect 10244 12220 10272 12260
rect 10502 12248 10508 12300
rect 10560 12288 10566 12300
rect 12820 12288 12848 12328
rect 12894 12316 12900 12368
rect 12952 12356 12958 12368
rect 15470 12356 15476 12368
rect 12952 12328 15332 12356
rect 15431 12328 15476 12356
rect 12952 12316 12958 12328
rect 10560 12260 12848 12288
rect 10560 12248 10566 12260
rect 10410 12229 10416 12232
rect 9493 12192 10272 12220
rect 9493 12189 9536 12192
rect 9456 12188 9536 12189
rect 9456 12183 9505 12188
rect 10408 12183 10416 12229
rect 10468 12220 10474 12232
rect 10594 12220 10600 12232
rect 10468 12192 10508 12220
rect 10555 12192 10600 12220
rect 9456 12180 9462 12183
rect 10410 12180 10416 12183
rect 10468 12180 10474 12192
rect 10594 12180 10600 12192
rect 10652 12180 10658 12232
rect 10796 12229 10824 12260
rect 12986 12248 12992 12300
rect 13044 12288 13050 12300
rect 15194 12288 15200 12300
rect 13044 12260 15200 12288
rect 13044 12248 13050 12260
rect 15194 12248 15200 12260
rect 15252 12248 15258 12300
rect 15304 12288 15332 12328
rect 15470 12316 15476 12328
rect 15528 12316 15534 12368
rect 17144 12288 17172 12387
rect 17770 12316 17776 12368
rect 17828 12356 17834 12368
rect 17957 12359 18015 12365
rect 17957 12356 17969 12359
rect 17828 12328 17969 12356
rect 17828 12316 17834 12328
rect 17957 12325 17969 12328
rect 18003 12325 18015 12359
rect 17957 12319 18015 12325
rect 17497 12291 17555 12297
rect 17497 12288 17509 12291
rect 15304 12260 17080 12288
rect 17144 12260 17509 12288
rect 10781 12223 10839 12229
rect 10781 12189 10793 12223
rect 10827 12189 10839 12223
rect 10781 12183 10839 12189
rect 11057 12223 11115 12229
rect 11057 12189 11069 12223
rect 11103 12220 11115 12223
rect 11146 12220 11152 12232
rect 11103 12192 11152 12220
rect 11103 12189 11115 12192
rect 11057 12183 11115 12189
rect 11146 12180 11152 12192
rect 11204 12180 11210 12232
rect 11238 12180 11244 12232
rect 11296 12220 11302 12232
rect 11477 12223 11535 12229
rect 11296 12192 11341 12220
rect 11296 12180 11302 12192
rect 11477 12189 11489 12223
rect 11523 12189 11535 12223
rect 12434 12220 12440 12232
rect 12395 12192 12440 12220
rect 11477 12183 11535 12189
rect 10318 12152 10324 12164
rect 9324 12124 10324 12152
rect 10318 12112 10324 12124
rect 10376 12112 10382 12164
rect 10505 12155 10563 12161
rect 10505 12121 10517 12155
rect 10551 12152 10563 12155
rect 10962 12152 10968 12164
rect 10551 12124 10968 12152
rect 10551 12121 10563 12124
rect 10505 12115 10563 12121
rect 10962 12112 10968 12124
rect 11020 12152 11026 12164
rect 11330 12155 11388 12161
rect 11330 12152 11342 12155
rect 11020 12124 11342 12152
rect 11020 12112 11026 12124
rect 11330 12121 11342 12124
rect 11376 12121 11388 12155
rect 11330 12115 11388 12121
rect 3326 12044 3332 12096
rect 3384 12084 3390 12096
rect 3973 12087 4031 12093
rect 3973 12084 3985 12087
rect 3384 12056 3985 12084
rect 3384 12044 3390 12056
rect 3973 12053 3985 12056
rect 4019 12053 4031 12087
rect 5810 12084 5816 12096
rect 5771 12056 5816 12084
rect 3973 12047 4031 12053
rect 5810 12044 5816 12056
rect 5868 12044 5874 12096
rect 7190 12044 7196 12096
rect 7248 12084 7254 12096
rect 7742 12084 7748 12096
rect 7248 12056 7748 12084
rect 7248 12044 7254 12056
rect 7742 12044 7748 12056
rect 7800 12044 7806 12096
rect 9582 12084 9588 12096
rect 9543 12056 9588 12084
rect 9582 12044 9588 12056
rect 9640 12044 9646 12096
rect 9674 12044 9680 12096
rect 9732 12084 9738 12096
rect 9732 12056 9777 12084
rect 9732 12044 9738 12056
rect 9858 12044 9864 12096
rect 9916 12084 9922 12096
rect 11492 12084 11520 12183
rect 12434 12180 12440 12192
rect 12492 12180 12498 12232
rect 12526 12180 12532 12232
rect 12584 12230 12590 12232
rect 12584 12220 12664 12230
rect 12894 12229 12900 12232
rect 12713 12223 12771 12229
rect 12713 12220 12725 12223
rect 12584 12202 12725 12220
rect 12584 12180 12590 12202
rect 12636 12192 12725 12202
rect 12713 12189 12725 12192
rect 12759 12189 12771 12223
rect 12713 12183 12771 12189
rect 12857 12223 12900 12229
rect 12857 12189 12869 12223
rect 12857 12183 12900 12189
rect 12894 12180 12900 12183
rect 12952 12180 12958 12232
rect 13078 12180 13084 12232
rect 13136 12220 13142 12232
rect 13449 12223 13507 12229
rect 13449 12220 13461 12223
rect 13136 12192 13461 12220
rect 13136 12180 13142 12192
rect 13449 12189 13461 12192
rect 13495 12189 13507 12223
rect 13630 12220 13636 12232
rect 13591 12192 13636 12220
rect 13449 12183 13507 12189
rect 13630 12180 13636 12192
rect 13688 12180 13694 12232
rect 14182 12220 14188 12232
rect 14143 12192 14188 12220
rect 14182 12180 14188 12192
rect 14240 12180 14246 12232
rect 15378 12220 15384 12232
rect 15339 12192 15384 12220
rect 15378 12180 15384 12192
rect 15436 12180 15442 12232
rect 16022 12180 16028 12232
rect 16080 12220 16086 12232
rect 16209 12223 16267 12229
rect 16209 12220 16221 12223
rect 16080 12192 16221 12220
rect 16080 12180 16086 12192
rect 16209 12189 16221 12192
rect 16255 12189 16267 12223
rect 16942 12220 16948 12232
rect 16903 12192 16948 12220
rect 16209 12183 16267 12189
rect 16942 12180 16948 12192
rect 17000 12180 17006 12232
rect 17052 12220 17080 12260
rect 17497 12257 17509 12260
rect 17543 12257 17555 12291
rect 17497 12251 17555 12257
rect 18049 12291 18107 12297
rect 18049 12257 18061 12291
rect 18095 12288 18107 12291
rect 18230 12288 18236 12300
rect 18095 12260 18236 12288
rect 18095 12257 18107 12260
rect 18049 12251 18107 12257
rect 18230 12248 18236 12260
rect 18288 12248 18294 12300
rect 18325 12223 18383 12229
rect 18325 12220 18337 12223
rect 17052 12192 18337 12220
rect 18325 12189 18337 12192
rect 18371 12189 18383 12223
rect 18325 12183 18383 12189
rect 12621 12155 12679 12161
rect 12621 12121 12633 12155
rect 12667 12152 12679 12155
rect 15286 12152 15292 12164
rect 12667 12124 15292 12152
rect 12667 12121 12679 12124
rect 12621 12115 12679 12121
rect 15286 12112 15292 12124
rect 15344 12112 15350 12164
rect 16669 12155 16727 12161
rect 16669 12152 16681 12155
rect 16040 12124 16681 12152
rect 16040 12096 16068 12124
rect 16669 12121 16681 12124
rect 16715 12121 16727 12155
rect 16669 12115 16727 12121
rect 9916 12056 11520 12084
rect 9916 12044 9922 12056
rect 11790 12044 11796 12096
rect 11848 12084 11854 12096
rect 11974 12084 11980 12096
rect 11848 12056 11980 12084
rect 11848 12044 11854 12056
rect 11974 12044 11980 12056
rect 12032 12044 12038 12096
rect 12802 12044 12808 12096
rect 12860 12084 12866 12096
rect 13633 12087 13691 12093
rect 13633 12084 13645 12087
rect 12860 12056 13645 12084
rect 12860 12044 12866 12056
rect 13633 12053 13645 12056
rect 13679 12084 13691 12087
rect 14826 12084 14832 12096
rect 13679 12056 14832 12084
rect 13679 12053 13691 12056
rect 13633 12047 13691 12053
rect 14826 12044 14832 12056
rect 14884 12044 14890 12096
rect 16022 12044 16028 12096
rect 16080 12044 16086 12096
rect 16114 12044 16120 12096
rect 16172 12084 16178 12096
rect 16301 12087 16359 12093
rect 16301 12084 16313 12087
rect 16172 12056 16313 12084
rect 16172 12044 16178 12056
rect 16301 12053 16313 12056
rect 16347 12053 16359 12087
rect 16758 12084 16764 12096
rect 16719 12056 16764 12084
rect 16301 12047 16359 12053
rect 16758 12044 16764 12056
rect 16816 12084 16822 12096
rect 17218 12084 17224 12096
rect 16816 12056 17224 12084
rect 16816 12044 16822 12056
rect 17218 12044 17224 12056
rect 17276 12044 17282 12096
rect 1104 11994 18860 12016
rect 1104 11942 8214 11994
rect 8266 11942 8278 11994
rect 8330 11942 8342 11994
rect 8394 11942 8406 11994
rect 8458 11942 8470 11994
rect 8522 11942 16214 11994
rect 16266 11942 16278 11994
rect 16330 11942 16342 11994
rect 16394 11942 16406 11994
rect 16458 11942 16470 11994
rect 16522 11942 18860 11994
rect 1104 11920 18860 11942
rect 2958 11880 2964 11892
rect 2919 11852 2964 11880
rect 2958 11840 2964 11852
rect 3016 11840 3022 11892
rect 5629 11883 5687 11889
rect 5629 11880 5641 11883
rect 3528 11852 5641 11880
rect 2314 11812 2320 11824
rect 2275 11784 2320 11812
rect 2314 11772 2320 11784
rect 2372 11772 2378 11824
rect 3418 11812 3424 11824
rect 3379 11784 3424 11812
rect 3418 11772 3424 11784
rect 3476 11772 3482 11824
rect 3053 11747 3111 11753
rect 3053 11713 3065 11747
rect 3099 11713 3111 11747
rect 3053 11707 3111 11713
rect 1486 11636 1492 11688
rect 1544 11676 1550 11688
rect 1765 11679 1823 11685
rect 1765 11676 1777 11679
rect 1544 11648 1777 11676
rect 1544 11636 1550 11648
rect 1765 11645 1777 11648
rect 1811 11645 1823 11679
rect 1765 11639 1823 11645
rect 2222 11608 2228 11620
rect 2183 11580 2228 11608
rect 2222 11568 2228 11580
rect 2280 11568 2286 11620
rect 3068 11608 3096 11707
rect 3326 11704 3332 11756
rect 3384 11744 3390 11756
rect 3528 11753 3556 11852
rect 5629 11849 5641 11852
rect 5675 11880 5687 11883
rect 6178 11880 6184 11892
rect 5675 11852 6184 11880
rect 5675 11849 5687 11852
rect 5629 11843 5687 11849
rect 6178 11840 6184 11852
rect 6236 11840 6242 11892
rect 6917 11883 6975 11889
rect 6917 11849 6929 11883
rect 6963 11880 6975 11883
rect 7006 11880 7012 11892
rect 6963 11852 7012 11880
rect 6963 11849 6975 11852
rect 6917 11843 6975 11849
rect 7006 11840 7012 11852
rect 7064 11840 7070 11892
rect 9125 11883 9183 11889
rect 7668 11852 8432 11880
rect 4062 11772 4068 11824
rect 4120 11812 4126 11824
rect 5166 11812 5172 11824
rect 4120 11784 5172 11812
rect 4120 11772 4126 11784
rect 5166 11772 5172 11784
rect 5224 11772 5230 11824
rect 5261 11815 5319 11821
rect 5261 11781 5273 11815
rect 5307 11812 5319 11815
rect 5902 11812 5908 11824
rect 5307 11784 5908 11812
rect 5307 11781 5319 11784
rect 5261 11775 5319 11781
rect 5902 11772 5908 11784
rect 5960 11772 5966 11824
rect 5997 11815 6055 11821
rect 5997 11781 6009 11815
rect 6043 11812 6055 11815
rect 6270 11812 6276 11824
rect 6043 11784 6276 11812
rect 6043 11781 6055 11784
rect 5997 11775 6055 11781
rect 6270 11772 6276 11784
rect 6328 11772 6334 11824
rect 6549 11815 6607 11821
rect 6549 11781 6561 11815
rect 6595 11812 6607 11815
rect 7668 11812 7696 11852
rect 6595 11784 7696 11812
rect 7745 11815 7803 11821
rect 6595 11781 6607 11784
rect 6549 11775 6607 11781
rect 7745 11781 7757 11815
rect 7791 11812 7803 11815
rect 8202 11812 8208 11824
rect 7791 11784 8208 11812
rect 7791 11781 7803 11784
rect 7745 11775 7803 11781
rect 8202 11772 8208 11784
rect 8260 11772 8266 11824
rect 3513 11747 3571 11753
rect 3513 11744 3525 11747
rect 3384 11716 3525 11744
rect 3384 11704 3390 11716
rect 3513 11713 3525 11716
rect 3559 11713 3571 11747
rect 3513 11707 3571 11713
rect 3697 11747 3755 11753
rect 3697 11713 3709 11747
rect 3743 11744 3755 11747
rect 4801 11747 4859 11753
rect 3743 11716 4752 11744
rect 3743 11713 3755 11716
rect 3697 11707 3755 11713
rect 3878 11676 3884 11688
rect 3791 11648 3884 11676
rect 3878 11636 3884 11648
rect 3936 11676 3942 11688
rect 4249 11679 4307 11685
rect 4249 11676 4261 11679
rect 3936 11648 4261 11676
rect 3936 11636 3942 11648
rect 4249 11645 4261 11648
rect 4295 11645 4307 11679
rect 4724 11676 4752 11716
rect 4801 11713 4813 11747
rect 4847 11744 4859 11747
rect 5077 11747 5135 11753
rect 5077 11744 5089 11747
rect 4847 11716 5089 11744
rect 4847 11713 4859 11716
rect 4801 11707 4859 11713
rect 5077 11713 5089 11716
rect 5123 11713 5135 11747
rect 5184 11744 5212 11772
rect 5537 11747 5595 11753
rect 5537 11744 5549 11747
rect 5184 11716 5549 11744
rect 5077 11707 5135 11713
rect 5537 11713 5549 11716
rect 5583 11713 5595 11747
rect 5537 11707 5595 11713
rect 5813 11747 5871 11753
rect 5813 11713 5825 11747
rect 5859 11744 5871 11747
rect 6086 11744 6092 11756
rect 5859 11716 6092 11744
rect 5859 11713 5871 11716
rect 5813 11707 5871 11713
rect 6086 11704 6092 11716
rect 6144 11704 6150 11756
rect 7006 11704 7012 11756
rect 7064 11744 7070 11756
rect 7101 11747 7159 11753
rect 7101 11744 7113 11747
rect 7064 11716 7113 11744
rect 7064 11704 7070 11716
rect 7101 11713 7113 11716
rect 7147 11713 7159 11747
rect 7101 11707 7159 11713
rect 7377 11747 7435 11753
rect 7377 11713 7389 11747
rect 7423 11744 7435 11747
rect 8018 11744 8024 11756
rect 7423 11716 8024 11744
rect 7423 11713 7435 11716
rect 7377 11707 7435 11713
rect 8018 11704 8024 11716
rect 8076 11704 8082 11756
rect 8297 11747 8355 11753
rect 8297 11713 8309 11747
rect 8343 11713 8355 11747
rect 8404 11744 8432 11852
rect 9125 11849 9137 11883
rect 9171 11880 9183 11883
rect 9398 11880 9404 11892
rect 9171 11852 9404 11880
rect 9171 11849 9183 11852
rect 9125 11843 9183 11849
rect 9398 11840 9404 11852
rect 9456 11840 9462 11892
rect 9493 11883 9551 11889
rect 9493 11849 9505 11883
rect 9539 11880 9551 11883
rect 9674 11880 9680 11892
rect 9539 11852 9680 11880
rect 9539 11849 9551 11852
rect 9493 11843 9551 11849
rect 9674 11840 9680 11852
rect 9732 11840 9738 11892
rect 9769 11883 9827 11889
rect 9769 11849 9781 11883
rect 9815 11880 9827 11883
rect 10502 11880 10508 11892
rect 9815 11852 10508 11880
rect 9815 11849 9827 11852
rect 9769 11843 9827 11849
rect 10502 11840 10508 11852
rect 10560 11840 10566 11892
rect 10594 11840 10600 11892
rect 10652 11880 10658 11892
rect 10873 11883 10931 11889
rect 10873 11880 10885 11883
rect 10652 11852 10885 11880
rect 10652 11840 10658 11852
rect 10873 11849 10885 11852
rect 10919 11849 10931 11883
rect 10873 11843 10931 11849
rect 11054 11840 11060 11892
rect 11112 11880 11118 11892
rect 11112 11852 11928 11880
rect 11112 11840 11118 11852
rect 8570 11772 8576 11824
rect 8628 11812 8634 11824
rect 9950 11812 9956 11824
rect 8628 11784 9956 11812
rect 8628 11772 8634 11784
rect 9950 11772 9956 11784
rect 10008 11772 10014 11824
rect 10134 11772 10140 11824
rect 10192 11812 10198 11824
rect 10612 11812 10640 11840
rect 10192 11784 10640 11812
rect 10192 11772 10198 11784
rect 11238 11772 11244 11824
rect 11296 11812 11302 11824
rect 11698 11812 11704 11824
rect 11296 11784 11704 11812
rect 11296 11772 11302 11784
rect 11698 11772 11704 11784
rect 11756 11772 11762 11824
rect 11900 11821 11928 11852
rect 12158 11840 12164 11892
rect 12216 11880 12222 11892
rect 13265 11883 13323 11889
rect 12216 11852 13124 11880
rect 12216 11840 12222 11852
rect 11885 11815 11943 11821
rect 11885 11781 11897 11815
rect 11931 11812 11943 11815
rect 12342 11812 12348 11824
rect 11931 11784 12348 11812
rect 11931 11781 11943 11784
rect 11885 11775 11943 11781
rect 12342 11772 12348 11784
rect 12400 11772 12406 11824
rect 13096 11821 13124 11852
rect 13265 11849 13277 11883
rect 13311 11880 13323 11883
rect 13814 11880 13820 11892
rect 13311 11852 13820 11880
rect 13311 11849 13323 11852
rect 13265 11843 13323 11849
rect 13814 11840 13820 11852
rect 13872 11840 13878 11892
rect 14090 11840 14096 11892
rect 14148 11880 14154 11892
rect 15378 11880 15384 11892
rect 14148 11852 15056 11880
rect 15339 11852 15384 11880
rect 14148 11840 14154 11852
rect 15028 11824 15056 11852
rect 15378 11840 15384 11852
rect 15436 11840 15442 11892
rect 13081 11815 13139 11821
rect 13081 11781 13093 11815
rect 13127 11781 13139 11815
rect 13906 11812 13912 11824
rect 13867 11784 13912 11812
rect 13081 11775 13139 11781
rect 13906 11772 13912 11784
rect 13964 11772 13970 11824
rect 14274 11812 14280 11824
rect 14235 11784 14280 11812
rect 14274 11772 14280 11784
rect 14332 11812 14338 11824
rect 14918 11812 14924 11824
rect 14332 11784 14924 11812
rect 14332 11772 14338 11784
rect 14918 11772 14924 11784
rect 14976 11772 14982 11824
rect 15010 11772 15016 11824
rect 15068 11812 15074 11824
rect 15068 11784 15161 11812
rect 15212 11784 16896 11812
rect 15068 11772 15074 11784
rect 8481 11747 8539 11753
rect 8481 11744 8493 11747
rect 8404 11716 8493 11744
rect 8297 11707 8355 11713
rect 8481 11713 8493 11716
rect 8527 11744 8539 11747
rect 9490 11744 9496 11756
rect 8527 11716 9496 11744
rect 8527 11713 8539 11716
rect 8481 11707 8539 11713
rect 4724 11648 5304 11676
rect 4249 11639 4307 11645
rect 4709 11611 4767 11617
rect 4709 11608 4721 11611
rect 3068 11580 4721 11608
rect 4709 11577 4721 11580
rect 4755 11608 4767 11611
rect 5166 11608 5172 11620
rect 4755 11580 5172 11608
rect 4755 11577 4767 11580
rect 4709 11571 4767 11577
rect 5166 11568 5172 11580
rect 5224 11568 5230 11620
rect 5276 11540 5304 11648
rect 5350 11636 5356 11688
rect 5408 11676 5414 11688
rect 8113 11679 8171 11685
rect 8113 11676 8125 11679
rect 5408 11648 8125 11676
rect 5408 11636 5414 11648
rect 8113 11645 8125 11648
rect 8159 11645 8171 11679
rect 8113 11639 8171 11645
rect 7285 11611 7343 11617
rect 7285 11577 7297 11611
rect 7331 11608 7343 11611
rect 8202 11608 8208 11620
rect 7331 11580 8208 11608
rect 7331 11577 7343 11580
rect 7285 11571 7343 11577
rect 8202 11568 8208 11580
rect 8260 11568 8266 11620
rect 8312 11608 8340 11707
rect 9490 11704 9496 11716
rect 9548 11704 9554 11756
rect 9858 11704 9864 11756
rect 9916 11744 9922 11756
rect 10045 11747 10103 11753
rect 10045 11744 10057 11747
rect 9916 11716 10057 11744
rect 9916 11704 9922 11716
rect 10045 11713 10057 11716
rect 10091 11713 10103 11747
rect 10226 11744 10232 11756
rect 10187 11716 10232 11744
rect 10045 11707 10103 11713
rect 10226 11704 10232 11716
rect 10284 11704 10290 11756
rect 10689 11747 10747 11753
rect 10689 11713 10701 11747
rect 10735 11744 10747 11747
rect 11256 11744 11284 11772
rect 10735 11716 11284 11744
rect 10735 11713 10747 11716
rect 10689 11707 10747 11713
rect 8662 11636 8668 11688
rect 8720 11676 8726 11688
rect 9677 11679 9735 11685
rect 9677 11676 9689 11679
rect 8720 11648 9689 11676
rect 8720 11636 8726 11648
rect 9677 11645 9689 11648
rect 9723 11645 9735 11679
rect 9950 11676 9956 11688
rect 9911 11648 9956 11676
rect 9677 11639 9735 11645
rect 9950 11636 9956 11648
rect 10008 11636 10014 11688
rect 10502 11676 10508 11688
rect 10463 11648 10508 11676
rect 10502 11636 10508 11648
rect 10560 11636 10566 11688
rect 8570 11608 8576 11620
rect 8312 11580 8576 11608
rect 8570 11568 8576 11580
rect 8628 11568 8634 11620
rect 9490 11568 9496 11620
rect 9548 11608 9554 11620
rect 10704 11608 10732 11707
rect 11514 11704 11520 11756
rect 11572 11744 11578 11756
rect 11609 11747 11667 11753
rect 11609 11744 11621 11747
rect 11572 11716 11621 11744
rect 11572 11704 11578 11716
rect 11609 11713 11621 11716
rect 11655 11713 11667 11747
rect 11609 11707 11667 11713
rect 11793 11747 11851 11753
rect 11793 11713 11805 11747
rect 11839 11713 11851 11747
rect 11974 11744 11980 11756
rect 12032 11753 12038 11756
rect 11940 11716 11980 11744
rect 11793 11707 11851 11713
rect 9548 11580 10732 11608
rect 9548 11568 9554 11580
rect 11606 11568 11612 11620
rect 11664 11608 11670 11620
rect 11808 11608 11836 11707
rect 11974 11704 11980 11716
rect 12032 11707 12040 11753
rect 12529 11747 12587 11753
rect 12529 11744 12541 11747
rect 12084 11716 12541 11744
rect 12032 11704 12038 11707
rect 12084 11688 12112 11716
rect 12529 11713 12541 11716
rect 12575 11713 12587 11747
rect 12529 11707 12587 11713
rect 13541 11747 13599 11753
rect 13541 11713 13553 11747
rect 13587 11744 13599 11747
rect 14090 11744 14096 11756
rect 13587 11716 14096 11744
rect 13587 11713 13599 11716
rect 13541 11707 13599 11713
rect 14090 11704 14096 11716
rect 14148 11704 14154 11756
rect 14366 11704 14372 11756
rect 14424 11744 14430 11756
rect 15212 11744 15240 11784
rect 14424 11716 14469 11744
rect 14844 11716 15240 11744
rect 15269 11747 15327 11753
rect 14424 11704 14430 11716
rect 12066 11636 12072 11688
rect 12124 11636 12130 11688
rect 14844 11676 14872 11716
rect 15269 11713 15281 11747
rect 15315 11744 15327 11747
rect 15746 11744 15752 11756
rect 15315 11716 15752 11744
rect 15315 11713 15327 11716
rect 15269 11707 15327 11713
rect 15746 11704 15752 11716
rect 15804 11704 15810 11756
rect 16114 11704 16120 11756
rect 16172 11744 16178 11756
rect 16868 11753 16896 11784
rect 16209 11747 16267 11753
rect 16209 11744 16221 11747
rect 16172 11716 16221 11744
rect 16172 11704 16178 11716
rect 16209 11713 16221 11716
rect 16255 11713 16267 11747
rect 16209 11707 16267 11713
rect 16853 11747 16911 11753
rect 16853 11713 16865 11747
rect 16899 11744 16911 11747
rect 17678 11744 17684 11756
rect 16899 11716 17684 11744
rect 16899 11713 16911 11716
rect 16853 11707 16911 11713
rect 15470 11676 15476 11688
rect 12176 11648 14872 11676
rect 15431 11648 15476 11676
rect 12176 11617 12204 11648
rect 15470 11636 15476 11648
rect 15528 11636 15534 11688
rect 15562 11636 15568 11688
rect 15620 11676 15626 11688
rect 16224 11676 16252 11707
rect 17678 11704 17684 11716
rect 17736 11704 17742 11756
rect 17773 11747 17831 11753
rect 17773 11713 17785 11747
rect 17819 11713 17831 11747
rect 17773 11707 17831 11713
rect 17788 11676 17816 11707
rect 15620 11648 15665 11676
rect 16224 11648 17816 11676
rect 15620 11636 15626 11648
rect 16868 11620 16896 11648
rect 11664 11580 11836 11608
rect 12161 11611 12219 11617
rect 11664 11568 11670 11580
rect 12161 11577 12173 11611
rect 12207 11577 12219 11611
rect 14829 11611 14887 11617
rect 14829 11608 14841 11611
rect 12161 11571 12219 11577
rect 12406 11580 14841 11608
rect 10870 11540 10876 11552
rect 5276 11512 10876 11540
rect 10870 11500 10876 11512
rect 10928 11500 10934 11552
rect 10962 11500 10968 11552
rect 11020 11540 11026 11552
rect 12406 11540 12434 11580
rect 14829 11577 14841 11580
rect 14875 11577 14887 11611
rect 14829 11571 14887 11577
rect 14918 11568 14924 11620
rect 14976 11608 14982 11620
rect 15841 11611 15899 11617
rect 15841 11608 15853 11611
rect 14976 11580 15853 11608
rect 14976 11568 14982 11580
rect 15841 11577 15853 11580
rect 15887 11608 15899 11611
rect 16758 11608 16764 11620
rect 15887 11580 16764 11608
rect 15887 11577 15899 11580
rect 15841 11571 15899 11577
rect 16758 11568 16764 11580
rect 16816 11568 16822 11620
rect 16850 11568 16856 11620
rect 16908 11568 16914 11620
rect 18138 11608 18144 11620
rect 18099 11580 18144 11608
rect 18138 11568 18144 11580
rect 18196 11568 18202 11620
rect 12618 11540 12624 11552
rect 11020 11512 12434 11540
rect 12579 11512 12624 11540
rect 11020 11500 11026 11512
rect 12618 11500 12624 11512
rect 12676 11500 12682 11552
rect 12802 11500 12808 11552
rect 12860 11540 12866 11552
rect 13265 11543 13323 11549
rect 13265 11540 13277 11543
rect 12860 11512 13277 11540
rect 12860 11500 12866 11512
rect 13265 11509 13277 11512
rect 13311 11540 13323 11543
rect 13354 11540 13360 11552
rect 13311 11512 13360 11540
rect 13311 11509 13323 11512
rect 13265 11503 13323 11509
rect 13354 11500 13360 11512
rect 13412 11500 13418 11552
rect 13538 11500 13544 11552
rect 13596 11540 13602 11552
rect 14642 11540 14648 11552
rect 13596 11512 14648 11540
rect 13596 11500 13602 11512
rect 14642 11500 14648 11512
rect 14700 11500 14706 11552
rect 16393 11543 16451 11549
rect 16393 11509 16405 11543
rect 16439 11540 16451 11543
rect 17126 11540 17132 11552
rect 16439 11512 17132 11540
rect 16439 11509 16451 11512
rect 16393 11503 16451 11509
rect 17126 11500 17132 11512
rect 17184 11500 17190 11552
rect 1104 11450 18860 11472
rect 1104 11398 4214 11450
rect 4266 11398 4278 11450
rect 4330 11398 4342 11450
rect 4394 11398 4406 11450
rect 4458 11398 4470 11450
rect 4522 11398 12214 11450
rect 12266 11398 12278 11450
rect 12330 11398 12342 11450
rect 12394 11398 12406 11450
rect 12458 11398 12470 11450
rect 12522 11398 18860 11450
rect 1104 11376 18860 11398
rect 3418 11336 3424 11348
rect 3379 11308 3424 11336
rect 3418 11296 3424 11308
rect 3476 11296 3482 11348
rect 7101 11339 7159 11345
rect 7101 11305 7113 11339
rect 7147 11336 7159 11339
rect 10962 11336 10968 11348
rect 7147 11308 10968 11336
rect 7147 11305 7159 11308
rect 7101 11299 7159 11305
rect 10962 11296 10968 11308
rect 11020 11296 11026 11348
rect 12986 11296 12992 11348
rect 13044 11336 13050 11348
rect 13630 11336 13636 11348
rect 13044 11308 13636 11336
rect 13044 11296 13050 11308
rect 13630 11296 13636 11308
rect 13688 11296 13694 11348
rect 13725 11339 13783 11345
rect 13725 11305 13737 11339
rect 13771 11336 13783 11339
rect 13814 11336 13820 11348
rect 13771 11308 13820 11336
rect 13771 11305 13783 11308
rect 13725 11299 13783 11305
rect 13814 11296 13820 11308
rect 13872 11296 13878 11348
rect 15286 11336 15292 11348
rect 15247 11308 15292 11336
rect 15286 11296 15292 11308
rect 15344 11296 15350 11348
rect 2222 11228 2228 11280
rect 2280 11268 2286 11280
rect 2777 11271 2835 11277
rect 2777 11268 2789 11271
rect 2280 11240 2789 11268
rect 2280 11228 2286 11240
rect 2777 11237 2789 11240
rect 2823 11237 2835 11271
rect 5166 11268 5172 11280
rect 5127 11240 5172 11268
rect 2777 11231 2835 11237
rect 5166 11228 5172 11240
rect 5224 11228 5230 11280
rect 6086 11228 6092 11280
rect 6144 11268 6150 11280
rect 7282 11268 7288 11280
rect 6144 11240 7288 11268
rect 6144 11228 6150 11240
rect 7282 11228 7288 11240
rect 7340 11268 7346 11280
rect 8662 11268 8668 11280
rect 7340 11240 8524 11268
rect 8623 11240 8668 11268
rect 7340 11228 7346 11240
rect 6730 11160 6736 11212
rect 6788 11200 6794 11212
rect 7576 11209 7604 11240
rect 7561 11203 7619 11209
rect 6788 11172 7488 11200
rect 6788 11160 6794 11172
rect 1486 11132 1492 11144
rect 1447 11104 1492 11132
rect 1486 11092 1492 11104
rect 1544 11092 1550 11144
rect 2958 11132 2964 11144
rect 2919 11104 2964 11132
rect 2958 11092 2964 11104
rect 3016 11092 3022 11144
rect 3878 11132 3884 11144
rect 3839 11104 3884 11132
rect 3878 11092 3884 11104
rect 3936 11092 3942 11144
rect 5353 11135 5411 11141
rect 5353 11101 5365 11135
rect 5399 11101 5411 11135
rect 5902 11132 5908 11144
rect 5863 11104 5908 11132
rect 5353 11095 5411 11101
rect 5368 11064 5396 11095
rect 5902 11092 5908 11104
rect 5960 11092 5966 11144
rect 6086 11092 6092 11144
rect 6144 11132 6150 11144
rect 6641 11135 6699 11141
rect 6641 11132 6653 11135
rect 6144 11104 6653 11132
rect 6144 11092 6150 11104
rect 6641 11101 6653 11104
rect 6687 11132 6699 11135
rect 6822 11132 6828 11144
rect 6687 11104 6828 11132
rect 6687 11101 6699 11104
rect 6641 11095 6699 11101
rect 6822 11092 6828 11104
rect 6880 11092 6886 11144
rect 7357 11135 7415 11141
rect 7357 11101 7369 11135
rect 7403 11132 7415 11135
rect 7460 11132 7488 11172
rect 7561 11169 7573 11203
rect 7607 11169 7619 11203
rect 7561 11163 7619 11169
rect 7653 11203 7711 11209
rect 7653 11169 7665 11203
rect 7699 11200 7711 11203
rect 8496 11200 8524 11240
rect 8662 11228 8668 11240
rect 8720 11228 8726 11280
rect 10042 11268 10048 11280
rect 10003 11240 10048 11268
rect 10042 11228 10048 11240
rect 10100 11228 10106 11280
rect 10502 11228 10508 11280
rect 10560 11268 10566 11280
rect 10597 11271 10655 11277
rect 10597 11268 10609 11271
rect 10560 11240 10609 11268
rect 10560 11228 10566 11240
rect 10597 11237 10609 11240
rect 10643 11237 10655 11271
rect 11146 11268 11152 11280
rect 10597 11231 10655 11237
rect 10704 11240 11152 11268
rect 9950 11200 9956 11212
rect 7699 11172 8156 11200
rect 8496 11172 9516 11200
rect 7699 11169 7711 11172
rect 7653 11163 7711 11169
rect 8128 11144 8156 11172
rect 9488 11144 9516 11172
rect 9692 11172 9956 11200
rect 7403 11104 7488 11132
rect 7403 11101 7415 11104
rect 7357 11095 7415 11101
rect 7834 11092 7840 11144
rect 7892 11132 7898 11144
rect 8021 11135 8079 11141
rect 8021 11132 8033 11135
rect 7892 11104 8033 11132
rect 7892 11092 7898 11104
rect 8021 11101 8033 11104
rect 8067 11101 8079 11135
rect 8021 11095 8079 11101
rect 8110 11092 8116 11144
rect 8168 11132 8174 11144
rect 8205 11135 8263 11141
rect 8205 11132 8217 11135
rect 8168 11104 8217 11132
rect 8168 11092 8174 11104
rect 8205 11101 8217 11104
rect 8251 11101 8263 11135
rect 8423 11135 8481 11141
rect 8205 11095 8263 11101
rect 8310 11113 8368 11119
rect 8310 11079 8322 11113
rect 8356 11079 8368 11113
rect 8423 11101 8435 11135
rect 8469 11132 8481 11135
rect 8754 11132 8760 11144
rect 8469 11104 8760 11132
rect 8469 11101 8481 11104
rect 8423 11095 8481 11101
rect 8754 11092 8760 11104
rect 8812 11132 8818 11144
rect 9275 11135 9333 11141
rect 9275 11132 9287 11135
rect 8812 11104 9287 11132
rect 8812 11092 8818 11104
rect 9275 11101 9287 11104
rect 9321 11101 9333 11135
rect 9275 11095 9333 11101
rect 9401 11135 9459 11141
rect 9401 11101 9413 11135
rect 9447 11101 9459 11135
rect 9488 11104 9496 11144
rect 9401 11095 9459 11101
rect 5721 11067 5779 11073
rect 5721 11064 5733 11067
rect 5368 11036 5733 11064
rect 5721 11033 5733 11036
rect 5767 11064 5779 11067
rect 5994 11064 6000 11076
rect 5767 11036 6000 11064
rect 5767 11033 5779 11036
rect 5721 11027 5779 11033
rect 5994 11024 6000 11036
rect 6052 11024 6058 11076
rect 7101 11067 7159 11073
rect 7101 11033 7113 11067
rect 7147 11064 7159 11067
rect 7190 11064 7196 11076
rect 7147 11036 7196 11064
rect 7147 11033 7159 11036
rect 7101 11027 7159 11033
rect 7190 11024 7196 11036
rect 7248 11024 7254 11076
rect 8310 11073 8368 11079
rect 2406 10956 2412 11008
rect 2464 10996 2470 11008
rect 7006 10996 7012 11008
rect 2464 10968 7012 10996
rect 2464 10956 2470 10968
rect 7006 10956 7012 10968
rect 7064 10956 7070 11008
rect 7466 10996 7472 11008
rect 7379 10968 7472 10996
rect 7466 10956 7472 10968
rect 7524 10996 7530 11008
rect 8312 10996 8340 11073
rect 9030 11024 9036 11076
rect 9088 11064 9094 11076
rect 9416 11064 9444 11095
rect 9490 11092 9496 11104
rect 9548 11132 9554 11144
rect 9692 11141 9720 11172
rect 9950 11160 9956 11172
rect 10008 11200 10014 11212
rect 10704 11200 10732 11240
rect 11146 11228 11152 11240
rect 11204 11228 11210 11280
rect 12618 11268 12624 11280
rect 12176 11240 12624 11268
rect 10008 11172 10732 11200
rect 10008 11160 10014 11172
rect 10870 11160 10876 11212
rect 10928 11200 10934 11212
rect 11057 11203 11115 11209
rect 11057 11200 11069 11203
rect 10928 11172 11069 11200
rect 10928 11160 10934 11172
rect 11057 11169 11069 11172
rect 11103 11169 11115 11203
rect 11057 11163 11115 11169
rect 11514 11160 11520 11212
rect 11572 11200 11578 11212
rect 11572 11172 11617 11200
rect 11572 11160 11578 11172
rect 9677 11135 9735 11141
rect 9548 11104 9592 11132
rect 9548 11092 9554 11104
rect 9677 11101 9689 11135
rect 9723 11101 9735 11135
rect 10410 11132 10416 11144
rect 10371 11104 10416 11132
rect 9677 11095 9735 11101
rect 10410 11092 10416 11104
rect 10468 11092 10474 11144
rect 10597 11135 10655 11141
rect 10597 11101 10609 11135
rect 10643 11132 10655 11135
rect 10778 11132 10784 11144
rect 10643 11104 10784 11132
rect 10643 11101 10655 11104
rect 10597 11095 10655 11101
rect 10778 11092 10784 11104
rect 10836 11092 10842 11144
rect 10962 11132 10968 11144
rect 10923 11104 10968 11132
rect 10962 11092 10968 11104
rect 11020 11092 11026 11144
rect 11241 11135 11299 11141
rect 11241 11128 11253 11135
rect 11164 11101 11253 11128
rect 11287 11101 11299 11135
rect 11164 11100 11299 11101
rect 10686 11064 10692 11076
rect 9088 11036 9133 11064
rect 9416 11036 10692 11064
rect 9088 11024 9094 11036
rect 9416 10996 9444 11036
rect 10686 11024 10692 11036
rect 10744 11024 10750 11076
rect 7524 10968 9444 10996
rect 7524 10956 7530 10968
rect 10226 10956 10232 11008
rect 10284 10996 10290 11008
rect 11164 10996 11192 11100
rect 11241 11095 11299 11100
rect 11333 11135 11391 11141
rect 11333 11101 11345 11135
rect 11379 11108 11391 11135
rect 11492 11110 11652 11132
rect 11440 11108 11652 11110
rect 11379 11104 11652 11108
rect 11379 11101 11520 11104
rect 11333 11095 11520 11101
rect 11348 11082 11520 11095
rect 11348 11080 11468 11082
rect 11624 11064 11652 11104
rect 11698 11092 11704 11144
rect 11756 11124 11762 11144
rect 12176 11141 12204 11240
rect 12618 11228 12624 11240
rect 12676 11268 12682 11280
rect 14921 11271 14979 11277
rect 12676 11240 14596 11268
rect 12676 11228 12682 11240
rect 12529 11203 12587 11209
rect 12529 11169 12541 11203
rect 12575 11200 12587 11203
rect 12894 11200 12900 11212
rect 12575 11172 12900 11200
rect 12575 11169 12587 11172
rect 12529 11163 12587 11169
rect 12894 11160 12900 11172
rect 12952 11160 12958 11212
rect 13262 11200 13268 11212
rect 13223 11172 13268 11200
rect 13262 11160 13268 11172
rect 13320 11160 13326 11212
rect 14568 11209 14596 11240
rect 14921 11237 14933 11271
rect 14967 11268 14979 11271
rect 15194 11268 15200 11280
rect 14967 11240 15200 11268
rect 14967 11237 14979 11240
rect 14921 11231 14979 11237
rect 15194 11228 15200 11240
rect 15252 11268 15258 11280
rect 15562 11268 15568 11280
rect 15252 11240 15568 11268
rect 15252 11228 15258 11240
rect 15562 11228 15568 11240
rect 15620 11228 15626 11280
rect 15948 11240 17264 11268
rect 14553 11203 14611 11209
rect 13740 11172 14320 11200
rect 11885 11135 11943 11141
rect 11885 11126 11897 11135
rect 11808 11124 11897 11126
rect 11756 11101 11897 11124
rect 11931 11101 11943 11135
rect 12069 11135 12127 11141
rect 12069 11126 12081 11135
rect 11756 11098 11943 11101
rect 11756 11096 11836 11098
rect 11756 11092 11762 11096
rect 11885 11095 11943 11098
rect 11992 11101 12081 11126
rect 12115 11101 12127 11135
rect 11992 11098 12127 11101
rect 11992 11064 12020 11098
rect 12069 11095 12127 11098
rect 12161 11135 12219 11141
rect 12161 11101 12173 11135
rect 12207 11101 12219 11135
rect 12161 11095 12219 11101
rect 12287 11135 12345 11141
rect 12287 11101 12299 11135
rect 12333 11132 12345 11135
rect 12434 11132 12440 11144
rect 12333 11104 12440 11132
rect 12333 11101 12345 11104
rect 12287 11095 12345 11101
rect 12434 11092 12440 11104
rect 12492 11092 12498 11144
rect 11624 11036 12020 11064
rect 12912 11064 12940 11160
rect 13740 11144 13768 11172
rect 13170 11132 13176 11144
rect 13131 11104 13176 11132
rect 13170 11092 13176 11104
rect 13228 11092 13234 11144
rect 13446 11132 13452 11144
rect 13407 11104 13452 11132
rect 13446 11092 13452 11104
rect 13504 11092 13510 11144
rect 13541 11135 13599 11141
rect 13541 11101 13553 11135
rect 13587 11132 13599 11135
rect 13722 11132 13728 11144
rect 13587 11104 13728 11132
rect 13587 11101 13599 11104
rect 13541 11095 13599 11101
rect 13722 11092 13728 11104
rect 13780 11092 13786 11144
rect 14185 11135 14243 11141
rect 14185 11132 14197 11135
rect 13924 11104 14197 11132
rect 13814 11064 13820 11076
rect 12912 11036 13820 11064
rect 10284 10968 11192 10996
rect 10284 10956 10290 10968
rect 11514 10956 11520 11008
rect 11572 10996 11578 11008
rect 11808 10996 11836 11036
rect 13814 11024 13820 11036
rect 13872 11024 13878 11076
rect 11572 10968 11836 10996
rect 11572 10956 11578 10968
rect 12342 10956 12348 11008
rect 12400 10996 12406 11008
rect 12805 10999 12863 11005
rect 12805 10996 12817 10999
rect 12400 10968 12817 10996
rect 12400 10956 12406 10968
rect 12805 10965 12817 10968
rect 12851 10965 12863 10999
rect 12805 10959 12863 10965
rect 13630 10956 13636 11008
rect 13688 10996 13694 11008
rect 13924 10996 13952 11104
rect 14185 11101 14197 11104
rect 14231 11101 14243 11135
rect 14292 11132 14320 11172
rect 14553 11169 14565 11203
rect 14599 11169 14611 11203
rect 14553 11163 14611 11169
rect 14642 11160 14648 11212
rect 14700 11200 14706 11212
rect 14700 11172 15424 11200
rect 14700 11160 14706 11172
rect 14350 11135 14408 11141
rect 14350 11132 14362 11135
rect 14292 11104 14362 11132
rect 14185 11095 14243 11101
rect 14350 11101 14362 11104
rect 14396 11101 14408 11135
rect 14350 11095 14408 11101
rect 14461 11135 14519 11141
rect 14461 11101 14473 11135
rect 14507 11101 14519 11135
rect 14461 11095 14519 11101
rect 14737 11135 14795 11141
rect 14737 11101 14749 11135
rect 14783 11101 14795 11135
rect 14737 11095 14795 11101
rect 14476 11064 14504 11095
rect 14292 11036 14504 11064
rect 14752 11064 14780 11095
rect 14826 11092 14832 11144
rect 14884 11132 14890 11144
rect 15396 11141 15424 11172
rect 15197 11135 15255 11141
rect 15197 11132 15209 11135
rect 14884 11104 15209 11132
rect 14884 11092 14890 11104
rect 15197 11101 15209 11104
rect 15243 11101 15255 11135
rect 15197 11095 15255 11101
rect 15381 11135 15439 11141
rect 15381 11101 15393 11135
rect 15427 11101 15439 11135
rect 15381 11095 15439 11101
rect 15838 11092 15844 11144
rect 15896 11132 15902 11144
rect 15948 11141 15976 11240
rect 17126 11200 17132 11212
rect 17087 11172 17132 11200
rect 17126 11160 17132 11172
rect 17184 11160 17190 11212
rect 17236 11200 17264 11240
rect 17494 11228 17500 11280
rect 17552 11268 17558 11280
rect 17957 11271 18015 11277
rect 17957 11268 17969 11271
rect 17552 11240 17969 11268
rect 17552 11228 17558 11240
rect 17957 11237 17969 11240
rect 18003 11237 18015 11271
rect 17957 11231 18015 11237
rect 17681 11203 17739 11209
rect 17681 11200 17693 11203
rect 17236 11172 17693 11200
rect 17681 11169 17693 11172
rect 17727 11169 17739 11203
rect 17681 11163 17739 11169
rect 15933 11135 15991 11141
rect 15933 11132 15945 11135
rect 15896 11104 15945 11132
rect 15896 11092 15902 11104
rect 15933 11101 15945 11104
rect 15979 11101 15991 11135
rect 16666 11132 16672 11144
rect 16579 11104 16672 11132
rect 15933 11095 15991 11101
rect 16666 11092 16672 11104
rect 16724 11132 16730 11144
rect 17221 11135 17279 11141
rect 17221 11132 17233 11135
rect 16724 11104 17233 11132
rect 16724 11092 16730 11104
rect 17221 11101 17233 11104
rect 17267 11101 17279 11135
rect 17221 11095 17279 11101
rect 18046 11092 18052 11144
rect 18104 11132 18110 11144
rect 18141 11135 18199 11141
rect 18141 11132 18153 11135
rect 18104 11104 18153 11132
rect 18104 11092 18110 11104
rect 18141 11101 18153 11104
rect 18187 11101 18199 11135
rect 18141 11095 18199 11101
rect 15562 11064 15568 11076
rect 14752 11036 15568 11064
rect 14292 11008 14320 11036
rect 15562 11024 15568 11036
rect 15620 11024 15626 11076
rect 16850 11064 16856 11076
rect 16811 11036 16856 11064
rect 16850 11024 16856 11036
rect 16908 11024 16914 11076
rect 13688 10968 13952 10996
rect 13688 10956 13694 10968
rect 14274 10956 14280 11008
rect 14332 10956 14338 11008
rect 1104 10906 18860 10928
rect 1104 10854 8214 10906
rect 8266 10854 8278 10906
rect 8330 10854 8342 10906
rect 8394 10854 8406 10906
rect 8458 10854 8470 10906
rect 8522 10854 16214 10906
rect 16266 10854 16278 10906
rect 16330 10854 16342 10906
rect 16394 10854 16406 10906
rect 16458 10854 16470 10906
rect 16522 10854 18860 10906
rect 1104 10832 18860 10854
rect 8481 10795 8539 10801
rect 5092 10764 8432 10792
rect 1486 10684 1492 10736
rect 1544 10724 1550 10736
rect 1857 10727 1915 10733
rect 1857 10724 1869 10727
rect 1544 10696 1869 10724
rect 1544 10684 1550 10696
rect 1857 10693 1869 10696
rect 1903 10693 1915 10727
rect 1857 10687 1915 10693
rect 2317 10727 2375 10733
rect 2317 10693 2329 10727
rect 2363 10724 2375 10727
rect 2593 10727 2651 10733
rect 2593 10724 2605 10727
rect 2363 10696 2605 10724
rect 2363 10693 2375 10696
rect 2317 10687 2375 10693
rect 2593 10693 2605 10696
rect 2639 10724 2651 10727
rect 2774 10724 2780 10736
rect 2639 10696 2780 10724
rect 2639 10693 2651 10696
rect 2593 10687 2651 10693
rect 2774 10684 2780 10696
rect 2832 10684 2838 10736
rect 3878 10684 3884 10736
rect 3936 10724 3942 10736
rect 5092 10733 5120 10764
rect 4893 10727 4951 10733
rect 4893 10724 4905 10727
rect 3936 10696 4905 10724
rect 3936 10684 3942 10696
rect 4893 10693 4905 10696
rect 4939 10693 4951 10727
rect 4893 10687 4951 10693
rect 5077 10727 5135 10733
rect 5077 10693 5089 10727
rect 5123 10693 5135 10727
rect 5077 10687 5135 10693
rect 5537 10727 5595 10733
rect 5537 10693 5549 10727
rect 5583 10724 5595 10727
rect 5810 10724 5816 10736
rect 5583 10696 5816 10724
rect 5583 10693 5595 10696
rect 5537 10687 5595 10693
rect 5810 10684 5816 10696
rect 5868 10684 5874 10736
rect 6730 10724 6736 10736
rect 6643 10696 6736 10724
rect 6730 10684 6736 10696
rect 6788 10724 6794 10736
rect 7098 10724 7104 10736
rect 6788 10696 7104 10724
rect 6788 10684 6794 10696
rect 7098 10684 7104 10696
rect 7156 10684 7162 10736
rect 8404 10724 8432 10764
rect 8481 10761 8493 10795
rect 8527 10792 8539 10795
rect 8570 10792 8576 10804
rect 8527 10764 8576 10792
rect 8527 10761 8539 10764
rect 8481 10755 8539 10761
rect 8570 10752 8576 10764
rect 8628 10752 8634 10804
rect 12250 10792 12256 10804
rect 8772 10764 12256 10792
rect 8772 10724 8800 10764
rect 12250 10752 12256 10764
rect 12308 10752 12314 10804
rect 14918 10792 14924 10804
rect 13188 10764 14924 10792
rect 13188 10736 13216 10764
rect 14918 10752 14924 10764
rect 14976 10752 14982 10804
rect 15194 10792 15200 10804
rect 15155 10764 15200 10792
rect 15194 10752 15200 10764
rect 15252 10752 15258 10804
rect 15289 10795 15347 10801
rect 15289 10761 15301 10795
rect 15335 10792 15347 10795
rect 15470 10792 15476 10804
rect 15335 10764 15476 10792
rect 15335 10761 15347 10764
rect 15289 10755 15347 10761
rect 10226 10724 10232 10736
rect 8404 10696 8800 10724
rect 9140 10696 10232 10724
rect 2038 10656 2044 10668
rect 1999 10628 2044 10656
rect 2038 10616 2044 10628
rect 2096 10616 2102 10668
rect 2225 10659 2283 10665
rect 2225 10625 2237 10659
rect 2271 10625 2283 10659
rect 2225 10619 2283 10625
rect 3697 10659 3755 10665
rect 3697 10625 3709 10659
rect 3743 10656 3755 10659
rect 4062 10656 4068 10668
rect 3743 10628 4068 10656
rect 3743 10625 3755 10628
rect 3697 10619 3755 10625
rect 2240 10588 2268 10619
rect 4062 10616 4068 10628
rect 4120 10616 4126 10668
rect 5629 10659 5687 10665
rect 5629 10625 5641 10659
rect 5675 10656 5687 10659
rect 5902 10656 5908 10668
rect 5675 10628 5908 10656
rect 5675 10625 5687 10628
rect 5629 10619 5687 10625
rect 5902 10616 5908 10628
rect 5960 10616 5966 10668
rect 6086 10656 6092 10668
rect 6047 10628 6092 10656
rect 6086 10616 6092 10628
rect 6144 10616 6150 10668
rect 7282 10656 7288 10668
rect 7243 10628 7288 10656
rect 7282 10616 7288 10628
rect 7340 10616 7346 10668
rect 7466 10656 7472 10668
rect 7427 10628 7472 10656
rect 7466 10616 7472 10628
rect 7524 10616 7530 10668
rect 7561 10659 7619 10665
rect 7561 10625 7573 10659
rect 7607 10656 7619 10659
rect 7926 10656 7932 10668
rect 7607 10628 7932 10656
rect 7607 10625 7619 10628
rect 7561 10619 7619 10625
rect 7926 10616 7932 10628
rect 7984 10656 7990 10668
rect 8021 10659 8079 10665
rect 8021 10656 8033 10659
rect 7984 10628 8033 10656
rect 7984 10616 7990 10628
rect 8021 10625 8033 10628
rect 8067 10625 8079 10659
rect 8021 10619 8079 10625
rect 8294 10616 8300 10668
rect 8352 10665 8358 10668
rect 8352 10659 8371 10665
rect 8359 10625 8371 10659
rect 8352 10619 8371 10625
rect 8352 10616 8358 10619
rect 8478 10616 8484 10668
rect 8536 10656 8542 10668
rect 9140 10665 9168 10696
rect 10226 10684 10232 10696
rect 10284 10684 10290 10736
rect 10781 10727 10839 10733
rect 10781 10693 10793 10727
rect 10827 10724 10839 10727
rect 11054 10724 11060 10736
rect 10827 10696 11060 10724
rect 10827 10693 10839 10696
rect 10781 10687 10839 10693
rect 11054 10684 11060 10696
rect 11112 10684 11118 10736
rect 12342 10724 12348 10736
rect 11440 10696 12348 10724
rect 11440 10668 11468 10696
rect 12342 10684 12348 10696
rect 12400 10684 12406 10736
rect 12526 10724 12532 10736
rect 12487 10696 12532 10724
rect 12526 10684 12532 10696
rect 12584 10724 12590 10736
rect 13170 10724 13176 10736
rect 12584 10696 13176 10724
rect 12584 10684 12590 10696
rect 13170 10684 13176 10696
rect 13228 10684 13234 10736
rect 13354 10684 13360 10736
rect 13412 10724 13418 10736
rect 13449 10727 13507 10733
rect 13449 10724 13461 10727
rect 13412 10696 13461 10724
rect 13412 10684 13418 10696
rect 13449 10693 13461 10696
rect 13495 10724 13507 10727
rect 13630 10724 13636 10736
rect 13495 10696 13636 10724
rect 13495 10693 13507 10696
rect 13449 10687 13507 10693
rect 13630 10684 13636 10696
rect 13688 10684 13694 10736
rect 13814 10684 13820 10736
rect 13872 10724 13878 10736
rect 14277 10727 14335 10733
rect 14277 10724 14289 10727
rect 13872 10696 14289 10724
rect 13872 10684 13878 10696
rect 14277 10693 14289 10696
rect 14323 10693 14335 10727
rect 14458 10724 14464 10736
rect 14419 10696 14464 10724
rect 14277 10687 14335 10693
rect 14458 10684 14464 10696
rect 14516 10684 14522 10736
rect 15304 10724 15332 10755
rect 15470 10752 15476 10764
rect 15528 10752 15534 10804
rect 16393 10795 16451 10801
rect 16393 10761 16405 10795
rect 16439 10792 16451 10795
rect 16666 10792 16672 10804
rect 16439 10764 16672 10792
rect 16439 10761 16451 10764
rect 16393 10755 16451 10761
rect 16666 10752 16672 10764
rect 16724 10752 16730 10804
rect 15838 10724 15844 10736
rect 14752 10696 15332 10724
rect 15799 10696 15844 10724
rect 8941 10659 8999 10665
rect 8941 10656 8953 10659
rect 8536 10628 8953 10656
rect 8536 10616 8542 10628
rect 8941 10625 8953 10628
rect 8987 10625 8999 10659
rect 8941 10619 8999 10625
rect 9125 10659 9183 10665
rect 9125 10625 9137 10659
rect 9171 10625 9183 10659
rect 9125 10619 9183 10625
rect 9309 10659 9367 10665
rect 9309 10625 9321 10659
rect 9355 10656 9367 10659
rect 9858 10656 9864 10668
rect 9355 10628 9864 10656
rect 9355 10625 9367 10628
rect 9309 10619 9367 10625
rect 9858 10616 9864 10628
rect 9916 10616 9922 10668
rect 9950 10616 9956 10668
rect 10008 10656 10014 10668
rect 10008 10628 10364 10656
rect 10008 10616 10014 10628
rect 2314 10588 2320 10600
rect 2240 10560 2320 10588
rect 2314 10548 2320 10560
rect 2372 10548 2378 10600
rect 3970 10588 3976 10600
rect 3931 10560 3976 10588
rect 3970 10548 3976 10560
rect 4028 10548 4034 10600
rect 4525 10591 4583 10597
rect 4525 10557 4537 10591
rect 4571 10588 4583 10591
rect 4798 10588 4804 10600
rect 4571 10560 4804 10588
rect 4571 10557 4583 10560
rect 4525 10551 4583 10557
rect 4798 10548 4804 10560
rect 4856 10588 4862 10600
rect 10137 10591 10195 10597
rect 4856 10560 7236 10588
rect 4856 10548 4862 10560
rect 3418 10480 3424 10532
rect 3476 10520 3482 10532
rect 3476 10492 4476 10520
rect 3476 10480 3482 10492
rect 3142 10452 3148 10464
rect 3103 10424 3148 10452
rect 3142 10412 3148 10424
rect 3200 10412 3206 10464
rect 3510 10412 3516 10464
rect 3568 10452 3574 10464
rect 3605 10455 3663 10461
rect 3605 10452 3617 10455
rect 3568 10424 3617 10452
rect 3568 10412 3574 10424
rect 3605 10421 3617 10424
rect 3651 10421 3663 10455
rect 4448 10452 4476 10492
rect 6914 10452 6920 10464
rect 4448 10424 6920 10452
rect 3605 10415 3663 10421
rect 6914 10412 6920 10424
rect 6972 10412 6978 10464
rect 7006 10412 7012 10464
rect 7064 10452 7070 10464
rect 7101 10455 7159 10461
rect 7101 10452 7113 10455
rect 7064 10424 7113 10452
rect 7064 10412 7070 10424
rect 7101 10421 7113 10424
rect 7147 10421 7159 10455
rect 7208 10452 7236 10560
rect 8496 10560 9904 10588
rect 8113 10523 8171 10529
rect 8113 10489 8125 10523
rect 8159 10520 8171 10523
rect 8202 10520 8208 10532
rect 8159 10492 8208 10520
rect 8159 10489 8171 10492
rect 8113 10483 8171 10489
rect 8202 10480 8208 10492
rect 8260 10480 8266 10532
rect 8496 10520 8524 10560
rect 8304 10492 8524 10520
rect 8304 10452 8332 10492
rect 9030 10480 9036 10532
rect 9088 10520 9094 10532
rect 9582 10520 9588 10532
rect 9088 10492 9588 10520
rect 9088 10480 9094 10492
rect 9582 10480 9588 10492
rect 9640 10480 9646 10532
rect 9766 10520 9772 10532
rect 9727 10492 9772 10520
rect 9766 10480 9772 10492
rect 9824 10480 9830 10532
rect 9876 10520 9904 10560
rect 10137 10557 10149 10591
rect 10183 10588 10195 10591
rect 10226 10588 10232 10600
rect 10183 10560 10232 10588
rect 10183 10557 10195 10560
rect 10137 10551 10195 10557
rect 10226 10548 10232 10560
rect 10284 10548 10290 10600
rect 10336 10588 10364 10628
rect 10502 10616 10508 10668
rect 10560 10656 10566 10668
rect 10689 10659 10747 10665
rect 10560 10628 10605 10656
rect 10560 10616 10566 10628
rect 10689 10625 10701 10659
rect 10735 10625 10747 10659
rect 10689 10619 10747 10625
rect 10925 10659 10983 10665
rect 10925 10625 10937 10659
rect 10971 10656 10983 10659
rect 11422 10656 11428 10668
rect 10971 10628 11428 10656
rect 10971 10625 10983 10628
rect 10925 10619 10983 10625
rect 10704 10588 10732 10619
rect 11422 10616 11428 10628
rect 11480 10616 11486 10668
rect 11882 10616 11888 10668
rect 11940 10656 11946 10668
rect 11977 10659 12035 10665
rect 11977 10656 11989 10659
rect 11940 10628 11989 10656
rect 11940 10616 11946 10628
rect 11977 10625 11989 10628
rect 12023 10625 12035 10659
rect 12158 10656 12164 10668
rect 12119 10628 12164 10656
rect 11977 10619 12035 10625
rect 12158 10616 12164 10628
rect 12216 10616 12222 10668
rect 12618 10656 12624 10668
rect 12579 10628 12624 10656
rect 12618 10616 12624 10628
rect 12676 10616 12682 10668
rect 12805 10659 12863 10665
rect 12805 10625 12817 10659
rect 12851 10656 12863 10659
rect 13078 10656 13084 10668
rect 12851 10628 13084 10656
rect 12851 10625 12863 10628
rect 12805 10619 12863 10625
rect 13078 10616 13084 10628
rect 13136 10616 13142 10668
rect 13262 10656 13268 10668
rect 13223 10628 13268 10656
rect 13262 10616 13268 10628
rect 13320 10616 13326 10668
rect 14752 10665 14780 10696
rect 15838 10684 15844 10696
rect 15896 10684 15902 10736
rect 17494 10724 17500 10736
rect 17455 10696 17500 10724
rect 17494 10684 17500 10696
rect 17552 10684 17558 10736
rect 18138 10684 18144 10736
rect 18196 10724 18202 10736
rect 18233 10727 18291 10733
rect 18233 10724 18245 10727
rect 18196 10696 18245 10724
rect 18196 10684 18202 10696
rect 18233 10693 18245 10696
rect 18279 10693 18291 10727
rect 18233 10687 18291 10693
rect 14737 10659 14795 10665
rect 14737 10625 14749 10659
rect 14783 10625 14795 10659
rect 14737 10619 14795 10625
rect 15105 10659 15163 10665
rect 15105 10625 15117 10659
rect 15151 10656 15163 10659
rect 15286 10656 15292 10668
rect 15151 10628 15292 10656
rect 15151 10625 15163 10628
rect 15105 10619 15163 10625
rect 15286 10616 15292 10628
rect 15344 10616 15350 10668
rect 15470 10665 15476 10668
rect 15427 10659 15476 10665
rect 15427 10625 15439 10659
rect 15473 10625 15476 10659
rect 15427 10619 15476 10625
rect 15470 10616 15476 10619
rect 15528 10616 15534 10668
rect 15657 10659 15715 10665
rect 15657 10656 15669 10659
rect 15580 10628 15669 10656
rect 11606 10588 11612 10600
rect 10336 10560 11612 10588
rect 11606 10548 11612 10560
rect 11664 10548 11670 10600
rect 11698 10548 11704 10600
rect 11756 10588 11762 10600
rect 13541 10591 13599 10597
rect 13541 10588 13553 10591
rect 11756 10560 13553 10588
rect 11756 10548 11762 10560
rect 13541 10557 13553 10560
rect 13587 10588 13599 10591
rect 14274 10588 14280 10600
rect 13587 10560 14280 10588
rect 13587 10557 13599 10560
rect 13541 10551 13599 10557
rect 14274 10548 14280 10560
rect 14332 10588 14338 10600
rect 14550 10588 14556 10600
rect 14332 10560 14556 10588
rect 14332 10548 14338 10560
rect 14550 10548 14556 10560
rect 14608 10548 14614 10600
rect 11057 10523 11115 10529
rect 11057 10520 11069 10523
rect 9876 10492 11069 10520
rect 11057 10489 11069 10492
rect 11103 10489 11115 10523
rect 11057 10483 11115 10489
rect 11146 10480 11152 10532
rect 11204 10520 11210 10532
rect 12161 10523 12219 10529
rect 12161 10520 12173 10523
rect 11204 10492 12173 10520
rect 11204 10480 11210 10492
rect 12161 10489 12173 10492
rect 12207 10489 12219 10523
rect 12161 10483 12219 10489
rect 12618 10480 12624 10532
rect 12676 10520 12682 10532
rect 12894 10520 12900 10532
rect 12676 10492 12900 10520
rect 12676 10480 12682 10492
rect 12894 10480 12900 10492
rect 12952 10480 12958 10532
rect 7208 10424 8332 10452
rect 7101 10415 7159 10421
rect 8386 10412 8392 10464
rect 8444 10452 8450 10464
rect 8846 10452 8852 10464
rect 8444 10424 8852 10452
rect 8444 10412 8450 10424
rect 8846 10412 8852 10424
rect 8904 10452 8910 10464
rect 9490 10452 9496 10464
rect 8904 10424 9496 10452
rect 8904 10412 8910 10424
rect 9490 10412 9496 10424
rect 9548 10412 9554 10464
rect 9677 10455 9735 10461
rect 9677 10421 9689 10455
rect 9723 10452 9735 10455
rect 9858 10452 9864 10464
rect 9723 10424 9864 10452
rect 9723 10421 9735 10424
rect 9677 10415 9735 10421
rect 9858 10412 9864 10424
rect 9916 10452 9922 10464
rect 10410 10452 10416 10464
rect 9916 10424 10416 10452
rect 9916 10412 9922 10424
rect 10410 10412 10416 10424
rect 10468 10412 10474 10464
rect 10870 10412 10876 10464
rect 10928 10452 10934 10464
rect 12802 10452 12808 10464
rect 10928 10424 12808 10452
rect 10928 10412 10934 10424
rect 12802 10412 12808 10424
rect 12860 10412 12866 10464
rect 13906 10412 13912 10464
rect 13964 10452 13970 10464
rect 14461 10455 14519 10461
rect 14461 10452 14473 10455
rect 13964 10424 14473 10452
rect 13964 10412 13970 10424
rect 14461 10421 14473 10424
rect 14507 10421 14519 10455
rect 14461 10415 14519 10421
rect 15010 10412 15016 10464
rect 15068 10452 15074 10464
rect 15580 10452 15608 10628
rect 15657 10625 15669 10628
rect 15703 10625 15715 10659
rect 15657 10619 15715 10625
rect 16301 10659 16359 10665
rect 16301 10625 16313 10659
rect 16347 10656 16359 10659
rect 18325 10659 18383 10665
rect 18325 10656 18337 10659
rect 16347 10628 18337 10656
rect 16347 10625 16359 10628
rect 16301 10619 16359 10625
rect 18325 10625 18337 10628
rect 18371 10625 18383 10659
rect 18325 10619 18383 10625
rect 16758 10548 16764 10600
rect 16816 10588 16822 10600
rect 16945 10591 17003 10597
rect 16945 10588 16957 10591
rect 16816 10560 16957 10588
rect 16816 10548 16822 10560
rect 16945 10557 16957 10560
rect 16991 10557 17003 10591
rect 16945 10551 17003 10557
rect 17678 10548 17684 10600
rect 17736 10588 17742 10600
rect 17773 10591 17831 10597
rect 17773 10588 17785 10591
rect 17736 10560 17785 10588
rect 17736 10548 17742 10560
rect 17773 10557 17785 10560
rect 17819 10557 17831 10591
rect 17773 10551 17831 10557
rect 17402 10520 17408 10532
rect 17363 10492 17408 10520
rect 17402 10480 17408 10492
rect 17460 10480 17466 10532
rect 15068 10424 15608 10452
rect 15068 10412 15074 10424
rect 1104 10362 18860 10384
rect 1104 10310 4214 10362
rect 4266 10310 4278 10362
rect 4330 10310 4342 10362
rect 4394 10310 4406 10362
rect 4458 10310 4470 10362
rect 4522 10310 12214 10362
rect 12266 10310 12278 10362
rect 12330 10310 12342 10362
rect 12394 10310 12406 10362
rect 12458 10310 12470 10362
rect 12522 10310 18860 10362
rect 1104 10288 18860 10310
rect 3970 10208 3976 10260
rect 4028 10248 4034 10260
rect 5077 10251 5135 10257
rect 5077 10248 5089 10251
rect 4028 10220 5089 10248
rect 4028 10208 4034 10220
rect 5077 10217 5089 10220
rect 5123 10217 5135 10251
rect 11885 10251 11943 10257
rect 5077 10211 5135 10217
rect 5184 10220 11560 10248
rect 3421 10183 3479 10189
rect 3421 10149 3433 10183
rect 3467 10180 3479 10183
rect 3878 10180 3884 10192
rect 3467 10152 3884 10180
rect 3467 10149 3479 10152
rect 3421 10143 3479 10149
rect 3878 10140 3884 10152
rect 3936 10140 3942 10192
rect 3510 10112 3516 10124
rect 3471 10084 3516 10112
rect 3510 10072 3516 10084
rect 3568 10072 3574 10124
rect 3786 10072 3792 10124
rect 3844 10112 3850 10124
rect 5184 10112 5212 10220
rect 7193 10183 7251 10189
rect 7193 10149 7205 10183
rect 7239 10180 7251 10183
rect 11422 10180 11428 10192
rect 7239 10152 11428 10180
rect 7239 10149 7251 10152
rect 7193 10143 7251 10149
rect 11422 10140 11428 10152
rect 11480 10140 11486 10192
rect 3844 10084 5212 10112
rect 3844 10072 3850 10084
rect 5902 10072 5908 10124
rect 5960 10112 5966 10124
rect 6457 10115 6515 10121
rect 5960 10084 6132 10112
rect 5960 10072 5966 10084
rect 2406 10044 2412 10056
rect 2367 10016 2412 10044
rect 2406 10004 2412 10016
rect 2464 10004 2470 10056
rect 2593 10047 2651 10053
rect 2593 10013 2605 10047
rect 2639 10044 2651 10047
rect 2774 10044 2780 10056
rect 2639 10016 2780 10044
rect 2639 10013 2651 10016
rect 2593 10007 2651 10013
rect 2774 10004 2780 10016
rect 2832 10044 2838 10056
rect 2961 10047 3019 10053
rect 2961 10044 2973 10047
rect 2832 10016 2973 10044
rect 2832 10004 2838 10016
rect 2961 10013 2973 10016
rect 3007 10013 3019 10047
rect 4062 10044 4068 10056
rect 4023 10016 4068 10044
rect 2961 10007 3019 10013
rect 4062 10004 4068 10016
rect 4120 10004 4126 10056
rect 4798 10044 4804 10056
rect 4759 10016 4804 10044
rect 4798 10004 4804 10016
rect 4856 10004 4862 10056
rect 5258 10044 5264 10056
rect 5219 10016 5264 10044
rect 5258 10004 5264 10016
rect 5316 10004 5322 10056
rect 5813 10047 5871 10053
rect 5813 10013 5825 10047
rect 5859 10044 5871 10047
rect 5994 10044 6000 10056
rect 5859 10016 6000 10044
rect 5859 10013 5871 10016
rect 5813 10007 5871 10013
rect 5994 10004 6000 10016
rect 6052 10004 6058 10056
rect 6104 10053 6132 10084
rect 6457 10081 6469 10115
rect 6503 10112 6515 10115
rect 7282 10112 7288 10124
rect 6503 10084 7288 10112
rect 6503 10081 6515 10084
rect 6457 10075 6515 10081
rect 7282 10072 7288 10084
rect 7340 10072 7346 10124
rect 7834 10072 7840 10124
rect 7892 10112 7898 10124
rect 7929 10115 7987 10121
rect 7929 10112 7941 10115
rect 7892 10084 7941 10112
rect 7892 10072 7898 10084
rect 7929 10081 7941 10084
rect 7975 10081 7987 10115
rect 8294 10112 8300 10124
rect 7929 10075 7987 10081
rect 8128 10084 8300 10112
rect 6089 10047 6147 10053
rect 6089 10013 6101 10047
rect 6135 10013 6147 10047
rect 6089 10007 6147 10013
rect 6365 10047 6423 10053
rect 6365 10013 6377 10047
rect 6411 10044 6423 10047
rect 7006 10044 7012 10056
rect 6411 10016 6868 10044
rect 6967 10016 7012 10044
rect 6411 10013 6423 10016
rect 6365 10007 6423 10013
rect 2133 9979 2191 9985
rect 2133 9976 2145 9979
rect 1780 9948 2145 9976
rect 1780 9920 1808 9948
rect 2133 9945 2145 9948
rect 2179 9945 2191 9979
rect 2133 9939 2191 9945
rect 3881 9979 3939 9985
rect 3881 9945 3893 9979
rect 3927 9976 3939 9979
rect 4246 9976 4252 9988
rect 3927 9948 4252 9976
rect 3927 9945 3939 9948
rect 3881 9939 3939 9945
rect 4246 9936 4252 9948
rect 4304 9936 4310 9988
rect 6730 9976 6736 9988
rect 5644 9948 6316 9976
rect 6691 9948 6736 9976
rect 1762 9908 1768 9920
rect 1723 9880 1768 9908
rect 1762 9868 1768 9880
rect 1820 9868 1826 9920
rect 2225 9911 2283 9917
rect 2225 9877 2237 9911
rect 2271 9908 2283 9911
rect 2314 9908 2320 9920
rect 2271 9880 2320 9908
rect 2271 9877 2283 9880
rect 2225 9871 2283 9877
rect 2314 9868 2320 9880
rect 2372 9908 2378 9920
rect 3326 9908 3332 9920
rect 2372 9880 3332 9908
rect 2372 9868 2378 9880
rect 3326 9868 3332 9880
rect 3384 9908 3390 9920
rect 5644 9917 5672 9948
rect 5629 9911 5687 9917
rect 5629 9908 5641 9911
rect 3384 9880 5641 9908
rect 3384 9868 3390 9880
rect 5629 9877 5641 9880
rect 5675 9877 5687 9911
rect 6288 9908 6316 9948
rect 6730 9936 6736 9948
rect 6788 9936 6794 9988
rect 6840 9976 6868 10016
rect 7006 10004 7012 10016
rect 7064 10004 7070 10056
rect 8128 10053 8156 10084
rect 8294 10072 8300 10084
rect 8352 10072 8358 10124
rect 8389 10115 8447 10121
rect 8389 10081 8401 10115
rect 8435 10112 8447 10115
rect 8662 10112 8668 10124
rect 8435 10084 8668 10112
rect 8435 10081 8447 10084
rect 8389 10075 8447 10081
rect 8662 10072 8668 10084
rect 8720 10072 8726 10124
rect 9766 10112 9772 10124
rect 9232 10084 9772 10112
rect 8095 10047 8156 10053
rect 8095 10013 8107 10047
rect 8141 10016 8156 10047
rect 8141 10013 8153 10016
rect 8095 10007 8153 10013
rect 8202 10004 8208 10056
rect 8260 10044 8266 10056
rect 8481 10047 8539 10053
rect 8260 10016 8305 10044
rect 8260 10004 8266 10016
rect 8481 10013 8493 10047
rect 8527 10044 8539 10047
rect 8754 10044 8760 10056
rect 8527 10016 8760 10044
rect 8527 10013 8539 10016
rect 8481 10007 8539 10013
rect 8754 10004 8760 10016
rect 8812 10004 8818 10056
rect 9232 10053 9260 10084
rect 9766 10072 9772 10084
rect 9824 10072 9830 10124
rect 10042 10112 10048 10124
rect 10003 10084 10048 10112
rect 10042 10072 10048 10084
rect 10100 10072 10106 10124
rect 10410 10072 10416 10124
rect 10468 10112 10474 10124
rect 10468 10084 10916 10112
rect 10468 10072 10474 10084
rect 9217 10047 9275 10053
rect 9217 10013 9229 10047
rect 9263 10013 9275 10047
rect 9217 10007 9275 10013
rect 9401 10047 9459 10053
rect 9401 10013 9413 10047
rect 9447 10013 9459 10047
rect 9858 10044 9864 10056
rect 9819 10016 9864 10044
rect 9401 10007 9459 10013
rect 8570 9976 8576 9988
rect 6840 9948 8576 9976
rect 8570 9936 8576 9948
rect 8628 9976 8634 9988
rect 9033 9979 9091 9985
rect 9033 9976 9045 9979
rect 8628 9948 9045 9976
rect 8628 9936 8634 9948
rect 9033 9945 9045 9948
rect 9079 9945 9091 9979
rect 9416 9976 9444 10007
rect 9858 10004 9864 10016
rect 9916 10004 9922 10056
rect 10428 10044 10456 10072
rect 10888 10056 10916 10084
rect 11072 10084 11468 10112
rect 9968 10016 10456 10044
rect 10689 10047 10747 10053
rect 9968 9976 9996 10016
rect 10689 10013 10701 10047
rect 10735 10044 10747 10047
rect 10778 10044 10784 10056
rect 10735 10016 10784 10044
rect 10735 10013 10747 10016
rect 10689 10007 10747 10013
rect 10778 10004 10784 10016
rect 10836 10004 10842 10056
rect 10870 10004 10876 10056
rect 10928 10044 10934 10056
rect 10928 10016 10973 10044
rect 10928 10004 10934 10016
rect 11072 9988 11100 10084
rect 11440 10053 11468 10084
rect 11149 10047 11207 10053
rect 11149 10013 11161 10047
rect 11195 10013 11207 10047
rect 11149 10007 11207 10013
rect 11333 10047 11391 10053
rect 11333 10013 11345 10047
rect 11379 10013 11391 10047
rect 11333 10007 11391 10013
rect 11425 10047 11483 10053
rect 11425 10013 11437 10047
rect 11471 10013 11483 10047
rect 11532 10044 11560 10220
rect 11885 10217 11897 10251
rect 11931 10248 11943 10251
rect 11974 10248 11980 10260
rect 11931 10220 11980 10248
rect 11931 10217 11943 10220
rect 11885 10211 11943 10217
rect 11974 10208 11980 10220
rect 12032 10208 12038 10260
rect 12069 10251 12127 10257
rect 12069 10217 12081 10251
rect 12115 10248 12127 10251
rect 13538 10248 13544 10260
rect 12115 10220 13544 10248
rect 12115 10217 12127 10220
rect 12069 10211 12127 10217
rect 13538 10208 13544 10220
rect 13596 10208 13602 10260
rect 14182 10208 14188 10260
rect 14240 10248 14246 10260
rect 14277 10251 14335 10257
rect 14277 10248 14289 10251
rect 14240 10220 14289 10248
rect 14240 10208 14246 10220
rect 14277 10217 14289 10220
rect 14323 10217 14335 10251
rect 18046 10248 18052 10260
rect 18007 10220 18052 10248
rect 14277 10211 14335 10217
rect 18046 10208 18052 10220
rect 18104 10208 18110 10260
rect 12802 10140 12808 10192
rect 12860 10180 12866 10192
rect 13262 10180 13268 10192
rect 12860 10152 13268 10180
rect 12860 10140 12866 10152
rect 13262 10140 13268 10152
rect 13320 10140 13326 10192
rect 14918 10140 14924 10192
rect 14976 10180 14982 10192
rect 14976 10152 15792 10180
rect 14976 10140 14982 10152
rect 14182 10112 14188 10124
rect 12636 10084 14188 10112
rect 12636 10044 12664 10084
rect 14182 10072 14188 10084
rect 14240 10112 14246 10124
rect 15010 10112 15016 10124
rect 14240 10084 14504 10112
rect 14240 10072 14246 10084
rect 11532 10016 12664 10044
rect 12713 10047 12771 10053
rect 11425 10007 11483 10013
rect 12713 10013 12725 10047
rect 12759 10044 12771 10047
rect 12802 10044 12808 10056
rect 12759 10016 12808 10044
rect 12759 10013 12771 10016
rect 12713 10007 12771 10013
rect 10134 9976 10140 9988
rect 9416 9948 9996 9976
rect 10095 9948 10140 9976
rect 9033 9939 9091 9945
rect 10134 9936 10140 9948
rect 10192 9936 10198 9988
rect 10229 9979 10287 9985
rect 10229 9945 10241 9979
rect 10275 9976 10287 9979
rect 11054 9976 11060 9988
rect 10275 9948 11060 9976
rect 10275 9945 10287 9948
rect 10229 9939 10287 9945
rect 11054 9936 11060 9948
rect 11112 9936 11118 9988
rect 6825 9911 6883 9917
rect 6825 9908 6837 9911
rect 6288 9880 6837 9908
rect 5629 9871 5687 9877
rect 6825 9877 6837 9880
rect 6871 9877 6883 9911
rect 6825 9871 6883 9877
rect 7926 9868 7932 9920
rect 7984 9908 7990 9920
rect 9490 9908 9496 9920
rect 7984 9880 9496 9908
rect 7984 9868 7990 9880
rect 9490 9868 9496 9880
rect 9548 9868 9554 9920
rect 9674 9868 9680 9920
rect 9732 9908 9738 9920
rect 10597 9911 10655 9917
rect 10597 9908 10609 9911
rect 9732 9880 10609 9908
rect 9732 9868 9738 9880
rect 10597 9877 10609 9880
rect 10643 9877 10655 9911
rect 10597 9871 10655 9877
rect 10686 9868 10692 9920
rect 10744 9908 10750 9920
rect 11164 9908 11192 10007
rect 11348 9976 11376 10007
rect 12802 10004 12808 10016
rect 12860 10004 12866 10056
rect 13081 10047 13139 10053
rect 13081 10044 13093 10047
rect 13004 10016 13093 10044
rect 11698 9976 11704 9988
rect 11348 9948 11704 9976
rect 11698 9936 11704 9948
rect 11756 9976 11762 9988
rect 12253 9979 12311 9985
rect 12253 9976 12265 9979
rect 11756 9948 12265 9976
rect 11756 9936 11762 9948
rect 12253 9945 12265 9948
rect 12299 9976 12311 9979
rect 12299 9948 12434 9976
rect 12299 9945 12311 9948
rect 12253 9939 12311 9945
rect 11514 9908 11520 9920
rect 10744 9880 11520 9908
rect 10744 9868 10750 9880
rect 11514 9868 11520 9880
rect 11572 9868 11578 9920
rect 12066 9908 12072 9920
rect 12027 9880 12072 9908
rect 12066 9868 12072 9880
rect 12124 9868 12130 9920
rect 12406 9908 12434 9948
rect 12618 9908 12624 9920
rect 12406 9880 12624 9908
rect 12618 9868 12624 9880
rect 12676 9868 12682 9920
rect 13004 9908 13032 10016
rect 13081 10013 13093 10016
rect 13127 10013 13139 10047
rect 13262 10044 13268 10056
rect 13223 10016 13268 10044
rect 13081 10007 13139 10013
rect 13262 10004 13268 10016
rect 13320 10004 13326 10056
rect 13449 10047 13507 10053
rect 13449 10013 13461 10047
rect 13495 10044 13507 10047
rect 13722 10044 13728 10056
rect 13495 10016 13728 10044
rect 13495 10013 13507 10016
rect 13449 10007 13507 10013
rect 13722 10004 13728 10016
rect 13780 10004 13786 10056
rect 14476 10053 14504 10084
rect 14568 10084 15016 10112
rect 14568 10053 14596 10084
rect 15010 10072 15016 10084
rect 15068 10072 15074 10124
rect 15378 10112 15384 10124
rect 15339 10084 15384 10112
rect 15378 10072 15384 10084
rect 15436 10072 15442 10124
rect 14461 10047 14519 10053
rect 14461 10013 14473 10047
rect 14507 10013 14519 10047
rect 14461 10007 14519 10013
rect 14553 10047 14611 10053
rect 14553 10013 14565 10047
rect 14599 10013 14611 10047
rect 14734 10044 14740 10056
rect 14695 10016 14740 10044
rect 14553 10007 14611 10013
rect 14734 10004 14740 10016
rect 14792 10004 14798 10056
rect 14826 10004 14832 10056
rect 14884 10044 14890 10056
rect 15102 10044 15108 10056
rect 14884 10016 14929 10044
rect 15063 10016 15108 10044
rect 14884 10004 14890 10016
rect 15102 10004 15108 10016
rect 15160 10004 15166 10056
rect 15289 10047 15347 10053
rect 15289 10013 15301 10047
rect 15335 10013 15347 10047
rect 15654 10044 15660 10056
rect 15615 10016 15660 10044
rect 15289 10007 15347 10013
rect 14642 9936 14648 9988
rect 14700 9976 14706 9988
rect 15304 9976 15332 10007
rect 15654 10004 15660 10016
rect 15712 10004 15718 10056
rect 15764 10044 15792 10152
rect 18064 10112 18092 10208
rect 17696 10084 18092 10112
rect 17696 10056 17724 10084
rect 16025 10047 16083 10053
rect 16025 10044 16037 10047
rect 15764 10016 16037 10044
rect 16025 10013 16037 10016
rect 16071 10013 16083 10047
rect 16758 10044 16764 10056
rect 16719 10016 16764 10044
rect 16025 10007 16083 10013
rect 16758 10004 16764 10016
rect 16816 10004 16822 10056
rect 17678 10044 17684 10056
rect 17591 10016 17684 10044
rect 17678 10004 17684 10016
rect 17736 10004 17742 10056
rect 18138 10044 18144 10056
rect 18099 10016 18144 10044
rect 18138 10004 18144 10016
rect 18196 10004 18202 10056
rect 14700 9948 16252 9976
rect 14700 9936 14706 9948
rect 13078 9908 13084 9920
rect 13004 9880 13084 9908
rect 13078 9868 13084 9880
rect 13136 9868 13142 9920
rect 13170 9868 13176 9920
rect 13228 9908 13234 9920
rect 16224 9917 16252 9948
rect 16666 9936 16672 9988
rect 16724 9976 16730 9988
rect 17402 9976 17408 9988
rect 16724 9948 17408 9976
rect 16724 9936 16730 9948
rect 17402 9936 17408 9948
rect 17460 9936 17466 9988
rect 13817 9911 13875 9917
rect 13817 9908 13829 9911
rect 13228 9880 13829 9908
rect 13228 9868 13234 9880
rect 13817 9877 13829 9880
rect 13863 9877 13875 9911
rect 13817 9871 13875 9877
rect 16209 9911 16267 9917
rect 16209 9877 16221 9911
rect 16255 9877 16267 9911
rect 16209 9871 16267 9877
rect 1104 9818 18860 9840
rect 1104 9766 8214 9818
rect 8266 9766 8278 9818
rect 8330 9766 8342 9818
rect 8394 9766 8406 9818
rect 8458 9766 8470 9818
rect 8522 9766 16214 9818
rect 16266 9766 16278 9818
rect 16330 9766 16342 9818
rect 16394 9766 16406 9818
rect 16458 9766 16470 9818
rect 16522 9766 18860 9818
rect 1104 9744 18860 9766
rect 2590 9664 2596 9716
rect 2648 9704 2654 9716
rect 3418 9704 3424 9716
rect 2648 9676 3424 9704
rect 2648 9664 2654 9676
rect 3418 9664 3424 9676
rect 3476 9664 3482 9716
rect 3694 9664 3700 9716
rect 3752 9704 3758 9716
rect 3752 9676 11008 9704
rect 3752 9664 3758 9676
rect 3142 9596 3148 9648
rect 3200 9636 3206 9648
rect 5902 9636 5908 9648
rect 3200 9608 5908 9636
rect 3200 9596 3206 9608
rect 5902 9596 5908 9608
rect 5960 9636 5966 9648
rect 8662 9636 8668 9648
rect 5960 9608 6500 9636
rect 5960 9596 5966 9608
rect 2222 9568 2228 9580
rect 2183 9540 2228 9568
rect 2222 9528 2228 9540
rect 2280 9528 2286 9580
rect 2774 9528 2780 9580
rect 2832 9568 2838 9580
rect 4246 9568 4252 9580
rect 2832 9540 2877 9568
rect 4159 9540 4252 9568
rect 2832 9528 2838 9540
rect 4246 9528 4252 9540
rect 4304 9528 4310 9580
rect 5074 9568 5080 9580
rect 5035 9540 5080 9568
rect 5074 9528 5080 9540
rect 5132 9528 5138 9580
rect 5629 9571 5687 9577
rect 5629 9537 5641 9571
rect 5675 9568 5687 9571
rect 5718 9568 5724 9580
rect 5675 9540 5724 9568
rect 5675 9537 5687 9540
rect 5629 9531 5687 9537
rect 5718 9528 5724 9540
rect 5776 9528 5782 9580
rect 6086 9568 6092 9580
rect 6047 9540 6092 9568
rect 6086 9528 6092 9540
rect 6144 9528 6150 9580
rect 6472 9577 6500 9608
rect 7300 9608 8668 9636
rect 6457 9571 6515 9577
rect 6457 9537 6469 9571
rect 6503 9537 6515 9571
rect 6457 9531 6515 9537
rect 7101 9571 7159 9577
rect 7101 9537 7113 9571
rect 7147 9537 7159 9571
rect 7101 9531 7159 9537
rect 4264 9500 4292 9528
rect 5258 9500 5264 9512
rect 4264 9472 5264 9500
rect 5258 9460 5264 9472
rect 5316 9460 5322 9512
rect 5997 9503 6055 9509
rect 5997 9469 6009 9503
rect 6043 9500 6055 9503
rect 7116 9500 7144 9531
rect 7190 9528 7196 9580
rect 7248 9528 7254 9580
rect 7300 9577 7328 9608
rect 8662 9596 8668 9608
rect 8720 9596 8726 9648
rect 9122 9636 9128 9648
rect 9083 9608 9128 9636
rect 9122 9596 9128 9608
rect 9180 9596 9186 9648
rect 10042 9636 10048 9648
rect 9324 9608 10048 9636
rect 7285 9571 7343 9577
rect 7285 9537 7297 9571
rect 7331 9537 7343 9571
rect 7285 9531 7343 9537
rect 7377 9571 7435 9577
rect 7377 9537 7389 9571
rect 7423 9537 7435 9571
rect 7377 9531 7435 9537
rect 8021 9571 8079 9577
rect 8021 9537 8033 9571
rect 8067 9568 8079 9571
rect 8294 9568 8300 9580
rect 8067 9540 8156 9568
rect 8255 9540 8300 9568
rect 8067 9537 8079 9540
rect 8021 9531 8079 9537
rect 6043 9472 7144 9500
rect 7208 9500 7236 9528
rect 7392 9500 7420 9531
rect 7926 9500 7932 9512
rect 7208 9472 7420 9500
rect 7887 9472 7932 9500
rect 6043 9469 6055 9472
rect 5997 9463 6055 9469
rect 3878 9392 3884 9444
rect 3936 9432 3942 9444
rect 4065 9435 4123 9441
rect 4065 9432 4077 9435
rect 3936 9404 4077 9432
rect 3936 9392 3942 9404
rect 4065 9401 4077 9404
rect 4111 9401 4123 9435
rect 7190 9432 7196 9444
rect 7151 9404 7196 9432
rect 4065 9395 4123 9401
rect 7190 9392 7196 9404
rect 7248 9392 7254 9444
rect 2038 9364 2044 9376
rect 1999 9336 2044 9364
rect 2038 9324 2044 9336
rect 2096 9324 2102 9376
rect 4890 9364 4896 9376
rect 4851 9336 4896 9364
rect 4890 9324 4896 9336
rect 4948 9324 4954 9376
rect 6641 9367 6699 9373
rect 6641 9333 6653 9367
rect 6687 9364 6699 9367
rect 6914 9364 6920 9376
rect 6687 9336 6920 9364
rect 6687 9333 6699 9336
rect 6641 9327 6699 9333
rect 6914 9324 6920 9336
rect 6972 9364 6978 9376
rect 7300 9364 7328 9472
rect 7926 9460 7932 9472
rect 7984 9460 7990 9512
rect 8128 9500 8156 9540
rect 8294 9528 8300 9540
rect 8352 9528 8358 9580
rect 8478 9568 8484 9580
rect 8439 9540 8484 9568
rect 8478 9528 8484 9540
rect 8536 9528 8542 9580
rect 8938 9568 8944 9580
rect 8588 9540 8944 9568
rect 8588 9500 8616 9540
rect 8938 9528 8944 9540
rect 8996 9528 9002 9580
rect 9324 9577 9352 9608
rect 10042 9596 10048 9608
rect 10100 9596 10106 9648
rect 10134 9596 10140 9648
rect 10192 9645 10198 9648
rect 10192 9636 10204 9645
rect 10980 9636 11008 9676
rect 11054 9664 11060 9716
rect 11112 9704 11118 9716
rect 11149 9707 11207 9713
rect 11149 9704 11161 9707
rect 11112 9676 11161 9704
rect 11112 9664 11118 9676
rect 11149 9673 11161 9676
rect 11195 9704 11207 9707
rect 11195 9676 12434 9704
rect 11195 9673 11207 9676
rect 11149 9667 11207 9673
rect 11790 9636 11796 9648
rect 10192 9608 10237 9636
rect 10980 9608 11796 9636
rect 10192 9599 10204 9608
rect 10192 9596 10198 9599
rect 11790 9596 11796 9608
rect 11848 9596 11854 9648
rect 12406 9636 12434 9676
rect 13446 9664 13452 9716
rect 13504 9704 13510 9716
rect 13504 9676 14412 9704
rect 13504 9664 13510 9676
rect 13998 9636 14004 9648
rect 12406 9608 14004 9636
rect 13998 9596 14004 9608
rect 14056 9596 14062 9648
rect 9309 9571 9367 9577
rect 9309 9537 9321 9571
rect 9355 9537 9367 9571
rect 9309 9531 9367 9537
rect 9493 9571 9551 9577
rect 9493 9537 9505 9571
rect 9539 9568 9551 9571
rect 9582 9568 9588 9580
rect 9539 9540 9588 9568
rect 9539 9537 9551 9540
rect 9493 9531 9551 9537
rect 9582 9528 9588 9540
rect 9640 9528 9646 9580
rect 9674 9528 9680 9580
rect 9732 9568 9738 9580
rect 9769 9571 9827 9577
rect 9769 9568 9781 9571
rect 9732 9540 9781 9568
rect 9732 9528 9738 9540
rect 9769 9537 9781 9540
rect 9815 9537 9827 9571
rect 9769 9531 9827 9537
rect 10413 9571 10471 9577
rect 10413 9537 10425 9571
rect 10459 9568 10471 9571
rect 10502 9568 10508 9580
rect 10459 9540 10508 9568
rect 10459 9537 10471 9540
rect 10413 9531 10471 9537
rect 10502 9528 10508 9540
rect 10560 9528 10566 9580
rect 10778 9568 10784 9580
rect 10739 9540 10784 9568
rect 10778 9528 10784 9540
rect 10836 9528 10842 9580
rect 10962 9568 10968 9580
rect 10923 9540 10968 9568
rect 10962 9528 10968 9540
rect 11020 9528 11026 9580
rect 11698 9568 11704 9580
rect 11659 9540 11704 9568
rect 11698 9528 11704 9540
rect 11756 9528 11762 9580
rect 11977 9571 12035 9577
rect 11977 9537 11989 9571
rect 12023 9568 12035 9571
rect 12437 9571 12495 9577
rect 12023 9540 12388 9568
rect 12023 9537 12035 9540
rect 11977 9531 12035 9537
rect 8128 9472 8616 9500
rect 8662 9460 8668 9512
rect 8720 9500 8726 9512
rect 11609 9503 11667 9509
rect 11609 9500 11621 9503
rect 8720 9472 11621 9500
rect 8720 9460 8726 9472
rect 11609 9469 11621 9472
rect 11655 9469 11667 9503
rect 11609 9463 11667 9469
rect 11882 9460 11888 9512
rect 11940 9500 11946 9512
rect 12253 9503 12311 9509
rect 12253 9500 12265 9503
rect 11940 9472 12265 9500
rect 11940 9460 11946 9472
rect 12253 9469 12265 9472
rect 12299 9469 12311 9503
rect 12360 9500 12388 9540
rect 12437 9537 12449 9571
rect 12483 9568 12495 9571
rect 12526 9568 12532 9580
rect 12483 9540 12532 9568
rect 12483 9537 12495 9540
rect 12437 9531 12495 9537
rect 12526 9528 12532 9540
rect 12584 9528 12590 9580
rect 12618 9528 12624 9580
rect 12676 9568 12682 9580
rect 12989 9571 13047 9577
rect 12989 9568 13001 9571
rect 12676 9540 13001 9568
rect 12676 9528 12682 9540
rect 12989 9537 13001 9540
rect 13035 9537 13047 9571
rect 13170 9568 13176 9580
rect 13131 9540 13176 9568
rect 12989 9531 13047 9537
rect 13170 9528 13176 9540
rect 13228 9528 13234 9580
rect 13446 9528 13452 9580
rect 13504 9568 13510 9580
rect 13633 9571 13691 9577
rect 13633 9568 13645 9571
rect 13504 9540 13645 9568
rect 13504 9528 13510 9540
rect 13633 9537 13645 9540
rect 13679 9537 13691 9571
rect 13633 9531 13691 9537
rect 13722 9528 13728 9580
rect 13780 9568 13786 9580
rect 14274 9568 14280 9580
rect 13780 9540 14280 9568
rect 13780 9528 13786 9540
rect 14274 9528 14280 9540
rect 14332 9528 14338 9580
rect 14384 9577 14412 9676
rect 14734 9664 14740 9716
rect 14792 9704 14798 9716
rect 14792 9676 15424 9704
rect 14792 9664 14798 9676
rect 15286 9636 15292 9648
rect 15247 9608 15292 9636
rect 15286 9596 15292 9608
rect 15344 9596 15350 9648
rect 15396 9636 15424 9676
rect 16393 9639 16451 9645
rect 15396 9608 15792 9636
rect 14369 9571 14427 9577
rect 14369 9537 14381 9571
rect 14415 9537 14427 9571
rect 14550 9568 14556 9580
rect 14511 9540 14556 9568
rect 14369 9531 14427 9537
rect 14550 9528 14556 9540
rect 14608 9528 14614 9580
rect 15194 9568 15200 9580
rect 15155 9540 15200 9568
rect 15194 9528 15200 9540
rect 15252 9528 15258 9580
rect 15378 9568 15384 9580
rect 15339 9540 15384 9568
rect 15378 9528 15384 9540
rect 15436 9528 15442 9580
rect 15654 9568 15660 9580
rect 15615 9540 15660 9568
rect 15654 9528 15660 9540
rect 15712 9528 15718 9580
rect 15764 9568 15792 9608
rect 16393 9605 16405 9639
rect 16439 9636 16451 9639
rect 16666 9636 16672 9648
rect 16439 9608 16672 9636
rect 16439 9605 16451 9608
rect 16393 9599 16451 9605
rect 16666 9596 16672 9608
rect 16724 9596 16730 9648
rect 16758 9596 16764 9648
rect 16816 9636 16822 9648
rect 16853 9639 16911 9645
rect 16853 9636 16865 9639
rect 16816 9608 16865 9636
rect 16816 9596 16822 9608
rect 16853 9605 16865 9608
rect 16899 9605 16911 9639
rect 17218 9636 17224 9648
rect 17179 9608 17224 9636
rect 16853 9599 16911 9605
rect 17218 9596 17224 9608
rect 17276 9596 17282 9648
rect 17037 9571 17095 9577
rect 17037 9568 17049 9571
rect 15764 9540 17049 9568
rect 17037 9537 17049 9540
rect 17083 9537 17095 9571
rect 17037 9531 17095 9537
rect 17313 9571 17371 9577
rect 17313 9537 17325 9571
rect 17359 9568 17371 9571
rect 17770 9568 17776 9580
rect 17359 9540 17776 9568
rect 17359 9537 17371 9540
rect 17313 9531 17371 9537
rect 17770 9528 17776 9540
rect 17828 9528 17834 9580
rect 13078 9500 13084 9512
rect 12360 9472 13084 9500
rect 12253 9463 12311 9469
rect 13078 9460 13084 9472
rect 13136 9460 13142 9512
rect 13357 9503 13415 9509
rect 13357 9469 13369 9503
rect 13403 9500 13415 9503
rect 13403 9472 14596 9500
rect 13403 9469 13415 9472
rect 13357 9463 13415 9469
rect 12621 9435 12679 9441
rect 8496 9404 12572 9432
rect 6972 9336 7328 9364
rect 7561 9367 7619 9373
rect 6972 9324 6978 9336
rect 7561 9333 7573 9367
rect 7607 9364 7619 9367
rect 8496 9364 8524 9404
rect 7607 9336 8524 9364
rect 7607 9333 7619 9336
rect 7561 9327 7619 9333
rect 8570 9324 8576 9376
rect 8628 9364 8634 9376
rect 8757 9367 8815 9373
rect 8757 9364 8769 9367
rect 8628 9336 8769 9364
rect 8628 9324 8634 9336
rect 8757 9333 8769 9336
rect 8803 9364 8815 9367
rect 9950 9364 9956 9376
rect 8803 9336 9956 9364
rect 8803 9333 8815 9336
rect 8757 9327 8815 9333
rect 9950 9324 9956 9336
rect 10008 9324 10014 9376
rect 10137 9367 10195 9373
rect 10137 9333 10149 9367
rect 10183 9364 10195 9367
rect 10502 9364 10508 9376
rect 10183 9336 10508 9364
rect 10183 9333 10195 9336
rect 10137 9327 10195 9333
rect 10502 9324 10508 9336
rect 10560 9324 10566 9376
rect 12544 9364 12572 9404
rect 12621 9401 12633 9435
rect 12667 9432 12679 9435
rect 12710 9432 12716 9444
rect 12667 9404 12716 9432
rect 12667 9401 12679 9404
rect 12621 9395 12679 9401
rect 12710 9392 12716 9404
rect 12768 9392 12774 9444
rect 12802 9392 12808 9444
rect 12860 9432 12866 9444
rect 13372 9432 13400 9463
rect 14458 9432 14464 9444
rect 12860 9404 13400 9432
rect 14419 9404 14464 9432
rect 12860 9392 12866 9404
rect 14458 9392 14464 9404
rect 14516 9392 14522 9444
rect 14568 9432 14596 9472
rect 16666 9460 16672 9512
rect 16724 9500 16730 9512
rect 17589 9503 17647 9509
rect 17589 9500 17601 9503
rect 16724 9472 17601 9500
rect 16724 9460 16730 9472
rect 17589 9469 17601 9472
rect 17635 9469 17647 9503
rect 18141 9503 18199 9509
rect 18141 9500 18153 9503
rect 17589 9463 17647 9469
rect 17696 9472 18153 9500
rect 14734 9432 14740 9444
rect 14568 9404 14740 9432
rect 14734 9392 14740 9404
rect 14792 9392 14798 9444
rect 15378 9392 15384 9444
rect 15436 9432 15442 9444
rect 15562 9432 15568 9444
rect 15436 9404 15568 9432
rect 15436 9392 15442 9404
rect 15562 9392 15568 9404
rect 15620 9392 15626 9444
rect 16301 9435 16359 9441
rect 16301 9401 16313 9435
rect 16347 9432 16359 9435
rect 17696 9432 17724 9472
rect 18141 9469 18153 9472
rect 18187 9469 18199 9503
rect 18141 9463 18199 9469
rect 18046 9432 18052 9444
rect 16347 9404 17724 9432
rect 18007 9404 18052 9432
rect 16347 9401 16359 9404
rect 16301 9395 16359 9401
rect 18046 9392 18052 9404
rect 18104 9392 18110 9444
rect 13538 9364 13544 9376
rect 12544 9336 13544 9364
rect 13538 9324 13544 9336
rect 13596 9324 13602 9376
rect 13630 9324 13636 9376
rect 13688 9364 13694 9376
rect 13725 9367 13783 9373
rect 13725 9364 13737 9367
rect 13688 9336 13737 9364
rect 13688 9324 13694 9336
rect 13725 9333 13737 9336
rect 13771 9333 13783 9367
rect 13725 9327 13783 9333
rect 13814 9324 13820 9376
rect 13872 9364 13878 9376
rect 16022 9364 16028 9376
rect 13872 9336 16028 9364
rect 13872 9324 13878 9336
rect 16022 9324 16028 9336
rect 16080 9324 16086 9376
rect 1104 9274 18860 9296
rect 1104 9222 4214 9274
rect 4266 9222 4278 9274
rect 4330 9222 4342 9274
rect 4394 9222 4406 9274
rect 4458 9222 4470 9274
rect 4522 9222 12214 9274
rect 12266 9222 12278 9274
rect 12330 9222 12342 9274
rect 12394 9222 12406 9274
rect 12458 9222 12470 9274
rect 12522 9222 18860 9274
rect 1104 9200 18860 9222
rect 3513 9163 3571 9169
rect 3513 9129 3525 9163
rect 3559 9160 3571 9163
rect 5718 9160 5724 9172
rect 3559 9132 5724 9160
rect 3559 9129 3571 9132
rect 3513 9123 3571 9129
rect 5718 9120 5724 9132
rect 5776 9120 5782 9172
rect 7282 9160 7288 9172
rect 7116 9132 7288 9160
rect 5077 9095 5135 9101
rect 5077 9061 5089 9095
rect 5123 9092 5135 9095
rect 5258 9092 5264 9104
rect 5123 9064 5264 9092
rect 5123 9061 5135 9064
rect 5077 9055 5135 9061
rect 5258 9052 5264 9064
rect 5316 9052 5322 9104
rect 6914 9092 6920 9104
rect 6196 9064 6920 9092
rect 2590 8984 2596 9036
rect 2648 9024 2654 9036
rect 6196 9033 6224 9064
rect 6914 9052 6920 9064
rect 6972 9052 6978 9104
rect 7116 9033 7144 9132
rect 7282 9120 7288 9132
rect 7340 9160 7346 9172
rect 9858 9160 9864 9172
rect 7340 9132 9864 9160
rect 7340 9120 7346 9132
rect 9858 9120 9864 9132
rect 9916 9120 9922 9172
rect 10502 9160 10508 9172
rect 10463 9132 10508 9160
rect 10502 9120 10508 9132
rect 10560 9120 10566 9172
rect 10778 9120 10784 9172
rect 10836 9160 10842 9172
rect 11701 9163 11759 9169
rect 11701 9160 11713 9163
rect 10836 9132 11713 9160
rect 10836 9120 10842 9132
rect 11701 9129 11713 9132
rect 11747 9160 11759 9163
rect 12434 9160 12440 9172
rect 11747 9132 12440 9160
rect 11747 9129 11759 9132
rect 11701 9123 11759 9129
rect 12434 9120 12440 9132
rect 12492 9120 12498 9172
rect 13538 9120 13544 9172
rect 13596 9160 13602 9172
rect 13596 9132 16252 9160
rect 13596 9120 13602 9132
rect 7926 9052 7932 9104
rect 7984 9092 7990 9104
rect 8570 9092 8576 9104
rect 7984 9064 8576 9092
rect 7984 9052 7990 9064
rect 8570 9052 8576 9064
rect 8628 9052 8634 9104
rect 9582 9092 9588 9104
rect 9543 9064 9588 9092
rect 9582 9052 9588 9064
rect 9640 9052 9646 9104
rect 9766 9052 9772 9104
rect 9824 9092 9830 9104
rect 10686 9092 10692 9104
rect 9824 9064 10692 9092
rect 9824 9052 9830 9064
rect 10686 9052 10692 9064
rect 10744 9052 10750 9104
rect 10962 9092 10968 9104
rect 10888 9064 10968 9092
rect 3973 9027 4031 9033
rect 3973 9024 3985 9027
rect 2648 8996 3985 9024
rect 2648 8984 2654 8996
rect 3973 8993 3985 8996
rect 4019 9024 4031 9027
rect 5721 9027 5779 9033
rect 5721 9024 5733 9027
rect 4019 8996 5733 9024
rect 4019 8993 4031 8996
rect 3973 8987 4031 8993
rect 5721 8993 5733 8996
rect 5767 8993 5779 9027
rect 5721 8987 5779 8993
rect 6181 9027 6239 9033
rect 6181 8993 6193 9027
rect 6227 8993 6239 9027
rect 6181 8987 6239 8993
rect 7101 9027 7159 9033
rect 7101 8993 7113 9027
rect 7147 8993 7159 9027
rect 8662 9024 8668 9036
rect 7101 8987 7159 8993
rect 8036 8996 8668 9024
rect 2038 8956 2044 8968
rect 1999 8928 2044 8956
rect 2038 8916 2044 8928
rect 2096 8916 2102 8968
rect 4893 8959 4951 8965
rect 4893 8956 4905 8959
rect 4448 8928 4905 8956
rect 1486 8888 1492 8900
rect 1447 8860 1492 8888
rect 1486 8848 1492 8860
rect 1544 8848 1550 8900
rect 4154 8848 4160 8900
rect 4212 8888 4218 8900
rect 4448 8897 4476 8928
rect 4893 8925 4905 8928
rect 4939 8925 4951 8959
rect 5994 8956 6000 8968
rect 5955 8928 6000 8956
rect 4893 8919 4951 8925
rect 5994 8916 6000 8928
rect 6052 8916 6058 8968
rect 6822 8956 6828 8968
rect 6783 8928 6828 8956
rect 6822 8916 6828 8928
rect 6880 8916 6886 8968
rect 7190 8916 7196 8968
rect 7248 8956 7254 8968
rect 7469 8959 7527 8965
rect 7248 8928 7293 8956
rect 7248 8916 7254 8928
rect 7469 8925 7481 8959
rect 7515 8956 7527 8959
rect 7650 8956 7656 8968
rect 7515 8928 7656 8956
rect 7515 8925 7527 8928
rect 7469 8919 7527 8925
rect 7650 8916 7656 8928
rect 7708 8916 7714 8968
rect 7742 8916 7748 8968
rect 7800 8956 7806 8968
rect 8036 8965 8064 8996
rect 8662 8984 8668 8996
rect 8720 8984 8726 9036
rect 10888 9024 10916 9064
rect 10962 9052 10968 9064
rect 11020 9052 11026 9104
rect 12161 9095 12219 9101
rect 12161 9061 12173 9095
rect 12207 9092 12219 9095
rect 12526 9092 12532 9104
rect 12207 9064 12532 9092
rect 12207 9061 12219 9064
rect 12161 9055 12219 9061
rect 12526 9052 12532 9064
rect 12584 9092 12590 9104
rect 13078 9092 13084 9104
rect 12584 9064 13084 9092
rect 12584 9052 12590 9064
rect 13078 9052 13084 9064
rect 13136 9052 13142 9104
rect 14274 9052 14280 9104
rect 14332 9092 14338 9104
rect 14369 9095 14427 9101
rect 14369 9092 14381 9095
rect 14332 9064 14381 9092
rect 14332 9052 14338 9064
rect 14369 9061 14381 9064
rect 14415 9061 14427 9095
rect 14369 9055 14427 9061
rect 14458 9052 14464 9104
rect 14516 9052 14522 9104
rect 14737 9095 14795 9101
rect 14737 9061 14749 9095
rect 14783 9092 14795 9095
rect 15657 9095 15715 9101
rect 14783 9064 15608 9092
rect 14783 9061 14795 9064
rect 14737 9055 14795 9061
rect 9416 8996 11008 9024
rect 9416 8968 9444 8996
rect 8021 8959 8079 8965
rect 7800 8928 7845 8956
rect 7800 8916 7806 8928
rect 8021 8925 8033 8959
rect 8067 8925 8079 8959
rect 8021 8919 8079 8925
rect 8481 8959 8539 8965
rect 8481 8925 8493 8959
rect 8527 8925 8539 8959
rect 9398 8956 9404 8968
rect 9359 8928 9404 8956
rect 8481 8919 8539 8925
rect 4433 8891 4491 8897
rect 4433 8888 4445 8891
rect 4212 8860 4445 8888
rect 4212 8848 4218 8860
rect 4433 8857 4445 8860
rect 4479 8857 4491 8891
rect 4433 8851 4491 8857
rect 4525 8891 4583 8897
rect 4525 8857 4537 8891
rect 4571 8888 4583 8891
rect 5442 8888 5448 8900
rect 4571 8860 5448 8888
rect 4571 8857 4583 8860
rect 4525 8851 4583 8857
rect 5442 8848 5448 8860
rect 5500 8848 5506 8900
rect 5626 8888 5632 8900
rect 5587 8860 5632 8888
rect 5626 8848 5632 8860
rect 5684 8848 5690 8900
rect 8496 8888 8524 8919
rect 9398 8916 9404 8928
rect 9456 8916 9462 8968
rect 9490 8916 9496 8968
rect 9548 8956 9554 8968
rect 9585 8959 9643 8965
rect 9585 8956 9597 8959
rect 9548 8928 9597 8956
rect 9548 8916 9554 8928
rect 9585 8925 9597 8928
rect 9631 8956 9643 8959
rect 10594 8956 10600 8968
rect 9631 8928 10600 8956
rect 9631 8925 9643 8928
rect 9585 8919 9643 8925
rect 10594 8916 10600 8928
rect 10652 8916 10658 8968
rect 10980 8965 11008 8996
rect 11808 8996 12388 9024
rect 10689 8959 10747 8965
rect 10689 8925 10701 8959
rect 10735 8925 10747 8959
rect 10689 8919 10747 8925
rect 10780 8959 10838 8965
rect 10780 8925 10792 8959
rect 10826 8925 10838 8959
rect 10780 8919 10838 8925
rect 10936 8959 11008 8965
rect 10936 8925 10948 8959
rect 10982 8928 11008 8959
rect 11069 8959 11127 8965
rect 10982 8925 10994 8928
rect 10936 8919 10994 8925
rect 11069 8925 11081 8959
rect 11115 8956 11127 8959
rect 11698 8956 11704 8968
rect 11115 8928 11704 8956
rect 11115 8925 11127 8928
rect 11069 8919 11127 8925
rect 9766 8888 9772 8900
rect 8496 8860 9772 8888
rect 9766 8848 9772 8860
rect 9824 8848 9830 8900
rect 9953 8891 10011 8897
rect 9953 8857 9965 8891
rect 9999 8857 10011 8891
rect 9953 8851 10011 8857
rect 6641 8823 6699 8829
rect 6641 8789 6653 8823
rect 6687 8820 6699 8823
rect 7558 8820 7564 8832
rect 6687 8792 7564 8820
rect 6687 8789 6699 8792
rect 6641 8783 6699 8789
rect 7558 8780 7564 8792
rect 7616 8780 7622 8832
rect 7834 8820 7840 8832
rect 7795 8792 7840 8820
rect 7834 8780 7840 8792
rect 7892 8780 7898 8832
rect 8570 8820 8576 8832
rect 8531 8792 8576 8820
rect 8570 8780 8576 8792
rect 8628 8780 8634 8832
rect 8662 8780 8668 8832
rect 8720 8820 8726 8832
rect 9582 8820 9588 8832
rect 8720 8792 9588 8820
rect 8720 8780 8726 8792
rect 9582 8780 9588 8792
rect 9640 8780 9646 8832
rect 9968 8820 9996 8851
rect 10502 8848 10508 8900
rect 10560 8888 10566 8900
rect 10704 8888 10732 8919
rect 10560 8860 10732 8888
rect 10560 8848 10566 8860
rect 10795 8820 10823 8919
rect 11698 8916 11704 8928
rect 11756 8916 11762 8968
rect 11808 8965 11836 8996
rect 11793 8959 11851 8965
rect 11793 8925 11805 8959
rect 11839 8925 11851 8959
rect 12158 8956 12164 8968
rect 12119 8928 12164 8956
rect 11793 8919 11851 8925
rect 11808 8820 11836 8919
rect 12158 8916 12164 8928
rect 12216 8916 12222 8968
rect 12360 8965 12388 8996
rect 12434 8984 12440 9036
rect 12492 9024 12498 9036
rect 12986 9024 12992 9036
rect 12492 8996 12992 9024
rect 12492 8984 12498 8996
rect 12986 8984 12992 8996
rect 13044 9024 13050 9036
rect 14476 9024 14504 9052
rect 15580 9024 15608 9064
rect 15657 9061 15669 9095
rect 15703 9092 15715 9095
rect 16114 9092 16120 9104
rect 15703 9064 16120 9092
rect 15703 9061 15715 9064
rect 15657 9055 15715 9061
rect 16114 9052 16120 9064
rect 16172 9052 16178 9104
rect 13044 8996 13400 9024
rect 14476 8996 15148 9024
rect 15580 8996 16160 9024
rect 13044 8984 13050 8996
rect 12345 8959 12403 8965
rect 12345 8925 12357 8959
rect 12391 8956 12403 8959
rect 12802 8956 12808 8968
rect 12391 8928 12808 8956
rect 12391 8925 12403 8928
rect 12345 8919 12403 8925
rect 12802 8916 12808 8928
rect 12860 8916 12866 8968
rect 13078 8956 13084 8968
rect 13039 8928 13084 8956
rect 13078 8916 13084 8928
rect 13136 8916 13142 8968
rect 13372 8965 13400 8996
rect 13173 8959 13231 8965
rect 13173 8925 13185 8959
rect 13219 8925 13231 8959
rect 13173 8919 13231 8925
rect 13265 8959 13323 8965
rect 13265 8925 13277 8959
rect 13311 8925 13323 8959
rect 13265 8919 13323 8925
rect 13357 8959 13415 8965
rect 13357 8925 13369 8959
rect 13403 8956 13415 8959
rect 13446 8956 13452 8968
rect 13403 8928 13452 8956
rect 13403 8925 13415 8928
rect 13357 8919 13415 8925
rect 11882 8848 11888 8900
rect 11940 8888 11946 8900
rect 13188 8888 13216 8919
rect 11940 8860 13216 8888
rect 11940 8848 11946 8860
rect 9968 8792 11836 8820
rect 12710 8780 12716 8832
rect 12768 8820 12774 8832
rect 13280 8820 13308 8919
rect 13446 8916 13452 8928
rect 13504 8956 13510 8968
rect 13998 8956 14004 8968
rect 13504 8928 14004 8956
rect 13504 8916 13510 8928
rect 13998 8916 14004 8928
rect 14056 8916 14062 8968
rect 14090 8916 14096 8968
rect 14148 8956 14154 8968
rect 14277 8959 14335 8965
rect 14277 8956 14289 8959
rect 14148 8928 14289 8956
rect 14148 8916 14154 8928
rect 14277 8925 14289 8928
rect 14323 8925 14335 8959
rect 14277 8919 14335 8925
rect 14461 8959 14519 8965
rect 14461 8925 14473 8959
rect 14507 8925 14519 8959
rect 14461 8919 14519 8925
rect 13630 8848 13636 8900
rect 13688 8888 13694 8900
rect 14476 8888 14504 8919
rect 14550 8916 14556 8968
rect 14608 8956 14614 8968
rect 15120 8965 15148 8996
rect 15562 8965 15568 8968
rect 15105 8959 15163 8965
rect 14608 8928 14653 8956
rect 14608 8916 14614 8928
rect 15105 8925 15117 8959
rect 15151 8925 15163 8959
rect 15105 8919 15163 8925
rect 15525 8959 15568 8965
rect 15525 8925 15537 8959
rect 15620 8956 15626 8968
rect 16025 8959 16083 8965
rect 16025 8956 16037 8959
rect 15620 8928 16037 8956
rect 15525 8919 15568 8925
rect 15562 8916 15568 8919
rect 15620 8916 15626 8928
rect 16025 8925 16037 8928
rect 16071 8925 16083 8959
rect 16025 8919 16083 8925
rect 15289 8891 15347 8897
rect 15289 8888 15301 8891
rect 13688 8860 14504 8888
rect 14568 8860 15301 8888
rect 13688 8848 13694 8860
rect 12768 8792 13308 8820
rect 13541 8823 13599 8829
rect 12768 8780 12774 8792
rect 13541 8789 13553 8823
rect 13587 8820 13599 8823
rect 13814 8820 13820 8832
rect 13587 8792 13820 8820
rect 13587 8789 13599 8792
rect 13541 8783 13599 8789
rect 13814 8780 13820 8792
rect 13872 8780 13878 8832
rect 14090 8780 14096 8832
rect 14148 8820 14154 8832
rect 14568 8820 14596 8860
rect 15289 8857 15301 8860
rect 15335 8857 15347 8891
rect 15289 8851 15347 8857
rect 15381 8891 15439 8897
rect 15381 8857 15393 8891
rect 15427 8857 15439 8891
rect 16132 8888 16160 8996
rect 16224 8956 16252 9132
rect 18046 9052 18052 9104
rect 18104 9092 18110 9104
rect 18141 9095 18199 9101
rect 18141 9092 18153 9095
rect 18104 9064 18153 9092
rect 18104 9052 18110 9064
rect 18141 9061 18153 9064
rect 18187 9061 18199 9095
rect 18141 9055 18199 9061
rect 16666 8956 16672 8968
rect 16224 8928 16672 8956
rect 16666 8916 16672 8928
rect 16724 8916 16730 8968
rect 17678 8956 17684 8968
rect 17639 8928 17684 8956
rect 17678 8916 17684 8928
rect 17736 8916 17742 8968
rect 16942 8888 16948 8900
rect 16132 8860 16948 8888
rect 15381 8851 15439 8857
rect 14148 8792 14596 8820
rect 14148 8780 14154 8792
rect 15010 8780 15016 8832
rect 15068 8820 15074 8832
rect 15396 8820 15424 8851
rect 16942 8848 16948 8860
rect 17000 8848 17006 8900
rect 15470 8820 15476 8832
rect 15068 8792 15476 8820
rect 15068 8780 15074 8792
rect 15470 8780 15476 8792
rect 15528 8780 15534 8832
rect 1104 8730 18860 8752
rect 1104 8678 8214 8730
rect 8266 8678 8278 8730
rect 8330 8678 8342 8730
rect 8394 8678 8406 8730
rect 8458 8678 8470 8730
rect 8522 8678 16214 8730
rect 16266 8678 16278 8730
rect 16330 8678 16342 8730
rect 16394 8678 16406 8730
rect 16458 8678 16470 8730
rect 16522 8678 18860 8730
rect 1104 8656 18860 8678
rect 6086 8616 6092 8628
rect 5999 8588 6092 8616
rect 4154 8548 4160 8560
rect 4115 8520 4160 8548
rect 4154 8508 4160 8520
rect 4212 8508 4218 8560
rect 4433 8551 4491 8557
rect 4433 8517 4445 8551
rect 4479 8548 4491 8551
rect 5074 8548 5080 8560
rect 4479 8520 5080 8548
rect 4479 8517 4491 8520
rect 4433 8511 4491 8517
rect 2590 8480 2596 8492
rect 2551 8452 2596 8480
rect 2590 8440 2596 8452
rect 2648 8440 2654 8492
rect 4065 8483 4123 8489
rect 4065 8449 4077 8483
rect 4111 8480 4123 8483
rect 4448 8480 4476 8511
rect 5074 8508 5080 8520
rect 5132 8508 5138 8560
rect 5626 8508 5632 8560
rect 5684 8548 5690 8560
rect 5721 8551 5779 8557
rect 5721 8548 5733 8551
rect 5684 8520 5733 8548
rect 5684 8508 5690 8520
rect 5721 8517 5733 8520
rect 5767 8517 5779 8551
rect 5721 8511 5779 8517
rect 4614 8480 4620 8492
rect 4111 8452 4476 8480
rect 4575 8452 4620 8480
rect 4111 8449 4123 8452
rect 4065 8443 4123 8449
rect 4614 8440 4620 8452
rect 4672 8440 4678 8492
rect 5350 8480 5356 8492
rect 5311 8452 5356 8480
rect 5350 8440 5356 8452
rect 5408 8440 5414 8492
rect 6012 8489 6040 8588
rect 6086 8576 6092 8588
rect 6144 8616 6150 8628
rect 6638 8616 6644 8628
rect 6144 8588 6644 8616
rect 6144 8576 6150 8588
rect 6638 8576 6644 8588
rect 6696 8576 6702 8628
rect 7745 8619 7803 8625
rect 7745 8616 7757 8619
rect 6748 8588 7757 8616
rect 6748 8548 6776 8588
rect 7745 8585 7757 8588
rect 7791 8616 7803 8619
rect 7926 8616 7932 8628
rect 7791 8588 7932 8616
rect 7791 8585 7803 8588
rect 7745 8579 7803 8585
rect 7926 8576 7932 8588
rect 7984 8576 7990 8628
rect 9398 8616 9404 8628
rect 9048 8588 9404 8616
rect 6472 8520 6776 8548
rect 6472 8489 6500 8520
rect 6822 8508 6828 8560
rect 6880 8548 6886 8560
rect 7650 8548 7656 8560
rect 6880 8520 7236 8548
rect 6880 8508 6886 8520
rect 5813 8483 5871 8489
rect 5813 8449 5825 8483
rect 5859 8449 5871 8483
rect 5813 8443 5871 8449
rect 5997 8483 6055 8489
rect 5997 8449 6009 8483
rect 6043 8449 6055 8483
rect 5997 8443 6055 8449
rect 6457 8483 6515 8489
rect 6457 8449 6469 8483
rect 6503 8449 6515 8483
rect 6457 8443 6515 8449
rect 7101 8483 7159 8489
rect 7101 8449 7113 8483
rect 7147 8449 7159 8483
rect 7101 8443 7159 8449
rect 3970 8372 3976 8424
rect 4028 8412 4034 8424
rect 5534 8412 5540 8424
rect 4028 8384 5540 8412
rect 4028 8372 4034 8384
rect 5534 8372 5540 8384
rect 5592 8412 5598 8424
rect 5828 8412 5856 8443
rect 5592 8384 5856 8412
rect 5592 8372 5598 8384
rect 5902 8372 5908 8424
rect 5960 8412 5966 8424
rect 6472 8412 6500 8443
rect 5960 8384 6500 8412
rect 5960 8372 5966 8384
rect 6638 8304 6644 8356
rect 6696 8344 6702 8356
rect 7116 8344 7144 8443
rect 7208 8412 7236 8520
rect 7484 8520 7656 8548
rect 7285 8483 7343 8489
rect 7285 8449 7297 8483
rect 7331 8480 7343 8483
rect 7484 8480 7512 8520
rect 7650 8508 7656 8520
rect 7708 8548 7714 8560
rect 8662 8548 8668 8560
rect 7708 8520 8668 8548
rect 7708 8508 7714 8520
rect 8662 8508 8668 8520
rect 8720 8508 8726 8560
rect 7331 8452 7512 8480
rect 7331 8449 7343 8452
rect 7285 8443 7343 8449
rect 7558 8440 7564 8492
rect 7616 8480 7622 8492
rect 8018 8480 8024 8492
rect 7616 8452 8024 8480
rect 7616 8440 7622 8452
rect 8018 8440 8024 8452
rect 8076 8480 8082 8492
rect 8297 8483 8355 8489
rect 8297 8480 8309 8483
rect 8076 8452 8309 8480
rect 8076 8440 8082 8452
rect 8297 8449 8309 8452
rect 8343 8449 8355 8483
rect 8297 8443 8355 8449
rect 8481 8483 8539 8489
rect 8481 8449 8493 8483
rect 8527 8480 8539 8483
rect 8846 8480 8852 8492
rect 8527 8452 8852 8480
rect 8527 8449 8539 8452
rect 8481 8443 8539 8449
rect 7469 8415 7527 8421
rect 7469 8412 7481 8415
rect 7208 8384 7481 8412
rect 7469 8381 7481 8384
rect 7515 8412 7527 8415
rect 7742 8412 7748 8424
rect 7515 8384 7748 8412
rect 7515 8381 7527 8384
rect 7469 8375 7527 8381
rect 7742 8372 7748 8384
rect 7800 8372 7806 8424
rect 8110 8412 8116 8424
rect 8071 8384 8116 8412
rect 8110 8372 8116 8384
rect 8168 8372 8174 8424
rect 8312 8412 8340 8443
rect 8846 8440 8852 8452
rect 8904 8440 8910 8492
rect 8938 8440 8944 8492
rect 8996 8480 9002 8492
rect 9048 8489 9076 8588
rect 9398 8576 9404 8588
rect 9456 8616 9462 8628
rect 9456 8588 9904 8616
rect 9456 8576 9462 8588
rect 9674 8548 9680 8560
rect 9324 8520 9680 8548
rect 9324 8489 9352 8520
rect 9674 8508 9680 8520
rect 9732 8508 9738 8560
rect 9033 8483 9091 8489
rect 9033 8480 9045 8483
rect 8996 8452 9045 8480
rect 8996 8440 9002 8452
rect 9033 8449 9045 8452
rect 9079 8449 9091 8483
rect 9033 8443 9091 8449
rect 9309 8483 9367 8489
rect 9309 8449 9321 8483
rect 9355 8449 9367 8483
rect 9309 8443 9367 8449
rect 9585 8483 9643 8489
rect 9585 8449 9597 8483
rect 9631 8449 9643 8483
rect 9766 8480 9772 8492
rect 9727 8452 9772 8480
rect 9585 8443 9643 8449
rect 9490 8412 9496 8424
rect 8312 8384 9496 8412
rect 9490 8372 9496 8384
rect 9548 8372 9554 8424
rect 9600 8412 9628 8443
rect 9766 8440 9772 8452
rect 9824 8440 9830 8492
rect 9876 8480 9904 8588
rect 10134 8576 10140 8628
rect 10192 8616 10198 8628
rect 12805 8619 12863 8625
rect 10192 8588 12756 8616
rect 10192 8576 10198 8588
rect 9950 8508 9956 8560
rect 10008 8548 10014 8560
rect 10873 8551 10931 8557
rect 10008 8520 10640 8548
rect 10008 8508 10014 8520
rect 10045 8483 10103 8489
rect 10045 8480 10057 8483
rect 9876 8452 10057 8480
rect 10045 8449 10057 8452
rect 10091 8449 10103 8483
rect 10318 8480 10324 8492
rect 10279 8452 10324 8480
rect 10045 8443 10103 8449
rect 10318 8440 10324 8452
rect 10376 8440 10382 8492
rect 10410 8440 10416 8492
rect 10468 8480 10474 8492
rect 10612 8480 10640 8520
rect 10873 8517 10885 8551
rect 10919 8548 10931 8551
rect 12250 8548 12256 8560
rect 10919 8520 12256 8548
rect 10919 8517 10931 8520
rect 10873 8511 10931 8517
rect 12250 8508 12256 8520
rect 12308 8508 12314 8560
rect 12728 8548 12756 8588
rect 12805 8585 12817 8619
rect 12851 8616 12863 8619
rect 15102 8616 15108 8628
rect 12851 8588 15108 8616
rect 12851 8585 12863 8588
rect 12805 8579 12863 8585
rect 15102 8576 15108 8588
rect 15160 8576 15166 8628
rect 15194 8576 15200 8628
rect 15252 8616 15258 8628
rect 15252 8588 16068 8616
rect 15252 8576 15258 8588
rect 12728 8520 13382 8548
rect 13354 8511 13382 8520
rect 13354 8505 13414 8511
rect 13906 8508 13912 8560
rect 13964 8548 13970 8560
rect 14369 8551 14427 8557
rect 13964 8520 14228 8548
rect 13964 8508 13970 8520
rect 11149 8483 11207 8489
rect 11149 8480 11161 8483
rect 10468 8452 10513 8480
rect 10612 8452 11161 8480
rect 10468 8440 10474 8452
rect 11149 8449 11161 8452
rect 11195 8480 11207 8483
rect 11885 8483 11943 8489
rect 11885 8480 11897 8483
rect 11195 8452 11897 8480
rect 11195 8449 11207 8452
rect 11149 8443 11207 8449
rect 11885 8449 11897 8452
rect 11931 8480 11943 8483
rect 12345 8483 12403 8489
rect 11931 8452 12296 8480
rect 11931 8449 11943 8452
rect 11885 8443 11943 8449
rect 9858 8412 9864 8424
rect 9600 8384 9864 8412
rect 9858 8372 9864 8384
rect 9916 8372 9922 8424
rect 10226 8372 10232 8424
rect 10284 8412 10290 8424
rect 12158 8412 12164 8424
rect 10284 8384 12164 8412
rect 10284 8372 10290 8384
rect 10428 8356 10456 8384
rect 12158 8372 12164 8384
rect 12216 8372 12222 8424
rect 12268 8412 12296 8452
rect 12345 8449 12357 8483
rect 12391 8480 12403 8483
rect 12434 8480 12440 8492
rect 12391 8452 12440 8480
rect 12391 8449 12403 8452
rect 12345 8443 12403 8449
rect 12434 8440 12440 8452
rect 12492 8440 12498 8492
rect 13170 8480 13176 8492
rect 12544 8452 13176 8480
rect 12544 8412 12572 8452
rect 13170 8440 13176 8452
rect 13228 8440 13234 8492
rect 13354 8474 13368 8505
rect 13356 8471 13368 8474
rect 13402 8471 13414 8505
rect 13541 8483 13599 8489
rect 13356 8465 13414 8471
rect 13448 8473 13506 8479
rect 12268 8384 12572 8412
rect 7190 8344 7196 8356
rect 6696 8316 7196 8344
rect 6696 8304 6702 8316
rect 7190 8304 7196 8316
rect 7248 8344 7254 8356
rect 10134 8344 10140 8356
rect 7248 8316 10140 8344
rect 7248 8304 7254 8316
rect 10134 8304 10140 8316
rect 10192 8304 10198 8356
rect 10410 8304 10416 8356
rect 10468 8304 10474 8356
rect 11146 8304 11152 8356
rect 11204 8344 11210 8356
rect 11698 8344 11704 8356
rect 11204 8316 11704 8344
rect 11204 8304 11210 8316
rect 11698 8304 11704 8316
rect 11756 8304 11762 8356
rect 12894 8304 12900 8356
rect 12952 8344 12958 8356
rect 13081 8347 13139 8353
rect 13081 8344 13093 8347
rect 12952 8316 13093 8344
rect 12952 8304 12958 8316
rect 13081 8313 13093 8316
rect 13127 8313 13139 8347
rect 13081 8307 13139 8313
rect 1854 8276 1860 8288
rect 1815 8248 1860 8276
rect 1854 8236 1860 8248
rect 1912 8236 1918 8288
rect 9214 8276 9220 8288
rect 9175 8248 9220 8276
rect 9214 8236 9220 8248
rect 9272 8236 9278 8288
rect 9582 8236 9588 8288
rect 9640 8276 9646 8288
rect 11514 8276 11520 8288
rect 9640 8248 11520 8276
rect 9640 8236 9646 8248
rect 11514 8236 11520 8248
rect 11572 8236 11578 8288
rect 11974 8236 11980 8288
rect 12032 8276 12038 8288
rect 12253 8279 12311 8285
rect 12253 8276 12265 8279
rect 12032 8248 12265 8276
rect 12032 8236 12038 8248
rect 12253 8245 12265 8248
rect 12299 8245 12311 8279
rect 13372 8276 13400 8465
rect 13448 8439 13460 8473
rect 13494 8439 13506 8473
rect 13541 8449 13553 8483
rect 13587 8449 13599 8483
rect 13541 8443 13599 8449
rect 13725 8483 13783 8489
rect 13725 8449 13737 8483
rect 13771 8480 13783 8483
rect 13814 8480 13820 8492
rect 13771 8452 13820 8480
rect 13771 8449 13783 8452
rect 13725 8443 13783 8449
rect 13448 8433 13506 8439
rect 13464 8356 13492 8433
rect 13556 8356 13584 8443
rect 13814 8440 13820 8452
rect 13872 8440 13878 8492
rect 14090 8480 14096 8492
rect 14051 8452 14096 8480
rect 14090 8440 14096 8452
rect 14148 8440 14154 8492
rect 14200 8489 14228 8520
rect 14369 8517 14381 8551
rect 14415 8548 14427 8551
rect 14826 8548 14832 8560
rect 14415 8520 14832 8548
rect 14415 8517 14427 8520
rect 14369 8511 14427 8517
rect 14826 8508 14832 8520
rect 14884 8548 14890 8560
rect 15381 8551 15439 8557
rect 15381 8548 15393 8551
rect 14884 8520 15393 8548
rect 14884 8508 14890 8520
rect 15381 8517 15393 8520
rect 15427 8517 15439 8551
rect 15381 8511 15439 8517
rect 15470 8508 15476 8560
rect 15528 8548 15534 8560
rect 15528 8520 15573 8548
rect 15528 8508 15534 8520
rect 16040 8492 16068 8588
rect 17957 8551 18015 8557
rect 17957 8517 17969 8551
rect 18003 8548 18015 8551
rect 18046 8548 18052 8560
rect 18003 8520 18052 8548
rect 18003 8517 18015 8520
rect 17957 8511 18015 8517
rect 18046 8508 18052 8520
rect 18104 8508 18110 8560
rect 14185 8483 14243 8489
rect 14185 8449 14197 8483
rect 14231 8449 14243 8483
rect 14185 8443 14243 8449
rect 14921 8483 14979 8489
rect 14921 8449 14933 8483
rect 14967 8480 14979 8483
rect 15102 8480 15108 8492
rect 14967 8452 15108 8480
rect 14967 8449 14979 8452
rect 14921 8443 14979 8449
rect 15102 8440 15108 8452
rect 15160 8440 15166 8492
rect 15197 8483 15255 8489
rect 15197 8449 15209 8483
rect 15243 8480 15255 8483
rect 15286 8480 15292 8492
rect 15243 8452 15292 8480
rect 15243 8449 15255 8452
rect 15197 8443 15255 8449
rect 15286 8440 15292 8452
rect 15344 8440 15350 8492
rect 15617 8483 15675 8489
rect 15617 8449 15629 8483
rect 15663 8480 15675 8483
rect 15663 8452 15976 8480
rect 15663 8449 15675 8452
rect 15617 8443 15675 8449
rect 15948 8412 15976 8452
rect 16022 8440 16028 8492
rect 16080 8480 16086 8492
rect 16301 8483 16359 8489
rect 16301 8480 16313 8483
rect 16080 8452 16313 8480
rect 16080 8440 16086 8452
rect 16301 8449 16313 8452
rect 16347 8449 16359 8483
rect 16301 8443 16359 8449
rect 16408 8452 18460 8480
rect 16408 8412 16436 8452
rect 16756 8415 16814 8421
rect 16756 8412 16768 8415
rect 15948 8384 16436 8412
rect 16684 8384 16768 8412
rect 16684 8356 16712 8384
rect 16756 8381 16768 8384
rect 16802 8381 16814 8415
rect 16756 8375 16814 8381
rect 17313 8415 17371 8421
rect 17313 8381 17325 8415
rect 17359 8412 17371 8415
rect 17954 8412 17960 8424
rect 17359 8384 17960 8412
rect 17359 8381 17371 8384
rect 17313 8375 17371 8381
rect 17954 8372 17960 8384
rect 18012 8372 18018 8424
rect 18432 8356 18460 8452
rect 13446 8304 13452 8356
rect 13504 8304 13510 8356
rect 13538 8304 13544 8356
rect 13596 8304 13602 8356
rect 14550 8304 14556 8356
rect 14608 8344 14614 8356
rect 14737 8347 14795 8353
rect 14737 8344 14749 8347
rect 14608 8316 14749 8344
rect 14608 8304 14614 8316
rect 14737 8313 14749 8316
rect 14783 8313 14795 8347
rect 14737 8307 14795 8313
rect 15749 8347 15807 8353
rect 15749 8313 15761 8347
rect 15795 8344 15807 8347
rect 16666 8344 16672 8356
rect 15795 8316 16672 8344
rect 15795 8313 15807 8316
rect 15749 8307 15807 8313
rect 16666 8304 16672 8316
rect 16724 8304 16730 8356
rect 17218 8344 17224 8356
rect 17179 8316 17224 8344
rect 17218 8304 17224 8316
rect 17276 8304 17282 8356
rect 18414 8344 18420 8356
rect 18375 8316 18420 8344
rect 18414 8304 18420 8316
rect 18472 8304 18478 8356
rect 13630 8276 13636 8288
rect 13372 8248 13636 8276
rect 12253 8239 12311 8245
rect 13630 8236 13636 8248
rect 13688 8236 13694 8288
rect 14826 8236 14832 8288
rect 14884 8276 14890 8288
rect 15378 8276 15384 8288
rect 14884 8248 15384 8276
rect 14884 8236 14890 8248
rect 15378 8236 15384 8248
rect 15436 8276 15442 8288
rect 16209 8279 16267 8285
rect 16209 8276 16221 8279
rect 15436 8248 16221 8276
rect 15436 8236 15442 8248
rect 16209 8245 16221 8248
rect 16255 8245 16267 8279
rect 17862 8276 17868 8288
rect 17823 8248 17868 8276
rect 16209 8239 16267 8245
rect 17862 8236 17868 8248
rect 17920 8236 17926 8288
rect 1104 8186 18860 8208
rect 1104 8134 4214 8186
rect 4266 8134 4278 8186
rect 4330 8134 4342 8186
rect 4394 8134 4406 8186
rect 4458 8134 4470 8186
rect 4522 8134 12214 8186
rect 12266 8134 12278 8186
rect 12330 8134 12342 8186
rect 12394 8134 12406 8186
rect 12458 8134 12470 8186
rect 12522 8134 18860 8186
rect 1104 8112 18860 8134
rect 5442 8072 5448 8084
rect 5403 8044 5448 8072
rect 5442 8032 5448 8044
rect 5500 8032 5506 8084
rect 5902 8072 5908 8084
rect 5863 8044 5908 8072
rect 5902 8032 5908 8044
rect 5960 8032 5966 8084
rect 8938 8032 8944 8084
rect 8996 8072 9002 8084
rect 10045 8075 10103 8081
rect 10045 8072 10057 8075
rect 8996 8044 10057 8072
rect 8996 8032 9002 8044
rect 10045 8041 10057 8044
rect 10091 8041 10103 8075
rect 10045 8035 10103 8041
rect 10597 8075 10655 8081
rect 10597 8041 10609 8075
rect 10643 8041 10655 8075
rect 10597 8035 10655 8041
rect 11609 8075 11667 8081
rect 11609 8041 11621 8075
rect 11655 8041 11667 8075
rect 11609 8035 11667 8041
rect 4614 8004 4620 8016
rect 4575 7976 4620 8004
rect 4614 7964 4620 7976
rect 4672 7964 4678 8016
rect 4982 7964 4988 8016
rect 5040 8004 5046 8016
rect 5040 7976 6408 8004
rect 5040 7964 5046 7976
rect 4632 7936 4660 7964
rect 6380 7945 6408 7976
rect 7834 7964 7840 8016
rect 7892 8004 7898 8016
rect 10612 8004 10640 8035
rect 7892 7976 10640 8004
rect 7892 7964 7898 7976
rect 6365 7939 6423 7945
rect 4632 7908 5396 7936
rect 1486 7868 1492 7880
rect 1447 7840 1492 7868
rect 1486 7828 1492 7840
rect 1544 7828 1550 7880
rect 4525 7871 4583 7877
rect 4525 7837 4537 7871
rect 4571 7868 4583 7871
rect 4890 7868 4896 7880
rect 4571 7840 4896 7868
rect 4571 7837 4583 7840
rect 4525 7831 4583 7837
rect 4890 7828 4896 7840
rect 4948 7828 4954 7880
rect 5077 7871 5135 7877
rect 5077 7837 5089 7871
rect 5123 7868 5135 7871
rect 5258 7868 5264 7880
rect 5123 7840 5264 7868
rect 5123 7837 5135 7840
rect 5077 7831 5135 7837
rect 5258 7828 5264 7840
rect 5316 7828 5322 7880
rect 5368 7877 5396 7908
rect 6365 7905 6377 7939
rect 6411 7905 6423 7939
rect 6365 7899 6423 7905
rect 7285 7939 7343 7945
rect 7285 7905 7297 7939
rect 7331 7936 7343 7939
rect 7331 7908 7880 7936
rect 7331 7905 7343 7908
rect 7285 7899 7343 7905
rect 7852 7880 7880 7908
rect 7926 7896 7932 7948
rect 7984 7936 7990 7948
rect 8113 7939 8171 7945
rect 8113 7936 8125 7939
rect 7984 7908 8125 7936
rect 7984 7896 7990 7908
rect 8113 7905 8125 7908
rect 8159 7936 8171 7939
rect 9493 7939 9551 7945
rect 9493 7936 9505 7939
rect 8159 7908 9505 7936
rect 8159 7905 8171 7908
rect 8113 7899 8171 7905
rect 9493 7905 9505 7908
rect 9539 7936 9551 7939
rect 11422 7936 11428 7948
rect 9539 7908 11428 7936
rect 9539 7905 9551 7908
rect 9493 7899 9551 7905
rect 11422 7896 11428 7908
rect 11480 7896 11486 7948
rect 11624 7936 11652 8035
rect 12894 8032 12900 8084
rect 12952 8072 12958 8084
rect 13817 8075 13875 8081
rect 12952 8044 13584 8072
rect 12952 8032 12958 8044
rect 11793 8007 11851 8013
rect 11793 7973 11805 8007
rect 11839 8004 11851 8007
rect 13078 8004 13084 8016
rect 11839 7976 13084 8004
rect 11839 7973 11851 7976
rect 11793 7967 11851 7973
rect 13078 7964 13084 7976
rect 13136 8004 13142 8016
rect 13262 8004 13268 8016
rect 13136 7976 13268 8004
rect 13136 7964 13142 7976
rect 13262 7964 13268 7976
rect 13320 7964 13326 8016
rect 13556 7936 13584 8044
rect 13817 8041 13829 8075
rect 13863 8072 13875 8075
rect 14366 8072 14372 8084
rect 13863 8044 14372 8072
rect 13863 8041 13875 8044
rect 13817 8035 13875 8041
rect 14366 8032 14372 8044
rect 14424 8032 14430 8084
rect 14182 8004 14188 8016
rect 14143 7976 14188 8004
rect 14182 7964 14188 7976
rect 14240 7964 14246 8016
rect 16485 8007 16543 8013
rect 16485 7973 16497 8007
rect 16531 8004 16543 8007
rect 18046 8004 18052 8016
rect 16531 7976 18052 8004
rect 16531 7973 16543 7976
rect 16485 7967 16543 7973
rect 18046 7964 18052 7976
rect 18104 8004 18110 8016
rect 18141 8007 18199 8013
rect 18141 8004 18153 8007
rect 18104 7976 18153 8004
rect 18104 7964 18110 7976
rect 18141 7973 18153 7976
rect 18187 7973 18199 8007
rect 18141 7967 18199 7973
rect 14737 7939 14795 7945
rect 14737 7936 14749 7939
rect 11624 7908 12572 7936
rect 13556 7908 14749 7936
rect 5353 7871 5411 7877
rect 5353 7837 5365 7871
rect 5399 7837 5411 7871
rect 6638 7868 6644 7880
rect 6599 7840 6644 7868
rect 5353 7831 5411 7837
rect 6638 7828 6644 7840
rect 6696 7828 6702 7880
rect 7834 7828 7840 7880
rect 7892 7868 7898 7880
rect 7892 7840 7985 7868
rect 7892 7828 7898 7840
rect 8570 7828 8576 7880
rect 8628 7868 8634 7880
rect 9033 7871 9091 7877
rect 9033 7868 9045 7871
rect 8628 7840 9045 7868
rect 8628 7828 8634 7840
rect 9033 7837 9045 7840
rect 9079 7837 9091 7871
rect 9033 7831 9091 7837
rect 9309 7871 9367 7877
rect 9309 7837 9321 7871
rect 9355 7868 9367 7871
rect 9858 7868 9864 7880
rect 9355 7840 9536 7868
rect 9819 7840 9864 7868
rect 9355 7837 9367 7840
rect 9309 7831 9367 7837
rect 9508 7812 9536 7840
rect 9858 7828 9864 7840
rect 9916 7828 9922 7880
rect 10873 7871 10931 7877
rect 10336 7840 10732 7868
rect 3050 7800 3056 7812
rect 3011 7772 3056 7800
rect 3050 7760 3056 7772
rect 3108 7760 3114 7812
rect 3418 7760 3424 7812
rect 3476 7800 3482 7812
rect 3476 7772 9260 7800
rect 3476 7760 3482 7772
rect 4249 7735 4307 7741
rect 4249 7701 4261 7735
rect 4295 7732 4307 7735
rect 4614 7732 4620 7744
rect 4295 7704 4620 7732
rect 4295 7701 4307 7704
rect 4249 7695 4307 7701
rect 4614 7692 4620 7704
rect 4672 7692 4678 7744
rect 8662 7732 8668 7744
rect 8623 7704 8668 7732
rect 8662 7692 8668 7704
rect 8720 7692 8726 7744
rect 9122 7732 9128 7744
rect 9083 7704 9128 7732
rect 9122 7692 9128 7704
rect 9180 7692 9186 7744
rect 9232 7732 9260 7772
rect 9490 7760 9496 7812
rect 9548 7760 9554 7812
rect 10336 7732 10364 7840
rect 10413 7803 10471 7809
rect 10413 7769 10425 7803
rect 10459 7769 10471 7803
rect 10704 7800 10732 7840
rect 10873 7837 10885 7871
rect 10919 7868 10931 7871
rect 11241 7871 11299 7877
rect 11241 7868 11253 7871
rect 10919 7840 11253 7868
rect 10919 7837 10931 7840
rect 10873 7831 10931 7837
rect 11241 7837 11253 7840
rect 11287 7837 11299 7871
rect 11241 7831 11299 7837
rect 11618 7803 11676 7809
rect 11618 7800 11630 7803
rect 10704 7772 11630 7800
rect 10413 7763 10471 7769
rect 11618 7769 11630 7772
rect 11664 7769 11676 7803
rect 12250 7800 12256 7812
rect 11618 7763 11676 7769
rect 11992 7772 12256 7800
rect 9232 7704 10364 7732
rect 10428 7732 10456 7763
rect 10502 7732 10508 7744
rect 10428 7704 10508 7732
rect 10502 7692 10508 7704
rect 10560 7692 10566 7744
rect 10597 7735 10655 7741
rect 10597 7701 10609 7735
rect 10643 7732 10655 7735
rect 10686 7732 10692 7744
rect 10643 7704 10692 7732
rect 10643 7701 10655 7704
rect 10597 7695 10655 7701
rect 10686 7692 10692 7704
rect 10744 7732 10750 7744
rect 11992 7732 12020 7772
rect 12250 7760 12256 7772
rect 12308 7760 12314 7812
rect 12544 7800 12572 7908
rect 14737 7905 14749 7908
rect 14783 7905 14795 7939
rect 14737 7899 14795 7905
rect 15930 7896 15936 7948
rect 15988 7936 15994 7948
rect 16025 7939 16083 7945
rect 16025 7936 16037 7939
rect 15988 7908 16037 7936
rect 15988 7896 15994 7908
rect 16025 7905 16037 7908
rect 16071 7905 16083 7939
rect 16025 7899 16083 7905
rect 12710 7828 12716 7880
rect 12768 7868 12774 7880
rect 12986 7868 12992 7880
rect 12768 7840 12813 7868
rect 12947 7840 12992 7868
rect 12768 7828 12774 7840
rect 12986 7828 12992 7840
rect 13044 7828 13050 7880
rect 14826 7868 14832 7880
rect 14787 7840 14832 7868
rect 14826 7828 14832 7840
rect 14884 7828 14890 7880
rect 16040 7868 16068 7899
rect 16853 7871 16911 7877
rect 16853 7868 16865 7871
rect 16040 7840 16865 7868
rect 16853 7837 16865 7840
rect 16899 7837 16911 7871
rect 17862 7868 17868 7880
rect 17823 7840 17868 7868
rect 16853 7831 16911 7837
rect 17862 7828 17868 7840
rect 17920 7828 17926 7880
rect 12544 7772 16528 7800
rect 12158 7732 12164 7744
rect 10744 7704 12020 7732
rect 12119 7704 12164 7732
rect 10744 7692 10750 7704
rect 12158 7692 12164 7704
rect 12216 7692 12222 7744
rect 15654 7732 15660 7744
rect 15615 7704 15660 7732
rect 15654 7692 15660 7704
rect 15712 7692 15718 7744
rect 16500 7732 16528 7772
rect 16574 7760 16580 7812
rect 16632 7800 16638 7812
rect 16632 7772 16677 7800
rect 16632 7760 16638 7772
rect 17402 7732 17408 7744
rect 16500 7704 17408 7732
rect 17402 7692 17408 7704
rect 17460 7692 17466 7744
rect 1104 7642 18860 7664
rect 1104 7590 8214 7642
rect 8266 7590 8278 7642
rect 8330 7590 8342 7642
rect 8394 7590 8406 7642
rect 8458 7590 8470 7642
rect 8522 7590 16214 7642
rect 16266 7590 16278 7642
rect 16330 7590 16342 7642
rect 16394 7590 16406 7642
rect 16458 7590 16470 7642
rect 16522 7590 18860 7642
rect 1104 7568 18860 7590
rect 2317 7531 2375 7537
rect 2317 7497 2329 7531
rect 2363 7528 2375 7531
rect 2590 7528 2596 7540
rect 2363 7500 2596 7528
rect 2363 7497 2375 7500
rect 2317 7491 2375 7497
rect 2590 7488 2596 7500
rect 2648 7488 2654 7540
rect 4341 7531 4399 7537
rect 4341 7497 4353 7531
rect 4387 7528 4399 7531
rect 5074 7528 5080 7540
rect 4387 7500 5080 7528
rect 4387 7497 4399 7500
rect 4341 7491 4399 7497
rect 5074 7488 5080 7500
rect 5132 7488 5138 7540
rect 5534 7528 5540 7540
rect 5495 7500 5540 7528
rect 5534 7488 5540 7500
rect 5592 7488 5598 7540
rect 5902 7488 5908 7540
rect 5960 7528 5966 7540
rect 5997 7531 6055 7537
rect 5997 7528 6009 7531
rect 5960 7500 6009 7528
rect 5960 7488 5966 7500
rect 5997 7497 6009 7500
rect 6043 7497 6055 7531
rect 5997 7491 6055 7497
rect 7377 7531 7435 7537
rect 7377 7497 7389 7531
rect 7423 7497 7435 7531
rect 7834 7528 7840 7540
rect 7795 7500 7840 7528
rect 7377 7491 7435 7497
rect 4982 7420 4988 7472
rect 5040 7460 5046 7472
rect 7392 7460 7420 7491
rect 7834 7488 7840 7500
rect 7892 7488 7898 7540
rect 7929 7531 7987 7537
rect 7929 7497 7941 7531
rect 7975 7528 7987 7531
rect 8110 7528 8116 7540
rect 7975 7500 8116 7528
rect 7975 7497 7987 7500
rect 7929 7491 7987 7497
rect 8110 7488 8116 7500
rect 8168 7488 8174 7540
rect 11793 7531 11851 7537
rect 8312 7500 10916 7528
rect 7466 7460 7472 7472
rect 5040 7432 7236 7460
rect 7379 7432 7472 7460
rect 5040 7420 5046 7432
rect 1581 7395 1639 7401
rect 1581 7361 1593 7395
rect 1627 7392 1639 7395
rect 1854 7392 1860 7404
rect 1627 7364 1860 7392
rect 1627 7361 1639 7364
rect 1581 7355 1639 7361
rect 1854 7352 1860 7364
rect 1912 7352 1918 7404
rect 2038 7392 2044 7404
rect 1999 7364 2044 7392
rect 2038 7352 2044 7364
rect 2096 7352 2102 7404
rect 3142 7392 3148 7404
rect 3103 7364 3148 7392
rect 3142 7352 3148 7364
rect 3200 7352 3206 7404
rect 3513 7395 3571 7401
rect 3513 7361 3525 7395
rect 3559 7392 3571 7395
rect 3602 7392 3608 7404
rect 3559 7364 3608 7392
rect 3559 7361 3571 7364
rect 3513 7355 3571 7361
rect 3602 7352 3608 7364
rect 3660 7352 3666 7404
rect 3789 7395 3847 7401
rect 3789 7361 3801 7395
rect 3835 7392 3847 7395
rect 3970 7392 3976 7404
rect 3835 7364 3976 7392
rect 3835 7361 3847 7364
rect 3789 7355 3847 7361
rect 3970 7352 3976 7364
rect 4028 7352 4034 7404
rect 4433 7395 4491 7401
rect 4433 7361 4445 7395
rect 4479 7392 4491 7395
rect 4614 7392 4620 7404
rect 4479 7364 4620 7392
rect 4479 7361 4491 7364
rect 4433 7355 4491 7361
rect 4614 7352 4620 7364
rect 4672 7352 4678 7404
rect 4706 7352 4712 7404
rect 4764 7392 4770 7404
rect 4801 7395 4859 7401
rect 4801 7392 4813 7395
rect 4764 7364 4813 7392
rect 4764 7352 4770 7364
rect 4801 7361 4813 7364
rect 4847 7361 4859 7395
rect 5074 7392 5080 7404
rect 5035 7364 5080 7392
rect 4801 7355 4859 7361
rect 5074 7352 5080 7364
rect 5132 7352 5138 7404
rect 5902 7352 5908 7404
rect 5960 7392 5966 7404
rect 7208 7401 7236 7432
rect 7466 7420 7472 7432
rect 7524 7460 7530 7472
rect 8312 7469 8340 7500
rect 8297 7463 8355 7469
rect 8297 7460 8309 7463
rect 7524 7432 8309 7460
rect 7524 7420 7530 7432
rect 8297 7429 8309 7432
rect 8343 7429 8355 7463
rect 8297 7423 8355 7429
rect 8662 7420 8668 7472
rect 8720 7460 8726 7472
rect 10888 7460 10916 7500
rect 11793 7497 11805 7531
rect 11839 7528 11851 7531
rect 11882 7528 11888 7540
rect 11839 7500 11888 7528
rect 11839 7497 11851 7500
rect 11793 7491 11851 7497
rect 11882 7488 11888 7500
rect 11940 7528 11946 7540
rect 12158 7528 12164 7540
rect 11940 7500 12164 7528
rect 11940 7488 11946 7500
rect 12158 7488 12164 7500
rect 12216 7488 12222 7540
rect 15286 7488 15292 7540
rect 15344 7528 15350 7540
rect 15565 7531 15623 7537
rect 15565 7528 15577 7531
rect 15344 7500 15577 7528
rect 15344 7488 15350 7500
rect 15565 7497 15577 7500
rect 15611 7497 15623 7531
rect 15565 7491 15623 7497
rect 16301 7531 16359 7537
rect 16301 7497 16313 7531
rect 16347 7528 16359 7531
rect 16574 7528 16580 7540
rect 16347 7500 16580 7528
rect 16347 7497 16359 7500
rect 16301 7491 16359 7497
rect 16574 7488 16580 7500
rect 16632 7488 16638 7540
rect 17954 7528 17960 7540
rect 17915 7500 17960 7528
rect 17954 7488 17960 7500
rect 18012 7488 18018 7540
rect 8720 7432 10824 7460
rect 10888 7432 12204 7460
rect 8720 7420 8726 7432
rect 6733 7395 6791 7401
rect 6733 7392 6745 7395
rect 5960 7364 6745 7392
rect 5960 7352 5966 7364
rect 6733 7361 6745 7364
rect 6779 7361 6791 7395
rect 6733 7355 6791 7361
rect 7193 7395 7251 7401
rect 7193 7361 7205 7395
rect 7239 7361 7251 7395
rect 7193 7355 7251 7361
rect 7745 7395 7803 7401
rect 7745 7361 7757 7395
rect 7791 7392 7803 7395
rect 7926 7392 7932 7404
rect 7791 7364 7932 7392
rect 7791 7361 7803 7364
rect 7745 7355 7803 7361
rect 2406 7324 2412 7336
rect 2367 7296 2412 7324
rect 2406 7284 2412 7296
rect 2464 7284 2470 7336
rect 2774 7284 2780 7336
rect 2832 7324 2838 7336
rect 3418 7324 3424 7336
rect 2832 7296 2877 7324
rect 3379 7296 3424 7324
rect 2832 7284 2838 7296
rect 3418 7284 3424 7296
rect 3476 7284 3482 7336
rect 5169 7327 5227 7333
rect 5169 7293 5181 7327
rect 5215 7324 5227 7327
rect 5350 7324 5356 7336
rect 5215 7296 5356 7324
rect 5215 7293 5227 7296
rect 5169 7287 5227 7293
rect 5350 7284 5356 7296
rect 5408 7284 5414 7336
rect 7208 7324 7236 7355
rect 7926 7352 7932 7364
rect 7984 7352 7990 7404
rect 8018 7352 8024 7404
rect 8076 7401 8082 7404
rect 8076 7395 8099 7401
rect 8087 7361 8099 7395
rect 8938 7392 8944 7404
rect 8899 7364 8944 7392
rect 8076 7355 8099 7361
rect 8076 7352 8082 7355
rect 8938 7352 8944 7364
rect 8996 7352 9002 7404
rect 9122 7352 9128 7404
rect 9180 7392 9186 7404
rect 9674 7392 9680 7404
rect 9180 7364 9680 7392
rect 9180 7352 9186 7364
rect 9674 7352 9680 7364
rect 9732 7352 9738 7404
rect 9769 7395 9827 7401
rect 9769 7361 9781 7395
rect 9815 7392 9827 7395
rect 9950 7392 9956 7404
rect 9815 7364 9956 7392
rect 9815 7361 9827 7364
rect 9769 7355 9827 7361
rect 9950 7352 9956 7364
rect 10008 7352 10014 7404
rect 10410 7392 10416 7404
rect 10371 7364 10416 7392
rect 10410 7352 10416 7364
rect 10468 7352 10474 7404
rect 10502 7352 10508 7404
rect 10560 7392 10566 7404
rect 10560 7364 10605 7392
rect 10560 7352 10566 7364
rect 9140 7324 9168 7352
rect 9582 7324 9588 7336
rect 7208 7296 9168 7324
rect 9543 7296 9588 7324
rect 9582 7284 9588 7296
rect 9640 7284 9646 7336
rect 9858 7284 9864 7336
rect 9916 7324 9922 7336
rect 10428 7324 10456 7352
rect 9916 7296 10456 7324
rect 9916 7284 9922 7296
rect 9217 7259 9275 7265
rect 9217 7225 9229 7259
rect 9263 7256 9275 7259
rect 10502 7256 10508 7268
rect 9263 7228 10508 7256
rect 9263 7225 9275 7228
rect 9217 7219 9275 7225
rect 10502 7216 10508 7228
rect 10560 7216 10566 7268
rect 6546 7188 6552 7200
rect 6507 7160 6552 7188
rect 6546 7148 6552 7160
rect 6604 7148 6610 7200
rect 8481 7191 8539 7197
rect 8481 7157 8493 7191
rect 8527 7188 8539 7191
rect 9674 7188 9680 7200
rect 8527 7160 9680 7188
rect 8527 7157 8539 7160
rect 8481 7151 8539 7157
rect 9674 7148 9680 7160
rect 9732 7148 9738 7200
rect 9858 7148 9864 7200
rect 9916 7188 9922 7200
rect 9953 7191 10011 7197
rect 9953 7188 9965 7191
rect 9916 7160 9965 7188
rect 9916 7148 9922 7160
rect 9953 7157 9965 7160
rect 9999 7157 10011 7191
rect 10686 7188 10692 7200
rect 10647 7160 10692 7188
rect 9953 7151 10011 7157
rect 10686 7148 10692 7160
rect 10744 7148 10750 7200
rect 10796 7188 10824 7432
rect 11054 7352 11060 7404
rect 11112 7392 11118 7404
rect 11974 7401 11980 7404
rect 11701 7395 11759 7401
rect 11701 7392 11713 7395
rect 11112 7364 11713 7392
rect 11112 7352 11118 7364
rect 11701 7361 11713 7364
rect 11747 7361 11759 7395
rect 11701 7355 11759 7361
rect 11931 7395 11980 7401
rect 11931 7361 11943 7395
rect 11977 7361 11980 7395
rect 11931 7355 11980 7361
rect 11974 7352 11980 7355
rect 12032 7352 12038 7404
rect 12176 7401 12204 7432
rect 12250 7420 12256 7472
rect 12308 7460 12314 7472
rect 13081 7463 13139 7469
rect 13081 7460 13093 7463
rect 12308 7432 13093 7460
rect 12308 7420 12314 7432
rect 13081 7429 13093 7432
rect 13127 7429 13139 7463
rect 13081 7423 13139 7429
rect 13170 7420 13176 7472
rect 13228 7460 13234 7472
rect 16393 7463 16451 7469
rect 13228 7432 15792 7460
rect 13228 7420 13234 7432
rect 12161 7395 12219 7401
rect 12161 7361 12173 7395
rect 12207 7361 12219 7395
rect 12161 7355 12219 7361
rect 12345 7395 12403 7401
rect 12345 7361 12357 7395
rect 12391 7392 12403 7395
rect 12391 7364 13768 7392
rect 12391 7361 12403 7364
rect 12345 7355 12403 7361
rect 10870 7284 10876 7336
rect 10928 7324 10934 7336
rect 11609 7327 11667 7333
rect 11609 7324 11621 7327
rect 10928 7296 11621 7324
rect 10928 7284 10934 7296
rect 11609 7293 11621 7296
rect 11655 7293 11667 7327
rect 12176 7324 12204 7355
rect 12710 7324 12716 7336
rect 12176 7296 12716 7324
rect 11609 7287 11667 7293
rect 12710 7284 12716 7296
rect 12768 7324 12774 7336
rect 12989 7327 13047 7333
rect 12989 7324 13001 7327
rect 12768 7296 13001 7324
rect 12768 7284 12774 7296
rect 12989 7293 13001 7296
rect 13035 7293 13047 7327
rect 12989 7287 13047 7293
rect 13173 7327 13231 7333
rect 13173 7293 13185 7327
rect 13219 7324 13231 7327
rect 13446 7324 13452 7336
rect 13219 7296 13452 7324
rect 13219 7293 13231 7296
rect 13173 7287 13231 7293
rect 13004 7256 13032 7287
rect 13446 7284 13452 7296
rect 13504 7284 13510 7336
rect 13740 7324 13768 7364
rect 13814 7352 13820 7404
rect 13872 7392 13878 7404
rect 13909 7395 13967 7401
rect 13909 7392 13921 7395
rect 13872 7364 13921 7392
rect 13872 7352 13878 7364
rect 13909 7361 13921 7364
rect 13955 7361 13967 7395
rect 13909 7355 13967 7361
rect 14090 7352 14096 7404
rect 14148 7392 14154 7404
rect 14645 7395 14703 7401
rect 14645 7392 14657 7395
rect 14148 7364 14657 7392
rect 14148 7352 14154 7364
rect 14645 7361 14657 7364
rect 14691 7361 14703 7395
rect 14645 7355 14703 7361
rect 15013 7395 15071 7401
rect 15013 7361 15025 7395
rect 15059 7392 15071 7395
rect 15194 7392 15200 7404
rect 15059 7364 15200 7392
rect 15059 7361 15071 7364
rect 15013 7355 15071 7361
rect 15194 7352 15200 7364
rect 15252 7352 15258 7404
rect 15764 7401 15792 7432
rect 16393 7429 16405 7463
rect 16439 7460 16451 7463
rect 17218 7460 17224 7472
rect 16439 7432 17224 7460
rect 16439 7429 16451 7432
rect 16393 7423 16451 7429
rect 17218 7420 17224 7432
rect 17276 7460 17282 7472
rect 17405 7463 17463 7469
rect 17405 7460 17417 7463
rect 17276 7432 17417 7460
rect 17276 7420 17282 7432
rect 17405 7429 17417 7432
rect 17451 7429 17463 7463
rect 17405 7423 17463 7429
rect 17681 7463 17739 7469
rect 17681 7429 17693 7463
rect 17727 7460 17739 7463
rect 17862 7460 17868 7472
rect 17727 7432 17868 7460
rect 17727 7429 17739 7432
rect 17681 7423 17739 7429
rect 17862 7420 17868 7432
rect 17920 7420 17926 7472
rect 15749 7395 15807 7401
rect 15749 7361 15761 7395
rect 15795 7392 15807 7395
rect 16206 7392 16212 7404
rect 15795 7364 16212 7392
rect 15795 7361 15807 7364
rect 15749 7355 15807 7361
rect 16206 7352 16212 7364
rect 16264 7352 16270 7404
rect 16666 7352 16672 7404
rect 16724 7392 16730 7404
rect 16761 7395 16819 7401
rect 16761 7392 16773 7395
rect 16724 7364 16773 7392
rect 16724 7352 16730 7364
rect 16761 7361 16773 7364
rect 16807 7361 16819 7395
rect 17880 7392 17908 7420
rect 18141 7395 18199 7401
rect 18141 7392 18153 7395
rect 17880 7364 18153 7392
rect 16761 7355 16819 7361
rect 18141 7361 18153 7364
rect 18187 7361 18199 7395
rect 18141 7355 18199 7361
rect 14829 7327 14887 7333
rect 14829 7324 14841 7327
rect 13740 7296 14841 7324
rect 14829 7293 14841 7296
rect 14875 7324 14887 7327
rect 15470 7324 15476 7336
rect 14875 7296 15476 7324
rect 14875 7293 14887 7296
rect 14829 7287 14887 7293
rect 15470 7284 15476 7296
rect 15528 7284 15534 7336
rect 13538 7256 13544 7268
rect 13004 7228 13216 7256
rect 13499 7228 13544 7256
rect 13078 7188 13084 7200
rect 10796 7160 13084 7188
rect 13078 7148 13084 7160
rect 13136 7148 13142 7200
rect 13188 7188 13216 7228
rect 13538 7216 13544 7228
rect 13596 7216 13602 7268
rect 15010 7256 15016 7268
rect 14971 7228 15016 7256
rect 15010 7216 15016 7228
rect 15068 7216 15074 7268
rect 13722 7188 13728 7200
rect 13188 7160 13728 7188
rect 13722 7148 13728 7160
rect 13780 7148 13786 7200
rect 14090 7188 14096 7200
rect 14051 7160 14096 7188
rect 14090 7148 14096 7160
rect 14148 7148 14154 7200
rect 1104 7098 18860 7120
rect 1104 7046 4214 7098
rect 4266 7046 4278 7098
rect 4330 7046 4342 7098
rect 4394 7046 4406 7098
rect 4458 7046 4470 7098
rect 4522 7046 12214 7098
rect 12266 7046 12278 7098
rect 12330 7046 12342 7098
rect 12394 7046 12406 7098
rect 12458 7046 12470 7098
rect 12522 7046 18860 7098
rect 1104 7024 18860 7046
rect 2774 6944 2780 6996
rect 2832 6984 2838 6996
rect 3145 6987 3203 6993
rect 3145 6984 3157 6987
rect 2832 6956 3157 6984
rect 2832 6944 2838 6956
rect 3145 6953 3157 6956
rect 3191 6953 3203 6987
rect 3145 6947 3203 6953
rect 9490 6944 9496 6996
rect 9548 6984 9554 6996
rect 9858 6984 9864 6996
rect 9548 6956 9864 6984
rect 9548 6944 9554 6956
rect 9858 6944 9864 6956
rect 9916 6944 9922 6996
rect 12406 6956 14596 6984
rect 2038 6876 2044 6928
rect 2096 6916 2102 6928
rect 2133 6919 2191 6925
rect 2133 6916 2145 6919
rect 2096 6888 2145 6916
rect 2096 6876 2102 6888
rect 2133 6885 2145 6888
rect 2179 6916 2191 6919
rect 2682 6916 2688 6928
rect 2179 6888 2688 6916
rect 2179 6885 2191 6888
rect 2133 6879 2191 6885
rect 2682 6876 2688 6888
rect 2740 6876 2746 6928
rect 4614 6876 4620 6928
rect 4672 6916 4678 6928
rect 12406 6916 12434 6956
rect 4672 6888 12434 6916
rect 4672 6876 4678 6888
rect 13262 6876 13268 6928
rect 13320 6916 13326 6928
rect 13449 6919 13507 6925
rect 13449 6916 13461 6919
rect 13320 6888 13461 6916
rect 13320 6876 13326 6888
rect 13449 6885 13461 6888
rect 13495 6885 13507 6919
rect 14568 6916 14596 6956
rect 17494 6916 17500 6928
rect 14568 6888 17500 6916
rect 13449 6879 13507 6885
rect 17494 6876 17500 6888
rect 17552 6876 17558 6928
rect 1670 6808 1676 6860
rect 1728 6848 1734 6860
rect 2501 6851 2559 6857
rect 2501 6848 2513 6851
rect 1728 6820 2513 6848
rect 1728 6808 1734 6820
rect 2501 6817 2513 6820
rect 2547 6817 2559 6851
rect 2501 6811 2559 6817
rect 3234 6808 3240 6860
rect 3292 6848 3298 6860
rect 4632 6848 4660 6876
rect 7466 6848 7472 6860
rect 3292 6820 4660 6848
rect 7427 6820 7472 6848
rect 3292 6808 3298 6820
rect 7466 6808 7472 6820
rect 7524 6808 7530 6860
rect 10597 6851 10655 6857
rect 9692 6820 10180 6848
rect 9692 6792 9720 6820
rect 1946 6780 1952 6792
rect 1907 6752 1952 6780
rect 1946 6740 1952 6752
rect 2004 6740 2010 6792
rect 2225 6783 2283 6789
rect 2225 6749 2237 6783
rect 2271 6780 2283 6783
rect 2406 6780 2412 6792
rect 2271 6752 2412 6780
rect 2271 6749 2283 6752
rect 2225 6743 2283 6749
rect 2406 6740 2412 6752
rect 2464 6740 2470 6792
rect 3329 6783 3387 6789
rect 3329 6749 3341 6783
rect 3375 6749 3387 6783
rect 3329 6743 3387 6749
rect 3513 6783 3571 6789
rect 3513 6749 3525 6783
rect 3559 6780 3571 6783
rect 3878 6780 3884 6792
rect 3559 6752 3884 6780
rect 3559 6749 3571 6752
rect 3513 6743 3571 6749
rect 3344 6712 3372 6743
rect 3878 6740 3884 6752
rect 3936 6740 3942 6792
rect 4706 6740 4712 6792
rect 4764 6780 4770 6792
rect 4801 6783 4859 6789
rect 4801 6780 4813 6783
rect 4764 6752 4813 6780
rect 4764 6740 4770 6752
rect 4801 6749 4813 6752
rect 4847 6749 4859 6783
rect 4801 6743 4859 6749
rect 5074 6740 5080 6792
rect 5132 6780 5138 6792
rect 5261 6783 5319 6789
rect 5261 6780 5273 6783
rect 5132 6752 5273 6780
rect 5132 6740 5138 6752
rect 5261 6749 5273 6752
rect 5307 6780 5319 6783
rect 5813 6783 5871 6789
rect 5813 6780 5825 6783
rect 5307 6752 5825 6780
rect 5307 6749 5319 6752
rect 5261 6743 5319 6749
rect 5813 6749 5825 6752
rect 5859 6749 5871 6783
rect 6825 6783 6883 6789
rect 5813 6743 5871 6749
rect 4433 6715 4491 6721
rect 4433 6712 4445 6715
rect 1596 6684 3280 6712
rect 3344 6684 4445 6712
rect 1596 6656 1624 6684
rect 1578 6644 1584 6656
rect 1539 6616 1584 6644
rect 1578 6604 1584 6616
rect 1636 6604 1642 6656
rect 2406 6644 2412 6656
rect 2367 6616 2412 6644
rect 2406 6604 2412 6616
rect 2464 6604 2470 6656
rect 2685 6647 2743 6653
rect 2685 6613 2697 6647
rect 2731 6644 2743 6647
rect 2774 6644 2780 6656
rect 2731 6616 2780 6644
rect 2731 6613 2743 6616
rect 2685 6607 2743 6613
rect 2774 6604 2780 6616
rect 2832 6604 2838 6656
rect 3252 6644 3280 6684
rect 4433 6681 4445 6684
rect 4479 6712 4491 6715
rect 4890 6712 4896 6724
rect 4479 6684 4896 6712
rect 4479 6681 4491 6684
rect 4433 6675 4491 6681
rect 4890 6672 4896 6684
rect 4948 6672 4954 6724
rect 6748 6712 6776 6766
rect 6825 6749 6837 6783
rect 6871 6780 6883 6783
rect 6914 6780 6920 6792
rect 6871 6752 6920 6780
rect 6871 6749 6883 6752
rect 6825 6743 6883 6749
rect 6914 6740 6920 6752
rect 6972 6740 6978 6792
rect 8110 6780 8116 6792
rect 7958 6752 8116 6780
rect 8110 6740 8116 6752
rect 8168 6740 8174 6792
rect 9674 6740 9680 6792
rect 9732 6740 9738 6792
rect 10045 6783 10103 6789
rect 10045 6749 10057 6783
rect 10091 6749 10103 6783
rect 10152 6780 10180 6820
rect 10597 6817 10609 6851
rect 10643 6848 10655 6851
rect 10686 6848 10692 6860
rect 10643 6820 10692 6848
rect 10643 6817 10655 6820
rect 10597 6811 10655 6817
rect 10686 6808 10692 6820
rect 10744 6808 10750 6860
rect 14090 6848 14096 6860
rect 13464 6820 14096 6848
rect 10870 6789 10876 6792
rect 10827 6783 10876 6789
rect 10827 6780 10839 6783
rect 10152 6752 10839 6780
rect 10045 6743 10103 6749
rect 10827 6749 10839 6752
rect 10873 6749 10876 6783
rect 10827 6743 10876 6749
rect 7006 6712 7012 6724
rect 6748 6684 7012 6712
rect 7006 6672 7012 6684
rect 7064 6672 7070 6724
rect 8297 6715 8355 6721
rect 8297 6681 8309 6715
rect 8343 6712 8355 6715
rect 8570 6712 8576 6724
rect 8343 6684 8576 6712
rect 8343 6681 8355 6684
rect 8297 6675 8355 6681
rect 8570 6672 8576 6684
rect 8628 6672 8634 6724
rect 9033 6715 9091 6721
rect 9033 6681 9045 6715
rect 9079 6712 9091 6715
rect 9122 6712 9128 6724
rect 9079 6684 9128 6712
rect 9079 6681 9091 6684
rect 9033 6675 9091 6681
rect 9122 6672 9128 6684
rect 9180 6672 9186 6724
rect 10060 6712 10088 6743
rect 10870 6740 10876 6743
rect 10928 6740 10934 6792
rect 10965 6783 11023 6789
rect 10965 6749 10977 6783
rect 11011 6780 11023 6783
rect 11054 6780 11060 6792
rect 11011 6752 11060 6780
rect 11011 6749 11023 6752
rect 10965 6743 11023 6749
rect 10980 6712 11008 6743
rect 11054 6740 11060 6752
rect 11112 6740 11118 6792
rect 11517 6783 11575 6789
rect 11517 6749 11529 6783
rect 11563 6749 11575 6783
rect 11882 6780 11888 6792
rect 11843 6752 11888 6780
rect 11517 6743 11575 6749
rect 10060 6684 11008 6712
rect 3878 6644 3884 6656
rect 3252 6616 3884 6644
rect 3878 6604 3884 6616
rect 3936 6644 3942 6656
rect 4065 6647 4123 6653
rect 4065 6644 4077 6647
rect 3936 6616 4077 6644
rect 3936 6604 3942 6616
rect 4065 6613 4077 6616
rect 4111 6613 4123 6647
rect 4065 6607 4123 6613
rect 10965 6647 11023 6653
rect 10965 6613 10977 6647
rect 11011 6644 11023 6647
rect 11532 6644 11560 6743
rect 11882 6740 11888 6752
rect 11940 6740 11946 6792
rect 12250 6740 12256 6792
rect 12308 6780 12314 6792
rect 13019 6783 13077 6789
rect 13019 6780 13031 6783
rect 12308 6752 13031 6780
rect 12308 6740 12314 6752
rect 13019 6749 13031 6752
rect 13065 6780 13077 6783
rect 13464 6780 13492 6820
rect 14090 6808 14096 6820
rect 14148 6808 14154 6860
rect 15194 6848 15200 6860
rect 15155 6820 15200 6848
rect 15194 6808 15200 6820
rect 15252 6848 15258 6860
rect 17310 6848 17316 6860
rect 15252 6820 15792 6848
rect 15252 6808 15258 6820
rect 13065 6752 13492 6780
rect 13065 6749 13077 6752
rect 13019 6743 13077 6749
rect 13538 6740 13544 6792
rect 13596 6780 13602 6792
rect 13596 6752 13641 6780
rect 13596 6740 13602 6752
rect 13722 6740 13728 6792
rect 13780 6780 13786 6792
rect 14277 6783 14335 6789
rect 14277 6780 14289 6783
rect 13780 6752 14289 6780
rect 13780 6740 13786 6752
rect 14277 6749 14289 6752
rect 14323 6749 14335 6783
rect 14277 6743 14335 6749
rect 14645 6783 14703 6789
rect 14645 6749 14657 6783
rect 14691 6780 14703 6783
rect 15286 6780 15292 6792
rect 14691 6752 15292 6780
rect 14691 6749 14703 6752
rect 14645 6743 14703 6749
rect 15286 6740 15292 6752
rect 15344 6740 15350 6792
rect 15470 6740 15476 6792
rect 15528 6780 15534 6792
rect 15764 6789 15792 6820
rect 17144 6820 17316 6848
rect 15565 6783 15623 6789
rect 15565 6780 15577 6783
rect 15528 6752 15577 6780
rect 15528 6740 15534 6752
rect 15565 6749 15577 6752
rect 15611 6749 15623 6783
rect 15565 6743 15623 6749
rect 15749 6783 15807 6789
rect 15749 6749 15761 6783
rect 15795 6749 15807 6783
rect 15749 6743 15807 6749
rect 16114 6740 16120 6792
rect 16172 6780 16178 6792
rect 17144 6789 17172 6820
rect 17310 6808 17316 6820
rect 17368 6848 17374 6860
rect 18049 6851 18107 6857
rect 18049 6848 18061 6851
rect 17368 6820 18061 6848
rect 17368 6808 17374 6820
rect 18049 6817 18061 6820
rect 18095 6817 18107 6851
rect 18049 6811 18107 6817
rect 16393 6783 16451 6789
rect 16393 6780 16405 6783
rect 16172 6752 16405 6780
rect 16172 6740 16178 6752
rect 16393 6749 16405 6752
rect 16439 6749 16451 6783
rect 16393 6743 16451 6749
rect 17129 6783 17187 6789
rect 17129 6749 17141 6783
rect 17175 6749 17187 6783
rect 17589 6783 17647 6789
rect 17589 6780 17601 6783
rect 17129 6743 17187 6749
rect 17236 6752 17601 6780
rect 16408 6712 16436 6743
rect 17236 6712 17264 6752
rect 17589 6749 17601 6752
rect 17635 6749 17647 6783
rect 17589 6743 17647 6749
rect 16408 6684 17264 6712
rect 17313 6715 17371 6721
rect 17313 6681 17325 6715
rect 17359 6712 17371 6715
rect 18046 6712 18052 6724
rect 17359 6684 18052 6712
rect 17359 6681 17371 6684
rect 17313 6675 17371 6681
rect 18046 6672 18052 6684
rect 18104 6672 18110 6724
rect 18138 6672 18144 6724
rect 18196 6712 18202 6724
rect 18196 6684 18241 6712
rect 18196 6672 18202 6684
rect 11011 6616 11560 6644
rect 11011 6613 11023 6616
rect 10965 6607 11023 6613
rect 12158 6604 12164 6656
rect 12216 6644 12222 6656
rect 12529 6647 12587 6653
rect 12529 6644 12541 6647
rect 12216 6616 12541 6644
rect 12216 6604 12222 6616
rect 12529 6613 12541 6616
rect 12575 6613 12587 6647
rect 12529 6607 12587 6613
rect 12710 6604 12716 6656
rect 12768 6644 12774 6656
rect 12897 6647 12955 6653
rect 12897 6644 12909 6647
rect 12768 6616 12909 6644
rect 12768 6604 12774 6616
rect 12897 6613 12909 6616
rect 12943 6613 12955 6647
rect 13078 6644 13084 6656
rect 13039 6616 13084 6644
rect 12897 6607 12955 6613
rect 13078 6604 13084 6616
rect 13136 6604 13142 6656
rect 15930 6644 15936 6656
rect 15891 6616 15936 6644
rect 15930 6604 15936 6616
rect 15988 6604 15994 6656
rect 1104 6554 18860 6576
rect 1104 6502 8214 6554
rect 8266 6502 8278 6554
rect 8330 6502 8342 6554
rect 8394 6502 8406 6554
rect 8458 6502 8470 6554
rect 8522 6502 16214 6554
rect 16266 6502 16278 6554
rect 16330 6502 16342 6554
rect 16394 6502 16406 6554
rect 16458 6502 16470 6554
rect 16522 6502 18860 6554
rect 1104 6480 18860 6502
rect 2682 6400 2688 6452
rect 2740 6440 2746 6452
rect 4341 6443 4399 6449
rect 4341 6440 4353 6443
rect 2740 6412 4353 6440
rect 2740 6400 2746 6412
rect 2406 6332 2412 6384
rect 2464 6372 2470 6384
rect 3528 6372 3556 6412
rect 4341 6409 4353 6412
rect 4387 6409 4399 6443
rect 4341 6403 4399 6409
rect 8481 6443 8539 6449
rect 8481 6409 8493 6443
rect 8527 6440 8539 6443
rect 8570 6440 8576 6452
rect 8527 6412 8576 6440
rect 8527 6409 8539 6412
rect 8481 6403 8539 6409
rect 8570 6400 8576 6412
rect 8628 6400 8634 6452
rect 9122 6440 9128 6452
rect 9083 6412 9128 6440
rect 9122 6400 9128 6412
rect 9180 6400 9186 6452
rect 12158 6440 12164 6452
rect 12119 6412 12164 6440
rect 12158 6400 12164 6412
rect 12216 6400 12222 6452
rect 15749 6443 15807 6449
rect 15749 6409 15761 6443
rect 15795 6440 15807 6443
rect 16574 6440 16580 6452
rect 15795 6412 16580 6440
rect 15795 6409 15807 6412
rect 15749 6403 15807 6409
rect 16574 6400 16580 6412
rect 16632 6440 16638 6452
rect 17034 6440 17040 6452
rect 16632 6412 17040 6440
rect 16632 6400 16638 6412
rect 17034 6400 17040 6412
rect 17092 6400 17098 6452
rect 3970 6372 3976 6384
rect 2464 6344 3372 6372
rect 3528 6344 3648 6372
rect 3931 6344 3976 6372
rect 2464 6332 2470 6344
rect 1946 6304 1952 6316
rect 1596 6276 1952 6304
rect 1596 6112 1624 6276
rect 1946 6264 1952 6276
rect 2004 6264 2010 6316
rect 2501 6307 2559 6313
rect 2501 6273 2513 6307
rect 2547 6273 2559 6307
rect 2501 6267 2559 6273
rect 2516 6168 2544 6267
rect 2590 6264 2596 6316
rect 2648 6304 2654 6316
rect 2648 6276 2693 6304
rect 2648 6264 2654 6276
rect 2774 6264 2780 6316
rect 2832 6304 2838 6316
rect 3344 6313 3372 6344
rect 3329 6307 3387 6313
rect 2832 6276 2877 6304
rect 2832 6264 2838 6276
rect 3329 6273 3341 6307
rect 3375 6273 3387 6307
rect 3510 6304 3516 6316
rect 3471 6276 3516 6304
rect 3329 6267 3387 6273
rect 3510 6264 3516 6276
rect 3568 6264 3574 6316
rect 3620 6313 3648 6344
rect 3970 6332 3976 6344
rect 4028 6332 4034 6384
rect 4614 6372 4620 6384
rect 4448 6344 4620 6372
rect 3605 6307 3663 6313
rect 3605 6273 3617 6307
rect 3651 6273 3663 6307
rect 3605 6267 3663 6273
rect 3694 6264 3700 6316
rect 3752 6304 3758 6316
rect 3752 6276 3797 6304
rect 3752 6264 3758 6276
rect 4062 6264 4068 6316
rect 4120 6304 4126 6316
rect 4448 6313 4476 6344
rect 4614 6332 4620 6344
rect 4672 6332 4678 6384
rect 4890 6332 4896 6384
rect 4948 6372 4954 6384
rect 4948 6344 5304 6372
rect 4948 6332 4954 6344
rect 5276 6313 5304 6344
rect 5442 6332 5448 6384
rect 5500 6372 5506 6384
rect 6914 6372 6920 6384
rect 5500 6344 5856 6372
rect 5500 6332 5506 6344
rect 4249 6307 4307 6313
rect 4249 6304 4261 6307
rect 4120 6276 4261 6304
rect 4120 6264 4126 6276
rect 4249 6273 4261 6276
rect 4295 6273 4307 6307
rect 4249 6267 4307 6273
rect 4433 6307 4491 6313
rect 4433 6273 4445 6307
rect 4479 6273 4491 6307
rect 5135 6307 5193 6313
rect 5135 6304 5147 6307
rect 4433 6267 4491 6273
rect 4540 6276 5147 6304
rect 2681 6239 2739 6245
rect 2681 6205 2693 6239
rect 2727 6236 2739 6239
rect 2866 6236 2872 6248
rect 2727 6208 2872 6236
rect 2727 6205 2739 6208
rect 2681 6199 2739 6205
rect 2866 6196 2872 6208
rect 2924 6196 2930 6248
rect 3878 6196 3884 6248
rect 3936 6236 3942 6248
rect 4540 6236 4568 6276
rect 5135 6273 5147 6276
rect 5181 6273 5193 6307
rect 5135 6267 5193 6273
rect 5261 6307 5319 6313
rect 5261 6273 5273 6307
rect 5307 6273 5319 6307
rect 5261 6267 5319 6273
rect 5350 6264 5356 6316
rect 5408 6304 5414 6316
rect 5828 6313 5856 6344
rect 6656 6344 6920 6372
rect 6656 6313 6684 6344
rect 6914 6332 6920 6344
rect 6972 6372 6978 6384
rect 7466 6372 7472 6384
rect 6972 6344 7472 6372
rect 6972 6332 6978 6344
rect 7466 6332 7472 6344
rect 7524 6332 7530 6384
rect 10873 6375 10931 6381
rect 9048 6344 10824 6372
rect 5537 6307 5595 6313
rect 5408 6276 5453 6304
rect 5408 6264 5414 6276
rect 5537 6273 5549 6307
rect 5583 6273 5595 6307
rect 5537 6267 5595 6273
rect 5813 6307 5871 6313
rect 5813 6273 5825 6307
rect 5859 6273 5871 6307
rect 5813 6267 5871 6273
rect 6641 6307 6699 6313
rect 6641 6273 6653 6307
rect 6687 6273 6699 6307
rect 6641 6267 6699 6273
rect 6825 6307 6883 6313
rect 6825 6273 6837 6307
rect 6871 6304 6883 6307
rect 7006 6304 7012 6316
rect 6871 6276 7012 6304
rect 6871 6273 6883 6276
rect 6825 6267 6883 6273
rect 3936 6208 4568 6236
rect 5552 6236 5580 6267
rect 7006 6264 7012 6276
rect 7064 6264 7070 6316
rect 9048 6313 9076 6344
rect 7653 6307 7711 6313
rect 7653 6273 7665 6307
rect 7699 6304 7711 6307
rect 8573 6307 8631 6313
rect 7699 6276 8064 6304
rect 7699 6273 7711 6276
rect 7653 6267 7711 6273
rect 6457 6239 6515 6245
rect 6457 6236 6469 6239
rect 5552 6208 6469 6236
rect 3936 6196 3942 6208
rect 6457 6205 6469 6208
rect 6503 6205 6515 6239
rect 6457 6199 6515 6205
rect 3602 6168 3608 6180
rect 2516 6140 3608 6168
rect 3602 6128 3608 6140
rect 3660 6168 3666 6180
rect 8036 6177 8064 6276
rect 8573 6273 8585 6307
rect 8619 6304 8631 6307
rect 9033 6307 9091 6313
rect 9033 6304 9045 6307
rect 8619 6276 9045 6304
rect 8619 6273 8631 6276
rect 8573 6267 8631 6273
rect 9033 6273 9045 6276
rect 9079 6273 9091 6307
rect 9953 6307 10011 6313
rect 9953 6304 9965 6307
rect 9033 6267 9091 6273
rect 9600 6276 9965 6304
rect 8478 6236 8484 6248
rect 8439 6208 8484 6236
rect 8478 6196 8484 6208
rect 8536 6196 8542 6248
rect 8938 6196 8944 6248
rect 8996 6236 9002 6248
rect 9125 6239 9183 6245
rect 9125 6236 9137 6239
rect 8996 6208 9137 6236
rect 8996 6196 9002 6208
rect 9125 6205 9137 6208
rect 9171 6205 9183 6239
rect 9125 6199 9183 6205
rect 9600 6177 9628 6276
rect 9953 6273 9965 6276
rect 9999 6273 10011 6307
rect 10502 6304 10508 6316
rect 10463 6276 10508 6304
rect 9953 6267 10011 6273
rect 10502 6264 10508 6276
rect 10560 6264 10566 6316
rect 10686 6304 10692 6316
rect 10647 6276 10692 6304
rect 10686 6264 10692 6276
rect 10744 6264 10750 6316
rect 10796 6304 10824 6344
rect 10873 6341 10885 6375
rect 10919 6372 10931 6375
rect 11054 6372 11060 6384
rect 10919 6344 11060 6372
rect 10919 6341 10931 6344
rect 10873 6335 10931 6341
rect 11054 6332 11060 6344
rect 11112 6332 11118 6384
rect 12250 6372 12256 6384
rect 12211 6344 12256 6372
rect 12250 6332 12256 6344
rect 12308 6332 12314 6384
rect 14826 6372 14832 6384
rect 14200 6344 14832 6372
rect 12268 6304 12296 6332
rect 14200 6313 14228 6344
rect 14826 6332 14832 6344
rect 14884 6332 14890 6384
rect 15838 6332 15844 6384
rect 15896 6372 15902 6384
rect 16025 6375 16083 6381
rect 16025 6372 16037 6375
rect 15896 6344 16037 6372
rect 15896 6332 15902 6344
rect 16025 6341 16037 6344
rect 16071 6341 16083 6375
rect 16025 6335 16083 6341
rect 16209 6375 16267 6381
rect 16209 6341 16221 6375
rect 16255 6372 16267 6375
rect 17126 6372 17132 6384
rect 16255 6344 17132 6372
rect 16255 6341 16267 6344
rect 16209 6335 16267 6341
rect 17126 6332 17132 6344
rect 17184 6332 17190 6384
rect 10796 6276 12296 6304
rect 13173 6307 13231 6313
rect 13173 6273 13185 6307
rect 13219 6304 13231 6307
rect 14185 6307 14243 6313
rect 14185 6304 14197 6307
rect 13219 6276 14197 6304
rect 13219 6273 13231 6276
rect 13173 6267 13231 6273
rect 14185 6273 14197 6276
rect 14231 6273 14243 6307
rect 14185 6267 14243 6273
rect 14277 6307 14335 6313
rect 14277 6273 14289 6307
rect 14323 6304 14335 6307
rect 15010 6304 15016 6316
rect 14323 6276 14872 6304
rect 14971 6276 15016 6304
rect 14323 6273 14335 6276
rect 14277 6267 14335 6273
rect 12161 6239 12219 6245
rect 12161 6205 12173 6239
rect 12207 6236 12219 6239
rect 12802 6236 12808 6248
rect 12207 6208 12808 6236
rect 12207 6205 12219 6208
rect 12161 6199 12219 6205
rect 12802 6196 12808 6208
rect 12860 6196 12866 6248
rect 4893 6171 4951 6177
rect 4893 6168 4905 6171
rect 3660 6140 4905 6168
rect 3660 6128 3666 6140
rect 4893 6137 4905 6140
rect 4939 6137 4951 6171
rect 4893 6131 4951 6137
rect 8021 6171 8079 6177
rect 8021 6137 8033 6171
rect 8067 6137 8079 6171
rect 8021 6131 8079 6137
rect 9585 6171 9643 6177
rect 9585 6137 9597 6171
rect 9631 6137 9643 6171
rect 9585 6131 9643 6137
rect 9950 6128 9956 6180
rect 10008 6168 10014 6180
rect 13188 6168 13216 6267
rect 13262 6196 13268 6248
rect 13320 6236 13326 6248
rect 13449 6239 13507 6245
rect 13320 6208 13365 6236
rect 13320 6196 13326 6208
rect 13449 6205 13461 6239
rect 13495 6236 13507 6239
rect 14001 6239 14059 6245
rect 14001 6236 14013 6239
rect 13495 6208 14013 6236
rect 13495 6205 13507 6208
rect 13449 6199 13507 6205
rect 14001 6205 14013 6208
rect 14047 6205 14059 6239
rect 14001 6199 14059 6205
rect 14090 6196 14096 6248
rect 14148 6236 14154 6248
rect 14292 6236 14320 6267
rect 14844 6245 14872 6276
rect 15010 6264 15016 6276
rect 15068 6264 15074 6316
rect 15105 6307 15163 6313
rect 15105 6273 15117 6307
rect 15151 6304 15163 6307
rect 15930 6304 15936 6316
rect 15151 6276 15936 6304
rect 15151 6273 15163 6276
rect 15105 6267 15163 6273
rect 15930 6264 15936 6276
rect 15988 6264 15994 6316
rect 16393 6307 16451 6313
rect 16393 6273 16405 6307
rect 16439 6304 16451 6307
rect 16853 6307 16911 6313
rect 16853 6304 16865 6307
rect 16439 6276 16865 6304
rect 16439 6273 16451 6276
rect 16393 6267 16451 6273
rect 16853 6273 16865 6276
rect 16899 6273 16911 6307
rect 18046 6304 18052 6316
rect 18007 6276 18052 6304
rect 16853 6267 16911 6273
rect 18046 6264 18052 6276
rect 18104 6264 18110 6316
rect 14148 6208 14320 6236
rect 14737 6239 14795 6245
rect 14148 6196 14154 6208
rect 14737 6205 14749 6239
rect 14783 6205 14795 6239
rect 14737 6199 14795 6205
rect 14829 6239 14887 6245
rect 14829 6205 14841 6239
rect 14875 6205 14887 6239
rect 14829 6199 14887 6205
rect 10008 6140 13216 6168
rect 14752 6168 14780 6199
rect 15286 6196 15292 6248
rect 15344 6196 15350 6248
rect 15304 6168 15332 6196
rect 14752 6140 15332 6168
rect 10008 6128 10014 6140
rect 17494 6128 17500 6180
rect 17552 6168 17558 6180
rect 18141 6171 18199 6177
rect 18141 6168 18153 6171
rect 17552 6140 18153 6168
rect 17552 6128 17558 6140
rect 18141 6137 18153 6140
rect 18187 6137 18199 6171
rect 18141 6131 18199 6137
rect 1578 6100 1584 6112
rect 1539 6072 1584 6100
rect 1578 6060 1584 6072
rect 1636 6060 1642 6112
rect 2041 6103 2099 6109
rect 2041 6069 2053 6103
rect 2087 6100 2099 6103
rect 2590 6100 2596 6112
rect 2087 6072 2596 6100
rect 2087 6069 2099 6072
rect 2041 6063 2099 6069
rect 2590 6060 2596 6072
rect 2648 6060 2654 6112
rect 2961 6103 3019 6109
rect 2961 6069 2973 6103
rect 3007 6100 3019 6103
rect 4982 6100 4988 6112
rect 3007 6072 4988 6100
rect 3007 6069 3019 6072
rect 2961 6063 3019 6069
rect 4982 6060 4988 6072
rect 5040 6060 5046 6112
rect 5074 6060 5080 6112
rect 5132 6100 5138 6112
rect 5905 6103 5963 6109
rect 5905 6100 5917 6103
rect 5132 6072 5917 6100
rect 5132 6060 5138 6072
rect 5905 6069 5917 6072
rect 5951 6069 5963 6103
rect 5905 6063 5963 6069
rect 7282 6060 7288 6112
rect 7340 6100 7346 6112
rect 7469 6103 7527 6109
rect 7469 6100 7481 6103
rect 7340 6072 7481 6100
rect 7340 6060 7346 6072
rect 7469 6069 7481 6072
rect 7515 6069 7527 6103
rect 7469 6063 7527 6069
rect 9674 6060 9680 6112
rect 9732 6100 9738 6112
rect 10137 6103 10195 6109
rect 10137 6100 10149 6103
rect 9732 6072 10149 6100
rect 9732 6060 9738 6072
rect 10137 6069 10149 6072
rect 10183 6069 10195 6103
rect 10137 6063 10195 6069
rect 11514 6060 11520 6112
rect 11572 6100 11578 6112
rect 11701 6103 11759 6109
rect 11701 6100 11713 6103
rect 11572 6072 11713 6100
rect 11572 6060 11578 6072
rect 11701 6069 11713 6072
rect 11747 6069 11759 6103
rect 11701 6063 11759 6069
rect 13633 6103 13691 6109
rect 13633 6069 13645 6103
rect 13679 6100 13691 6103
rect 13998 6100 14004 6112
rect 13679 6072 14004 6100
rect 13679 6069 13691 6072
rect 13633 6063 13691 6069
rect 13998 6060 14004 6072
rect 14056 6060 14062 6112
rect 15286 6100 15292 6112
rect 15247 6072 15292 6100
rect 15286 6060 15292 6072
rect 15344 6060 15350 6112
rect 1104 6010 18860 6032
rect 1104 5958 4214 6010
rect 4266 5958 4278 6010
rect 4330 5958 4342 6010
rect 4394 5958 4406 6010
rect 4458 5958 4470 6010
rect 4522 5958 12214 6010
rect 12266 5958 12278 6010
rect 12330 5958 12342 6010
rect 12394 5958 12406 6010
rect 12458 5958 12470 6010
rect 12522 5958 18860 6010
rect 1104 5936 18860 5958
rect 2133 5899 2191 5905
rect 2133 5865 2145 5899
rect 2179 5896 2191 5899
rect 2406 5896 2412 5908
rect 2179 5868 2412 5896
rect 2179 5865 2191 5868
rect 2133 5859 2191 5865
rect 2406 5856 2412 5868
rect 2464 5856 2470 5908
rect 2498 5856 2504 5908
rect 2556 5896 2562 5908
rect 3145 5899 3203 5905
rect 3145 5896 3157 5899
rect 2556 5868 3157 5896
rect 2556 5856 2562 5868
rect 3145 5865 3157 5868
rect 3191 5896 3203 5899
rect 3510 5896 3516 5908
rect 3191 5868 3516 5896
rect 3191 5865 3203 5868
rect 3145 5859 3203 5865
rect 3510 5856 3516 5868
rect 3568 5856 3574 5908
rect 4062 5896 4068 5908
rect 4023 5868 4068 5896
rect 4062 5856 4068 5868
rect 4120 5856 4126 5908
rect 4249 5899 4307 5905
rect 4249 5865 4261 5899
rect 4295 5896 4307 5899
rect 4798 5896 4804 5908
rect 4295 5868 4804 5896
rect 4295 5865 4307 5868
rect 4249 5859 4307 5865
rect 4798 5856 4804 5868
rect 4856 5856 4862 5908
rect 8478 5856 8484 5908
rect 8536 5896 8542 5908
rect 8754 5896 8760 5908
rect 8536 5868 8760 5896
rect 8536 5856 8542 5868
rect 8754 5856 8760 5868
rect 8812 5896 8818 5908
rect 9582 5896 9588 5908
rect 8812 5868 9588 5896
rect 8812 5856 8818 5868
rect 9582 5856 9588 5868
rect 9640 5856 9646 5908
rect 13357 5899 13415 5905
rect 13357 5865 13369 5899
rect 13403 5896 13415 5899
rect 16574 5896 16580 5908
rect 13403 5868 16580 5896
rect 13403 5865 13415 5868
rect 13357 5859 13415 5865
rect 16574 5856 16580 5868
rect 16632 5856 16638 5908
rect 18049 5899 18107 5905
rect 18049 5865 18061 5899
rect 18095 5896 18107 5899
rect 18138 5896 18144 5908
rect 18095 5868 18144 5896
rect 18095 5865 18107 5868
rect 18049 5859 18107 5865
rect 18138 5856 18144 5868
rect 18196 5856 18202 5908
rect 2774 5828 2780 5840
rect 2240 5800 2780 5828
rect 2240 5701 2268 5800
rect 2774 5788 2780 5800
rect 2832 5828 2838 5840
rect 3878 5828 3884 5840
rect 2832 5800 3884 5828
rect 2832 5788 2838 5800
rect 3878 5788 3884 5800
rect 3936 5788 3942 5840
rect 2590 5720 2596 5772
rect 2648 5760 2654 5772
rect 2961 5763 3019 5769
rect 2961 5760 2973 5763
rect 2648 5732 2973 5760
rect 2648 5720 2654 5732
rect 2961 5729 2973 5732
rect 3007 5729 3019 5763
rect 2961 5723 3019 5729
rect 2041 5695 2099 5701
rect 2041 5661 2053 5695
rect 2087 5661 2099 5695
rect 2041 5655 2099 5661
rect 2225 5695 2283 5701
rect 2225 5661 2237 5695
rect 2271 5661 2283 5695
rect 2498 5692 2504 5704
rect 2459 5664 2504 5692
rect 2225 5655 2283 5661
rect 2056 5624 2084 5655
rect 2498 5652 2504 5664
rect 2556 5652 2562 5704
rect 2682 5692 2688 5704
rect 2643 5664 2688 5692
rect 2682 5652 2688 5664
rect 2740 5652 2746 5704
rect 2777 5695 2835 5701
rect 2777 5661 2789 5695
rect 2823 5661 2835 5695
rect 2777 5655 2835 5661
rect 2869 5695 2927 5701
rect 2869 5661 2881 5695
rect 2915 5692 2927 5695
rect 4080 5692 4108 5856
rect 4706 5828 4712 5840
rect 4667 5800 4712 5828
rect 4706 5788 4712 5800
rect 4764 5788 4770 5840
rect 6914 5788 6920 5840
rect 6972 5828 6978 5840
rect 7193 5831 7251 5837
rect 7193 5828 7205 5831
rect 6972 5800 7205 5828
rect 6972 5788 6978 5800
rect 7193 5797 7205 5800
rect 7239 5797 7251 5831
rect 17494 5828 17500 5840
rect 17455 5800 17500 5828
rect 7193 5791 7251 5797
rect 17494 5788 17500 5800
rect 17552 5788 17558 5840
rect 17770 5788 17776 5840
rect 17828 5828 17834 5840
rect 18325 5831 18383 5837
rect 18325 5828 18337 5831
rect 17828 5800 18337 5828
rect 17828 5788 17834 5800
rect 18325 5797 18337 5800
rect 18371 5797 18383 5831
rect 18325 5791 18383 5797
rect 5629 5763 5687 5769
rect 5629 5760 5641 5763
rect 2915 5664 4108 5692
rect 4356 5732 5641 5760
rect 2915 5661 2927 5664
rect 2869 5655 2927 5661
rect 2516 5624 2544 5652
rect 2056 5596 2544 5624
rect 2792 5624 2820 5655
rect 4356 5636 4384 5732
rect 5629 5729 5641 5732
rect 5675 5729 5687 5763
rect 8110 5760 8116 5772
rect 8071 5732 8116 5760
rect 5629 5723 5687 5729
rect 8110 5720 8116 5732
rect 8168 5720 8174 5772
rect 9490 5760 9496 5772
rect 8312 5732 9496 5760
rect 5534 5692 5540 5704
rect 5495 5664 5540 5692
rect 5534 5652 5540 5664
rect 5592 5652 5598 5704
rect 5997 5695 6055 5701
rect 5997 5661 6009 5695
rect 6043 5661 6055 5695
rect 6362 5692 6368 5704
rect 6323 5664 6368 5692
rect 5997 5655 6055 5661
rect 4249 5627 4307 5633
rect 2792 5596 2912 5624
rect 1581 5559 1639 5565
rect 1581 5525 1593 5559
rect 1627 5556 1639 5559
rect 2774 5556 2780 5568
rect 1627 5528 2780 5556
rect 1627 5525 1639 5528
rect 1581 5519 1639 5525
rect 2774 5516 2780 5528
rect 2832 5516 2838 5568
rect 2884 5556 2912 5596
rect 4249 5593 4261 5627
rect 4295 5624 4307 5627
rect 4338 5624 4344 5636
rect 4295 5596 4344 5624
rect 4295 5593 4307 5596
rect 4249 5587 4307 5593
rect 4338 5584 4344 5596
rect 4396 5584 4402 5636
rect 4433 5627 4491 5633
rect 4433 5593 4445 5627
rect 4479 5624 4491 5627
rect 4479 5596 4752 5624
rect 4479 5593 4491 5596
rect 4433 5587 4491 5593
rect 4724 5568 4752 5596
rect 4798 5584 4804 5636
rect 4856 5624 4862 5636
rect 4893 5627 4951 5633
rect 4893 5624 4905 5627
rect 4856 5596 4905 5624
rect 4856 5584 4862 5596
rect 4893 5593 4905 5596
rect 4939 5593 4951 5627
rect 5258 5624 5264 5636
rect 5219 5596 5264 5624
rect 4893 5587 4951 5593
rect 5258 5584 5264 5596
rect 5316 5584 5322 5636
rect 5442 5584 5448 5636
rect 5500 5624 5506 5636
rect 6012 5624 6040 5655
rect 6362 5652 6368 5664
rect 6420 5652 6426 5704
rect 7466 5692 7472 5704
rect 7427 5664 7472 5692
rect 7466 5652 7472 5664
rect 7524 5692 7530 5704
rect 8018 5692 8024 5704
rect 7524 5664 8024 5692
rect 7524 5652 7530 5664
rect 8018 5652 8024 5664
rect 8076 5652 8082 5704
rect 8312 5701 8340 5732
rect 9490 5720 9496 5732
rect 9548 5720 9554 5772
rect 10045 5763 10103 5769
rect 10045 5729 10057 5763
rect 10091 5760 10103 5763
rect 10594 5760 10600 5772
rect 10091 5732 10600 5760
rect 10091 5729 10103 5732
rect 10045 5723 10103 5729
rect 8297 5695 8355 5701
rect 8297 5661 8309 5695
rect 8343 5661 8355 5695
rect 8297 5655 8355 5661
rect 8481 5695 8539 5701
rect 8481 5661 8493 5695
rect 8527 5692 8539 5695
rect 8527 5664 9536 5692
rect 8527 5661 8539 5664
rect 8481 5655 8539 5661
rect 5500 5596 6040 5624
rect 7745 5627 7803 5633
rect 5500 5584 5506 5596
rect 7745 5593 7757 5627
rect 7791 5624 7803 5627
rect 9398 5624 9404 5636
rect 7791 5596 9404 5624
rect 7791 5593 7803 5596
rect 7745 5587 7803 5593
rect 9398 5584 9404 5596
rect 9456 5584 9462 5636
rect 9508 5624 9536 5664
rect 9582 5652 9588 5704
rect 9640 5692 9646 5704
rect 9677 5695 9735 5701
rect 9677 5692 9689 5695
rect 9640 5664 9689 5692
rect 9640 5652 9646 5664
rect 9677 5661 9689 5664
rect 9723 5661 9735 5695
rect 9950 5692 9956 5704
rect 9911 5664 9956 5692
rect 9677 5655 9735 5661
rect 9950 5652 9956 5664
rect 10008 5652 10014 5704
rect 10060 5624 10088 5723
rect 10594 5720 10600 5732
rect 10652 5720 10658 5772
rect 15197 5763 15255 5769
rect 15197 5729 15209 5763
rect 15243 5760 15255 5763
rect 15654 5760 15660 5772
rect 15243 5732 15660 5760
rect 15243 5729 15255 5732
rect 15197 5723 15255 5729
rect 15654 5720 15660 5732
rect 15712 5720 15718 5772
rect 15838 5720 15844 5772
rect 15896 5760 15902 5772
rect 17037 5763 17095 5769
rect 17037 5760 17049 5763
rect 15896 5732 17049 5760
rect 15896 5720 15902 5732
rect 17037 5729 17049 5732
rect 17083 5729 17095 5763
rect 17037 5723 17095 5729
rect 11514 5692 11520 5704
rect 11475 5664 11520 5692
rect 11514 5652 11520 5664
rect 11572 5652 11578 5704
rect 13173 5695 13231 5701
rect 13173 5661 13185 5695
rect 13219 5692 13231 5695
rect 13906 5692 13912 5704
rect 13219 5664 13912 5692
rect 13219 5661 13231 5664
rect 13173 5655 13231 5661
rect 13906 5652 13912 5664
rect 13964 5652 13970 5704
rect 14182 5692 14188 5704
rect 14143 5664 14188 5692
rect 14182 5652 14188 5664
rect 14240 5652 14246 5704
rect 14369 5695 14427 5701
rect 14369 5661 14381 5695
rect 14415 5661 14427 5695
rect 14369 5655 14427 5661
rect 9508 5596 10088 5624
rect 13722 5584 13728 5636
rect 13780 5624 13786 5636
rect 14384 5624 14412 5655
rect 14734 5652 14740 5704
rect 14792 5692 14798 5704
rect 14921 5695 14979 5701
rect 14921 5692 14933 5695
rect 14792 5664 14933 5692
rect 14792 5652 14798 5664
rect 14921 5661 14933 5664
rect 14967 5661 14979 5695
rect 14921 5655 14979 5661
rect 17865 5695 17923 5701
rect 17865 5661 17877 5695
rect 17911 5692 17923 5695
rect 18046 5692 18052 5704
rect 17911 5664 18052 5692
rect 17911 5661 17923 5664
rect 17865 5655 17923 5661
rect 18046 5652 18052 5664
rect 18104 5652 18110 5704
rect 13780 5596 14412 5624
rect 15304 5596 15686 5624
rect 13780 5584 13786 5596
rect 4614 5556 4620 5568
rect 2884 5528 4620 5556
rect 4614 5516 4620 5528
rect 4672 5516 4678 5568
rect 4706 5516 4712 5568
rect 4764 5556 4770 5568
rect 4985 5559 5043 5565
rect 4985 5556 4997 5559
rect 4764 5528 4997 5556
rect 4764 5516 4770 5528
rect 4985 5525 4997 5528
rect 5031 5525 5043 5559
rect 4985 5519 5043 5525
rect 5074 5516 5080 5568
rect 5132 5556 5138 5568
rect 6549 5559 6607 5565
rect 5132 5528 5177 5556
rect 5132 5516 5138 5528
rect 6549 5525 6561 5559
rect 6595 5556 6607 5559
rect 6730 5556 6736 5568
rect 6595 5528 6736 5556
rect 6595 5525 6607 5528
rect 6549 5519 6607 5525
rect 6730 5516 6736 5528
rect 6788 5516 6794 5568
rect 7006 5516 7012 5568
rect 7064 5556 7070 5568
rect 7653 5559 7711 5565
rect 7653 5556 7665 5559
rect 7064 5528 7665 5556
rect 7064 5516 7070 5528
rect 7653 5525 7665 5528
rect 7699 5556 7711 5559
rect 7926 5556 7932 5568
rect 7699 5528 7932 5556
rect 7699 5525 7711 5528
rect 7653 5519 7711 5525
rect 7926 5516 7932 5528
rect 7984 5516 7990 5568
rect 11330 5556 11336 5568
rect 11291 5528 11336 5556
rect 11330 5516 11336 5528
rect 11388 5516 11394 5568
rect 14461 5559 14519 5565
rect 14461 5525 14473 5559
rect 14507 5556 14519 5559
rect 15304 5556 15332 5596
rect 17586 5584 17592 5636
rect 17644 5624 17650 5636
rect 17644 5596 17689 5624
rect 17644 5584 17650 5596
rect 14507 5528 15332 5556
rect 14507 5525 14519 5528
rect 14461 5519 14519 5525
rect 16022 5516 16028 5568
rect 16080 5556 16086 5568
rect 16669 5559 16727 5565
rect 16669 5556 16681 5559
rect 16080 5528 16681 5556
rect 16080 5516 16086 5528
rect 16669 5525 16681 5528
rect 16715 5525 16727 5559
rect 16669 5519 16727 5525
rect 1104 5466 18860 5488
rect 1104 5414 8214 5466
rect 8266 5414 8278 5466
rect 8330 5414 8342 5466
rect 8394 5414 8406 5466
rect 8458 5414 8470 5466
rect 8522 5414 16214 5466
rect 16266 5414 16278 5466
rect 16330 5414 16342 5466
rect 16394 5414 16406 5466
rect 16458 5414 16470 5466
rect 16522 5414 18860 5466
rect 1104 5392 18860 5414
rect 3513 5355 3571 5361
rect 3513 5321 3525 5355
rect 3559 5352 3571 5355
rect 3694 5352 3700 5364
rect 3559 5324 3700 5352
rect 3559 5321 3571 5324
rect 3513 5315 3571 5321
rect 3694 5312 3700 5324
rect 3752 5312 3758 5364
rect 4065 5355 4123 5361
rect 4065 5321 4077 5355
rect 4111 5321 4123 5355
rect 4065 5315 4123 5321
rect 4525 5355 4583 5361
rect 4525 5321 4537 5355
rect 4571 5352 4583 5355
rect 4614 5352 4620 5364
rect 4571 5324 4620 5352
rect 4571 5321 4583 5324
rect 4525 5315 4583 5321
rect 2774 5244 2780 5296
rect 2832 5284 2838 5296
rect 4080 5284 4108 5315
rect 4614 5312 4620 5324
rect 4672 5312 4678 5364
rect 5258 5312 5264 5364
rect 5316 5352 5322 5364
rect 5353 5355 5411 5361
rect 5353 5352 5365 5355
rect 5316 5324 5365 5352
rect 5316 5312 5322 5324
rect 5353 5321 5365 5324
rect 5399 5321 5411 5355
rect 8754 5352 8760 5364
rect 8715 5324 8760 5352
rect 5353 5315 5411 5321
rect 8754 5312 8760 5324
rect 8812 5312 8818 5364
rect 10410 5312 10416 5364
rect 10468 5352 10474 5364
rect 10873 5355 10931 5361
rect 10873 5352 10885 5355
rect 10468 5324 10885 5352
rect 10468 5312 10474 5324
rect 10873 5321 10885 5324
rect 10919 5321 10931 5355
rect 10873 5315 10931 5321
rect 12802 5312 12808 5364
rect 12860 5352 12866 5364
rect 13357 5355 13415 5361
rect 13357 5352 13369 5355
rect 12860 5324 13369 5352
rect 12860 5312 12866 5324
rect 13357 5321 13369 5324
rect 13403 5321 13415 5355
rect 13357 5315 13415 5321
rect 14826 5312 14832 5364
rect 14884 5352 14890 5364
rect 15473 5355 15531 5361
rect 15473 5352 15485 5355
rect 14884 5324 15485 5352
rect 14884 5312 14890 5324
rect 15473 5321 15485 5324
rect 15519 5321 15531 5355
rect 15473 5315 15531 5321
rect 15746 5312 15752 5364
rect 15804 5352 15810 5364
rect 15841 5355 15899 5361
rect 15841 5352 15853 5355
rect 15804 5324 15853 5352
rect 15804 5312 15810 5324
rect 15841 5321 15853 5324
rect 15887 5321 15899 5355
rect 15841 5315 15899 5321
rect 16393 5355 16451 5361
rect 16393 5321 16405 5355
rect 16439 5352 16451 5355
rect 16574 5352 16580 5364
rect 16439 5324 16580 5352
rect 16439 5321 16451 5324
rect 16393 5315 16451 5321
rect 16574 5312 16580 5324
rect 16632 5352 16638 5364
rect 16761 5355 16819 5361
rect 16761 5352 16773 5355
rect 16632 5324 16773 5352
rect 16632 5312 16638 5324
rect 16761 5321 16773 5324
rect 16807 5321 16819 5355
rect 17310 5352 17316 5364
rect 17271 5324 17316 5352
rect 16761 5315 16819 5321
rect 5442 5284 5448 5296
rect 2832 5256 3188 5284
rect 4080 5256 5448 5284
rect 2832 5244 2838 5256
rect 3160 5225 3188 5256
rect 5442 5244 5448 5256
rect 5500 5244 5506 5296
rect 7282 5284 7288 5296
rect 7243 5256 7288 5284
rect 7282 5244 7288 5256
rect 7340 5244 7346 5296
rect 9122 5284 9128 5296
rect 8510 5256 9128 5284
rect 9122 5244 9128 5256
rect 9180 5244 9186 5296
rect 9401 5287 9459 5293
rect 9401 5253 9413 5287
rect 9447 5284 9459 5287
rect 9674 5284 9680 5296
rect 9447 5256 9680 5284
rect 9447 5253 9459 5256
rect 9401 5247 9459 5253
rect 9674 5244 9680 5256
rect 9732 5244 9738 5296
rect 10134 5244 10140 5296
rect 10192 5244 10198 5296
rect 11330 5244 11336 5296
rect 11388 5284 11394 5296
rect 11885 5287 11943 5293
rect 11885 5284 11897 5287
rect 11388 5256 11897 5284
rect 11388 5244 11394 5256
rect 11885 5253 11897 5256
rect 11931 5253 11943 5287
rect 11885 5247 11943 5253
rect 12618 5244 12624 5296
rect 12676 5244 12682 5296
rect 13998 5284 14004 5296
rect 13959 5256 14004 5284
rect 13998 5244 14004 5256
rect 14056 5244 14062 5296
rect 14458 5244 14464 5296
rect 14516 5244 14522 5296
rect 16776 5284 16804 5315
rect 17310 5312 17316 5324
rect 17368 5312 17374 5364
rect 17218 5284 17224 5296
rect 16776 5256 17224 5284
rect 17218 5244 17224 5256
rect 17276 5244 17282 5296
rect 17497 5287 17555 5293
rect 17497 5253 17509 5287
rect 17543 5284 17555 5287
rect 17586 5284 17592 5296
rect 17543 5256 17592 5284
rect 17543 5253 17555 5256
rect 17497 5247 17555 5253
rect 17586 5244 17592 5256
rect 17644 5244 17650 5296
rect 2501 5219 2559 5225
rect 2501 5185 2513 5219
rect 2547 5216 2559 5219
rect 2869 5219 2927 5225
rect 2869 5216 2881 5219
rect 2547 5188 2881 5216
rect 2547 5185 2559 5188
rect 2501 5179 2559 5185
rect 2869 5185 2881 5188
rect 2915 5185 2927 5219
rect 2869 5179 2927 5185
rect 3145 5219 3203 5225
rect 3145 5185 3157 5219
rect 3191 5216 3203 5219
rect 3234 5216 3240 5228
rect 3191 5188 3240 5216
rect 3191 5185 3203 5188
rect 3145 5179 3203 5185
rect 3234 5176 3240 5188
rect 3292 5176 3298 5228
rect 3973 5219 4031 5225
rect 3973 5185 3985 5219
rect 4019 5185 4031 5219
rect 4154 5216 4160 5228
rect 4115 5188 4160 5216
rect 3973 5179 4031 5185
rect 3988 5148 4016 5179
rect 4154 5176 4160 5188
rect 4212 5176 4218 5228
rect 4338 5176 4344 5228
rect 4396 5216 4402 5228
rect 4433 5219 4491 5225
rect 4433 5216 4445 5219
rect 4396 5188 4445 5216
rect 4396 5176 4402 5188
rect 4433 5185 4445 5188
rect 4479 5185 4491 5219
rect 4433 5179 4491 5185
rect 4614 5176 4620 5228
rect 4672 5216 4678 5228
rect 4801 5219 4859 5225
rect 4801 5216 4813 5219
rect 4672 5188 4813 5216
rect 4672 5176 4678 5188
rect 4801 5185 4813 5188
rect 4847 5185 4859 5219
rect 4801 5179 4859 5185
rect 4890 5176 4896 5228
rect 4948 5216 4954 5228
rect 5537 5219 5595 5225
rect 5537 5216 5549 5219
rect 4948 5188 5549 5216
rect 4948 5176 4954 5188
rect 5537 5185 5549 5188
rect 5583 5185 5595 5219
rect 5537 5179 5595 5185
rect 6733 5219 6791 5225
rect 6733 5185 6745 5219
rect 6779 5216 6791 5219
rect 6914 5216 6920 5228
rect 6779 5188 6920 5216
rect 6779 5185 6791 5188
rect 6733 5179 6791 5185
rect 6914 5176 6920 5188
rect 6972 5176 6978 5228
rect 13725 5219 13783 5225
rect 13725 5185 13737 5219
rect 13771 5185 13783 5219
rect 13725 5179 13783 5185
rect 4908 5148 4936 5176
rect 3988 5120 4936 5148
rect 4985 5151 5043 5157
rect 4985 5117 4997 5151
rect 5031 5117 5043 5151
rect 4985 5111 5043 5117
rect 4154 5040 4160 5092
rect 4212 5080 4218 5092
rect 4706 5080 4712 5092
rect 4212 5052 4712 5080
rect 4212 5040 4218 5052
rect 4706 5040 4712 5052
rect 4764 5040 4770 5092
rect 4798 5040 4804 5092
rect 4856 5080 4862 5092
rect 5000 5080 5028 5111
rect 5074 5108 5080 5160
rect 5132 5148 5138 5160
rect 5721 5151 5779 5157
rect 5721 5148 5733 5151
rect 5132 5120 5733 5148
rect 5132 5108 5138 5120
rect 5721 5117 5733 5120
rect 5767 5117 5779 5151
rect 5721 5111 5779 5117
rect 6178 5108 6184 5160
rect 6236 5148 6242 5160
rect 7009 5151 7067 5157
rect 7009 5148 7021 5151
rect 6236 5120 7021 5148
rect 6236 5108 6242 5120
rect 7009 5117 7021 5120
rect 7055 5148 7067 5151
rect 9125 5151 9183 5157
rect 9125 5148 9137 5151
rect 7055 5120 9137 5148
rect 7055 5117 7067 5120
rect 7009 5111 7067 5117
rect 9125 5117 9137 5120
rect 9171 5148 9183 5151
rect 9766 5148 9772 5160
rect 9171 5120 9772 5148
rect 9171 5117 9183 5120
rect 9125 5111 9183 5117
rect 9766 5108 9772 5120
rect 9824 5148 9830 5160
rect 11609 5151 11667 5157
rect 11609 5148 11621 5151
rect 9824 5120 11621 5148
rect 9824 5108 9830 5120
rect 11609 5117 11621 5120
rect 11655 5148 11667 5151
rect 11974 5148 11980 5160
rect 11655 5120 11980 5148
rect 11655 5117 11667 5120
rect 11609 5111 11667 5117
rect 11974 5108 11980 5120
rect 12032 5108 12038 5160
rect 13740 5148 13768 5179
rect 14734 5148 14740 5160
rect 13740 5120 14740 5148
rect 14734 5108 14740 5120
rect 14792 5108 14798 5160
rect 17678 5108 17684 5160
rect 17736 5148 17742 5160
rect 17957 5151 18015 5157
rect 17957 5148 17969 5151
rect 17736 5120 17969 5148
rect 17736 5108 17742 5120
rect 17957 5117 17969 5120
rect 18003 5117 18015 5151
rect 17957 5111 18015 5117
rect 4856 5052 5028 5080
rect 4856 5040 4862 5052
rect 2406 4972 2412 5024
rect 2464 5012 2470 5024
rect 2501 5015 2559 5021
rect 2501 5012 2513 5015
rect 2464 4984 2513 5012
rect 2464 4972 2470 4984
rect 2501 4981 2513 4984
rect 2547 4981 2559 5015
rect 2501 4975 2559 4981
rect 4062 4972 4068 5024
rect 4120 5012 4126 5024
rect 5997 5015 6055 5021
rect 5997 5012 6009 5015
rect 4120 4984 6009 5012
rect 4120 4972 4126 4984
rect 5997 4981 6009 4984
rect 6043 4981 6055 5015
rect 5997 4975 6055 4981
rect 6454 4972 6460 5024
rect 6512 5012 6518 5024
rect 6549 5015 6607 5021
rect 6549 5012 6561 5015
rect 6512 4984 6561 5012
rect 6512 4972 6518 4984
rect 6549 4981 6561 4984
rect 6595 4981 6607 5015
rect 6549 4975 6607 4981
rect 1104 4922 18860 4944
rect 1104 4870 4214 4922
rect 4266 4870 4278 4922
rect 4330 4870 4342 4922
rect 4394 4870 4406 4922
rect 4458 4870 4470 4922
rect 4522 4870 12214 4922
rect 12266 4870 12278 4922
rect 12330 4870 12342 4922
rect 12394 4870 12406 4922
rect 12458 4870 12470 4922
rect 12522 4870 18860 4922
rect 1104 4848 18860 4870
rect 2498 4808 2504 4820
rect 2459 4780 2504 4808
rect 2498 4768 2504 4780
rect 2556 4768 2562 4820
rect 2958 4808 2964 4820
rect 2919 4780 2964 4808
rect 2958 4768 2964 4780
rect 3016 4768 3022 4820
rect 4706 4768 4712 4820
rect 4764 4808 4770 4820
rect 5074 4808 5080 4820
rect 4764 4780 5080 4808
rect 4764 4768 4770 4780
rect 5074 4768 5080 4780
rect 5132 4768 5138 4820
rect 6546 4808 6552 4820
rect 6012 4780 6552 4808
rect 2976 4740 3004 4768
rect 2976 4712 4476 4740
rect 1673 4675 1731 4681
rect 1673 4641 1685 4675
rect 1719 4672 1731 4675
rect 1762 4672 1768 4684
rect 1719 4644 1768 4672
rect 1719 4641 1731 4644
rect 1673 4635 1731 4641
rect 1762 4632 1768 4644
rect 1820 4672 1826 4684
rect 4062 4672 4068 4684
rect 1820 4644 4068 4672
rect 1820 4632 1826 4644
rect 4062 4632 4068 4644
rect 4120 4632 4126 4684
rect 1857 4607 1915 4613
rect 1857 4573 1869 4607
rect 1903 4604 1915 4607
rect 2130 4604 2136 4616
rect 1903 4576 2136 4604
rect 1903 4573 1915 4576
rect 1857 4567 1915 4573
rect 2130 4564 2136 4576
rect 2188 4564 2194 4616
rect 2590 4604 2596 4616
rect 2551 4576 2596 4604
rect 2590 4564 2596 4576
rect 2648 4564 2654 4616
rect 3513 4607 3571 4613
rect 3513 4573 3525 4607
rect 3559 4573 3571 4607
rect 4246 4604 4252 4616
rect 4207 4576 4252 4604
rect 3513 4567 3571 4573
rect 3528 4536 3556 4567
rect 4246 4564 4252 4576
rect 4304 4564 4310 4616
rect 4448 4613 4476 4712
rect 5261 4675 5319 4681
rect 5261 4641 5273 4675
rect 5307 4672 5319 4675
rect 5534 4672 5540 4684
rect 5307 4644 5540 4672
rect 5307 4641 5319 4644
rect 5261 4635 5319 4641
rect 5534 4632 5540 4644
rect 5592 4632 5598 4684
rect 6012 4616 6040 4780
rect 6546 4768 6552 4780
rect 6604 4808 6610 4820
rect 7926 4808 7932 4820
rect 6604 4780 7512 4808
rect 7887 4780 7932 4808
rect 6604 4768 6610 4780
rect 7484 4740 7512 4780
rect 7926 4768 7932 4780
rect 7984 4768 7990 4820
rect 11241 4811 11299 4817
rect 11241 4777 11253 4811
rect 11287 4808 11299 4811
rect 13538 4808 13544 4820
rect 11287 4780 13544 4808
rect 11287 4777 11299 4780
rect 11241 4771 11299 4777
rect 13538 4768 13544 4780
rect 13596 4768 13602 4820
rect 13814 4808 13820 4820
rect 13648 4780 13820 4808
rect 10134 4740 10140 4752
rect 7484 4712 7880 4740
rect 10095 4712 10140 4740
rect 7852 4684 7880 4712
rect 10134 4700 10140 4712
rect 10192 4700 10198 4752
rect 6454 4672 6460 4684
rect 6415 4644 6460 4672
rect 6454 4632 6460 4644
rect 6512 4632 6518 4684
rect 7834 4632 7840 4684
rect 7892 4672 7898 4684
rect 7892 4644 8708 4672
rect 7892 4632 7898 4644
rect 4433 4607 4491 4613
rect 4433 4573 4445 4607
rect 4479 4573 4491 4607
rect 4890 4604 4896 4616
rect 4851 4576 4896 4604
rect 4433 4567 4491 4573
rect 4890 4564 4896 4576
rect 4948 4564 4954 4616
rect 5074 4604 5080 4616
rect 5035 4576 5080 4604
rect 5074 4564 5080 4576
rect 5132 4564 5138 4616
rect 5629 4607 5687 4613
rect 5629 4573 5641 4607
rect 5675 4573 5687 4607
rect 5629 4567 5687 4573
rect 5905 4607 5963 4613
rect 5905 4573 5917 4607
rect 5951 4604 5963 4607
rect 5994 4604 6000 4616
rect 5951 4576 6000 4604
rect 5951 4573 5963 4576
rect 5905 4567 5963 4573
rect 4522 4536 4528 4548
rect 3528 4508 4528 4536
rect 4522 4496 4528 4508
rect 4580 4496 4586 4548
rect 4617 4539 4675 4545
rect 4617 4505 4629 4539
rect 4663 4536 4675 4539
rect 5644 4536 5672 4567
rect 5994 4564 6000 4576
rect 6052 4564 6058 4616
rect 6178 4604 6184 4616
rect 6139 4576 6184 4604
rect 6178 4564 6184 4576
rect 6236 4564 6242 4616
rect 8680 4613 8708 4644
rect 9122 4632 9128 4684
rect 9180 4672 9186 4684
rect 9217 4675 9275 4681
rect 9217 4672 9229 4675
rect 9180 4644 9229 4672
rect 9180 4632 9186 4644
rect 9217 4641 9229 4644
rect 9263 4641 9275 4675
rect 9217 4635 9275 4641
rect 9324 4644 10088 4672
rect 9324 4616 9352 4644
rect 8389 4607 8447 4613
rect 8389 4573 8401 4607
rect 8435 4573 8447 4607
rect 8389 4567 8447 4573
rect 8665 4607 8723 4613
rect 8665 4573 8677 4607
rect 8711 4573 8723 4607
rect 9306 4604 9312 4616
rect 9267 4576 9312 4604
rect 8665 4567 8723 4573
rect 8297 4539 8355 4545
rect 8297 4536 8309 4539
rect 4663 4508 6868 4536
rect 7682 4508 8309 4536
rect 4663 4505 4675 4508
rect 4617 4499 4675 4505
rect 1854 4428 1860 4480
rect 1912 4468 1918 4480
rect 2041 4471 2099 4477
rect 2041 4468 2053 4471
rect 1912 4440 2053 4468
rect 1912 4428 1918 4440
rect 2041 4437 2053 4440
rect 2087 4437 2099 4471
rect 3326 4468 3332 4480
rect 3287 4440 3332 4468
rect 2041 4431 2099 4437
rect 3326 4428 3332 4440
rect 3384 4428 3390 4480
rect 3973 4471 4031 4477
rect 3973 4437 3985 4471
rect 4019 4468 4031 4471
rect 4246 4468 4252 4480
rect 4019 4440 4252 4468
rect 4019 4437 4031 4440
rect 3973 4431 4031 4437
rect 4246 4428 4252 4440
rect 4304 4468 4310 4480
rect 4706 4468 4712 4480
rect 4304 4440 4712 4468
rect 4304 4428 4310 4440
rect 4706 4428 4712 4440
rect 4764 4428 4770 4480
rect 4982 4428 4988 4480
rect 5040 4468 5046 4480
rect 5629 4471 5687 4477
rect 5629 4468 5641 4471
rect 5040 4440 5641 4468
rect 5040 4428 5046 4440
rect 5629 4437 5641 4440
rect 5675 4437 5687 4471
rect 6840 4468 6868 4508
rect 8297 4505 8309 4508
rect 8343 4505 8355 4539
rect 8297 4499 8355 4505
rect 8404 4468 8432 4567
rect 8570 4468 8576 4480
rect 6840 4440 8576 4468
rect 5629 4431 5687 4437
rect 8570 4428 8576 4440
rect 8628 4428 8634 4480
rect 8680 4468 8708 4567
rect 9306 4564 9312 4576
rect 9364 4564 9370 4616
rect 10060 4613 10088 4644
rect 11974 4632 11980 4684
rect 12032 4672 12038 4684
rect 12989 4675 13047 4681
rect 12989 4672 13001 4675
rect 12032 4644 13001 4672
rect 12032 4632 12038 4644
rect 12989 4641 13001 4644
rect 13035 4672 13047 4675
rect 13648 4672 13676 4780
rect 13814 4768 13820 4780
rect 13872 4808 13878 4820
rect 14369 4811 14427 4817
rect 14369 4808 14381 4811
rect 13872 4780 14381 4808
rect 13872 4768 13878 4780
rect 14369 4777 14381 4780
rect 14415 4777 14427 4811
rect 14369 4771 14427 4777
rect 16114 4768 16120 4820
rect 16172 4808 16178 4820
rect 16485 4811 16543 4817
rect 16485 4808 16497 4811
rect 16172 4780 16497 4808
rect 16172 4768 16178 4780
rect 16485 4777 16497 4780
rect 16531 4777 16543 4811
rect 16485 4771 16543 4777
rect 13725 4743 13783 4749
rect 13725 4709 13737 4743
rect 13771 4740 13783 4743
rect 14458 4740 14464 4752
rect 13771 4712 14464 4740
rect 13771 4709 13783 4712
rect 13725 4703 13783 4709
rect 14458 4700 14464 4712
rect 14516 4700 14522 4752
rect 14734 4672 14740 4684
rect 13035 4644 13492 4672
rect 13035 4641 13047 4644
rect 12989 4635 13047 4641
rect 9585 4607 9643 4613
rect 9585 4573 9597 4607
rect 9631 4604 9643 4607
rect 9953 4607 10011 4613
rect 9953 4604 9965 4607
rect 9631 4576 9965 4604
rect 9631 4573 9643 4576
rect 9585 4567 9643 4573
rect 9953 4573 9965 4576
rect 9999 4573 10011 4607
rect 9953 4567 10011 4573
rect 10045 4607 10103 4613
rect 10045 4573 10057 4607
rect 10091 4573 10103 4607
rect 10045 4567 10103 4573
rect 9968 4536 9996 4567
rect 10870 4536 10876 4548
rect 9968 4508 10876 4536
rect 10870 4496 10876 4508
rect 10928 4496 10934 4548
rect 11974 4496 11980 4548
rect 12032 4496 12038 4548
rect 12710 4536 12716 4548
rect 12671 4508 12716 4536
rect 12710 4496 12716 4508
rect 12768 4496 12774 4548
rect 13464 4536 13492 4644
rect 13556 4644 13676 4672
rect 14695 4644 14740 4672
rect 13556 4613 13584 4644
rect 14734 4632 14740 4644
rect 14792 4632 14798 4684
rect 16850 4632 16856 4684
rect 16908 4672 16914 4684
rect 17681 4675 17739 4681
rect 17681 4672 17693 4675
rect 16908 4644 17693 4672
rect 16908 4632 16914 4644
rect 17681 4641 17693 4644
rect 17727 4641 17739 4675
rect 17681 4635 17739 4641
rect 13541 4607 13599 4613
rect 13541 4573 13553 4607
rect 13587 4573 13599 4607
rect 13722 4604 13728 4616
rect 13683 4576 13728 4604
rect 13541 4567 13599 4573
rect 13722 4564 13728 4576
rect 13780 4564 13786 4616
rect 13906 4564 13912 4616
rect 13964 4604 13970 4616
rect 14185 4607 14243 4613
rect 14185 4604 14197 4607
rect 13964 4576 14197 4604
rect 13964 4564 13970 4576
rect 14185 4573 14197 4576
rect 14231 4573 14243 4607
rect 14185 4567 14243 4573
rect 14752 4536 14780 4632
rect 17126 4604 17132 4616
rect 17087 4576 17132 4604
rect 17126 4564 17132 4576
rect 17184 4564 17190 4616
rect 17218 4564 17224 4616
rect 17276 4604 17282 4616
rect 17589 4607 17647 4613
rect 17276 4576 17321 4604
rect 17276 4564 17282 4576
rect 17589 4573 17601 4607
rect 17635 4573 17647 4607
rect 18046 4604 18052 4616
rect 18007 4576 18052 4604
rect 17589 4567 17647 4573
rect 13464 4508 14780 4536
rect 15013 4539 15071 4545
rect 15013 4505 15025 4539
rect 15059 4536 15071 4539
rect 15286 4536 15292 4548
rect 15059 4508 15292 4536
rect 15059 4505 15071 4508
rect 15013 4499 15071 4505
rect 15286 4496 15292 4508
rect 15344 4496 15350 4548
rect 15470 4496 15476 4548
rect 15528 4496 15534 4548
rect 16942 4536 16948 4548
rect 16903 4508 16948 4536
rect 16942 4496 16948 4508
rect 17000 4496 17006 4548
rect 17034 4496 17040 4548
rect 17092 4536 17098 4548
rect 17604 4536 17632 4567
rect 18046 4564 18052 4576
rect 18104 4564 18110 4616
rect 17092 4508 17632 4536
rect 17092 4496 17098 4508
rect 16022 4468 16028 4480
rect 8680 4440 16028 4468
rect 16022 4428 16028 4440
rect 16080 4428 16086 4480
rect 1104 4378 18860 4400
rect 1104 4326 8214 4378
rect 8266 4326 8278 4378
rect 8330 4326 8342 4378
rect 8394 4326 8406 4378
rect 8458 4326 8470 4378
rect 8522 4326 16214 4378
rect 16266 4326 16278 4378
rect 16330 4326 16342 4378
rect 16394 4326 16406 4378
rect 16458 4326 16470 4378
rect 16522 4326 18860 4378
rect 1104 4304 18860 4326
rect 2498 4224 2504 4276
rect 2556 4224 2562 4276
rect 4157 4267 4215 4273
rect 4157 4233 4169 4267
rect 4203 4264 4215 4267
rect 4890 4264 4896 4276
rect 4203 4236 4896 4264
rect 4203 4233 4215 4236
rect 4157 4227 4215 4233
rect 4890 4224 4896 4236
rect 4948 4264 4954 4276
rect 5077 4267 5135 4273
rect 5077 4264 5089 4267
rect 4948 4236 5089 4264
rect 4948 4224 4954 4236
rect 5077 4233 5089 4236
rect 5123 4233 5135 4267
rect 11974 4264 11980 4276
rect 11935 4236 11980 4264
rect 5077 4227 5135 4233
rect 11974 4224 11980 4236
rect 12032 4224 12038 4276
rect 12618 4264 12624 4276
rect 12579 4236 12624 4264
rect 12618 4224 12624 4236
rect 12676 4224 12682 4276
rect 14185 4267 14243 4273
rect 14185 4233 14197 4267
rect 14231 4264 14243 4267
rect 15470 4264 15476 4276
rect 14231 4236 15476 4264
rect 14231 4233 14243 4236
rect 14185 4227 14243 4233
rect 15470 4224 15476 4236
rect 15528 4224 15534 4276
rect 16853 4267 16911 4273
rect 16853 4233 16865 4267
rect 16899 4264 16911 4267
rect 17034 4264 17040 4276
rect 16899 4236 17040 4264
rect 16899 4233 16911 4236
rect 16853 4227 16911 4233
rect 17034 4224 17040 4236
rect 17092 4224 17098 4276
rect 17218 4224 17224 4276
rect 17276 4264 17282 4276
rect 17276 4236 18092 4264
rect 17276 4224 17282 4236
rect 1670 4196 1676 4208
rect 1631 4168 1676 4196
rect 1670 4156 1676 4168
rect 1728 4156 1734 4208
rect 2133 4199 2191 4205
rect 2133 4165 2145 4199
rect 2179 4196 2191 4199
rect 2516 4196 2544 4224
rect 4982 4196 4988 4208
rect 2179 4168 2544 4196
rect 3910 4168 4988 4196
rect 2179 4165 2191 4168
rect 2133 4159 2191 4165
rect 4982 4156 4988 4168
rect 5040 4156 5046 4208
rect 7466 4156 7472 4208
rect 7524 4156 7530 4208
rect 9306 4156 9312 4208
rect 9364 4196 9370 4208
rect 13722 4196 13728 4208
rect 9364 4168 13728 4196
rect 9364 4156 9370 4168
rect 1854 4128 1860 4140
rect 1815 4100 1860 4128
rect 1854 4088 1860 4100
rect 1912 4088 1918 4140
rect 2041 4131 2099 4137
rect 2041 4097 2053 4131
rect 2087 4128 2099 4131
rect 2222 4128 2228 4140
rect 2087 4100 2228 4128
rect 2087 4097 2099 4100
rect 2041 4091 2099 4097
rect 2222 4088 2228 4100
rect 2280 4088 2286 4140
rect 2406 4128 2412 4140
rect 2367 4100 2412 4128
rect 2406 4088 2412 4100
rect 2464 4088 2470 4140
rect 5626 4128 5632 4140
rect 5587 4100 5632 4128
rect 5626 4088 5632 4100
rect 5684 4088 5690 4140
rect 5810 4128 5816 4140
rect 5771 4100 5816 4128
rect 5810 4088 5816 4100
rect 5868 4088 5874 4140
rect 8570 4128 8576 4140
rect 8531 4100 8576 4128
rect 8570 4088 8576 4100
rect 8628 4128 8634 4140
rect 9125 4131 9183 4137
rect 9125 4128 9137 4131
rect 8628 4100 9137 4128
rect 8628 4088 8634 4100
rect 9125 4097 9137 4100
rect 9171 4097 9183 4131
rect 9858 4128 9864 4140
rect 9819 4100 9864 4128
rect 9125 4091 9183 4097
rect 9858 4088 9864 4100
rect 9916 4088 9922 4140
rect 10045 4131 10103 4137
rect 10045 4097 10057 4131
rect 10091 4128 10103 4131
rect 10410 4128 10416 4140
rect 10091 4100 10416 4128
rect 10091 4097 10103 4100
rect 10045 4091 10103 4097
rect 10410 4088 10416 4100
rect 10468 4088 10474 4140
rect 10594 4128 10600 4140
rect 10555 4100 10600 4128
rect 10594 4088 10600 4100
rect 10652 4088 10658 4140
rect 11808 4137 11836 4168
rect 11793 4131 11851 4137
rect 11793 4097 11805 4131
rect 11839 4097 11851 4131
rect 11793 4091 11851 4097
rect 12069 4131 12127 4137
rect 12069 4097 12081 4131
rect 12115 4128 12127 4131
rect 12434 4128 12440 4140
rect 12115 4100 12440 4128
rect 12115 4097 12127 4100
rect 12406 4098 12440 4100
rect 12069 4091 12127 4097
rect 2685 4063 2743 4069
rect 2685 4029 2697 4063
rect 2731 4060 2743 4063
rect 3326 4060 3332 4072
rect 2731 4032 3332 4060
rect 2731 4029 2743 4032
rect 2685 4023 2743 4029
rect 3326 4020 3332 4032
rect 3384 4020 3390 4072
rect 4985 4063 5043 4069
rect 4985 4029 4997 4063
rect 5031 4029 5043 4063
rect 5166 4060 5172 4072
rect 5127 4032 5172 4060
rect 4985 4023 5043 4029
rect 4522 3952 4528 4004
rect 4580 3992 4586 4004
rect 4617 3995 4675 4001
rect 4617 3992 4629 3995
rect 4580 3964 4629 3992
rect 4580 3952 4586 3964
rect 4617 3961 4629 3964
rect 4663 3961 4675 3995
rect 5000 3992 5028 4023
rect 5166 4020 5172 4032
rect 5224 4020 5230 4072
rect 5534 4060 5540 4072
rect 5495 4032 5540 4060
rect 5534 4020 5540 4032
rect 5592 4020 5598 4072
rect 5718 4020 5724 4072
rect 5776 4060 5782 4072
rect 6178 4060 6184 4072
rect 5776 4032 6184 4060
rect 5776 4020 5782 4032
rect 6178 4020 6184 4032
rect 6236 4060 6242 4072
rect 6457 4063 6515 4069
rect 6457 4060 6469 4063
rect 6236 4032 6469 4060
rect 6236 4020 6242 4032
rect 6457 4029 6469 4032
rect 6503 4029 6515 4063
rect 6730 4060 6736 4072
rect 6691 4032 6736 4060
rect 6457 4023 6515 4029
rect 6730 4020 6736 4032
rect 6788 4020 6794 4072
rect 7742 4020 7748 4072
rect 7800 4060 7806 4072
rect 9674 4060 9680 4072
rect 7800 4032 9444 4060
rect 9635 4032 9680 4060
rect 7800 4020 7806 4032
rect 5074 3992 5080 4004
rect 4987 3964 5080 3992
rect 4617 3955 4675 3961
rect 5074 3952 5080 3964
rect 5132 3992 5138 4004
rect 5132 3964 6500 3992
rect 5132 3952 5138 3964
rect 6472 3936 6500 3964
rect 8478 3952 8484 4004
rect 8536 3992 8542 4004
rect 9306 3992 9312 4004
rect 8536 3964 9312 3992
rect 8536 3952 8542 3964
rect 9306 3952 9312 3964
rect 9364 3952 9370 4004
rect 9416 3992 9444 4032
rect 9674 4020 9680 4032
rect 9732 4020 9738 4072
rect 10778 4060 10784 4072
rect 10739 4032 10784 4060
rect 10778 4020 10784 4032
rect 10836 4020 10842 4072
rect 10870 4020 10876 4072
rect 10928 4060 10934 4072
rect 12084 4060 12112 4091
rect 12434 4088 12440 4098
rect 12492 4128 12498 4140
rect 13188 4137 13216 4168
rect 13722 4156 13728 4168
rect 13780 4156 13786 4208
rect 16666 4196 16672 4208
rect 16054 4168 16672 4196
rect 16666 4156 16672 4168
rect 16724 4156 16730 4208
rect 17126 4156 17132 4208
rect 17184 4196 17190 4208
rect 17954 4196 17960 4208
rect 17184 4168 17816 4196
rect 17915 4168 17960 4196
rect 17184 4156 17190 4168
rect 12621 4131 12679 4137
rect 12492 4100 12537 4128
rect 12492 4088 12498 4100
rect 12621 4097 12633 4131
rect 12667 4128 12679 4131
rect 13173 4131 13231 4137
rect 12667 4100 13124 4128
rect 12667 4097 12679 4100
rect 12621 4091 12679 4097
rect 12636 4060 12664 4091
rect 12986 4060 12992 4072
rect 10928 4032 12112 4060
rect 12360 4032 12664 4060
rect 12947 4032 12992 4060
rect 10928 4020 10934 4032
rect 12360 3992 12388 4032
rect 12986 4020 12992 4032
rect 13044 4020 13050 4072
rect 13096 4060 13124 4100
rect 13173 4097 13185 4131
rect 13219 4097 13231 4131
rect 13173 4091 13231 4097
rect 13357 4131 13415 4137
rect 13357 4097 13369 4131
rect 13403 4128 13415 4131
rect 13814 4128 13820 4140
rect 13403 4100 13820 4128
rect 13403 4097 13415 4100
rect 13357 4091 13415 4097
rect 13814 4088 13820 4100
rect 13872 4088 13878 4140
rect 14001 4131 14059 4137
rect 14001 4097 14013 4131
rect 14047 4128 14059 4131
rect 14090 4128 14096 4140
rect 14047 4100 14096 4128
rect 14047 4097 14059 4100
rect 14001 4091 14059 4097
rect 14090 4088 14096 4100
rect 14148 4088 14154 4140
rect 14185 4131 14243 4137
rect 14185 4097 14197 4131
rect 14231 4097 14243 4131
rect 14185 4091 14243 4097
rect 17037 4131 17095 4137
rect 17037 4097 17049 4131
rect 17083 4128 17095 4131
rect 17678 4128 17684 4140
rect 17083 4100 17540 4128
rect 17639 4100 17684 4128
rect 17083 4097 17095 4100
rect 17037 4091 17095 4097
rect 14200 4060 14228 4091
rect 14366 4060 14372 4072
rect 13096 4032 14372 4060
rect 14366 4020 14372 4032
rect 14424 4020 14430 4072
rect 14550 4060 14556 4072
rect 14511 4032 14556 4060
rect 14550 4020 14556 4032
rect 14608 4020 14614 4072
rect 14829 4063 14887 4069
rect 14829 4029 14841 4063
rect 14875 4060 14887 4063
rect 16574 4060 16580 4072
rect 14875 4032 16580 4060
rect 14875 4029 14887 4032
rect 14829 4023 14887 4029
rect 16574 4020 16580 4032
rect 16632 4020 16638 4072
rect 17313 4063 17371 4069
rect 17313 4029 17325 4063
rect 17359 4029 17371 4063
rect 17512 4060 17540 4100
rect 17678 4088 17684 4100
rect 17736 4088 17742 4140
rect 17788 4128 17816 4168
rect 17954 4156 17960 4168
rect 18012 4156 18018 4208
rect 18064 4196 18092 4236
rect 18064 4168 18184 4196
rect 18049 4131 18107 4137
rect 18049 4128 18061 4131
rect 17788 4100 18061 4128
rect 18049 4097 18061 4100
rect 18095 4097 18107 4131
rect 18156 4128 18184 4168
rect 18230 4128 18236 4140
rect 18156 4100 18236 4128
rect 18049 4091 18107 4097
rect 18230 4088 18236 4100
rect 18288 4128 18294 4140
rect 18288 4100 18381 4128
rect 18288 4088 18294 4100
rect 18322 4060 18328 4072
rect 17512 4032 18328 4060
rect 17313 4023 17371 4029
rect 9416 3964 12388 3992
rect 16114 3952 16120 4004
rect 16172 3992 16178 4004
rect 17126 3992 17132 4004
rect 16172 3964 17132 3992
rect 16172 3952 16178 3964
rect 17126 3952 17132 3964
rect 17184 3992 17190 4004
rect 17328 3992 17356 4023
rect 18322 4020 18328 4032
rect 18380 4020 18386 4072
rect 17184 3964 17356 3992
rect 17184 3952 17190 3964
rect 6454 3884 6460 3936
rect 6512 3884 6518 3936
rect 6730 3884 6736 3936
rect 6788 3924 6794 3936
rect 8205 3927 8263 3933
rect 8205 3924 8217 3927
rect 6788 3896 8217 3924
rect 6788 3884 6794 3896
rect 8205 3893 8217 3896
rect 8251 3893 8263 3927
rect 8205 3887 8263 3893
rect 8757 3927 8815 3933
rect 8757 3893 8769 3927
rect 8803 3924 8815 3927
rect 9214 3924 9220 3936
rect 8803 3896 9220 3924
rect 8803 3893 8815 3896
rect 8757 3887 8815 3893
rect 9214 3884 9220 3896
rect 9272 3884 9278 3936
rect 10410 3924 10416 3936
rect 10371 3896 10416 3924
rect 10410 3884 10416 3896
rect 10468 3884 10474 3936
rect 12434 3884 12440 3936
rect 12492 3924 12498 3936
rect 14182 3924 14188 3936
rect 12492 3896 14188 3924
rect 12492 3884 12498 3896
rect 14182 3884 14188 3896
rect 14240 3884 14246 3936
rect 16301 3927 16359 3933
rect 16301 3893 16313 3927
rect 16347 3924 16359 3927
rect 16758 3924 16764 3936
rect 16347 3896 16764 3924
rect 16347 3893 16359 3896
rect 16301 3887 16359 3893
rect 16758 3884 16764 3896
rect 16816 3884 16822 3936
rect 17494 3884 17500 3936
rect 17552 3924 17558 3936
rect 17681 3927 17739 3933
rect 17681 3924 17693 3927
rect 17552 3896 17693 3924
rect 17552 3884 17558 3896
rect 17681 3893 17693 3896
rect 17727 3893 17739 3927
rect 17681 3887 17739 3893
rect 1104 3834 18860 3856
rect 1104 3782 4214 3834
rect 4266 3782 4278 3834
rect 4330 3782 4342 3834
rect 4394 3782 4406 3834
rect 4458 3782 4470 3834
rect 4522 3782 12214 3834
rect 12266 3782 12278 3834
rect 12330 3782 12342 3834
rect 12394 3782 12406 3834
rect 12458 3782 12470 3834
rect 12522 3782 18860 3834
rect 1104 3760 18860 3782
rect 2777 3723 2835 3729
rect 2777 3689 2789 3723
rect 2823 3720 2835 3723
rect 3142 3720 3148 3732
rect 2823 3692 3148 3720
rect 2823 3689 2835 3692
rect 2777 3683 2835 3689
rect 3142 3680 3148 3692
rect 3200 3680 3206 3732
rect 6273 3723 6331 3729
rect 6273 3689 6285 3723
rect 6319 3720 6331 3723
rect 6362 3720 6368 3732
rect 6319 3692 6368 3720
rect 6319 3689 6331 3692
rect 6273 3683 6331 3689
rect 6362 3680 6368 3692
rect 6420 3680 6426 3732
rect 6454 3680 6460 3732
rect 6512 3720 6518 3732
rect 10778 3720 10784 3732
rect 6512 3692 10784 3720
rect 6512 3680 6518 3692
rect 10778 3680 10784 3692
rect 10836 3720 10842 3732
rect 13357 3723 13415 3729
rect 13357 3720 13369 3723
rect 10836 3692 13369 3720
rect 10836 3680 10842 3692
rect 4614 3612 4620 3664
rect 4672 3652 4678 3664
rect 6733 3655 6791 3661
rect 6733 3652 6745 3655
rect 4672 3624 6745 3652
rect 4672 3612 4678 3624
rect 6733 3621 6745 3624
rect 6779 3621 6791 3655
rect 6733 3615 6791 3621
rect 9398 3612 9404 3664
rect 9456 3652 9462 3664
rect 9456 3624 10732 3652
rect 9456 3612 9462 3624
rect 1854 3544 1860 3596
rect 1912 3584 1918 3596
rect 2133 3587 2191 3593
rect 2133 3584 2145 3587
rect 1912 3556 2145 3584
rect 1912 3544 1918 3556
rect 2133 3553 2145 3556
rect 2179 3553 2191 3587
rect 2133 3547 2191 3553
rect 2222 3544 2228 3596
rect 2280 3584 2286 3596
rect 2409 3587 2467 3593
rect 2409 3584 2421 3587
rect 2280 3556 2421 3584
rect 2280 3544 2286 3556
rect 2409 3553 2421 3556
rect 2455 3553 2467 3587
rect 3878 3584 3884 3596
rect 3839 3556 3884 3584
rect 2409 3547 2467 3553
rect 3878 3544 3884 3556
rect 3936 3544 3942 3596
rect 5166 3544 5172 3596
rect 5224 3584 5230 3596
rect 5442 3584 5448 3596
rect 5224 3556 5448 3584
rect 5224 3544 5230 3556
rect 5442 3544 5448 3556
rect 5500 3584 5506 3596
rect 5721 3587 5779 3593
rect 5721 3584 5733 3587
rect 5500 3556 5733 3584
rect 5500 3544 5506 3556
rect 5721 3553 5733 3556
rect 5767 3553 5779 3587
rect 7466 3584 7472 3596
rect 7427 3556 7472 3584
rect 5721 3547 5779 3553
rect 7466 3544 7472 3556
rect 7524 3544 7530 3596
rect 8570 3584 8576 3596
rect 7668 3556 8576 3584
rect 7668 3528 7696 3556
rect 8570 3544 8576 3556
rect 8628 3544 8634 3596
rect 9048 3556 9720 3584
rect 1673 3519 1731 3525
rect 1673 3485 1685 3519
rect 1719 3516 1731 3519
rect 1762 3516 1768 3528
rect 1719 3488 1768 3516
rect 1719 3485 1731 3488
rect 1673 3479 1731 3485
rect 1762 3476 1768 3488
rect 1820 3476 1826 3528
rect 3234 3476 3240 3528
rect 3292 3516 3298 3528
rect 3329 3519 3387 3525
rect 3329 3516 3341 3519
rect 3292 3488 3341 3516
rect 3292 3476 3298 3488
rect 3329 3485 3341 3488
rect 3375 3485 3387 3519
rect 4614 3516 4620 3528
rect 4575 3488 4620 3516
rect 3329 3479 3387 3485
rect 4614 3476 4620 3488
rect 4672 3476 4678 3528
rect 4893 3519 4951 3525
rect 4893 3485 4905 3519
rect 4939 3516 4951 3519
rect 5534 3516 5540 3528
rect 4939 3488 5540 3516
rect 4939 3485 4951 3488
rect 4893 3479 4951 3485
rect 5534 3476 5540 3488
rect 5592 3476 5598 3528
rect 6638 3516 6644 3528
rect 6599 3488 6644 3516
rect 6638 3476 6644 3488
rect 6696 3476 6702 3528
rect 7098 3516 7104 3528
rect 7059 3488 7104 3516
rect 7098 3476 7104 3488
rect 7156 3476 7162 3528
rect 7650 3516 7656 3528
rect 7563 3488 7656 3516
rect 7650 3476 7656 3488
rect 7708 3476 7714 3528
rect 7834 3516 7840 3528
rect 7795 3488 7840 3516
rect 7834 3476 7840 3488
rect 7892 3476 7898 3528
rect 8478 3516 8484 3528
rect 8439 3488 8484 3516
rect 8478 3476 8484 3488
rect 8536 3476 8542 3528
rect 8662 3516 8668 3528
rect 8623 3488 8668 3516
rect 8662 3476 8668 3488
rect 8720 3476 8726 3528
rect 9048 3525 9076 3556
rect 9033 3519 9091 3525
rect 9033 3485 9045 3519
rect 9079 3485 9091 3519
rect 9033 3479 9091 3485
rect 9125 3519 9183 3525
rect 9125 3485 9137 3519
rect 9171 3485 9183 3519
rect 9125 3479 9183 3485
rect 9309 3519 9367 3525
rect 9309 3485 9321 3519
rect 9355 3516 9367 3519
rect 9398 3516 9404 3528
rect 9355 3488 9404 3516
rect 9355 3485 9367 3488
rect 9309 3479 9367 3485
rect 2590 3448 2596 3460
rect 2551 3420 2596 3448
rect 2590 3408 2596 3420
rect 2648 3408 2654 3460
rect 2774 3408 2780 3460
rect 2832 3448 2838 3460
rect 5261 3451 5319 3457
rect 5261 3448 5273 3451
rect 2832 3420 5273 3448
rect 2832 3408 2838 3420
rect 5261 3417 5273 3420
rect 5307 3417 5319 3451
rect 5261 3411 5319 3417
rect 5997 3451 6055 3457
rect 5997 3417 6009 3451
rect 6043 3448 6055 3451
rect 7116 3448 7144 3476
rect 6043 3420 7144 3448
rect 6043 3417 6055 3420
rect 5997 3411 6055 3417
rect 8018 3408 8024 3460
rect 8076 3448 8082 3460
rect 9048 3448 9076 3479
rect 8076 3420 9076 3448
rect 9140 3448 9168 3479
rect 9398 3476 9404 3488
rect 9456 3476 9462 3528
rect 9692 3516 9720 3556
rect 10704 3528 10732 3624
rect 9858 3516 9864 3528
rect 9692 3488 9864 3516
rect 9858 3476 9864 3488
rect 9916 3516 9922 3528
rect 9953 3519 10011 3525
rect 9953 3516 9965 3519
rect 9916 3488 9965 3516
rect 9916 3476 9922 3488
rect 9953 3485 9965 3488
rect 9999 3485 10011 3519
rect 10229 3519 10287 3525
rect 10229 3516 10241 3519
rect 9953 3479 10011 3485
rect 10060 3488 10241 3516
rect 10060 3448 10088 3488
rect 10229 3485 10241 3488
rect 10275 3516 10287 3519
rect 10410 3516 10416 3528
rect 10275 3488 10416 3516
rect 10275 3485 10287 3488
rect 10229 3479 10287 3485
rect 10410 3476 10416 3488
rect 10468 3476 10474 3528
rect 10686 3516 10692 3528
rect 10647 3488 10692 3516
rect 10686 3476 10692 3488
rect 10744 3476 10750 3528
rect 10873 3519 10931 3525
rect 10873 3485 10885 3519
rect 10919 3485 10931 3519
rect 10873 3479 10931 3485
rect 10965 3519 11023 3525
rect 10965 3485 10977 3519
rect 11011 3485 11023 3519
rect 10965 3479 11023 3485
rect 11074 3519 11132 3525
rect 11074 3485 11086 3519
rect 11120 3516 11132 3519
rect 11164 3516 11192 3692
rect 13357 3689 13369 3692
rect 13403 3689 13415 3723
rect 13357 3683 13415 3689
rect 16853 3723 16911 3729
rect 16853 3689 16865 3723
rect 16899 3720 16911 3723
rect 16899 3692 17908 3720
rect 16899 3689 16911 3692
rect 16853 3683 16911 3689
rect 11514 3544 11520 3596
rect 11572 3584 11578 3596
rect 11609 3587 11667 3593
rect 11609 3584 11621 3587
rect 11572 3556 11621 3584
rect 11572 3544 11578 3556
rect 11609 3553 11621 3556
rect 11655 3553 11667 3587
rect 11609 3547 11667 3553
rect 15381 3587 15439 3593
rect 15381 3553 15393 3587
rect 15427 3584 15439 3587
rect 16850 3584 16856 3596
rect 15427 3556 16856 3584
rect 15427 3553 15439 3556
rect 15381 3547 15439 3553
rect 16850 3544 16856 3556
rect 16908 3544 16914 3596
rect 17880 3593 17908 3692
rect 18230 3680 18236 3732
rect 18288 3720 18294 3732
rect 18325 3723 18383 3729
rect 18325 3720 18337 3723
rect 18288 3692 18337 3720
rect 18288 3680 18294 3692
rect 18325 3689 18337 3692
rect 18371 3689 18383 3723
rect 18325 3683 18383 3689
rect 17865 3587 17923 3593
rect 17865 3553 17877 3587
rect 17911 3584 17923 3587
rect 18046 3584 18052 3596
rect 17911 3556 18052 3584
rect 17911 3553 17923 3556
rect 17865 3547 17923 3553
rect 18046 3544 18052 3556
rect 18104 3544 18110 3596
rect 11120 3488 11192 3516
rect 11120 3485 11132 3488
rect 11074 3479 11132 3485
rect 9140 3420 10088 3448
rect 10137 3451 10195 3457
rect 8076 3408 8082 3420
rect 10137 3417 10149 3451
rect 10183 3448 10195 3451
rect 10888 3448 10916 3479
rect 10183 3420 10916 3448
rect 10183 3417 10195 3420
rect 10137 3411 10195 3417
rect 1762 3380 1768 3392
rect 1723 3352 1768 3380
rect 1762 3340 1768 3352
rect 1820 3340 1826 3392
rect 2498 3340 2504 3392
rect 2556 3380 2562 3392
rect 2556 3352 2601 3380
rect 2556 3340 2562 3352
rect 2866 3340 2872 3392
rect 2924 3380 2930 3392
rect 3237 3383 3295 3389
rect 3237 3380 3249 3383
rect 2924 3352 3249 3380
rect 2924 3340 2930 3352
rect 3237 3349 3249 3352
rect 3283 3349 3295 3383
rect 3237 3343 3295 3349
rect 5813 3383 5871 3389
rect 5813 3349 5825 3383
rect 5859 3380 5871 3383
rect 5902 3380 5908 3392
rect 5859 3352 5908 3380
rect 5859 3349 5871 3352
rect 5813 3343 5871 3349
rect 5902 3340 5908 3352
rect 5960 3340 5966 3392
rect 8573 3383 8631 3389
rect 8573 3349 8585 3383
rect 8619 3380 8631 3383
rect 8754 3380 8760 3392
rect 8619 3352 8760 3380
rect 8619 3349 8631 3352
rect 8573 3343 8631 3349
rect 8754 3340 8760 3352
rect 8812 3340 8818 3392
rect 9490 3380 9496 3392
rect 9451 3352 9496 3380
rect 9490 3340 9496 3352
rect 9548 3340 9554 3392
rect 10594 3340 10600 3392
rect 10652 3380 10658 3392
rect 10980 3380 11008 3479
rect 12986 3476 12992 3528
rect 13044 3476 13050 3528
rect 14182 3516 14188 3528
rect 14143 3488 14188 3516
rect 14182 3476 14188 3488
rect 14240 3476 14246 3528
rect 14366 3516 14372 3528
rect 14327 3488 14372 3516
rect 14366 3476 14372 3488
rect 14424 3476 14430 3528
rect 14550 3476 14556 3528
rect 14608 3516 14614 3528
rect 15105 3519 15163 3525
rect 15105 3516 15117 3519
rect 14608 3488 15117 3516
rect 14608 3476 14614 3488
rect 15105 3485 15117 3488
rect 15151 3485 15163 3519
rect 15105 3479 15163 3485
rect 17957 3519 18015 3525
rect 17957 3485 17969 3519
rect 18003 3516 18015 3519
rect 18322 3516 18328 3528
rect 18003 3488 18328 3516
rect 18003 3485 18015 3488
rect 17957 3479 18015 3485
rect 18322 3476 18328 3488
rect 18380 3476 18386 3528
rect 11333 3451 11391 3457
rect 11333 3417 11345 3451
rect 11379 3448 11391 3451
rect 11885 3451 11943 3457
rect 11885 3448 11897 3451
rect 11379 3420 11897 3448
rect 11379 3417 11391 3420
rect 11333 3411 11391 3417
rect 11885 3417 11897 3420
rect 11931 3417 11943 3451
rect 14384 3448 14412 3476
rect 15654 3448 15660 3460
rect 14384 3420 15660 3448
rect 11885 3411 11943 3417
rect 15654 3408 15660 3420
rect 15712 3408 15718 3460
rect 16942 3448 16948 3460
rect 16606 3420 16948 3448
rect 16942 3408 16948 3420
rect 17000 3408 17006 3460
rect 14274 3380 14280 3392
rect 10652 3352 11008 3380
rect 14235 3352 14280 3380
rect 10652 3340 10658 3352
rect 14274 3340 14280 3352
rect 14332 3340 14338 3392
rect 17218 3340 17224 3392
rect 17276 3380 17282 3392
rect 17387 3383 17445 3389
rect 17387 3380 17399 3383
rect 17276 3352 17399 3380
rect 17276 3340 17282 3352
rect 17387 3349 17399 3352
rect 17433 3349 17445 3383
rect 17387 3343 17445 3349
rect 17770 3340 17776 3392
rect 17828 3380 17834 3392
rect 17865 3383 17923 3389
rect 17865 3380 17877 3383
rect 17828 3352 17877 3380
rect 17828 3340 17834 3352
rect 17865 3349 17877 3352
rect 17911 3349 17923 3383
rect 17865 3343 17923 3349
rect 1104 3290 18860 3312
rect 1104 3238 8214 3290
rect 8266 3238 8278 3290
rect 8330 3238 8342 3290
rect 8394 3238 8406 3290
rect 8458 3238 8470 3290
rect 8522 3238 16214 3290
rect 16266 3238 16278 3290
rect 16330 3238 16342 3290
rect 16394 3238 16406 3290
rect 16458 3238 16470 3290
rect 16522 3238 18860 3290
rect 1104 3216 18860 3238
rect 2222 3136 2228 3188
rect 2280 3136 2286 3188
rect 2682 3176 2688 3188
rect 2643 3148 2688 3176
rect 2682 3136 2688 3148
rect 2740 3136 2746 3188
rect 4062 3136 4068 3188
rect 4120 3176 4126 3188
rect 4341 3179 4399 3185
rect 4341 3176 4353 3179
rect 4120 3148 4353 3176
rect 4120 3136 4126 3148
rect 4341 3145 4353 3148
rect 4387 3145 4399 3179
rect 4798 3176 4804 3188
rect 4759 3148 4804 3176
rect 4341 3139 4399 3145
rect 4798 3136 4804 3148
rect 4856 3136 4862 3188
rect 5810 3176 5816 3188
rect 5771 3148 5816 3176
rect 5810 3136 5816 3148
rect 5868 3136 5874 3188
rect 7374 3136 7380 3188
rect 7432 3176 7438 3188
rect 7469 3179 7527 3185
rect 7469 3176 7481 3179
rect 7432 3148 7481 3176
rect 7432 3136 7438 3148
rect 7469 3145 7481 3148
rect 7515 3176 7527 3179
rect 7742 3176 7748 3188
rect 7515 3148 7748 3176
rect 7515 3145 7527 3148
rect 7469 3139 7527 3145
rect 7742 3136 7748 3148
rect 7800 3136 7806 3188
rect 8018 3176 8024 3188
rect 7979 3148 8024 3176
rect 8018 3136 8024 3148
rect 8076 3136 8082 3188
rect 9214 3136 9220 3188
rect 9272 3176 9278 3188
rect 16114 3176 16120 3188
rect 9272 3148 12434 3176
rect 9272 3136 9278 3148
rect 2041 3111 2099 3117
rect 2041 3077 2053 3111
rect 2087 3108 2099 3111
rect 2240 3108 2268 3136
rect 2087 3080 2268 3108
rect 6012 3080 6776 3108
rect 2087 3077 2099 3080
rect 2041 3071 2099 3077
rect 1762 3040 1768 3052
rect 1723 3012 1768 3040
rect 1762 3000 1768 3012
rect 1820 3000 1826 3052
rect 2130 3000 2136 3052
rect 2188 3040 2194 3052
rect 2225 3043 2283 3049
rect 2225 3040 2237 3043
rect 2188 3012 2237 3040
rect 2188 3000 2194 3012
rect 2225 3009 2237 3012
rect 2271 3040 2283 3043
rect 2961 3043 3019 3049
rect 2961 3040 2973 3043
rect 2271 3012 2973 3040
rect 2271 3009 2283 3012
rect 2225 3003 2283 3009
rect 2961 3009 2973 3012
rect 3007 3009 3019 3043
rect 2961 3003 3019 3009
rect 3789 3043 3847 3049
rect 3789 3009 3801 3043
rect 3835 3009 3847 3043
rect 3789 3003 3847 3009
rect 3973 3043 4031 3049
rect 3973 3009 3985 3043
rect 4019 3040 4031 3043
rect 4982 3040 4988 3052
rect 4019 3012 4988 3040
rect 4019 3009 4031 3012
rect 3973 3003 4031 3009
rect 3804 2972 3832 3003
rect 4982 3000 4988 3012
rect 5040 3000 5046 3052
rect 5077 3043 5135 3049
rect 5077 3009 5089 3043
rect 5123 3009 5135 3043
rect 5077 3003 5135 3009
rect 5261 3043 5319 3049
rect 5261 3009 5273 3043
rect 5307 3009 5319 3043
rect 5261 3003 5319 3009
rect 4154 2972 4160 2984
rect 3804 2944 4160 2972
rect 4154 2932 4160 2944
rect 4212 2972 4218 2984
rect 5092 2972 5120 3003
rect 4212 2944 5120 2972
rect 5276 2972 5304 3003
rect 5350 3000 5356 3052
rect 5408 3040 5414 3052
rect 5813 3043 5871 3049
rect 5408 3012 5453 3040
rect 5408 3000 5414 3012
rect 5813 3009 5825 3043
rect 5859 3040 5871 3043
rect 5902 3040 5908 3052
rect 5859 3012 5908 3040
rect 5859 3009 5871 3012
rect 5813 3003 5871 3009
rect 5902 3000 5908 3012
rect 5960 3038 5966 3052
rect 6012 3038 6040 3080
rect 6748 3052 6776 3080
rect 8754 3068 8760 3120
rect 8812 3068 8818 3120
rect 9490 3108 9496 3120
rect 9451 3080 9496 3108
rect 9490 3068 9496 3080
rect 9548 3068 9554 3120
rect 11514 3108 11520 3120
rect 9784 3080 11520 3108
rect 9784 3052 9812 3080
rect 11514 3068 11520 3080
rect 11572 3068 11578 3120
rect 12406 3108 12434 3148
rect 14108 3148 16120 3176
rect 14108 3108 14136 3148
rect 16114 3136 16120 3148
rect 16172 3136 16178 3188
rect 16301 3179 16359 3185
rect 16301 3145 16313 3179
rect 16347 3176 16359 3179
rect 17862 3176 17868 3188
rect 16347 3148 17868 3176
rect 16347 3145 16359 3148
rect 16301 3139 16359 3145
rect 17862 3136 17868 3148
rect 17920 3136 17926 3188
rect 17957 3179 18015 3185
rect 17957 3145 17969 3179
rect 18003 3176 18015 3179
rect 18046 3176 18052 3188
rect 18003 3148 18052 3176
rect 18003 3145 18015 3148
rect 17957 3139 18015 3145
rect 18046 3136 18052 3148
rect 18104 3136 18110 3188
rect 12406 3080 14136 3108
rect 5960 3010 6040 3038
rect 6089 3043 6147 3049
rect 5960 3000 5966 3010
rect 6089 3009 6101 3043
rect 6135 3040 6147 3043
rect 6135 3012 6684 3040
rect 6135 3009 6147 3012
rect 6089 3003 6147 3009
rect 5626 2972 5632 2984
rect 5276 2944 5632 2972
rect 4212 2932 4218 2944
rect 5626 2932 5632 2944
rect 5684 2972 5690 2984
rect 6549 2975 6607 2981
rect 6549 2972 6561 2975
rect 5684 2944 6561 2972
rect 5684 2932 5690 2944
rect 6549 2941 6561 2944
rect 6595 2941 6607 2975
rect 6656 2972 6684 3012
rect 6730 3000 6736 3052
rect 6788 3040 6794 3052
rect 7650 3040 7656 3052
rect 6788 3012 6833 3040
rect 7611 3012 7656 3040
rect 6788 3000 6794 3012
rect 7650 3000 7656 3012
rect 7708 3000 7714 3052
rect 9766 3000 9772 3052
rect 9824 3040 9830 3052
rect 9824 3012 9869 3040
rect 9824 3000 9830 3012
rect 10502 3000 10508 3052
rect 10560 3040 10566 3052
rect 10781 3043 10839 3049
rect 10781 3040 10793 3043
rect 10560 3012 10793 3040
rect 10560 3000 10566 3012
rect 10781 3009 10793 3012
rect 10827 3009 10839 3043
rect 11606 3040 11612 3052
rect 11567 3012 11612 3040
rect 10781 3003 10839 3009
rect 11606 3000 11612 3012
rect 11664 3000 11670 3052
rect 11790 3040 11796 3052
rect 11751 3012 11796 3040
rect 11790 3000 11796 3012
rect 11848 3000 11854 3052
rect 12452 3049 12480 3080
rect 13372 3049 13400 3080
rect 12437 3043 12495 3049
rect 12437 3009 12449 3043
rect 12483 3009 12495 3043
rect 12437 3003 12495 3009
rect 12713 3043 12771 3049
rect 12713 3009 12725 3043
rect 12759 3009 12771 3043
rect 12713 3003 12771 3009
rect 13357 3043 13415 3049
rect 13357 3009 13369 3043
rect 13403 3009 13415 3043
rect 13357 3003 13415 3009
rect 13633 3043 13691 3049
rect 13633 3009 13645 3043
rect 13679 3040 13691 3043
rect 13814 3040 13820 3052
rect 13679 3012 13820 3040
rect 13679 3009 13691 3012
rect 13633 3003 13691 3009
rect 6917 2975 6975 2981
rect 6917 2972 6929 2975
rect 6656 2944 6929 2972
rect 6549 2935 6607 2941
rect 6917 2941 6929 2944
rect 6963 2972 6975 2975
rect 7098 2972 7104 2984
rect 6963 2944 7104 2972
rect 6963 2941 6975 2944
rect 6917 2935 6975 2941
rect 7098 2932 7104 2944
rect 7156 2972 7162 2984
rect 7156 2944 9720 2972
rect 7156 2932 7162 2944
rect 2406 2864 2412 2916
rect 2464 2904 2470 2916
rect 3326 2904 3332 2916
rect 2464 2876 3332 2904
rect 2464 2864 2470 2876
rect 3326 2864 3332 2876
rect 3384 2904 3390 2916
rect 5718 2904 5724 2916
rect 3384 2876 5724 2904
rect 3384 2864 3390 2876
rect 5718 2864 5724 2876
rect 5776 2864 5782 2916
rect 9692 2904 9720 2944
rect 10226 2932 10232 2984
rect 10284 2972 10290 2984
rect 10597 2975 10655 2981
rect 10597 2972 10609 2975
rect 10284 2944 10609 2972
rect 10284 2932 10290 2944
rect 10597 2941 10609 2944
rect 10643 2941 10655 2975
rect 11146 2972 11152 2984
rect 10597 2935 10655 2941
rect 10704 2944 11152 2972
rect 10704 2904 10732 2944
rect 11146 2932 11152 2944
rect 11204 2932 11210 2984
rect 12728 2972 12756 3003
rect 13648 2972 13676 3003
rect 13814 3000 13820 3012
rect 13872 3040 13878 3052
rect 14108 3049 14136 3080
rect 14277 3111 14335 3117
rect 14277 3077 14289 3111
rect 14323 3108 14335 3111
rect 14323 3080 15318 3108
rect 14323 3077 14335 3080
rect 14277 3071 14335 3077
rect 17402 3068 17408 3120
rect 17460 3108 17466 3120
rect 17497 3111 17555 3117
rect 17497 3108 17509 3111
rect 17460 3080 17509 3108
rect 17460 3068 17466 3080
rect 17497 3077 17509 3080
rect 17543 3077 17555 3111
rect 17497 3071 17555 3077
rect 13909 3043 13967 3049
rect 13909 3040 13921 3043
rect 13872 3012 13921 3040
rect 13872 3000 13878 3012
rect 13909 3009 13921 3012
rect 13955 3009 13967 3043
rect 13909 3003 13967 3009
rect 14093 3043 14151 3049
rect 14093 3009 14105 3043
rect 14139 3009 14151 3043
rect 17218 3040 17224 3052
rect 17179 3012 17224 3040
rect 14093 3003 14151 3009
rect 17218 3000 17224 3012
rect 17276 3000 17282 3052
rect 14550 2972 14556 2984
rect 11808 2944 13676 2972
rect 14511 2944 14556 2972
rect 11054 2904 11060 2916
rect 9692 2876 10732 2904
rect 11015 2876 11060 2904
rect 11054 2864 11060 2876
rect 11112 2864 11118 2916
rect 8754 2796 8760 2848
rect 8812 2836 8818 2848
rect 11808 2836 11836 2944
rect 14550 2932 14556 2944
rect 14608 2932 14614 2984
rect 14829 2975 14887 2981
rect 14829 2941 14841 2975
rect 14875 2972 14887 2975
rect 17494 2972 17500 2984
rect 14875 2944 17500 2972
rect 14875 2941 14887 2944
rect 14829 2935 14887 2941
rect 17494 2932 17500 2944
rect 17552 2932 17558 2984
rect 17770 2972 17776 2984
rect 17731 2944 17776 2972
rect 17770 2932 17776 2944
rect 17828 2932 17834 2984
rect 18230 2972 18236 2984
rect 18191 2944 18236 2972
rect 18230 2932 18236 2944
rect 18288 2932 18294 2984
rect 12437 2907 12495 2913
rect 12437 2873 12449 2907
rect 12483 2904 12495 2907
rect 12618 2904 12624 2916
rect 12483 2876 12624 2904
rect 12483 2873 12495 2876
rect 12437 2867 12495 2873
rect 12618 2864 12624 2876
rect 12676 2864 12682 2916
rect 13354 2904 13360 2916
rect 13315 2876 13360 2904
rect 13354 2864 13360 2876
rect 13412 2864 13418 2916
rect 8812 2808 11836 2836
rect 8812 2796 8818 2808
rect 11882 2796 11888 2848
rect 11940 2836 11946 2848
rect 11977 2839 12035 2845
rect 11977 2836 11989 2839
rect 11940 2808 11989 2836
rect 11940 2796 11946 2808
rect 11977 2805 11989 2808
rect 12023 2805 12035 2839
rect 17034 2836 17040 2848
rect 16995 2808 17040 2836
rect 11977 2799 12035 2805
rect 17034 2796 17040 2808
rect 17092 2796 17098 2848
rect 1104 2746 18860 2768
rect 1104 2694 4214 2746
rect 4266 2694 4278 2746
rect 4330 2694 4342 2746
rect 4394 2694 4406 2746
rect 4458 2694 4470 2746
rect 4522 2694 12214 2746
rect 12266 2694 12278 2746
rect 12330 2694 12342 2746
rect 12394 2694 12406 2746
rect 12458 2694 12470 2746
rect 12522 2694 18860 2746
rect 1104 2672 18860 2694
rect 2498 2632 2504 2644
rect 2459 2604 2504 2632
rect 2498 2592 2504 2604
rect 2556 2592 2562 2644
rect 5350 2592 5356 2644
rect 5408 2632 5414 2644
rect 7929 2635 7987 2641
rect 7929 2632 7941 2635
rect 5408 2604 7941 2632
rect 5408 2592 5414 2604
rect 7929 2601 7941 2604
rect 7975 2601 7987 2635
rect 10229 2635 10287 2641
rect 10229 2632 10241 2635
rect 7929 2595 7987 2601
rect 8220 2604 10241 2632
rect 3234 2564 3240 2576
rect 3195 2536 3240 2564
rect 3234 2524 3240 2536
rect 3292 2524 3298 2576
rect 4433 2567 4491 2573
rect 4433 2533 4445 2567
rect 4479 2564 4491 2567
rect 4614 2564 4620 2576
rect 4479 2536 4620 2564
rect 4479 2533 4491 2536
rect 4433 2527 4491 2533
rect 4614 2524 4620 2536
rect 4672 2524 4678 2576
rect 2866 2496 2872 2508
rect 2700 2468 2872 2496
rect 1857 2431 1915 2437
rect 1857 2397 1869 2431
rect 1903 2397 1915 2431
rect 1857 2391 1915 2397
rect 1872 2360 1900 2391
rect 2038 2388 2044 2440
rect 2096 2428 2102 2440
rect 2700 2437 2728 2468
rect 2866 2456 2872 2468
rect 2924 2456 2930 2508
rect 4525 2499 4583 2505
rect 4525 2465 4537 2499
rect 4571 2496 4583 2499
rect 5368 2496 5396 2592
rect 5718 2496 5724 2508
rect 4571 2468 5396 2496
rect 5679 2468 5724 2496
rect 4571 2465 4583 2468
rect 4525 2459 4583 2465
rect 5718 2456 5724 2468
rect 5776 2456 5782 2508
rect 7469 2499 7527 2505
rect 7469 2465 7481 2499
rect 7515 2465 7527 2499
rect 7469 2459 7527 2465
rect 2317 2431 2375 2437
rect 2317 2428 2329 2431
rect 2096 2400 2329 2428
rect 2096 2388 2102 2400
rect 2317 2397 2329 2400
rect 2363 2397 2375 2431
rect 2317 2391 2375 2397
rect 2685 2431 2743 2437
rect 2685 2397 2697 2431
rect 2731 2397 2743 2431
rect 2685 2391 2743 2397
rect 2774 2388 2780 2440
rect 2832 2428 2838 2440
rect 2832 2400 2877 2428
rect 2832 2388 2838 2400
rect 3142 2388 3148 2440
rect 3200 2428 3206 2440
rect 3237 2431 3295 2437
rect 3237 2428 3249 2431
rect 3200 2400 3249 2428
rect 3200 2388 3206 2400
rect 3237 2397 3249 2400
rect 3283 2397 3295 2431
rect 3237 2391 3295 2397
rect 3513 2431 3571 2437
rect 3513 2397 3525 2431
rect 3559 2428 3571 2431
rect 3973 2431 4031 2437
rect 3559 2400 3924 2428
rect 3559 2397 3571 2400
rect 3513 2391 3571 2397
rect 2866 2360 2872 2372
rect 1872 2332 2872 2360
rect 2866 2320 2872 2332
rect 2924 2320 2930 2372
rect 1673 2295 1731 2301
rect 1673 2261 1685 2295
rect 1719 2292 1731 2295
rect 3602 2292 3608 2304
rect 1719 2264 3608 2292
rect 1719 2261 1731 2264
rect 1673 2255 1731 2261
rect 3602 2252 3608 2264
rect 3660 2252 3666 2304
rect 3896 2292 3924 2400
rect 3973 2397 3985 2431
rect 4019 2397 4031 2431
rect 4154 2428 4160 2440
rect 4115 2400 4160 2428
rect 3973 2391 4031 2397
rect 3988 2360 4016 2391
rect 4154 2388 4160 2400
rect 4212 2428 4218 2440
rect 5077 2431 5135 2437
rect 5077 2428 5089 2431
rect 4212 2400 5089 2428
rect 4212 2388 4218 2400
rect 5077 2397 5089 2400
rect 5123 2397 5135 2431
rect 5258 2428 5264 2440
rect 5219 2400 5264 2428
rect 5077 2391 5135 2397
rect 5258 2388 5264 2400
rect 5316 2388 5322 2440
rect 5445 2431 5503 2437
rect 5445 2397 5457 2431
rect 5491 2397 5503 2431
rect 7484 2428 7512 2459
rect 7558 2428 7564 2440
rect 7471 2400 7564 2428
rect 5445 2391 5503 2397
rect 4982 2360 4988 2372
rect 3988 2332 4988 2360
rect 4982 2320 4988 2332
rect 5040 2320 5046 2372
rect 4798 2292 4804 2304
rect 3896 2264 4804 2292
rect 4798 2252 4804 2264
rect 4856 2252 4862 2304
rect 5460 2292 5488 2391
rect 7558 2388 7564 2400
rect 7616 2428 7622 2440
rect 8220 2437 8248 2604
rect 10229 2601 10241 2604
rect 10275 2632 10287 2635
rect 10502 2632 10508 2644
rect 10275 2604 10508 2632
rect 10275 2601 10287 2604
rect 10229 2595 10287 2601
rect 10502 2592 10508 2604
rect 10560 2592 10566 2644
rect 11241 2635 11299 2641
rect 11241 2601 11253 2635
rect 11287 2632 11299 2635
rect 11790 2632 11796 2644
rect 11287 2604 11796 2632
rect 11287 2601 11299 2604
rect 11241 2595 11299 2601
rect 11790 2592 11796 2604
rect 11848 2592 11854 2644
rect 13725 2635 13783 2641
rect 13725 2632 13737 2635
rect 11900 2604 13737 2632
rect 11146 2524 11152 2576
rect 11204 2564 11210 2576
rect 11900 2564 11928 2604
rect 13725 2601 13737 2604
rect 13771 2601 13783 2635
rect 13725 2595 13783 2601
rect 14182 2592 14188 2644
rect 14240 2632 14246 2644
rect 14369 2635 14427 2641
rect 14369 2632 14381 2635
rect 14240 2604 14381 2632
rect 14240 2592 14246 2604
rect 14369 2601 14381 2604
rect 14415 2601 14427 2635
rect 14369 2595 14427 2601
rect 17586 2564 17592 2576
rect 11204 2536 11928 2564
rect 17547 2536 17592 2564
rect 11204 2524 11210 2536
rect 17586 2524 17592 2536
rect 17644 2524 17650 2576
rect 10594 2496 10600 2508
rect 10520 2468 10600 2496
rect 8113 2431 8171 2437
rect 8113 2428 8125 2431
rect 7616 2400 8125 2428
rect 7616 2388 7622 2400
rect 8113 2397 8125 2400
rect 8159 2397 8171 2431
rect 8113 2391 8171 2397
rect 8205 2431 8263 2437
rect 8205 2397 8217 2431
rect 8251 2397 8263 2431
rect 8205 2391 8263 2397
rect 5994 2360 6000 2372
rect 5955 2332 6000 2360
rect 5994 2320 6000 2332
rect 6052 2320 6058 2372
rect 6454 2320 6460 2372
rect 6512 2320 6518 2372
rect 7742 2320 7748 2372
rect 7800 2360 7806 2372
rect 8220 2360 8248 2391
rect 8662 2388 8668 2440
rect 8720 2428 8726 2440
rect 9125 2431 9183 2437
rect 9125 2428 9137 2431
rect 8720 2400 9137 2428
rect 8720 2388 8726 2400
rect 9125 2397 9137 2400
rect 9171 2397 9183 2431
rect 9125 2391 9183 2397
rect 9214 2388 9220 2440
rect 9272 2428 9278 2440
rect 10520 2437 10548 2468
rect 10594 2456 10600 2468
rect 10652 2496 10658 2508
rect 10781 2499 10839 2505
rect 10781 2496 10793 2499
rect 10652 2468 10793 2496
rect 10652 2456 10658 2468
rect 10781 2465 10793 2468
rect 10827 2465 10839 2499
rect 10781 2459 10839 2465
rect 11606 2456 11612 2508
rect 11664 2496 11670 2508
rect 11977 2499 12035 2505
rect 11977 2496 11989 2499
rect 11664 2468 11989 2496
rect 11664 2456 11670 2468
rect 11977 2465 11989 2468
rect 12023 2465 12035 2499
rect 11977 2459 12035 2465
rect 14550 2456 14556 2508
rect 14608 2496 14614 2508
rect 15105 2499 15163 2505
rect 15105 2496 15117 2499
rect 14608 2468 15117 2496
rect 14608 2456 14614 2468
rect 15105 2465 15117 2468
rect 15151 2465 15163 2499
rect 15105 2459 15163 2465
rect 15381 2499 15439 2505
rect 15381 2465 15393 2499
rect 15427 2496 15439 2499
rect 17034 2496 17040 2508
rect 15427 2468 17040 2496
rect 15427 2465 15439 2468
rect 15381 2459 15439 2465
rect 17034 2456 17040 2468
rect 17092 2456 17098 2508
rect 17954 2456 17960 2508
rect 18012 2456 18018 2508
rect 9309 2431 9367 2437
rect 9309 2428 9321 2431
rect 9272 2400 9321 2428
rect 9272 2388 9278 2400
rect 9309 2397 9321 2400
rect 9355 2397 9367 2431
rect 9309 2391 9367 2397
rect 10505 2431 10563 2437
rect 10505 2397 10517 2431
rect 10551 2397 10563 2431
rect 10505 2391 10563 2397
rect 10965 2431 11023 2437
rect 10965 2397 10977 2431
rect 11011 2428 11023 2431
rect 11054 2428 11060 2440
rect 11011 2400 11060 2428
rect 11011 2397 11023 2400
rect 10965 2391 11023 2397
rect 11054 2388 11060 2400
rect 11112 2388 11118 2440
rect 13354 2388 13360 2440
rect 13412 2388 13418 2440
rect 13906 2388 13912 2440
rect 13964 2428 13970 2440
rect 14185 2431 14243 2437
rect 14185 2428 14197 2431
rect 13964 2400 14197 2428
rect 13964 2388 13970 2400
rect 14185 2397 14197 2400
rect 14231 2397 14243 2431
rect 17972 2428 18000 2456
rect 16514 2400 18000 2428
rect 14185 2391 14243 2397
rect 7800 2332 8248 2360
rect 10045 2363 10103 2369
rect 7800 2320 7806 2332
rect 10045 2329 10057 2363
rect 10091 2360 10103 2363
rect 11146 2360 11152 2372
rect 10091 2332 11152 2360
rect 10091 2329 10103 2332
rect 10045 2323 10103 2329
rect 11146 2320 11152 2332
rect 11204 2320 11210 2372
rect 11333 2363 11391 2369
rect 11333 2329 11345 2363
rect 11379 2329 11391 2363
rect 11333 2323 11391 2329
rect 8570 2292 8576 2304
rect 5460 2264 8576 2292
rect 8570 2252 8576 2264
rect 8628 2252 8634 2304
rect 9214 2292 9220 2304
rect 9175 2264 9220 2292
rect 9214 2252 9220 2264
rect 9272 2252 9278 2304
rect 10226 2292 10232 2304
rect 10187 2264 10232 2292
rect 10226 2252 10232 2264
rect 10284 2252 10290 2304
rect 11054 2252 11060 2304
rect 11112 2292 11118 2304
rect 11348 2292 11376 2323
rect 11974 2320 11980 2372
rect 12032 2360 12038 2372
rect 12253 2363 12311 2369
rect 12253 2360 12265 2363
rect 12032 2332 12265 2360
rect 12032 2320 12038 2332
rect 12253 2329 12265 2332
rect 12299 2329 12311 2363
rect 12253 2323 12311 2329
rect 17865 2363 17923 2369
rect 17865 2329 17877 2363
rect 17911 2329 17923 2363
rect 17865 2323 17923 2329
rect 11112 2264 11376 2292
rect 14829 2295 14887 2301
rect 11112 2252 11118 2264
rect 14829 2261 14841 2295
rect 14875 2292 14887 2295
rect 14918 2292 14924 2304
rect 14875 2264 14924 2292
rect 14875 2261 14887 2264
rect 14829 2255 14887 2261
rect 14918 2252 14924 2264
rect 14976 2252 14982 2304
rect 16853 2295 16911 2301
rect 16853 2261 16865 2295
rect 16899 2292 16911 2295
rect 17770 2292 17776 2304
rect 16899 2264 17776 2292
rect 16899 2261 16911 2264
rect 16853 2255 16911 2261
rect 17770 2252 17776 2264
rect 17828 2292 17834 2304
rect 17880 2292 17908 2323
rect 17954 2320 17960 2372
rect 18012 2360 18018 2372
rect 18049 2363 18107 2369
rect 18049 2360 18061 2363
rect 18012 2332 18061 2360
rect 18012 2320 18018 2332
rect 18049 2329 18061 2332
rect 18095 2329 18107 2363
rect 18049 2323 18107 2329
rect 18141 2363 18199 2369
rect 18141 2329 18153 2363
rect 18187 2360 18199 2363
rect 18322 2360 18328 2372
rect 18187 2332 18328 2360
rect 18187 2329 18199 2332
rect 18141 2323 18199 2329
rect 18322 2320 18328 2332
rect 18380 2320 18386 2372
rect 17828 2264 17908 2292
rect 17828 2252 17834 2264
rect 1104 2202 18860 2224
rect 1104 2150 8214 2202
rect 8266 2150 8278 2202
rect 8330 2150 8342 2202
rect 8394 2150 8406 2202
rect 8458 2150 8470 2202
rect 8522 2150 16214 2202
rect 16266 2150 16278 2202
rect 16330 2150 16342 2202
rect 16394 2150 16406 2202
rect 16458 2150 16470 2202
rect 16522 2150 18860 2202
rect 1104 2128 18860 2150
rect 3142 2088 3148 2100
rect 2240 2060 3148 2088
rect 1673 2023 1731 2029
rect 1673 1989 1685 2023
rect 1719 2020 1731 2023
rect 2038 2020 2044 2032
rect 1719 1992 2044 2020
rect 1719 1989 1731 1992
rect 1673 1983 1731 1989
rect 2038 1980 2044 1992
rect 2096 1980 2102 2032
rect 1857 1955 1915 1961
rect 1857 1921 1869 1955
rect 1903 1921 1915 1955
rect 1857 1915 1915 1921
rect 1949 1955 2007 1961
rect 1949 1921 1961 1955
rect 1995 1952 2007 1955
rect 2240 1952 2268 2060
rect 3142 2048 3148 2060
rect 3200 2088 3206 2100
rect 4614 2088 4620 2100
rect 3200 2060 4620 2088
rect 3200 2048 3206 2060
rect 4614 2048 4620 2060
rect 4672 2088 4678 2100
rect 5077 2091 5135 2097
rect 5077 2088 5089 2091
rect 4672 2060 5089 2088
rect 4672 2048 4678 2060
rect 5077 2057 5089 2060
rect 5123 2088 5135 2091
rect 5258 2088 5264 2100
rect 5123 2060 5264 2088
rect 5123 2057 5135 2060
rect 5077 2051 5135 2057
rect 5258 2048 5264 2060
rect 5316 2048 5322 2100
rect 5997 2091 6055 2097
rect 5997 2057 6009 2091
rect 6043 2088 6055 2091
rect 6454 2088 6460 2100
rect 6043 2060 6460 2088
rect 6043 2057 6055 2060
rect 5997 2051 6055 2057
rect 6454 2048 6460 2060
rect 6512 2048 6518 2100
rect 6549 2091 6607 2097
rect 6549 2057 6561 2091
rect 6595 2088 6607 2091
rect 6638 2088 6644 2100
rect 6595 2060 6644 2088
rect 6595 2057 6607 2060
rect 6549 2051 6607 2057
rect 6638 2048 6644 2060
rect 6696 2048 6702 2100
rect 8389 2091 8447 2097
rect 8389 2057 8401 2091
rect 8435 2088 8447 2091
rect 8570 2088 8576 2100
rect 8435 2060 8576 2088
rect 8435 2057 8447 2060
rect 8389 2051 8447 2057
rect 8570 2048 8576 2060
rect 8628 2048 8634 2100
rect 14550 2088 14556 2100
rect 11624 2060 14556 2088
rect 11624 2032 11652 2060
rect 2409 2023 2467 2029
rect 2409 1989 2421 2023
rect 2455 2020 2467 2023
rect 2590 2020 2596 2032
rect 2455 1992 2596 2020
rect 2455 1989 2467 1992
rect 2409 1983 2467 1989
rect 2590 1980 2596 1992
rect 2648 1980 2654 2032
rect 3234 2020 3240 2032
rect 2700 1992 3240 2020
rect 2700 1961 2728 1992
rect 3234 1980 3240 1992
rect 3292 1980 3298 2032
rect 3602 2020 3608 2032
rect 3563 1992 3608 2020
rect 3602 1980 3608 1992
rect 3660 1980 3666 2032
rect 5166 2020 5172 2032
rect 4830 1992 5172 2020
rect 5166 1980 5172 1992
rect 5224 1980 5230 2032
rect 7374 2020 7380 2032
rect 6012 1992 7380 2020
rect 1995 1924 2268 1952
rect 2317 1955 2375 1961
rect 1995 1921 2007 1924
rect 1949 1915 2007 1921
rect 2317 1921 2329 1955
rect 2363 1921 2375 1955
rect 2317 1915 2375 1921
rect 2685 1955 2743 1961
rect 2685 1921 2697 1955
rect 2731 1921 2743 1955
rect 3326 1952 3332 1964
rect 3287 1924 3332 1952
rect 2685 1915 2743 1921
rect 1872 1884 1900 1915
rect 2332 1884 2360 1915
rect 3326 1912 3332 1924
rect 3384 1912 3390 1964
rect 5813 1955 5871 1961
rect 5813 1921 5825 1955
rect 5859 1952 5871 1955
rect 5902 1952 5908 1964
rect 5859 1924 5908 1952
rect 5859 1921 5871 1924
rect 5813 1915 5871 1921
rect 5902 1912 5908 1924
rect 5960 1912 5966 1964
rect 6012 1961 6040 1992
rect 7374 1980 7380 1992
rect 7432 1980 7438 2032
rect 9214 1980 9220 2032
rect 9272 1980 9278 2032
rect 11606 2020 11612 2032
rect 10152 1992 11612 2020
rect 5997 1955 6055 1961
rect 5997 1921 6009 1955
rect 6043 1921 6055 1955
rect 5997 1915 6055 1921
rect 6457 1955 6515 1961
rect 6457 1921 6469 1955
rect 6503 1952 6515 1955
rect 6730 1952 6736 1964
rect 6503 1924 6736 1952
rect 6503 1921 6515 1924
rect 6457 1915 6515 1921
rect 2774 1884 2780 1896
rect 1872 1856 1992 1884
rect 2332 1856 2780 1884
rect 1964 1748 1992 1856
rect 2774 1844 2780 1856
rect 2832 1844 2838 1896
rect 2869 1887 2927 1893
rect 2869 1853 2881 1887
rect 2915 1884 2927 1887
rect 4154 1884 4160 1896
rect 2915 1856 4160 1884
rect 2915 1853 2927 1856
rect 2869 1847 2927 1853
rect 4154 1844 4160 1856
rect 4212 1844 4218 1896
rect 5350 1844 5356 1896
rect 5408 1884 5414 1896
rect 6012 1884 6040 1915
rect 6730 1912 6736 1924
rect 6788 1912 6794 1964
rect 7558 1912 7564 1964
rect 7616 1912 7622 1964
rect 10152 1961 10180 1992
rect 11606 1980 11612 1992
rect 11664 1980 11670 2032
rect 12618 1980 12624 2032
rect 12676 1980 12682 2032
rect 10137 1955 10195 1961
rect 10137 1921 10149 1955
rect 10183 1921 10195 1955
rect 10137 1915 10195 1921
rect 10505 1955 10563 1961
rect 10505 1921 10517 1955
rect 10551 1952 10563 1955
rect 10686 1952 10692 1964
rect 10551 1924 10692 1952
rect 10551 1921 10563 1924
rect 10505 1915 10563 1921
rect 6917 1887 6975 1893
rect 6917 1884 6929 1887
rect 5408 1856 6040 1884
rect 6104 1856 6929 1884
rect 5408 1844 5414 1856
rect 4982 1776 4988 1828
rect 5040 1816 5046 1828
rect 6104 1816 6132 1856
rect 6917 1853 6929 1856
rect 6963 1853 6975 1887
rect 7742 1884 7748 1896
rect 7703 1856 7748 1884
rect 6917 1847 6975 1853
rect 7742 1844 7748 1856
rect 7800 1844 7806 1896
rect 9398 1844 9404 1896
rect 9456 1884 9462 1896
rect 9861 1887 9919 1893
rect 9861 1884 9873 1887
rect 9456 1856 9873 1884
rect 9456 1844 9462 1856
rect 9861 1853 9873 1856
rect 9907 1853 9919 1887
rect 9861 1847 9919 1853
rect 10520 1816 10548 1915
rect 10686 1912 10692 1924
rect 10744 1912 10750 1964
rect 11054 1952 11060 1964
rect 11015 1924 11060 1952
rect 11054 1912 11060 1924
rect 11112 1912 11118 1964
rect 13464 1961 13492 2060
rect 14550 2048 14556 2060
rect 14608 2088 14614 2100
rect 18141 2091 18199 2097
rect 14608 2060 15608 2088
rect 14608 2048 14614 2060
rect 14274 1980 14280 2032
rect 14332 1980 14338 2032
rect 15580 1961 15608 2060
rect 18141 2057 18153 2091
rect 18187 2088 18199 2091
rect 18230 2088 18236 2100
rect 18187 2060 18236 2088
rect 18187 2057 18199 2060
rect 18141 2051 18199 2057
rect 18230 2048 18236 2060
rect 18288 2048 18294 2100
rect 16942 2020 16948 2032
rect 15948 1992 16948 2020
rect 13449 1955 13507 1961
rect 13449 1921 13461 1955
rect 13495 1921 13507 1955
rect 13449 1915 13507 1921
rect 15565 1955 15623 1961
rect 15565 1921 15577 1955
rect 15611 1921 15623 1955
rect 15565 1915 15623 1921
rect 15654 1912 15660 1964
rect 15712 1952 15718 1964
rect 15948 1961 15976 1992
rect 16942 1980 16948 1992
rect 17000 1980 17006 2032
rect 15933 1955 15991 1961
rect 15933 1952 15945 1955
rect 15712 1924 15945 1952
rect 15712 1912 15718 1924
rect 15933 1921 15945 1924
rect 15979 1921 15991 1955
rect 16114 1952 16120 1964
rect 16075 1924 16120 1952
rect 15933 1915 15991 1921
rect 16114 1912 16120 1924
rect 16172 1912 16178 1964
rect 16758 1912 16764 1964
rect 16816 1952 16822 1964
rect 17129 1955 17187 1961
rect 17129 1952 17141 1955
rect 16816 1924 17141 1952
rect 16816 1912 16822 1924
rect 17129 1921 17141 1924
rect 17175 1921 17187 1955
rect 17129 1915 17187 1921
rect 17313 1955 17371 1961
rect 17313 1921 17325 1955
rect 17359 1921 17371 1955
rect 17313 1915 17371 1921
rect 11146 1884 11152 1896
rect 11107 1856 11152 1884
rect 11146 1844 11152 1856
rect 11204 1844 11210 1896
rect 13173 1887 13231 1893
rect 13173 1884 13185 1887
rect 11992 1856 13185 1884
rect 5040 1788 6132 1816
rect 10428 1788 10548 1816
rect 10781 1819 10839 1825
rect 5040 1776 5046 1788
rect 4798 1748 4804 1760
rect 1964 1720 4804 1748
rect 4798 1708 4804 1720
rect 4856 1708 4862 1760
rect 9214 1708 9220 1760
rect 9272 1748 9278 1760
rect 10428 1748 10456 1788
rect 10781 1785 10793 1819
rect 10827 1816 10839 1819
rect 11992 1816 12020 1856
rect 13173 1853 13185 1856
rect 13219 1853 13231 1887
rect 13173 1847 13231 1853
rect 14918 1844 14924 1896
rect 14976 1884 14982 1896
rect 15289 1887 15347 1893
rect 15289 1884 15301 1887
rect 14976 1856 15301 1884
rect 14976 1844 14982 1856
rect 15289 1853 15301 1856
rect 15335 1853 15347 1887
rect 15289 1847 15347 1853
rect 16574 1844 16580 1896
rect 16632 1884 16638 1896
rect 17328 1884 17356 1915
rect 16632 1856 17356 1884
rect 16632 1844 16638 1856
rect 15930 1816 15936 1828
rect 10827 1788 12020 1816
rect 15891 1788 15936 1816
rect 10827 1785 10839 1788
rect 10781 1779 10839 1785
rect 15930 1776 15936 1788
rect 15988 1776 15994 1828
rect 9272 1720 10456 1748
rect 9272 1708 9278 1720
rect 10502 1708 10508 1760
rect 10560 1748 10566 1760
rect 11701 1751 11759 1757
rect 11701 1748 11713 1751
rect 10560 1720 11713 1748
rect 10560 1708 10566 1720
rect 11701 1717 11713 1720
rect 11747 1717 11759 1751
rect 11701 1711 11759 1717
rect 13817 1751 13875 1757
rect 13817 1717 13829 1751
rect 13863 1748 13875 1751
rect 14826 1748 14832 1760
rect 13863 1720 14832 1748
rect 13863 1717 13875 1720
rect 13817 1711 13875 1717
rect 14826 1708 14832 1720
rect 14884 1708 14890 1760
rect 1104 1658 18860 1680
rect 1104 1606 4214 1658
rect 4266 1606 4278 1658
rect 4330 1606 4342 1658
rect 4394 1606 4406 1658
rect 4458 1606 4470 1658
rect 4522 1606 12214 1658
rect 12266 1606 12278 1658
rect 12330 1606 12342 1658
rect 12394 1606 12406 1658
rect 12458 1606 12470 1658
rect 12522 1606 18860 1658
rect 1104 1584 18860 1606
rect 2866 1504 2872 1556
rect 2924 1544 2930 1556
rect 3973 1547 4031 1553
rect 3973 1544 3985 1547
rect 2924 1516 3985 1544
rect 2924 1504 2930 1516
rect 3973 1513 3985 1516
rect 4019 1513 4031 1547
rect 3973 1507 4031 1513
rect 5905 1547 5963 1553
rect 5905 1513 5917 1547
rect 5951 1544 5963 1547
rect 5994 1544 6000 1556
rect 5951 1516 6000 1544
rect 5951 1513 5963 1516
rect 5905 1507 5963 1513
rect 5994 1504 6000 1516
rect 6052 1504 6058 1556
rect 11974 1504 11980 1556
rect 12032 1544 12038 1556
rect 12161 1547 12219 1553
rect 12161 1544 12173 1547
rect 12032 1516 12173 1544
rect 12032 1504 12038 1516
rect 12161 1513 12173 1516
rect 12207 1513 12219 1547
rect 12161 1507 12219 1513
rect 1486 1408 1492 1420
rect 1447 1380 1492 1408
rect 1486 1368 1492 1380
rect 1544 1368 1550 1420
rect 4433 1411 4491 1417
rect 4433 1377 4445 1411
rect 4479 1408 4491 1411
rect 4798 1408 4804 1420
rect 4479 1380 4804 1408
rect 4479 1377 4491 1380
rect 4433 1371 4491 1377
rect 4798 1368 4804 1380
rect 4856 1408 4862 1420
rect 7469 1411 7527 1417
rect 4856 1380 4936 1408
rect 4856 1368 4862 1380
rect 3237 1343 3295 1349
rect 3237 1309 3249 1343
rect 3283 1340 3295 1343
rect 3326 1340 3332 1352
rect 3283 1312 3332 1340
rect 3283 1309 3295 1312
rect 3237 1303 3295 1309
rect 3326 1300 3332 1312
rect 3384 1300 3390 1352
rect 4522 1272 4528 1284
rect 4483 1244 4528 1272
rect 4522 1232 4528 1244
rect 4580 1232 4586 1284
rect 4908 1272 4936 1380
rect 7469 1377 7481 1411
rect 7515 1408 7527 1411
rect 7742 1408 7748 1420
rect 7515 1380 7748 1408
rect 7515 1377 7527 1380
rect 7469 1371 7527 1377
rect 7742 1368 7748 1380
rect 7800 1368 7806 1420
rect 9398 1408 9404 1420
rect 9359 1380 9404 1408
rect 9398 1368 9404 1380
rect 9456 1368 9462 1420
rect 10226 1408 10232 1420
rect 9508 1380 10232 1408
rect 5166 1340 5172 1352
rect 5127 1312 5172 1340
rect 5166 1300 5172 1312
rect 5224 1300 5230 1352
rect 5350 1340 5356 1352
rect 5311 1312 5356 1340
rect 5350 1300 5356 1312
rect 5408 1300 5414 1352
rect 5537 1343 5595 1349
rect 5537 1309 5549 1343
rect 5583 1340 5595 1343
rect 5902 1340 5908 1352
rect 5583 1312 5908 1340
rect 5583 1309 5595 1312
rect 5537 1303 5595 1309
rect 5902 1300 5908 1312
rect 5960 1300 5966 1352
rect 6089 1343 6147 1349
rect 6089 1309 6101 1343
rect 6135 1340 6147 1343
rect 6991 1343 7049 1349
rect 6991 1340 7003 1343
rect 6135 1312 7003 1340
rect 6135 1309 6147 1312
rect 6089 1303 6147 1309
rect 6991 1309 7003 1312
rect 7037 1309 7049 1343
rect 6991 1303 7049 1309
rect 8389 1343 8447 1349
rect 8389 1309 8401 1343
rect 8435 1340 8447 1343
rect 8570 1340 8576 1352
rect 8435 1312 8576 1340
rect 8435 1309 8447 1312
rect 8389 1303 8447 1309
rect 8570 1300 8576 1312
rect 8628 1300 8634 1352
rect 9033 1343 9091 1349
rect 9033 1309 9045 1343
rect 9079 1309 9091 1343
rect 9214 1340 9220 1352
rect 9175 1312 9220 1340
rect 9033 1303 9091 1309
rect 7466 1272 7472 1284
rect 4908 1244 6914 1272
rect 7427 1244 7472 1272
rect 4433 1207 4491 1213
rect 4433 1173 4445 1207
rect 4479 1204 4491 1207
rect 4614 1204 4620 1216
rect 4479 1176 4620 1204
rect 4479 1173 4491 1176
rect 4433 1167 4491 1173
rect 4614 1164 4620 1176
rect 4672 1164 4678 1216
rect 6454 1204 6460 1216
rect 6415 1176 6460 1204
rect 6454 1164 6460 1176
rect 6512 1164 6518 1216
rect 6886 1204 6914 1244
rect 7466 1232 7472 1244
rect 7524 1232 7530 1284
rect 7558 1232 7564 1284
rect 7616 1272 7622 1284
rect 9048 1272 9076 1303
rect 9214 1300 9220 1312
rect 9272 1300 9278 1352
rect 9508 1340 9536 1380
rect 10226 1368 10232 1380
rect 10284 1408 10290 1420
rect 10321 1411 10379 1417
rect 10321 1408 10333 1411
rect 10284 1380 10333 1408
rect 10284 1368 10290 1380
rect 10321 1377 10333 1380
rect 10367 1377 10379 1411
rect 11146 1408 11152 1420
rect 11107 1380 11152 1408
rect 10321 1371 10379 1377
rect 11146 1368 11152 1380
rect 11204 1368 11210 1420
rect 14550 1408 14556 1420
rect 14511 1380 14556 1408
rect 14550 1368 14556 1380
rect 14608 1368 14614 1420
rect 14826 1408 14832 1420
rect 14787 1380 14832 1408
rect 14826 1368 14832 1380
rect 14884 1368 14890 1420
rect 16114 1368 16120 1420
rect 16172 1408 16178 1420
rect 16172 1380 16574 1408
rect 16172 1368 16178 1380
rect 9324 1312 9536 1340
rect 9585 1343 9643 1349
rect 9324 1272 9352 1312
rect 9585 1309 9597 1343
rect 9631 1340 9643 1343
rect 9674 1340 9680 1352
rect 9631 1312 9680 1340
rect 9631 1309 9643 1312
rect 9585 1303 9643 1309
rect 9674 1300 9680 1312
rect 9732 1300 9738 1352
rect 10502 1340 10508 1352
rect 10463 1312 10508 1340
rect 10502 1300 10508 1312
rect 10560 1300 10566 1352
rect 11882 1300 11888 1352
rect 11940 1340 11946 1352
rect 11977 1343 12035 1349
rect 11977 1340 11989 1343
rect 11940 1312 11989 1340
rect 11940 1300 11946 1312
rect 11977 1309 11989 1312
rect 12023 1309 12035 1343
rect 11977 1303 12035 1309
rect 15930 1300 15936 1352
rect 15988 1300 15994 1352
rect 16546 1340 16574 1380
rect 16761 1343 16819 1349
rect 16761 1340 16773 1343
rect 16546 1312 16773 1340
rect 16761 1309 16773 1312
rect 16807 1309 16819 1343
rect 16942 1340 16948 1352
rect 16903 1312 16948 1340
rect 16761 1303 16819 1309
rect 16942 1300 16948 1312
rect 17000 1300 17006 1352
rect 17586 1340 17592 1352
rect 17547 1312 17592 1340
rect 17586 1300 17592 1312
rect 17644 1300 17650 1352
rect 18141 1343 18199 1349
rect 18141 1309 18153 1343
rect 18187 1340 18199 1343
rect 18230 1340 18236 1352
rect 18187 1312 18236 1340
rect 18187 1309 18199 1312
rect 18141 1303 18199 1309
rect 18230 1300 18236 1312
rect 18288 1300 18294 1352
rect 7616 1244 7661 1272
rect 8588 1244 9352 1272
rect 9692 1272 9720 1300
rect 11054 1272 11060 1284
rect 9692 1244 11060 1272
rect 7616 1232 7622 1244
rect 8588 1213 8616 1244
rect 11054 1232 11060 1244
rect 11112 1232 11118 1284
rect 8573 1207 8631 1213
rect 8573 1204 8585 1207
rect 6886 1176 8585 1204
rect 8573 1173 8585 1176
rect 8619 1173 8631 1207
rect 8573 1167 8631 1173
rect 16301 1207 16359 1213
rect 16301 1173 16313 1207
rect 16347 1204 16359 1207
rect 16574 1204 16580 1216
rect 16347 1176 16580 1204
rect 16347 1173 16359 1176
rect 16301 1167 16359 1173
rect 16574 1164 16580 1176
rect 16632 1164 16638 1216
rect 16666 1164 16672 1216
rect 16724 1204 16730 1216
rect 16853 1207 16911 1213
rect 16853 1204 16865 1207
rect 16724 1176 16865 1204
rect 16724 1164 16730 1176
rect 16853 1173 16865 1176
rect 16899 1173 16911 1207
rect 16853 1167 16911 1173
rect 17494 1164 17500 1216
rect 17552 1204 17558 1216
rect 17773 1207 17831 1213
rect 17773 1204 17785 1207
rect 17552 1176 17785 1204
rect 17552 1164 17558 1176
rect 17773 1173 17785 1176
rect 17819 1173 17831 1207
rect 18322 1204 18328 1216
rect 18283 1176 18328 1204
rect 17773 1167 17831 1173
rect 18322 1164 18328 1176
rect 18380 1164 18386 1216
rect 1104 1114 18860 1136
rect 1104 1062 8214 1114
rect 8266 1062 8278 1114
rect 8330 1062 8342 1114
rect 8394 1062 8406 1114
rect 8458 1062 8470 1114
rect 8522 1062 16214 1114
rect 16266 1062 16278 1114
rect 16330 1062 16342 1114
rect 16394 1062 16406 1114
rect 16458 1062 16470 1114
rect 16522 1062 18860 1114
rect 1104 1040 18860 1062
rect 2774 960 2780 1012
rect 2832 1000 2838 1012
rect 6454 1000 6460 1012
rect 2832 972 6460 1000
rect 2832 960 2838 972
rect 6454 960 6460 972
rect 6512 960 6518 1012
rect 4522 892 4528 944
rect 4580 932 4586 944
rect 5442 932 5448 944
rect 4580 904 5448 932
rect 4580 892 4586 904
rect 5442 892 5448 904
rect 5500 932 5506 944
rect 7558 932 7564 944
rect 5500 904 7564 932
rect 5500 892 5506 904
rect 7558 892 7564 904
rect 7616 932 7622 944
rect 18322 932 18328 944
rect 7616 904 18328 932
rect 7616 892 7622 904
rect 18322 892 18328 904
rect 18380 892 18386 944
<< via1 >>
rect 12716 13676 12768 13728
rect 17316 13676 17368 13728
rect 4214 13574 4266 13626
rect 4278 13574 4330 13626
rect 4342 13574 4394 13626
rect 4406 13574 4458 13626
rect 4470 13574 4522 13626
rect 12214 13574 12266 13626
rect 12278 13574 12330 13626
rect 12342 13574 12394 13626
rect 12406 13574 12458 13626
rect 12470 13574 12522 13626
rect 1308 13472 1360 13524
rect 7104 13472 7156 13524
rect 8484 13472 8536 13524
rect 5540 13404 5592 13456
rect 13820 13404 13872 13456
rect 2964 13268 3016 13320
rect 4436 13268 4488 13320
rect 4528 13268 4580 13320
rect 6552 13336 6604 13388
rect 7012 13268 7064 13320
rect 8944 13336 8996 13388
rect 9312 13268 9364 13320
rect 10140 13311 10192 13320
rect 10140 13277 10149 13311
rect 10149 13277 10183 13311
rect 10183 13277 10192 13311
rect 10140 13268 10192 13277
rect 11612 13268 11664 13320
rect 12624 13268 12676 13320
rect 13084 13268 13136 13320
rect 14188 13311 14240 13320
rect 14188 13277 14197 13311
rect 14197 13277 14231 13311
rect 14231 13277 14240 13311
rect 14188 13268 14240 13277
rect 4344 13243 4396 13252
rect 4344 13209 4353 13243
rect 4353 13209 4387 13243
rect 4387 13209 4396 13243
rect 4344 13200 4396 13209
rect 6000 13200 6052 13252
rect 2228 13175 2280 13184
rect 2228 13141 2237 13175
rect 2237 13141 2271 13175
rect 2271 13141 2280 13175
rect 2228 13132 2280 13141
rect 2320 13175 2372 13184
rect 2320 13141 2329 13175
rect 2329 13141 2363 13175
rect 2363 13141 2372 13175
rect 2688 13175 2740 13184
rect 2320 13132 2372 13141
rect 2688 13141 2697 13175
rect 2697 13141 2731 13175
rect 2731 13141 2740 13175
rect 2688 13132 2740 13141
rect 5172 13175 5224 13184
rect 5172 13141 5181 13175
rect 5181 13141 5215 13175
rect 5215 13141 5224 13175
rect 5172 13132 5224 13141
rect 5632 13175 5684 13184
rect 5632 13141 5641 13175
rect 5641 13141 5675 13175
rect 5675 13141 5684 13175
rect 5632 13132 5684 13141
rect 6092 13175 6144 13184
rect 6092 13141 6101 13175
rect 6101 13141 6135 13175
rect 6135 13141 6144 13175
rect 6092 13132 6144 13141
rect 6184 13132 6236 13184
rect 7288 13200 7340 13252
rect 7564 13200 7616 13252
rect 9588 13243 9640 13252
rect 9588 13209 9597 13243
rect 9597 13209 9631 13243
rect 9631 13209 9640 13243
rect 9588 13200 9640 13209
rect 8576 13175 8628 13184
rect 8576 13141 8585 13175
rect 8585 13141 8619 13175
rect 8619 13141 8628 13175
rect 8576 13132 8628 13141
rect 9772 13200 9824 13252
rect 11336 13200 11388 13252
rect 12256 13243 12308 13252
rect 10600 13175 10652 13184
rect 10600 13141 10609 13175
rect 10609 13141 10643 13175
rect 10643 13141 10652 13175
rect 10600 13132 10652 13141
rect 10784 13132 10836 13184
rect 11060 13132 11112 13184
rect 12256 13209 12265 13243
rect 12265 13209 12299 13243
rect 12299 13209 12308 13243
rect 12256 13200 12308 13209
rect 12716 13243 12768 13252
rect 12716 13209 12725 13243
rect 12725 13209 12759 13243
rect 12759 13209 12768 13243
rect 12716 13200 12768 13209
rect 14648 13243 14700 13252
rect 13728 13132 13780 13184
rect 14648 13209 14657 13243
rect 14657 13209 14691 13243
rect 14691 13209 14700 13243
rect 14648 13200 14700 13209
rect 15384 13268 15436 13320
rect 17224 13336 17276 13388
rect 16764 13311 16816 13320
rect 16764 13277 16773 13311
rect 16773 13277 16807 13311
rect 16807 13277 16816 13311
rect 16764 13268 16816 13277
rect 16028 13200 16080 13252
rect 15752 13175 15804 13184
rect 15752 13141 15761 13175
rect 15761 13141 15795 13175
rect 15795 13141 15804 13175
rect 15752 13132 15804 13141
rect 17776 13175 17828 13184
rect 17776 13141 17785 13175
rect 17785 13141 17819 13175
rect 17819 13141 17828 13175
rect 17776 13132 17828 13141
rect 8214 13030 8266 13082
rect 8278 13030 8330 13082
rect 8342 13030 8394 13082
rect 8406 13030 8458 13082
rect 8470 13030 8522 13082
rect 16214 13030 16266 13082
rect 16278 13030 16330 13082
rect 16342 13030 16394 13082
rect 16406 13030 16458 13082
rect 16470 13030 16522 13082
rect 6092 12928 6144 12980
rect 6920 12928 6972 12980
rect 2228 12860 2280 12912
rect 4436 12860 4488 12912
rect 4896 12860 4948 12912
rect 5632 12860 5684 12912
rect 10600 12928 10652 12980
rect 11612 12928 11664 12980
rect 2964 12792 3016 12844
rect 4528 12835 4580 12844
rect 3148 12724 3200 12776
rect 4528 12801 4537 12835
rect 4537 12801 4571 12835
rect 4571 12801 4580 12835
rect 4528 12792 4580 12801
rect 5908 12792 5960 12844
rect 6828 12792 6880 12844
rect 7380 12792 7432 12844
rect 9312 12835 9364 12844
rect 9312 12801 9321 12835
rect 9321 12801 9355 12835
rect 9355 12801 9364 12835
rect 9312 12792 9364 12801
rect 9588 12860 9640 12912
rect 11060 12860 11112 12912
rect 10140 12792 10192 12844
rect 10784 12835 10836 12844
rect 10784 12801 10793 12835
rect 10793 12801 10827 12835
rect 10827 12801 10836 12835
rect 13820 12903 13872 12912
rect 11612 12835 11664 12844
rect 10784 12792 10836 12801
rect 11612 12801 11621 12835
rect 11621 12801 11655 12835
rect 11655 12801 11664 12835
rect 11612 12792 11664 12801
rect 4344 12656 4396 12708
rect 6276 12724 6328 12776
rect 6920 12724 6972 12776
rect 6552 12656 6604 12708
rect 7564 12656 7616 12708
rect 8944 12699 8996 12708
rect 8944 12665 8953 12699
rect 8953 12665 8987 12699
rect 8987 12665 8996 12699
rect 8944 12656 8996 12665
rect 13084 12835 13136 12844
rect 13084 12801 13093 12835
rect 13093 12801 13127 12835
rect 13127 12801 13136 12835
rect 13084 12792 13136 12801
rect 13820 12869 13829 12903
rect 13829 12869 13863 12903
rect 13863 12869 13872 12903
rect 13820 12860 13872 12869
rect 14648 12860 14700 12912
rect 15476 12860 15528 12912
rect 13912 12792 13964 12844
rect 14004 12835 14056 12844
rect 14004 12801 14013 12835
rect 14013 12801 14047 12835
rect 14047 12801 14056 12835
rect 14004 12792 14056 12801
rect 16764 12928 16816 12980
rect 15752 12835 15804 12844
rect 12072 12724 12124 12776
rect 15752 12801 15761 12835
rect 15761 12801 15795 12835
rect 15795 12801 15804 12835
rect 17040 12835 17092 12844
rect 15752 12792 15804 12801
rect 17040 12801 17049 12835
rect 17049 12801 17083 12835
rect 17083 12801 17092 12835
rect 17040 12792 17092 12801
rect 17776 12835 17828 12844
rect 17776 12801 17785 12835
rect 17785 12801 17819 12835
rect 17819 12801 17828 12835
rect 17776 12792 17828 12801
rect 12716 12656 12768 12708
rect 16028 12656 16080 12708
rect 1768 12588 1820 12640
rect 12256 12588 12308 12640
rect 14004 12588 14056 12640
rect 15384 12588 15436 12640
rect 18236 12631 18288 12640
rect 18236 12597 18245 12631
rect 18245 12597 18279 12631
rect 18279 12597 18288 12631
rect 18236 12588 18288 12597
rect 4214 12486 4266 12538
rect 4278 12486 4330 12538
rect 4342 12486 4394 12538
rect 4406 12486 4458 12538
rect 4470 12486 4522 12538
rect 12214 12486 12266 12538
rect 12278 12486 12330 12538
rect 12342 12486 12394 12538
rect 12406 12486 12458 12538
rect 12470 12486 12522 12538
rect 3424 12427 3476 12436
rect 3424 12393 3433 12427
rect 3433 12393 3467 12427
rect 3467 12393 3476 12427
rect 3424 12384 3476 12393
rect 4620 12384 4672 12436
rect 2228 12359 2280 12368
rect 2228 12325 2237 12359
rect 2237 12325 2271 12359
rect 2271 12325 2280 12359
rect 2228 12316 2280 12325
rect 3148 12359 3200 12368
rect 3148 12325 3157 12359
rect 3157 12325 3191 12359
rect 3191 12325 3200 12359
rect 3148 12316 3200 12325
rect 4896 12359 4948 12368
rect 4896 12325 4905 12359
rect 4905 12325 4939 12359
rect 4939 12325 4948 12359
rect 4896 12316 4948 12325
rect 1768 12291 1820 12300
rect 1768 12257 1777 12291
rect 1777 12257 1811 12291
rect 1811 12257 1820 12291
rect 1768 12248 1820 12257
rect 2688 12248 2740 12300
rect 5540 12248 5592 12300
rect 3424 12180 3476 12232
rect 5908 12248 5960 12300
rect 7564 12359 7616 12368
rect 7564 12325 7573 12359
rect 7573 12325 7607 12359
rect 7607 12325 7616 12359
rect 7564 12316 7616 12325
rect 7748 12384 7800 12436
rect 9128 12384 9180 12436
rect 9312 12384 9364 12436
rect 9496 12384 9548 12436
rect 11336 12384 11388 12436
rect 12072 12384 12124 12436
rect 7380 12248 7432 12300
rect 8576 12248 8628 12300
rect 9128 12248 9180 12300
rect 11796 12316 11848 12368
rect 11888 12316 11940 12368
rect 12808 12384 12860 12436
rect 13084 12384 13136 12436
rect 13728 12384 13780 12436
rect 14280 12384 14332 12436
rect 17040 12384 17092 12436
rect 12716 12316 12768 12368
rect 6000 12223 6052 12232
rect 2228 12112 2280 12164
rect 6000 12189 6009 12223
rect 6009 12189 6043 12223
rect 6043 12189 6052 12223
rect 6000 12180 6052 12189
rect 6276 12223 6328 12232
rect 6276 12189 6285 12223
rect 6285 12189 6319 12223
rect 6319 12189 6328 12223
rect 6276 12180 6328 12189
rect 8484 12112 8536 12164
rect 8944 12112 8996 12164
rect 9220 12155 9272 12164
rect 9220 12121 9229 12155
rect 9229 12121 9263 12155
rect 9263 12121 9272 12155
rect 9220 12112 9272 12121
rect 9404 12180 9456 12232
rect 10508 12248 10560 12300
rect 12900 12316 12952 12368
rect 15476 12359 15528 12368
rect 10416 12223 10468 12232
rect 10416 12189 10420 12223
rect 10420 12189 10454 12223
rect 10454 12189 10468 12223
rect 10600 12223 10652 12232
rect 10416 12180 10468 12189
rect 10600 12189 10609 12223
rect 10609 12189 10643 12223
rect 10643 12189 10652 12223
rect 10600 12180 10652 12189
rect 12992 12248 13044 12300
rect 15200 12248 15252 12300
rect 15476 12325 15485 12359
rect 15485 12325 15519 12359
rect 15519 12325 15528 12359
rect 15476 12316 15528 12325
rect 17776 12316 17828 12368
rect 11152 12180 11204 12232
rect 11244 12223 11296 12232
rect 11244 12189 11253 12223
rect 11253 12189 11287 12223
rect 11287 12189 11296 12223
rect 11244 12180 11296 12189
rect 12440 12223 12492 12232
rect 10324 12112 10376 12164
rect 10968 12112 11020 12164
rect 3332 12044 3384 12096
rect 5816 12087 5868 12096
rect 5816 12053 5825 12087
rect 5825 12053 5859 12087
rect 5859 12053 5868 12087
rect 5816 12044 5868 12053
rect 7196 12044 7248 12096
rect 7748 12044 7800 12096
rect 9588 12087 9640 12096
rect 9588 12053 9597 12087
rect 9597 12053 9631 12087
rect 9631 12053 9640 12087
rect 9588 12044 9640 12053
rect 9680 12087 9732 12096
rect 9680 12053 9689 12087
rect 9689 12053 9723 12087
rect 9723 12053 9732 12087
rect 9680 12044 9732 12053
rect 9864 12044 9916 12096
rect 12440 12189 12449 12223
rect 12449 12189 12483 12223
rect 12483 12189 12492 12223
rect 12440 12180 12492 12189
rect 12532 12180 12584 12232
rect 12900 12223 12952 12232
rect 12900 12189 12903 12223
rect 12903 12189 12952 12223
rect 12900 12180 12952 12189
rect 13084 12180 13136 12232
rect 13636 12223 13688 12232
rect 13636 12189 13645 12223
rect 13645 12189 13679 12223
rect 13679 12189 13688 12223
rect 13636 12180 13688 12189
rect 14188 12223 14240 12232
rect 14188 12189 14197 12223
rect 14197 12189 14231 12223
rect 14231 12189 14240 12223
rect 14188 12180 14240 12189
rect 15384 12223 15436 12232
rect 15384 12189 15393 12223
rect 15393 12189 15427 12223
rect 15427 12189 15436 12223
rect 15384 12180 15436 12189
rect 16028 12180 16080 12232
rect 16948 12223 17000 12232
rect 16948 12189 16957 12223
rect 16957 12189 16991 12223
rect 16991 12189 17000 12223
rect 16948 12180 17000 12189
rect 18236 12248 18288 12300
rect 15292 12112 15344 12164
rect 11796 12044 11848 12096
rect 11980 12087 12032 12096
rect 11980 12053 11989 12087
rect 11989 12053 12023 12087
rect 12023 12053 12032 12087
rect 11980 12044 12032 12053
rect 12808 12044 12860 12096
rect 14832 12044 14884 12096
rect 16028 12044 16080 12096
rect 16120 12044 16172 12096
rect 16764 12087 16816 12096
rect 16764 12053 16773 12087
rect 16773 12053 16807 12087
rect 16807 12053 16816 12087
rect 16764 12044 16816 12053
rect 17224 12044 17276 12096
rect 8214 11942 8266 11994
rect 8278 11942 8330 11994
rect 8342 11942 8394 11994
rect 8406 11942 8458 11994
rect 8470 11942 8522 11994
rect 16214 11942 16266 11994
rect 16278 11942 16330 11994
rect 16342 11942 16394 11994
rect 16406 11942 16458 11994
rect 16470 11942 16522 11994
rect 2964 11883 3016 11892
rect 2964 11849 2973 11883
rect 2973 11849 3007 11883
rect 3007 11849 3016 11883
rect 2964 11840 3016 11849
rect 2320 11815 2372 11824
rect 2320 11781 2329 11815
rect 2329 11781 2363 11815
rect 2363 11781 2372 11815
rect 2320 11772 2372 11781
rect 3424 11815 3476 11824
rect 3424 11781 3433 11815
rect 3433 11781 3467 11815
rect 3467 11781 3476 11815
rect 3424 11772 3476 11781
rect 1492 11636 1544 11688
rect 2228 11611 2280 11620
rect 2228 11577 2237 11611
rect 2237 11577 2271 11611
rect 2271 11577 2280 11611
rect 2228 11568 2280 11577
rect 3332 11704 3384 11756
rect 6184 11840 6236 11892
rect 7012 11840 7064 11892
rect 4068 11772 4120 11824
rect 5172 11772 5224 11824
rect 5908 11772 5960 11824
rect 6276 11772 6328 11824
rect 8208 11772 8260 11824
rect 3884 11679 3936 11688
rect 3884 11645 3893 11679
rect 3893 11645 3927 11679
rect 3927 11645 3936 11679
rect 3884 11636 3936 11645
rect 6092 11704 6144 11756
rect 7012 11704 7064 11756
rect 8024 11704 8076 11756
rect 9404 11840 9456 11892
rect 9680 11840 9732 11892
rect 10508 11840 10560 11892
rect 10600 11840 10652 11892
rect 11060 11840 11112 11892
rect 8576 11815 8628 11824
rect 8576 11781 8585 11815
rect 8585 11781 8619 11815
rect 8619 11781 8628 11815
rect 8576 11772 8628 11781
rect 9956 11772 10008 11824
rect 10140 11772 10192 11824
rect 11244 11772 11296 11824
rect 11704 11772 11756 11824
rect 12164 11840 12216 11892
rect 12348 11772 12400 11824
rect 13820 11840 13872 11892
rect 14096 11840 14148 11892
rect 15384 11883 15436 11892
rect 15384 11849 15393 11883
rect 15393 11849 15427 11883
rect 15427 11849 15436 11883
rect 15384 11840 15436 11849
rect 13912 11815 13964 11824
rect 13912 11781 13921 11815
rect 13921 11781 13955 11815
rect 13955 11781 13964 11815
rect 13912 11772 13964 11781
rect 14280 11815 14332 11824
rect 14280 11781 14289 11815
rect 14289 11781 14323 11815
rect 14323 11781 14332 11815
rect 14280 11772 14332 11781
rect 14924 11772 14976 11824
rect 15016 11815 15068 11824
rect 15016 11781 15025 11815
rect 15025 11781 15059 11815
rect 15059 11781 15068 11815
rect 15016 11772 15068 11781
rect 5172 11568 5224 11620
rect 5356 11636 5408 11688
rect 8208 11568 8260 11620
rect 9496 11704 9548 11756
rect 9864 11704 9916 11756
rect 10232 11747 10284 11756
rect 10232 11713 10241 11747
rect 10241 11713 10275 11747
rect 10275 11713 10284 11747
rect 10232 11704 10284 11713
rect 8668 11636 8720 11688
rect 9956 11679 10008 11688
rect 9956 11645 9965 11679
rect 9965 11645 9999 11679
rect 9999 11645 10008 11679
rect 9956 11636 10008 11645
rect 10508 11679 10560 11688
rect 10508 11645 10517 11679
rect 10517 11645 10551 11679
rect 10551 11645 10560 11679
rect 10508 11636 10560 11645
rect 8576 11568 8628 11620
rect 9496 11568 9548 11620
rect 11520 11704 11572 11756
rect 11980 11747 12032 11756
rect 11612 11568 11664 11620
rect 11980 11713 11994 11747
rect 11994 11713 12028 11747
rect 12028 11713 12032 11747
rect 11980 11704 12032 11713
rect 14096 11747 14148 11756
rect 14096 11713 14105 11747
rect 14105 11713 14139 11747
rect 14139 11713 14148 11747
rect 14096 11704 14148 11713
rect 14372 11747 14424 11756
rect 14372 11713 14381 11747
rect 14381 11713 14415 11747
rect 14415 11713 14424 11747
rect 14372 11704 14424 11713
rect 12072 11636 12124 11688
rect 15752 11704 15804 11756
rect 16120 11704 16172 11756
rect 15476 11679 15528 11688
rect 15476 11645 15485 11679
rect 15485 11645 15519 11679
rect 15519 11645 15528 11679
rect 15476 11636 15528 11645
rect 15568 11679 15620 11688
rect 15568 11645 15577 11679
rect 15577 11645 15611 11679
rect 15611 11645 15620 11679
rect 17684 11704 17736 11756
rect 15568 11636 15620 11645
rect 10876 11500 10928 11552
rect 10968 11500 11020 11552
rect 14924 11568 14976 11620
rect 16764 11568 16816 11620
rect 16856 11568 16908 11620
rect 18144 11611 18196 11620
rect 18144 11577 18153 11611
rect 18153 11577 18187 11611
rect 18187 11577 18196 11611
rect 18144 11568 18196 11577
rect 12624 11543 12676 11552
rect 12624 11509 12633 11543
rect 12633 11509 12667 11543
rect 12667 11509 12676 11543
rect 12624 11500 12676 11509
rect 12808 11500 12860 11552
rect 13360 11500 13412 11552
rect 13544 11500 13596 11552
rect 14648 11500 14700 11552
rect 17132 11500 17184 11552
rect 4214 11398 4266 11450
rect 4278 11398 4330 11450
rect 4342 11398 4394 11450
rect 4406 11398 4458 11450
rect 4470 11398 4522 11450
rect 12214 11398 12266 11450
rect 12278 11398 12330 11450
rect 12342 11398 12394 11450
rect 12406 11398 12458 11450
rect 12470 11398 12522 11450
rect 3424 11339 3476 11348
rect 3424 11305 3433 11339
rect 3433 11305 3467 11339
rect 3467 11305 3476 11339
rect 3424 11296 3476 11305
rect 10968 11296 11020 11348
rect 12992 11296 13044 11348
rect 13636 11296 13688 11348
rect 13820 11296 13872 11348
rect 15292 11339 15344 11348
rect 15292 11305 15301 11339
rect 15301 11305 15335 11339
rect 15335 11305 15344 11339
rect 15292 11296 15344 11305
rect 2228 11228 2280 11280
rect 5172 11271 5224 11280
rect 5172 11237 5181 11271
rect 5181 11237 5215 11271
rect 5215 11237 5224 11271
rect 5172 11228 5224 11237
rect 6092 11228 6144 11280
rect 7288 11228 7340 11280
rect 8668 11271 8720 11280
rect 6736 11160 6788 11212
rect 1492 11135 1544 11144
rect 1492 11101 1501 11135
rect 1501 11101 1535 11135
rect 1535 11101 1544 11135
rect 1492 11092 1544 11101
rect 2964 11135 3016 11144
rect 2964 11101 2973 11135
rect 2973 11101 3007 11135
rect 3007 11101 3016 11135
rect 2964 11092 3016 11101
rect 3884 11135 3936 11144
rect 3884 11101 3893 11135
rect 3893 11101 3927 11135
rect 3927 11101 3936 11135
rect 3884 11092 3936 11101
rect 5908 11135 5960 11144
rect 5908 11101 5917 11135
rect 5917 11101 5951 11135
rect 5951 11101 5960 11135
rect 5908 11092 5960 11101
rect 6092 11092 6144 11144
rect 6828 11092 6880 11144
rect 8668 11237 8677 11271
rect 8677 11237 8711 11271
rect 8711 11237 8720 11271
rect 8668 11228 8720 11237
rect 10048 11271 10100 11280
rect 10048 11237 10057 11271
rect 10057 11237 10091 11271
rect 10091 11237 10100 11271
rect 10048 11228 10100 11237
rect 10508 11228 10560 11280
rect 7840 11092 7892 11144
rect 8116 11092 8168 11144
rect 8760 11092 8812 11144
rect 9496 11135 9548 11144
rect 6000 11024 6052 11076
rect 7196 11024 7248 11076
rect 2412 10956 2464 11008
rect 7012 10956 7064 11008
rect 7472 10999 7524 11008
rect 7472 10965 7481 10999
rect 7481 10965 7515 10999
rect 7515 10965 7524 10999
rect 9036 11067 9088 11076
rect 9036 11033 9045 11067
rect 9045 11033 9079 11067
rect 9079 11033 9088 11067
rect 9496 11101 9504 11135
rect 9504 11101 9538 11135
rect 9538 11101 9548 11135
rect 9956 11160 10008 11212
rect 11152 11228 11204 11280
rect 10876 11160 10928 11212
rect 11520 11203 11572 11212
rect 11520 11169 11529 11203
rect 11529 11169 11563 11203
rect 11563 11169 11572 11203
rect 11520 11160 11572 11169
rect 9496 11092 9548 11101
rect 10416 11135 10468 11144
rect 10416 11101 10425 11135
rect 10425 11101 10459 11135
rect 10459 11101 10468 11135
rect 10416 11092 10468 11101
rect 10784 11092 10836 11144
rect 10968 11135 11020 11144
rect 10968 11101 10977 11135
rect 10977 11101 11011 11135
rect 11011 11101 11020 11135
rect 10968 11092 11020 11101
rect 9036 11024 9088 11033
rect 10692 11024 10744 11076
rect 7472 10956 7524 10965
rect 10232 10956 10284 11008
rect 11704 11092 11756 11144
rect 12624 11228 12676 11280
rect 12900 11160 12952 11212
rect 13268 11203 13320 11212
rect 13268 11169 13277 11203
rect 13277 11169 13311 11203
rect 13311 11169 13320 11203
rect 13268 11160 13320 11169
rect 15200 11228 15252 11280
rect 15568 11228 15620 11280
rect 12440 11092 12492 11144
rect 13176 11135 13228 11144
rect 13176 11101 13185 11135
rect 13185 11101 13219 11135
rect 13219 11101 13228 11135
rect 13176 11092 13228 11101
rect 13452 11135 13504 11144
rect 13452 11101 13461 11135
rect 13461 11101 13495 11135
rect 13495 11101 13504 11135
rect 13452 11092 13504 11101
rect 13728 11092 13780 11144
rect 11520 10956 11572 11008
rect 13820 11024 13872 11076
rect 12348 10956 12400 11008
rect 13636 10956 13688 11008
rect 14648 11160 14700 11212
rect 14832 11092 14884 11144
rect 15844 11092 15896 11144
rect 17132 11203 17184 11212
rect 17132 11169 17141 11203
rect 17141 11169 17175 11203
rect 17175 11169 17184 11203
rect 17132 11160 17184 11169
rect 17500 11228 17552 11280
rect 16672 11135 16724 11144
rect 16672 11101 16681 11135
rect 16681 11101 16715 11135
rect 16715 11101 16724 11135
rect 16672 11092 16724 11101
rect 18052 11092 18104 11144
rect 15568 11024 15620 11076
rect 16856 11067 16908 11076
rect 16856 11033 16865 11067
rect 16865 11033 16899 11067
rect 16899 11033 16908 11067
rect 16856 11024 16908 11033
rect 14280 10956 14332 11008
rect 8214 10854 8266 10906
rect 8278 10854 8330 10906
rect 8342 10854 8394 10906
rect 8406 10854 8458 10906
rect 8470 10854 8522 10906
rect 16214 10854 16266 10906
rect 16278 10854 16330 10906
rect 16342 10854 16394 10906
rect 16406 10854 16458 10906
rect 16470 10854 16522 10906
rect 1492 10684 1544 10736
rect 2780 10684 2832 10736
rect 3884 10684 3936 10736
rect 5816 10684 5868 10736
rect 6736 10727 6788 10736
rect 6736 10693 6745 10727
rect 6745 10693 6779 10727
rect 6779 10693 6788 10727
rect 6736 10684 6788 10693
rect 7104 10684 7156 10736
rect 8576 10752 8628 10804
rect 12256 10752 12308 10804
rect 14924 10752 14976 10804
rect 15200 10795 15252 10804
rect 15200 10761 15209 10795
rect 15209 10761 15243 10795
rect 15243 10761 15252 10795
rect 15200 10752 15252 10761
rect 2044 10659 2096 10668
rect 2044 10625 2053 10659
rect 2053 10625 2087 10659
rect 2087 10625 2096 10659
rect 2044 10616 2096 10625
rect 4068 10659 4120 10668
rect 4068 10625 4077 10659
rect 4077 10625 4111 10659
rect 4111 10625 4120 10659
rect 4068 10616 4120 10625
rect 5908 10616 5960 10668
rect 6092 10659 6144 10668
rect 6092 10625 6101 10659
rect 6101 10625 6135 10659
rect 6135 10625 6144 10659
rect 6092 10616 6144 10625
rect 7288 10659 7340 10668
rect 7288 10625 7297 10659
rect 7297 10625 7331 10659
rect 7331 10625 7340 10659
rect 7288 10616 7340 10625
rect 7472 10659 7524 10668
rect 7472 10625 7481 10659
rect 7481 10625 7515 10659
rect 7515 10625 7524 10659
rect 7472 10616 7524 10625
rect 7932 10616 7984 10668
rect 8300 10659 8352 10668
rect 8300 10625 8325 10659
rect 8325 10625 8352 10659
rect 8300 10616 8352 10625
rect 8484 10616 8536 10668
rect 10232 10684 10284 10736
rect 11060 10684 11112 10736
rect 12348 10684 12400 10736
rect 12532 10727 12584 10736
rect 12532 10693 12541 10727
rect 12541 10693 12575 10727
rect 12575 10693 12584 10727
rect 12532 10684 12584 10693
rect 13176 10684 13228 10736
rect 13360 10684 13412 10736
rect 13636 10684 13688 10736
rect 13820 10684 13872 10736
rect 14464 10727 14516 10736
rect 14464 10693 14473 10727
rect 14473 10693 14507 10727
rect 14507 10693 14516 10727
rect 14464 10684 14516 10693
rect 15476 10752 15528 10804
rect 16672 10752 16724 10804
rect 15844 10727 15896 10736
rect 9864 10616 9916 10668
rect 9956 10616 10008 10668
rect 2320 10548 2372 10600
rect 3976 10591 4028 10600
rect 3976 10557 3985 10591
rect 3985 10557 4019 10591
rect 4019 10557 4028 10591
rect 3976 10548 4028 10557
rect 4804 10548 4856 10600
rect 3424 10480 3476 10532
rect 3148 10455 3200 10464
rect 3148 10421 3157 10455
rect 3157 10421 3191 10455
rect 3191 10421 3200 10455
rect 3148 10412 3200 10421
rect 3516 10412 3568 10464
rect 6920 10412 6972 10464
rect 7012 10412 7064 10464
rect 8208 10480 8260 10532
rect 9036 10480 9088 10532
rect 9588 10480 9640 10532
rect 9772 10523 9824 10532
rect 9772 10489 9781 10523
rect 9781 10489 9815 10523
rect 9815 10489 9824 10523
rect 9772 10480 9824 10489
rect 10232 10548 10284 10600
rect 10508 10659 10560 10668
rect 10508 10625 10517 10659
rect 10517 10625 10551 10659
rect 10551 10625 10560 10659
rect 10508 10616 10560 10625
rect 11428 10616 11480 10668
rect 11888 10616 11940 10668
rect 12164 10659 12216 10668
rect 12164 10625 12173 10659
rect 12173 10625 12207 10659
rect 12207 10625 12216 10659
rect 12164 10616 12216 10625
rect 12624 10659 12676 10668
rect 12624 10625 12633 10659
rect 12633 10625 12667 10659
rect 12667 10625 12676 10659
rect 12624 10616 12676 10625
rect 13084 10616 13136 10668
rect 13268 10659 13320 10668
rect 13268 10625 13277 10659
rect 13277 10625 13311 10659
rect 13311 10625 13320 10659
rect 13268 10616 13320 10625
rect 15844 10693 15853 10727
rect 15853 10693 15887 10727
rect 15887 10693 15896 10727
rect 15844 10684 15896 10693
rect 17500 10727 17552 10736
rect 17500 10693 17509 10727
rect 17509 10693 17543 10727
rect 17543 10693 17552 10727
rect 17500 10684 17552 10693
rect 18144 10684 18196 10736
rect 15292 10616 15344 10668
rect 15476 10616 15528 10668
rect 11612 10548 11664 10600
rect 11704 10548 11756 10600
rect 14280 10548 14332 10600
rect 14556 10548 14608 10600
rect 11152 10480 11204 10532
rect 12624 10480 12676 10532
rect 12900 10480 12952 10532
rect 8392 10412 8444 10464
rect 8852 10412 8904 10464
rect 9496 10412 9548 10464
rect 9864 10412 9916 10464
rect 10416 10412 10468 10464
rect 10876 10412 10928 10464
rect 12808 10412 12860 10464
rect 13912 10412 13964 10464
rect 15016 10412 15068 10464
rect 16764 10548 16816 10600
rect 17684 10548 17736 10600
rect 17408 10523 17460 10532
rect 17408 10489 17417 10523
rect 17417 10489 17451 10523
rect 17451 10489 17460 10523
rect 17408 10480 17460 10489
rect 4214 10310 4266 10362
rect 4278 10310 4330 10362
rect 4342 10310 4394 10362
rect 4406 10310 4458 10362
rect 4470 10310 4522 10362
rect 12214 10310 12266 10362
rect 12278 10310 12330 10362
rect 12342 10310 12394 10362
rect 12406 10310 12458 10362
rect 12470 10310 12522 10362
rect 3976 10208 4028 10260
rect 3884 10140 3936 10192
rect 3516 10115 3568 10124
rect 3516 10081 3525 10115
rect 3525 10081 3559 10115
rect 3559 10081 3568 10115
rect 3516 10072 3568 10081
rect 3792 10072 3844 10124
rect 11428 10140 11480 10192
rect 5908 10072 5960 10124
rect 2412 10047 2464 10056
rect 2412 10013 2421 10047
rect 2421 10013 2455 10047
rect 2455 10013 2464 10047
rect 2412 10004 2464 10013
rect 2780 10004 2832 10056
rect 4068 10047 4120 10056
rect 4068 10013 4077 10047
rect 4077 10013 4111 10047
rect 4111 10013 4120 10047
rect 4068 10004 4120 10013
rect 4804 10047 4856 10056
rect 4804 10013 4813 10047
rect 4813 10013 4847 10047
rect 4847 10013 4856 10047
rect 4804 10004 4856 10013
rect 5264 10047 5316 10056
rect 5264 10013 5273 10047
rect 5273 10013 5307 10047
rect 5307 10013 5316 10047
rect 5264 10004 5316 10013
rect 6000 10004 6052 10056
rect 7288 10072 7340 10124
rect 7840 10072 7892 10124
rect 7012 10047 7064 10056
rect 4252 9936 4304 9988
rect 6736 9979 6788 9988
rect 1768 9911 1820 9920
rect 1768 9877 1777 9911
rect 1777 9877 1811 9911
rect 1811 9877 1820 9911
rect 1768 9868 1820 9877
rect 2320 9868 2372 9920
rect 3332 9868 3384 9920
rect 6736 9945 6745 9979
rect 6745 9945 6779 9979
rect 6779 9945 6788 9979
rect 6736 9936 6788 9945
rect 7012 10013 7021 10047
rect 7021 10013 7055 10047
rect 7055 10013 7064 10047
rect 7012 10004 7064 10013
rect 8300 10072 8352 10124
rect 8668 10072 8720 10124
rect 8208 10047 8260 10056
rect 8208 10013 8217 10047
rect 8217 10013 8251 10047
rect 8251 10013 8260 10047
rect 8208 10004 8260 10013
rect 8760 10004 8812 10056
rect 9772 10072 9824 10124
rect 10048 10115 10100 10124
rect 10048 10081 10057 10115
rect 10057 10081 10091 10115
rect 10091 10081 10100 10115
rect 10048 10072 10100 10081
rect 10416 10072 10468 10124
rect 9864 10047 9916 10056
rect 8576 9936 8628 9988
rect 9864 10013 9873 10047
rect 9873 10013 9907 10047
rect 9907 10013 9916 10047
rect 9864 10004 9916 10013
rect 10784 10004 10836 10056
rect 10876 10047 10928 10056
rect 10876 10013 10885 10047
rect 10885 10013 10919 10047
rect 10919 10013 10928 10047
rect 10876 10004 10928 10013
rect 11980 10208 12032 10260
rect 13544 10208 13596 10260
rect 14188 10208 14240 10260
rect 18052 10251 18104 10260
rect 18052 10217 18061 10251
rect 18061 10217 18095 10251
rect 18095 10217 18104 10251
rect 18052 10208 18104 10217
rect 12808 10140 12860 10192
rect 13268 10140 13320 10192
rect 14924 10140 14976 10192
rect 14188 10072 14240 10124
rect 10140 9979 10192 9988
rect 10140 9945 10149 9979
rect 10149 9945 10183 9979
rect 10183 9945 10192 9979
rect 10140 9936 10192 9945
rect 11060 9936 11112 9988
rect 7932 9868 7984 9920
rect 9496 9868 9548 9920
rect 9680 9868 9732 9920
rect 10692 9868 10744 9920
rect 12808 10004 12860 10056
rect 11704 9936 11756 9988
rect 11520 9868 11572 9920
rect 12072 9911 12124 9920
rect 12072 9877 12081 9911
rect 12081 9877 12115 9911
rect 12115 9877 12124 9911
rect 12072 9868 12124 9877
rect 12624 9911 12676 9920
rect 12624 9877 12633 9911
rect 12633 9877 12667 9911
rect 12667 9877 12676 9911
rect 12624 9868 12676 9877
rect 13268 10047 13320 10056
rect 13268 10013 13277 10047
rect 13277 10013 13311 10047
rect 13311 10013 13320 10047
rect 13268 10004 13320 10013
rect 13728 10004 13780 10056
rect 15016 10072 15068 10124
rect 15384 10115 15436 10124
rect 15384 10081 15393 10115
rect 15393 10081 15427 10115
rect 15427 10081 15436 10115
rect 15384 10072 15436 10081
rect 14740 10047 14792 10056
rect 14740 10013 14749 10047
rect 14749 10013 14783 10047
rect 14783 10013 14792 10047
rect 14740 10004 14792 10013
rect 14832 10047 14884 10056
rect 14832 10013 14841 10047
rect 14841 10013 14875 10047
rect 14875 10013 14884 10047
rect 15108 10047 15160 10056
rect 14832 10004 14884 10013
rect 15108 10013 15117 10047
rect 15117 10013 15151 10047
rect 15151 10013 15160 10047
rect 15108 10004 15160 10013
rect 15660 10047 15712 10056
rect 14648 9936 14700 9988
rect 15660 10013 15669 10047
rect 15669 10013 15703 10047
rect 15703 10013 15712 10047
rect 15660 10004 15712 10013
rect 16764 10047 16816 10056
rect 16764 10013 16773 10047
rect 16773 10013 16807 10047
rect 16807 10013 16816 10047
rect 16764 10004 16816 10013
rect 17684 10047 17736 10056
rect 17684 10013 17693 10047
rect 17693 10013 17727 10047
rect 17727 10013 17736 10047
rect 17684 10004 17736 10013
rect 18144 10047 18196 10056
rect 18144 10013 18153 10047
rect 18153 10013 18187 10047
rect 18187 10013 18196 10047
rect 18144 10004 18196 10013
rect 13084 9868 13136 9920
rect 13176 9868 13228 9920
rect 16672 9936 16724 9988
rect 17408 9979 17460 9988
rect 17408 9945 17417 9979
rect 17417 9945 17451 9979
rect 17451 9945 17460 9979
rect 17408 9936 17460 9945
rect 8214 9766 8266 9818
rect 8278 9766 8330 9818
rect 8342 9766 8394 9818
rect 8406 9766 8458 9818
rect 8470 9766 8522 9818
rect 16214 9766 16266 9818
rect 16278 9766 16330 9818
rect 16342 9766 16394 9818
rect 16406 9766 16458 9818
rect 16470 9766 16522 9818
rect 2596 9664 2648 9716
rect 3424 9664 3476 9716
rect 3700 9664 3752 9716
rect 3148 9596 3200 9648
rect 5908 9596 5960 9648
rect 2228 9571 2280 9580
rect 2228 9537 2237 9571
rect 2237 9537 2271 9571
rect 2271 9537 2280 9571
rect 2228 9528 2280 9537
rect 2780 9571 2832 9580
rect 2780 9537 2789 9571
rect 2789 9537 2823 9571
rect 2823 9537 2832 9571
rect 4252 9571 4304 9580
rect 2780 9528 2832 9537
rect 4252 9537 4261 9571
rect 4261 9537 4295 9571
rect 4295 9537 4304 9571
rect 4252 9528 4304 9537
rect 5080 9571 5132 9580
rect 5080 9537 5089 9571
rect 5089 9537 5123 9571
rect 5123 9537 5132 9571
rect 5080 9528 5132 9537
rect 5724 9528 5776 9580
rect 6092 9571 6144 9580
rect 6092 9537 6101 9571
rect 6101 9537 6135 9571
rect 6135 9537 6144 9571
rect 6092 9528 6144 9537
rect 5264 9460 5316 9512
rect 7196 9528 7248 9580
rect 8668 9596 8720 9648
rect 9128 9639 9180 9648
rect 9128 9605 9137 9639
rect 9137 9605 9171 9639
rect 9171 9605 9180 9639
rect 9128 9596 9180 9605
rect 8300 9571 8352 9580
rect 7932 9503 7984 9512
rect 3884 9392 3936 9444
rect 7196 9435 7248 9444
rect 7196 9401 7205 9435
rect 7205 9401 7239 9435
rect 7239 9401 7248 9435
rect 7196 9392 7248 9401
rect 2044 9367 2096 9376
rect 2044 9333 2053 9367
rect 2053 9333 2087 9367
rect 2087 9333 2096 9367
rect 2044 9324 2096 9333
rect 4896 9367 4948 9376
rect 4896 9333 4905 9367
rect 4905 9333 4939 9367
rect 4939 9333 4948 9367
rect 4896 9324 4948 9333
rect 6920 9324 6972 9376
rect 7932 9469 7941 9503
rect 7941 9469 7975 9503
rect 7975 9469 7984 9503
rect 7932 9460 7984 9469
rect 8300 9537 8309 9571
rect 8309 9537 8343 9571
rect 8343 9537 8352 9571
rect 8300 9528 8352 9537
rect 8484 9571 8536 9580
rect 8484 9537 8493 9571
rect 8493 9537 8527 9571
rect 8527 9537 8536 9571
rect 8484 9528 8536 9537
rect 8944 9528 8996 9580
rect 10048 9596 10100 9648
rect 10140 9639 10192 9648
rect 10140 9605 10158 9639
rect 10158 9605 10192 9639
rect 11060 9664 11112 9716
rect 10140 9596 10192 9605
rect 11796 9596 11848 9648
rect 13452 9664 13504 9716
rect 14004 9596 14056 9648
rect 9588 9528 9640 9580
rect 9680 9528 9732 9580
rect 10508 9528 10560 9580
rect 10784 9571 10836 9580
rect 10784 9537 10793 9571
rect 10793 9537 10827 9571
rect 10827 9537 10836 9571
rect 10784 9528 10836 9537
rect 10968 9571 11020 9580
rect 10968 9537 10977 9571
rect 10977 9537 11011 9571
rect 11011 9537 11020 9571
rect 10968 9528 11020 9537
rect 11704 9571 11756 9580
rect 11704 9537 11713 9571
rect 11713 9537 11747 9571
rect 11747 9537 11756 9571
rect 11704 9528 11756 9537
rect 8668 9460 8720 9512
rect 11888 9460 11940 9512
rect 12532 9528 12584 9580
rect 12624 9528 12676 9580
rect 13176 9571 13228 9580
rect 13176 9537 13185 9571
rect 13185 9537 13219 9571
rect 13219 9537 13228 9571
rect 13176 9528 13228 9537
rect 13452 9528 13504 9580
rect 13728 9528 13780 9580
rect 14280 9571 14332 9580
rect 14280 9537 14289 9571
rect 14289 9537 14323 9571
rect 14323 9537 14332 9571
rect 14280 9528 14332 9537
rect 14740 9664 14792 9716
rect 15292 9639 15344 9648
rect 15292 9605 15301 9639
rect 15301 9605 15335 9639
rect 15335 9605 15344 9639
rect 15292 9596 15344 9605
rect 14556 9571 14608 9580
rect 14556 9537 14565 9571
rect 14565 9537 14599 9571
rect 14599 9537 14608 9571
rect 14556 9528 14608 9537
rect 15200 9571 15252 9580
rect 15200 9537 15209 9571
rect 15209 9537 15243 9571
rect 15243 9537 15252 9571
rect 15200 9528 15252 9537
rect 15384 9571 15436 9580
rect 15384 9537 15393 9571
rect 15393 9537 15427 9571
rect 15427 9537 15436 9571
rect 15384 9528 15436 9537
rect 15660 9571 15712 9580
rect 15660 9537 15669 9571
rect 15669 9537 15703 9571
rect 15703 9537 15712 9571
rect 15660 9528 15712 9537
rect 16672 9596 16724 9648
rect 16764 9596 16816 9648
rect 17224 9639 17276 9648
rect 17224 9605 17233 9639
rect 17233 9605 17267 9639
rect 17267 9605 17276 9639
rect 17224 9596 17276 9605
rect 17776 9528 17828 9580
rect 13084 9460 13136 9512
rect 8576 9324 8628 9376
rect 9956 9324 10008 9376
rect 10508 9324 10560 9376
rect 12716 9392 12768 9444
rect 12808 9392 12860 9444
rect 14464 9435 14516 9444
rect 14464 9401 14473 9435
rect 14473 9401 14507 9435
rect 14507 9401 14516 9435
rect 14464 9392 14516 9401
rect 16672 9460 16724 9512
rect 14740 9392 14792 9444
rect 15384 9392 15436 9444
rect 15568 9392 15620 9444
rect 18052 9435 18104 9444
rect 18052 9401 18061 9435
rect 18061 9401 18095 9435
rect 18095 9401 18104 9435
rect 18052 9392 18104 9401
rect 13544 9324 13596 9376
rect 13636 9324 13688 9376
rect 13820 9324 13872 9376
rect 16028 9324 16080 9376
rect 4214 9222 4266 9274
rect 4278 9222 4330 9274
rect 4342 9222 4394 9274
rect 4406 9222 4458 9274
rect 4470 9222 4522 9274
rect 12214 9222 12266 9274
rect 12278 9222 12330 9274
rect 12342 9222 12394 9274
rect 12406 9222 12458 9274
rect 12470 9222 12522 9274
rect 5724 9120 5776 9172
rect 5264 9052 5316 9104
rect 2596 8984 2648 9036
rect 6920 9052 6972 9104
rect 7288 9120 7340 9172
rect 9864 9120 9916 9172
rect 10508 9163 10560 9172
rect 10508 9129 10517 9163
rect 10517 9129 10551 9163
rect 10551 9129 10560 9163
rect 10508 9120 10560 9129
rect 10784 9120 10836 9172
rect 12440 9120 12492 9172
rect 13544 9120 13596 9172
rect 7932 9052 7984 9104
rect 8576 9052 8628 9104
rect 9588 9095 9640 9104
rect 9588 9061 9597 9095
rect 9597 9061 9631 9095
rect 9631 9061 9640 9095
rect 9588 9052 9640 9061
rect 9772 9052 9824 9104
rect 10692 9052 10744 9104
rect 2044 8959 2096 8968
rect 2044 8925 2053 8959
rect 2053 8925 2087 8959
rect 2087 8925 2096 8959
rect 2044 8916 2096 8925
rect 1492 8891 1544 8900
rect 1492 8857 1501 8891
rect 1501 8857 1535 8891
rect 1535 8857 1544 8891
rect 1492 8848 1544 8857
rect 4160 8848 4212 8900
rect 6000 8959 6052 8968
rect 6000 8925 6009 8959
rect 6009 8925 6043 8959
rect 6043 8925 6052 8959
rect 6000 8916 6052 8925
rect 6828 8959 6880 8968
rect 6828 8925 6837 8959
rect 6837 8925 6871 8959
rect 6871 8925 6880 8959
rect 6828 8916 6880 8925
rect 7196 8959 7248 8968
rect 7196 8925 7205 8959
rect 7205 8925 7239 8959
rect 7239 8925 7248 8959
rect 7196 8916 7248 8925
rect 7656 8916 7708 8968
rect 7748 8959 7800 8968
rect 7748 8925 7757 8959
rect 7757 8925 7791 8959
rect 7791 8925 7800 8959
rect 8668 8984 8720 9036
rect 10968 9052 11020 9104
rect 12532 9052 12584 9104
rect 13084 9052 13136 9104
rect 14280 9052 14332 9104
rect 14464 9052 14516 9104
rect 7748 8916 7800 8925
rect 9404 8959 9456 8968
rect 5448 8848 5500 8900
rect 5632 8891 5684 8900
rect 5632 8857 5641 8891
rect 5641 8857 5675 8891
rect 5675 8857 5684 8891
rect 5632 8848 5684 8857
rect 9404 8925 9413 8959
rect 9413 8925 9447 8959
rect 9447 8925 9456 8959
rect 9404 8916 9456 8925
rect 9496 8916 9548 8968
rect 10600 8916 10652 8968
rect 9772 8848 9824 8900
rect 7564 8780 7616 8832
rect 7840 8823 7892 8832
rect 7840 8789 7849 8823
rect 7849 8789 7883 8823
rect 7883 8789 7892 8823
rect 7840 8780 7892 8789
rect 8576 8823 8628 8832
rect 8576 8789 8585 8823
rect 8585 8789 8619 8823
rect 8619 8789 8628 8823
rect 8576 8780 8628 8789
rect 8668 8780 8720 8832
rect 9588 8780 9640 8832
rect 10508 8848 10560 8900
rect 11704 8916 11756 8968
rect 12164 8959 12216 8968
rect 12164 8925 12173 8959
rect 12173 8925 12207 8959
rect 12207 8925 12216 8959
rect 12164 8916 12216 8925
rect 12440 8984 12492 9036
rect 12992 8984 13044 9036
rect 16120 9052 16172 9104
rect 12808 8916 12860 8968
rect 13084 8959 13136 8968
rect 13084 8925 13093 8959
rect 13093 8925 13127 8959
rect 13127 8925 13136 8959
rect 13084 8916 13136 8925
rect 11888 8848 11940 8900
rect 12716 8780 12768 8832
rect 13452 8916 13504 8968
rect 14004 8916 14056 8968
rect 14096 8916 14148 8968
rect 13636 8848 13688 8900
rect 14556 8959 14608 8968
rect 14556 8925 14565 8959
rect 14565 8925 14599 8959
rect 14599 8925 14608 8959
rect 14556 8916 14608 8925
rect 15568 8959 15620 8968
rect 15568 8925 15571 8959
rect 15571 8925 15620 8959
rect 15568 8916 15620 8925
rect 13820 8780 13872 8832
rect 14096 8780 14148 8832
rect 18052 9052 18104 9104
rect 16672 8959 16724 8968
rect 16672 8925 16681 8959
rect 16681 8925 16715 8959
rect 16715 8925 16724 8959
rect 16672 8916 16724 8925
rect 17684 8959 17736 8968
rect 17684 8925 17693 8959
rect 17693 8925 17727 8959
rect 17727 8925 17736 8959
rect 17684 8916 17736 8925
rect 15016 8780 15068 8832
rect 16948 8848 17000 8900
rect 15476 8780 15528 8832
rect 8214 8678 8266 8730
rect 8278 8678 8330 8730
rect 8342 8678 8394 8730
rect 8406 8678 8458 8730
rect 8470 8678 8522 8730
rect 16214 8678 16266 8730
rect 16278 8678 16330 8730
rect 16342 8678 16394 8730
rect 16406 8678 16458 8730
rect 16470 8678 16522 8730
rect 4160 8551 4212 8560
rect 4160 8517 4169 8551
rect 4169 8517 4203 8551
rect 4203 8517 4212 8551
rect 4160 8508 4212 8517
rect 2596 8483 2648 8492
rect 2596 8449 2605 8483
rect 2605 8449 2639 8483
rect 2639 8449 2648 8483
rect 2596 8440 2648 8449
rect 5080 8508 5132 8560
rect 5632 8508 5684 8560
rect 4620 8483 4672 8492
rect 4620 8449 4629 8483
rect 4629 8449 4663 8483
rect 4663 8449 4672 8483
rect 4620 8440 4672 8449
rect 5356 8483 5408 8492
rect 5356 8449 5365 8483
rect 5365 8449 5399 8483
rect 5399 8449 5408 8483
rect 5356 8440 5408 8449
rect 6092 8576 6144 8628
rect 6644 8619 6696 8628
rect 6644 8585 6653 8619
rect 6653 8585 6687 8619
rect 6687 8585 6696 8619
rect 6644 8576 6696 8585
rect 7932 8576 7984 8628
rect 6828 8508 6880 8560
rect 3976 8372 4028 8424
rect 5540 8372 5592 8424
rect 5908 8372 5960 8424
rect 6644 8304 6696 8356
rect 7656 8508 7708 8560
rect 8668 8508 8720 8560
rect 7564 8440 7616 8492
rect 8024 8440 8076 8492
rect 7748 8372 7800 8424
rect 8116 8415 8168 8424
rect 8116 8381 8125 8415
rect 8125 8381 8159 8415
rect 8159 8381 8168 8415
rect 8116 8372 8168 8381
rect 8852 8440 8904 8492
rect 8944 8440 8996 8492
rect 9404 8576 9456 8628
rect 9680 8508 9732 8560
rect 9772 8483 9824 8492
rect 9496 8372 9548 8424
rect 9772 8449 9781 8483
rect 9781 8449 9815 8483
rect 9815 8449 9824 8483
rect 9772 8440 9824 8449
rect 10140 8576 10192 8628
rect 9956 8508 10008 8560
rect 10324 8483 10376 8492
rect 10324 8449 10333 8483
rect 10333 8449 10367 8483
rect 10367 8449 10376 8483
rect 10324 8440 10376 8449
rect 10416 8483 10468 8492
rect 10416 8449 10425 8483
rect 10425 8449 10459 8483
rect 10459 8449 10468 8483
rect 12256 8508 12308 8560
rect 15108 8576 15160 8628
rect 15200 8576 15252 8628
rect 13912 8508 13964 8560
rect 10416 8440 10468 8449
rect 9864 8372 9916 8424
rect 10232 8372 10284 8424
rect 12164 8372 12216 8424
rect 12440 8440 12492 8492
rect 13176 8440 13228 8492
rect 7196 8304 7248 8356
rect 10140 8304 10192 8356
rect 10416 8304 10468 8356
rect 11152 8304 11204 8356
rect 11704 8347 11756 8356
rect 11704 8313 11713 8347
rect 11713 8313 11747 8347
rect 11747 8313 11756 8347
rect 11704 8304 11756 8313
rect 12900 8304 12952 8356
rect 1860 8279 1912 8288
rect 1860 8245 1869 8279
rect 1869 8245 1903 8279
rect 1903 8245 1912 8279
rect 1860 8236 1912 8245
rect 9220 8279 9272 8288
rect 9220 8245 9229 8279
rect 9229 8245 9263 8279
rect 9263 8245 9272 8279
rect 9220 8236 9272 8245
rect 9588 8236 9640 8288
rect 11520 8236 11572 8288
rect 11980 8236 12032 8288
rect 13820 8440 13872 8492
rect 14096 8483 14148 8492
rect 14096 8449 14105 8483
rect 14105 8449 14139 8483
rect 14139 8449 14148 8483
rect 14096 8440 14148 8449
rect 14832 8508 14884 8560
rect 15476 8551 15528 8560
rect 15476 8517 15485 8551
rect 15485 8517 15519 8551
rect 15519 8517 15528 8551
rect 15476 8508 15528 8517
rect 18052 8508 18104 8560
rect 15108 8440 15160 8492
rect 15292 8440 15344 8492
rect 16028 8440 16080 8492
rect 17960 8372 18012 8424
rect 13452 8304 13504 8356
rect 13544 8304 13596 8356
rect 14556 8304 14608 8356
rect 16672 8304 16724 8356
rect 17224 8347 17276 8356
rect 17224 8313 17233 8347
rect 17233 8313 17267 8347
rect 17267 8313 17276 8347
rect 17224 8304 17276 8313
rect 18420 8347 18472 8356
rect 18420 8313 18429 8347
rect 18429 8313 18463 8347
rect 18463 8313 18472 8347
rect 18420 8304 18472 8313
rect 13636 8236 13688 8288
rect 14832 8236 14884 8288
rect 15384 8236 15436 8288
rect 17868 8279 17920 8288
rect 17868 8245 17877 8279
rect 17877 8245 17911 8279
rect 17911 8245 17920 8279
rect 17868 8236 17920 8245
rect 4214 8134 4266 8186
rect 4278 8134 4330 8186
rect 4342 8134 4394 8186
rect 4406 8134 4458 8186
rect 4470 8134 4522 8186
rect 12214 8134 12266 8186
rect 12278 8134 12330 8186
rect 12342 8134 12394 8186
rect 12406 8134 12458 8186
rect 12470 8134 12522 8186
rect 5448 8075 5500 8084
rect 5448 8041 5457 8075
rect 5457 8041 5491 8075
rect 5491 8041 5500 8075
rect 5448 8032 5500 8041
rect 5908 8075 5960 8084
rect 5908 8041 5917 8075
rect 5917 8041 5951 8075
rect 5951 8041 5960 8075
rect 5908 8032 5960 8041
rect 8944 8032 8996 8084
rect 4620 8007 4672 8016
rect 4620 7973 4629 8007
rect 4629 7973 4663 8007
rect 4663 7973 4672 8007
rect 4620 7964 4672 7973
rect 4988 7964 5040 8016
rect 7840 7964 7892 8016
rect 1492 7871 1544 7880
rect 1492 7837 1501 7871
rect 1501 7837 1535 7871
rect 1535 7837 1544 7871
rect 1492 7828 1544 7837
rect 4896 7828 4948 7880
rect 5264 7828 5316 7880
rect 7932 7896 7984 7948
rect 11428 7896 11480 7948
rect 12900 8032 12952 8084
rect 13084 7964 13136 8016
rect 13268 7964 13320 8016
rect 14372 8032 14424 8084
rect 14188 8007 14240 8016
rect 14188 7973 14197 8007
rect 14197 7973 14231 8007
rect 14231 7973 14240 8007
rect 14188 7964 14240 7973
rect 18052 7964 18104 8016
rect 6644 7871 6696 7880
rect 6644 7837 6653 7871
rect 6653 7837 6687 7871
rect 6687 7837 6696 7871
rect 6644 7828 6696 7837
rect 7840 7871 7892 7880
rect 7840 7837 7849 7871
rect 7849 7837 7883 7871
rect 7883 7837 7892 7871
rect 7840 7828 7892 7837
rect 8576 7828 8628 7880
rect 9864 7871 9916 7880
rect 9864 7837 9873 7871
rect 9873 7837 9907 7871
rect 9907 7837 9916 7871
rect 9864 7828 9916 7837
rect 3056 7803 3108 7812
rect 3056 7769 3065 7803
rect 3065 7769 3099 7803
rect 3099 7769 3108 7803
rect 3056 7760 3108 7769
rect 3424 7760 3476 7812
rect 4620 7692 4672 7744
rect 8668 7735 8720 7744
rect 8668 7701 8677 7735
rect 8677 7701 8711 7735
rect 8711 7701 8720 7735
rect 8668 7692 8720 7701
rect 9128 7735 9180 7744
rect 9128 7701 9137 7735
rect 9137 7701 9171 7735
rect 9171 7701 9180 7735
rect 9128 7692 9180 7701
rect 9496 7760 9548 7812
rect 10508 7692 10560 7744
rect 10692 7692 10744 7744
rect 12256 7760 12308 7812
rect 15936 7896 15988 7948
rect 12716 7871 12768 7880
rect 12716 7837 12725 7871
rect 12725 7837 12759 7871
rect 12759 7837 12768 7871
rect 12992 7871 13044 7880
rect 12716 7828 12768 7837
rect 12992 7837 13001 7871
rect 13001 7837 13035 7871
rect 13035 7837 13044 7871
rect 12992 7828 13044 7837
rect 14832 7871 14884 7880
rect 14832 7837 14841 7871
rect 14841 7837 14875 7871
rect 14875 7837 14884 7871
rect 14832 7828 14884 7837
rect 17868 7871 17920 7880
rect 17868 7837 17877 7871
rect 17877 7837 17911 7871
rect 17911 7837 17920 7871
rect 17868 7828 17920 7837
rect 12164 7735 12216 7744
rect 12164 7701 12173 7735
rect 12173 7701 12207 7735
rect 12207 7701 12216 7735
rect 12164 7692 12216 7701
rect 15660 7735 15712 7744
rect 15660 7701 15669 7735
rect 15669 7701 15703 7735
rect 15703 7701 15712 7735
rect 15660 7692 15712 7701
rect 16580 7803 16632 7812
rect 16580 7769 16589 7803
rect 16589 7769 16623 7803
rect 16623 7769 16632 7803
rect 16580 7760 16632 7769
rect 17408 7692 17460 7744
rect 8214 7590 8266 7642
rect 8278 7590 8330 7642
rect 8342 7590 8394 7642
rect 8406 7590 8458 7642
rect 8470 7590 8522 7642
rect 16214 7590 16266 7642
rect 16278 7590 16330 7642
rect 16342 7590 16394 7642
rect 16406 7590 16458 7642
rect 16470 7590 16522 7642
rect 2596 7488 2648 7540
rect 5080 7488 5132 7540
rect 5540 7531 5592 7540
rect 5540 7497 5549 7531
rect 5549 7497 5583 7531
rect 5583 7497 5592 7531
rect 5540 7488 5592 7497
rect 5908 7488 5960 7540
rect 7840 7531 7892 7540
rect 4988 7420 5040 7472
rect 7840 7497 7849 7531
rect 7849 7497 7883 7531
rect 7883 7497 7892 7531
rect 7840 7488 7892 7497
rect 8116 7488 8168 7540
rect 1860 7395 1912 7404
rect 1860 7361 1869 7395
rect 1869 7361 1903 7395
rect 1903 7361 1912 7395
rect 1860 7352 1912 7361
rect 2044 7395 2096 7404
rect 2044 7361 2053 7395
rect 2053 7361 2087 7395
rect 2087 7361 2096 7395
rect 2044 7352 2096 7361
rect 3148 7395 3200 7404
rect 3148 7361 3157 7395
rect 3157 7361 3191 7395
rect 3191 7361 3200 7395
rect 3148 7352 3200 7361
rect 3608 7352 3660 7404
rect 3976 7352 4028 7404
rect 4620 7352 4672 7404
rect 4712 7352 4764 7404
rect 5080 7395 5132 7404
rect 5080 7361 5089 7395
rect 5089 7361 5123 7395
rect 5123 7361 5132 7395
rect 5080 7352 5132 7361
rect 5908 7352 5960 7404
rect 7472 7420 7524 7472
rect 8668 7420 8720 7472
rect 11888 7488 11940 7540
rect 12164 7488 12216 7540
rect 15292 7488 15344 7540
rect 16580 7488 16632 7540
rect 17960 7531 18012 7540
rect 17960 7497 17969 7531
rect 17969 7497 18003 7531
rect 18003 7497 18012 7531
rect 17960 7488 18012 7497
rect 2412 7327 2464 7336
rect 2412 7293 2421 7327
rect 2421 7293 2455 7327
rect 2455 7293 2464 7327
rect 2412 7284 2464 7293
rect 2780 7327 2832 7336
rect 2780 7293 2789 7327
rect 2789 7293 2823 7327
rect 2823 7293 2832 7327
rect 3424 7327 3476 7336
rect 2780 7284 2832 7293
rect 3424 7293 3433 7327
rect 3433 7293 3467 7327
rect 3467 7293 3476 7327
rect 3424 7284 3476 7293
rect 5356 7284 5408 7336
rect 7932 7352 7984 7404
rect 8024 7395 8076 7404
rect 8024 7361 8053 7395
rect 8053 7361 8076 7395
rect 8944 7395 8996 7404
rect 8024 7352 8076 7361
rect 8944 7361 8953 7395
rect 8953 7361 8987 7395
rect 8987 7361 8996 7395
rect 8944 7352 8996 7361
rect 9128 7395 9180 7404
rect 9128 7361 9137 7395
rect 9137 7361 9171 7395
rect 9171 7361 9180 7395
rect 9128 7352 9180 7361
rect 9680 7352 9732 7404
rect 9956 7352 10008 7404
rect 10416 7395 10468 7404
rect 10416 7361 10425 7395
rect 10425 7361 10459 7395
rect 10459 7361 10468 7395
rect 10416 7352 10468 7361
rect 10508 7395 10560 7404
rect 10508 7361 10517 7395
rect 10517 7361 10551 7395
rect 10551 7361 10560 7395
rect 10508 7352 10560 7361
rect 9588 7327 9640 7336
rect 9588 7293 9597 7327
rect 9597 7293 9631 7327
rect 9631 7293 9640 7327
rect 9588 7284 9640 7293
rect 9864 7284 9916 7336
rect 10508 7216 10560 7268
rect 6552 7191 6604 7200
rect 6552 7157 6561 7191
rect 6561 7157 6595 7191
rect 6595 7157 6604 7191
rect 6552 7148 6604 7157
rect 9680 7148 9732 7200
rect 9864 7148 9916 7200
rect 10692 7191 10744 7200
rect 10692 7157 10701 7191
rect 10701 7157 10735 7191
rect 10735 7157 10744 7191
rect 10692 7148 10744 7157
rect 11060 7352 11112 7404
rect 11980 7352 12032 7404
rect 12256 7420 12308 7472
rect 13176 7420 13228 7472
rect 10876 7284 10928 7336
rect 12716 7284 12768 7336
rect 13452 7284 13504 7336
rect 13820 7352 13872 7404
rect 14096 7352 14148 7404
rect 15200 7352 15252 7404
rect 17224 7420 17276 7472
rect 17868 7420 17920 7472
rect 16212 7352 16264 7404
rect 16672 7352 16724 7404
rect 15476 7284 15528 7336
rect 13544 7259 13596 7268
rect 13084 7148 13136 7200
rect 13544 7225 13553 7259
rect 13553 7225 13587 7259
rect 13587 7225 13596 7259
rect 13544 7216 13596 7225
rect 15016 7259 15068 7268
rect 15016 7225 15025 7259
rect 15025 7225 15059 7259
rect 15059 7225 15068 7259
rect 15016 7216 15068 7225
rect 13728 7148 13780 7200
rect 14096 7191 14148 7200
rect 14096 7157 14105 7191
rect 14105 7157 14139 7191
rect 14139 7157 14148 7191
rect 14096 7148 14148 7157
rect 4214 7046 4266 7098
rect 4278 7046 4330 7098
rect 4342 7046 4394 7098
rect 4406 7046 4458 7098
rect 4470 7046 4522 7098
rect 12214 7046 12266 7098
rect 12278 7046 12330 7098
rect 12342 7046 12394 7098
rect 12406 7046 12458 7098
rect 12470 7046 12522 7098
rect 2780 6944 2832 6996
rect 9496 6944 9548 6996
rect 9864 6944 9916 6996
rect 2044 6876 2096 6928
rect 2688 6876 2740 6928
rect 4620 6876 4672 6928
rect 13268 6876 13320 6928
rect 17500 6876 17552 6928
rect 1676 6808 1728 6860
rect 3240 6808 3292 6860
rect 7472 6851 7524 6860
rect 7472 6817 7481 6851
rect 7481 6817 7515 6851
rect 7515 6817 7524 6851
rect 7472 6808 7524 6817
rect 1952 6783 2004 6792
rect 1952 6749 1961 6783
rect 1961 6749 1995 6783
rect 1995 6749 2004 6783
rect 1952 6740 2004 6749
rect 2412 6740 2464 6792
rect 3884 6740 3936 6792
rect 4712 6740 4764 6792
rect 5080 6740 5132 6792
rect 1584 6647 1636 6656
rect 1584 6613 1593 6647
rect 1593 6613 1627 6647
rect 1627 6613 1636 6647
rect 1584 6604 1636 6613
rect 2412 6647 2464 6656
rect 2412 6613 2421 6647
rect 2421 6613 2455 6647
rect 2455 6613 2464 6647
rect 2412 6604 2464 6613
rect 2780 6604 2832 6656
rect 4896 6672 4948 6724
rect 6920 6740 6972 6792
rect 8116 6740 8168 6792
rect 9680 6740 9732 6792
rect 10692 6808 10744 6860
rect 7012 6672 7064 6724
rect 8576 6672 8628 6724
rect 9128 6672 9180 6724
rect 10876 6740 10928 6792
rect 11060 6740 11112 6792
rect 11888 6783 11940 6792
rect 3884 6604 3936 6656
rect 11888 6749 11897 6783
rect 11897 6749 11931 6783
rect 11931 6749 11940 6783
rect 11888 6740 11940 6749
rect 12256 6740 12308 6792
rect 14096 6808 14148 6860
rect 15200 6851 15252 6860
rect 15200 6817 15209 6851
rect 15209 6817 15243 6851
rect 15243 6817 15252 6851
rect 15200 6808 15252 6817
rect 13544 6783 13596 6792
rect 13544 6749 13553 6783
rect 13553 6749 13587 6783
rect 13587 6749 13596 6783
rect 13544 6740 13596 6749
rect 13728 6740 13780 6792
rect 15292 6740 15344 6792
rect 15476 6740 15528 6792
rect 16120 6740 16172 6792
rect 17316 6808 17368 6860
rect 18052 6672 18104 6724
rect 18144 6715 18196 6724
rect 18144 6681 18153 6715
rect 18153 6681 18187 6715
rect 18187 6681 18196 6715
rect 18144 6672 18196 6681
rect 12164 6604 12216 6656
rect 12716 6604 12768 6656
rect 13084 6647 13136 6656
rect 13084 6613 13093 6647
rect 13093 6613 13127 6647
rect 13127 6613 13136 6647
rect 13084 6604 13136 6613
rect 15936 6647 15988 6656
rect 15936 6613 15945 6647
rect 15945 6613 15979 6647
rect 15979 6613 15988 6647
rect 15936 6604 15988 6613
rect 8214 6502 8266 6554
rect 8278 6502 8330 6554
rect 8342 6502 8394 6554
rect 8406 6502 8458 6554
rect 8470 6502 8522 6554
rect 16214 6502 16266 6554
rect 16278 6502 16330 6554
rect 16342 6502 16394 6554
rect 16406 6502 16458 6554
rect 16470 6502 16522 6554
rect 2688 6400 2740 6452
rect 2412 6332 2464 6384
rect 8576 6400 8628 6452
rect 9128 6443 9180 6452
rect 9128 6409 9137 6443
rect 9137 6409 9171 6443
rect 9171 6409 9180 6443
rect 9128 6400 9180 6409
rect 12164 6443 12216 6452
rect 12164 6409 12173 6443
rect 12173 6409 12207 6443
rect 12207 6409 12216 6443
rect 12164 6400 12216 6409
rect 16580 6400 16632 6452
rect 17040 6400 17092 6452
rect 3976 6375 4028 6384
rect 1952 6307 2004 6316
rect 1952 6273 1961 6307
rect 1961 6273 1995 6307
rect 1995 6273 2004 6307
rect 1952 6264 2004 6273
rect 2596 6307 2648 6316
rect 2596 6273 2605 6307
rect 2605 6273 2639 6307
rect 2639 6273 2648 6307
rect 2596 6264 2648 6273
rect 2780 6307 2832 6316
rect 2780 6273 2789 6307
rect 2789 6273 2823 6307
rect 2823 6273 2832 6307
rect 2780 6264 2832 6273
rect 3516 6307 3568 6316
rect 3516 6273 3525 6307
rect 3525 6273 3559 6307
rect 3559 6273 3568 6307
rect 3516 6264 3568 6273
rect 3976 6341 3985 6375
rect 3985 6341 4019 6375
rect 4019 6341 4028 6375
rect 3976 6332 4028 6341
rect 3700 6307 3752 6316
rect 3700 6273 3710 6307
rect 3710 6273 3744 6307
rect 3744 6273 3752 6307
rect 3700 6264 3752 6273
rect 4068 6264 4120 6316
rect 4620 6332 4672 6384
rect 4896 6332 4948 6384
rect 5448 6332 5500 6384
rect 2872 6196 2924 6248
rect 3884 6196 3936 6248
rect 5356 6307 5408 6316
rect 5356 6273 5365 6307
rect 5365 6273 5399 6307
rect 5399 6273 5408 6307
rect 6920 6332 6972 6384
rect 7472 6332 7524 6384
rect 5356 6264 5408 6273
rect 7012 6264 7064 6316
rect 3608 6128 3660 6180
rect 8484 6239 8536 6248
rect 8484 6205 8493 6239
rect 8493 6205 8527 6239
rect 8527 6205 8536 6239
rect 8484 6196 8536 6205
rect 8944 6196 8996 6248
rect 10508 6307 10560 6316
rect 10508 6273 10517 6307
rect 10517 6273 10551 6307
rect 10551 6273 10560 6307
rect 10508 6264 10560 6273
rect 10692 6307 10744 6316
rect 10692 6273 10701 6307
rect 10701 6273 10735 6307
rect 10735 6273 10744 6307
rect 10692 6264 10744 6273
rect 11060 6332 11112 6384
rect 12256 6375 12308 6384
rect 12256 6341 12265 6375
rect 12265 6341 12299 6375
rect 12299 6341 12308 6375
rect 12256 6332 12308 6341
rect 14832 6332 14884 6384
rect 15844 6332 15896 6384
rect 17132 6332 17184 6384
rect 15016 6307 15068 6316
rect 12808 6196 12860 6248
rect 9956 6128 10008 6180
rect 13268 6239 13320 6248
rect 13268 6205 13277 6239
rect 13277 6205 13311 6239
rect 13311 6205 13320 6239
rect 13268 6196 13320 6205
rect 14096 6196 14148 6248
rect 15016 6273 15025 6307
rect 15025 6273 15059 6307
rect 15059 6273 15068 6307
rect 15016 6264 15068 6273
rect 15936 6264 15988 6316
rect 18052 6307 18104 6316
rect 18052 6273 18061 6307
rect 18061 6273 18095 6307
rect 18095 6273 18104 6307
rect 18052 6264 18104 6273
rect 15292 6196 15344 6248
rect 17500 6128 17552 6180
rect 1584 6103 1636 6112
rect 1584 6069 1593 6103
rect 1593 6069 1627 6103
rect 1627 6069 1636 6103
rect 1584 6060 1636 6069
rect 2596 6060 2648 6112
rect 4988 6060 5040 6112
rect 5080 6060 5132 6112
rect 7288 6060 7340 6112
rect 9680 6060 9732 6112
rect 11520 6060 11572 6112
rect 14004 6060 14056 6112
rect 15292 6103 15344 6112
rect 15292 6069 15301 6103
rect 15301 6069 15335 6103
rect 15335 6069 15344 6103
rect 15292 6060 15344 6069
rect 4214 5958 4266 6010
rect 4278 5958 4330 6010
rect 4342 5958 4394 6010
rect 4406 5958 4458 6010
rect 4470 5958 4522 6010
rect 12214 5958 12266 6010
rect 12278 5958 12330 6010
rect 12342 5958 12394 6010
rect 12406 5958 12458 6010
rect 12470 5958 12522 6010
rect 2412 5856 2464 5908
rect 2504 5856 2556 5908
rect 3516 5856 3568 5908
rect 4068 5899 4120 5908
rect 4068 5865 4077 5899
rect 4077 5865 4111 5899
rect 4111 5865 4120 5899
rect 4068 5856 4120 5865
rect 4804 5856 4856 5908
rect 8484 5856 8536 5908
rect 8760 5856 8812 5908
rect 9588 5856 9640 5908
rect 16580 5856 16632 5908
rect 18144 5856 18196 5908
rect 2780 5788 2832 5840
rect 3884 5788 3936 5840
rect 2596 5720 2648 5772
rect 2504 5695 2556 5704
rect 2504 5661 2513 5695
rect 2513 5661 2547 5695
rect 2547 5661 2556 5695
rect 2504 5652 2556 5661
rect 2688 5695 2740 5704
rect 2688 5661 2697 5695
rect 2697 5661 2731 5695
rect 2731 5661 2740 5695
rect 2688 5652 2740 5661
rect 4712 5831 4764 5840
rect 4712 5797 4721 5831
rect 4721 5797 4755 5831
rect 4755 5797 4764 5831
rect 4712 5788 4764 5797
rect 6920 5788 6972 5840
rect 17500 5831 17552 5840
rect 17500 5797 17509 5831
rect 17509 5797 17543 5831
rect 17543 5797 17552 5831
rect 17500 5788 17552 5797
rect 17776 5788 17828 5840
rect 8116 5763 8168 5772
rect 8116 5729 8125 5763
rect 8125 5729 8159 5763
rect 8159 5729 8168 5763
rect 8116 5720 8168 5729
rect 5540 5695 5592 5704
rect 5540 5661 5549 5695
rect 5549 5661 5583 5695
rect 5583 5661 5592 5695
rect 5540 5652 5592 5661
rect 6368 5695 6420 5704
rect 2780 5516 2832 5568
rect 4344 5584 4396 5636
rect 4804 5584 4856 5636
rect 5264 5627 5316 5636
rect 5264 5593 5273 5627
rect 5273 5593 5307 5627
rect 5307 5593 5316 5627
rect 5264 5584 5316 5593
rect 5448 5584 5500 5636
rect 6368 5661 6377 5695
rect 6377 5661 6411 5695
rect 6411 5661 6420 5695
rect 6368 5652 6420 5661
rect 7472 5695 7524 5704
rect 7472 5661 7481 5695
rect 7481 5661 7515 5695
rect 7515 5661 7524 5695
rect 7472 5652 7524 5661
rect 8024 5652 8076 5704
rect 9496 5720 9548 5772
rect 9404 5584 9456 5636
rect 9588 5652 9640 5704
rect 9956 5695 10008 5704
rect 9956 5661 9965 5695
rect 9965 5661 9999 5695
rect 9999 5661 10008 5695
rect 9956 5652 10008 5661
rect 10600 5720 10652 5772
rect 15660 5720 15712 5772
rect 15844 5720 15896 5772
rect 11520 5695 11572 5704
rect 11520 5661 11529 5695
rect 11529 5661 11563 5695
rect 11563 5661 11572 5695
rect 11520 5652 11572 5661
rect 13912 5652 13964 5704
rect 14188 5695 14240 5704
rect 14188 5661 14197 5695
rect 14197 5661 14231 5695
rect 14231 5661 14240 5695
rect 14188 5652 14240 5661
rect 13728 5584 13780 5636
rect 14740 5652 14792 5704
rect 18052 5652 18104 5704
rect 4620 5516 4672 5568
rect 4712 5516 4764 5568
rect 5080 5559 5132 5568
rect 5080 5525 5089 5559
rect 5089 5525 5123 5559
rect 5123 5525 5132 5559
rect 5080 5516 5132 5525
rect 6736 5516 6788 5568
rect 7012 5516 7064 5568
rect 7932 5516 7984 5568
rect 11336 5559 11388 5568
rect 11336 5525 11345 5559
rect 11345 5525 11379 5559
rect 11379 5525 11388 5559
rect 11336 5516 11388 5525
rect 17592 5627 17644 5636
rect 17592 5593 17601 5627
rect 17601 5593 17635 5627
rect 17635 5593 17644 5627
rect 17592 5584 17644 5593
rect 16028 5516 16080 5568
rect 8214 5414 8266 5466
rect 8278 5414 8330 5466
rect 8342 5414 8394 5466
rect 8406 5414 8458 5466
rect 8470 5414 8522 5466
rect 16214 5414 16266 5466
rect 16278 5414 16330 5466
rect 16342 5414 16394 5466
rect 16406 5414 16458 5466
rect 16470 5414 16522 5466
rect 3700 5312 3752 5364
rect 2780 5244 2832 5296
rect 4620 5312 4672 5364
rect 5264 5312 5316 5364
rect 8760 5355 8812 5364
rect 8760 5321 8769 5355
rect 8769 5321 8803 5355
rect 8803 5321 8812 5355
rect 8760 5312 8812 5321
rect 10416 5312 10468 5364
rect 12808 5312 12860 5364
rect 14832 5312 14884 5364
rect 15752 5312 15804 5364
rect 16580 5312 16632 5364
rect 17316 5355 17368 5364
rect 5448 5244 5500 5296
rect 7288 5287 7340 5296
rect 7288 5253 7297 5287
rect 7297 5253 7331 5287
rect 7331 5253 7340 5287
rect 7288 5244 7340 5253
rect 9128 5244 9180 5296
rect 9680 5244 9732 5296
rect 10140 5244 10192 5296
rect 11336 5244 11388 5296
rect 12624 5244 12676 5296
rect 14004 5287 14056 5296
rect 14004 5253 14013 5287
rect 14013 5253 14047 5287
rect 14047 5253 14056 5287
rect 14004 5244 14056 5253
rect 14464 5244 14516 5296
rect 17316 5321 17325 5355
rect 17325 5321 17359 5355
rect 17359 5321 17368 5355
rect 17316 5312 17368 5321
rect 17224 5244 17276 5296
rect 17592 5244 17644 5296
rect 3240 5176 3292 5228
rect 4160 5219 4212 5228
rect 4160 5185 4169 5219
rect 4169 5185 4203 5219
rect 4203 5185 4212 5219
rect 4160 5176 4212 5185
rect 4344 5176 4396 5228
rect 4620 5176 4672 5228
rect 4896 5176 4948 5228
rect 6920 5176 6972 5228
rect 4160 5040 4212 5092
rect 4712 5040 4764 5092
rect 4804 5040 4856 5092
rect 5080 5108 5132 5160
rect 6184 5108 6236 5160
rect 9772 5108 9824 5160
rect 11980 5108 12032 5160
rect 14740 5108 14792 5160
rect 17684 5108 17736 5160
rect 2412 4972 2464 5024
rect 4068 4972 4120 5024
rect 6460 4972 6512 5024
rect 4214 4870 4266 4922
rect 4278 4870 4330 4922
rect 4342 4870 4394 4922
rect 4406 4870 4458 4922
rect 4470 4870 4522 4922
rect 12214 4870 12266 4922
rect 12278 4870 12330 4922
rect 12342 4870 12394 4922
rect 12406 4870 12458 4922
rect 12470 4870 12522 4922
rect 2504 4811 2556 4820
rect 2504 4777 2513 4811
rect 2513 4777 2547 4811
rect 2547 4777 2556 4811
rect 2504 4768 2556 4777
rect 2964 4811 3016 4820
rect 2964 4777 2973 4811
rect 2973 4777 3007 4811
rect 3007 4777 3016 4811
rect 2964 4768 3016 4777
rect 4712 4768 4764 4820
rect 5080 4768 5132 4820
rect 1768 4632 1820 4684
rect 4068 4632 4120 4684
rect 2136 4564 2188 4616
rect 2596 4607 2648 4616
rect 2596 4573 2605 4607
rect 2605 4573 2639 4607
rect 2639 4573 2648 4607
rect 2596 4564 2648 4573
rect 4252 4607 4304 4616
rect 4252 4573 4261 4607
rect 4261 4573 4295 4607
rect 4295 4573 4304 4607
rect 4252 4564 4304 4573
rect 5540 4632 5592 4684
rect 6552 4768 6604 4820
rect 7932 4811 7984 4820
rect 7932 4777 7941 4811
rect 7941 4777 7975 4811
rect 7975 4777 7984 4811
rect 7932 4768 7984 4777
rect 13544 4768 13596 4820
rect 10140 4743 10192 4752
rect 10140 4709 10149 4743
rect 10149 4709 10183 4743
rect 10183 4709 10192 4743
rect 10140 4700 10192 4709
rect 6460 4675 6512 4684
rect 6460 4641 6469 4675
rect 6469 4641 6503 4675
rect 6503 4641 6512 4675
rect 6460 4632 6512 4641
rect 7840 4632 7892 4684
rect 4896 4607 4948 4616
rect 4896 4573 4905 4607
rect 4905 4573 4939 4607
rect 4939 4573 4948 4607
rect 4896 4564 4948 4573
rect 5080 4607 5132 4616
rect 5080 4573 5089 4607
rect 5089 4573 5123 4607
rect 5123 4573 5132 4607
rect 5080 4564 5132 4573
rect 4528 4496 4580 4548
rect 6000 4564 6052 4616
rect 6184 4607 6236 4616
rect 6184 4573 6193 4607
rect 6193 4573 6227 4607
rect 6227 4573 6236 4607
rect 6184 4564 6236 4573
rect 9128 4632 9180 4684
rect 9312 4607 9364 4616
rect 1860 4428 1912 4480
rect 3332 4471 3384 4480
rect 3332 4437 3341 4471
rect 3341 4437 3375 4471
rect 3375 4437 3384 4471
rect 3332 4428 3384 4437
rect 4252 4428 4304 4480
rect 4712 4428 4764 4480
rect 4988 4428 5040 4480
rect 8576 4428 8628 4480
rect 9312 4573 9321 4607
rect 9321 4573 9355 4607
rect 9355 4573 9364 4607
rect 9312 4564 9364 4573
rect 11980 4632 12032 4684
rect 13820 4768 13872 4820
rect 16120 4768 16172 4820
rect 14464 4700 14516 4752
rect 14740 4675 14792 4684
rect 10876 4496 10928 4548
rect 11980 4496 12032 4548
rect 12716 4539 12768 4548
rect 12716 4505 12725 4539
rect 12725 4505 12759 4539
rect 12759 4505 12768 4539
rect 12716 4496 12768 4505
rect 14740 4641 14749 4675
rect 14749 4641 14783 4675
rect 14783 4641 14792 4675
rect 14740 4632 14792 4641
rect 16856 4632 16908 4684
rect 13728 4607 13780 4616
rect 13728 4573 13737 4607
rect 13737 4573 13771 4607
rect 13771 4573 13780 4607
rect 13728 4564 13780 4573
rect 13912 4564 13964 4616
rect 17132 4607 17184 4616
rect 17132 4573 17141 4607
rect 17141 4573 17175 4607
rect 17175 4573 17184 4607
rect 17132 4564 17184 4573
rect 17224 4607 17276 4616
rect 17224 4573 17233 4607
rect 17233 4573 17267 4607
rect 17267 4573 17276 4607
rect 17224 4564 17276 4573
rect 18052 4607 18104 4616
rect 15292 4496 15344 4548
rect 15476 4496 15528 4548
rect 16948 4539 17000 4548
rect 16948 4505 16957 4539
rect 16957 4505 16991 4539
rect 16991 4505 17000 4539
rect 16948 4496 17000 4505
rect 17040 4496 17092 4548
rect 18052 4573 18061 4607
rect 18061 4573 18095 4607
rect 18095 4573 18104 4607
rect 18052 4564 18104 4573
rect 16028 4428 16080 4480
rect 8214 4326 8266 4378
rect 8278 4326 8330 4378
rect 8342 4326 8394 4378
rect 8406 4326 8458 4378
rect 8470 4326 8522 4378
rect 16214 4326 16266 4378
rect 16278 4326 16330 4378
rect 16342 4326 16394 4378
rect 16406 4326 16458 4378
rect 16470 4326 16522 4378
rect 2504 4224 2556 4276
rect 4896 4224 4948 4276
rect 11980 4267 12032 4276
rect 11980 4233 11989 4267
rect 11989 4233 12023 4267
rect 12023 4233 12032 4267
rect 11980 4224 12032 4233
rect 12624 4267 12676 4276
rect 12624 4233 12633 4267
rect 12633 4233 12667 4267
rect 12667 4233 12676 4267
rect 12624 4224 12676 4233
rect 15476 4224 15528 4276
rect 17040 4224 17092 4276
rect 17224 4224 17276 4276
rect 1676 4199 1728 4208
rect 1676 4165 1685 4199
rect 1685 4165 1719 4199
rect 1719 4165 1728 4199
rect 1676 4156 1728 4165
rect 4988 4156 5040 4208
rect 7472 4156 7524 4208
rect 9312 4156 9364 4208
rect 1860 4131 1912 4140
rect 1860 4097 1869 4131
rect 1869 4097 1903 4131
rect 1903 4097 1912 4131
rect 1860 4088 1912 4097
rect 2228 4088 2280 4140
rect 2412 4131 2464 4140
rect 2412 4097 2421 4131
rect 2421 4097 2455 4131
rect 2455 4097 2464 4131
rect 2412 4088 2464 4097
rect 5632 4131 5684 4140
rect 5632 4097 5641 4131
rect 5641 4097 5675 4131
rect 5675 4097 5684 4131
rect 5632 4088 5684 4097
rect 5816 4131 5868 4140
rect 5816 4097 5825 4131
rect 5825 4097 5859 4131
rect 5859 4097 5868 4131
rect 5816 4088 5868 4097
rect 8576 4131 8628 4140
rect 8576 4097 8585 4131
rect 8585 4097 8619 4131
rect 8619 4097 8628 4131
rect 8576 4088 8628 4097
rect 9864 4131 9916 4140
rect 9864 4097 9873 4131
rect 9873 4097 9907 4131
rect 9907 4097 9916 4131
rect 9864 4088 9916 4097
rect 10416 4088 10468 4140
rect 10600 4131 10652 4140
rect 10600 4097 10609 4131
rect 10609 4097 10643 4131
rect 10643 4097 10652 4131
rect 10600 4088 10652 4097
rect 12440 4131 12492 4140
rect 3332 4020 3384 4072
rect 5172 4063 5224 4072
rect 4528 3952 4580 4004
rect 5172 4029 5181 4063
rect 5181 4029 5215 4063
rect 5215 4029 5224 4063
rect 5172 4020 5224 4029
rect 5540 4063 5592 4072
rect 5540 4029 5549 4063
rect 5549 4029 5583 4063
rect 5583 4029 5592 4063
rect 5540 4020 5592 4029
rect 5724 4020 5776 4072
rect 6184 4020 6236 4072
rect 6736 4063 6788 4072
rect 6736 4029 6745 4063
rect 6745 4029 6779 4063
rect 6779 4029 6788 4063
rect 6736 4020 6788 4029
rect 7748 4020 7800 4072
rect 9680 4063 9732 4072
rect 5080 3952 5132 4004
rect 8484 3952 8536 4004
rect 9312 3995 9364 4004
rect 9312 3961 9321 3995
rect 9321 3961 9355 3995
rect 9355 3961 9364 3995
rect 9312 3952 9364 3961
rect 9680 4029 9689 4063
rect 9689 4029 9723 4063
rect 9723 4029 9732 4063
rect 9680 4020 9732 4029
rect 10784 4063 10836 4072
rect 10784 4029 10793 4063
rect 10793 4029 10827 4063
rect 10827 4029 10836 4063
rect 10784 4020 10836 4029
rect 10876 4020 10928 4072
rect 12440 4097 12449 4131
rect 12449 4097 12483 4131
rect 12483 4097 12492 4131
rect 13728 4156 13780 4208
rect 16672 4156 16724 4208
rect 17132 4156 17184 4208
rect 17960 4199 18012 4208
rect 12440 4088 12492 4097
rect 12992 4063 13044 4072
rect 12992 4029 13001 4063
rect 13001 4029 13035 4063
rect 13035 4029 13044 4063
rect 12992 4020 13044 4029
rect 13820 4088 13872 4140
rect 14096 4088 14148 4140
rect 17684 4131 17736 4140
rect 14372 4020 14424 4072
rect 14556 4063 14608 4072
rect 14556 4029 14565 4063
rect 14565 4029 14599 4063
rect 14599 4029 14608 4063
rect 14556 4020 14608 4029
rect 16580 4020 16632 4072
rect 17684 4097 17693 4131
rect 17693 4097 17727 4131
rect 17727 4097 17736 4131
rect 17684 4088 17736 4097
rect 17960 4165 17969 4199
rect 17969 4165 18003 4199
rect 18003 4165 18012 4199
rect 17960 4156 18012 4165
rect 18236 4131 18288 4140
rect 18236 4097 18245 4131
rect 18245 4097 18279 4131
rect 18279 4097 18288 4131
rect 18236 4088 18288 4097
rect 16120 3952 16172 4004
rect 17132 3952 17184 4004
rect 18328 4020 18380 4072
rect 6460 3884 6512 3936
rect 6736 3884 6788 3936
rect 9220 3884 9272 3936
rect 10416 3927 10468 3936
rect 10416 3893 10425 3927
rect 10425 3893 10459 3927
rect 10459 3893 10468 3927
rect 10416 3884 10468 3893
rect 12440 3884 12492 3936
rect 14188 3884 14240 3936
rect 16764 3884 16816 3936
rect 17500 3884 17552 3936
rect 4214 3782 4266 3834
rect 4278 3782 4330 3834
rect 4342 3782 4394 3834
rect 4406 3782 4458 3834
rect 4470 3782 4522 3834
rect 12214 3782 12266 3834
rect 12278 3782 12330 3834
rect 12342 3782 12394 3834
rect 12406 3782 12458 3834
rect 12470 3782 12522 3834
rect 3148 3680 3200 3732
rect 6368 3680 6420 3732
rect 6460 3680 6512 3732
rect 10784 3680 10836 3732
rect 4620 3612 4672 3664
rect 9404 3612 9456 3664
rect 1860 3544 1912 3596
rect 2228 3544 2280 3596
rect 3884 3587 3936 3596
rect 3884 3553 3893 3587
rect 3893 3553 3927 3587
rect 3927 3553 3936 3587
rect 3884 3544 3936 3553
rect 5172 3544 5224 3596
rect 5448 3544 5500 3596
rect 7472 3587 7524 3596
rect 7472 3553 7481 3587
rect 7481 3553 7515 3587
rect 7515 3553 7524 3587
rect 7472 3544 7524 3553
rect 8576 3544 8628 3596
rect 1768 3476 1820 3528
rect 3240 3476 3292 3528
rect 4620 3519 4672 3528
rect 4620 3485 4629 3519
rect 4629 3485 4663 3519
rect 4663 3485 4672 3519
rect 4620 3476 4672 3485
rect 5540 3476 5592 3528
rect 6644 3519 6696 3528
rect 6644 3485 6653 3519
rect 6653 3485 6687 3519
rect 6687 3485 6696 3519
rect 6644 3476 6696 3485
rect 7104 3519 7156 3528
rect 7104 3485 7113 3519
rect 7113 3485 7147 3519
rect 7147 3485 7156 3519
rect 7104 3476 7156 3485
rect 7656 3519 7708 3528
rect 7656 3485 7665 3519
rect 7665 3485 7699 3519
rect 7699 3485 7708 3519
rect 7656 3476 7708 3485
rect 7840 3519 7892 3528
rect 7840 3485 7849 3519
rect 7849 3485 7883 3519
rect 7883 3485 7892 3519
rect 7840 3476 7892 3485
rect 8484 3519 8536 3528
rect 8484 3485 8493 3519
rect 8493 3485 8527 3519
rect 8527 3485 8536 3519
rect 8484 3476 8536 3485
rect 8668 3519 8720 3528
rect 8668 3485 8677 3519
rect 8677 3485 8711 3519
rect 8711 3485 8720 3519
rect 8668 3476 8720 3485
rect 2596 3451 2648 3460
rect 2596 3417 2605 3451
rect 2605 3417 2639 3451
rect 2639 3417 2648 3451
rect 2596 3408 2648 3417
rect 2780 3408 2832 3460
rect 8024 3408 8076 3460
rect 9404 3476 9456 3528
rect 9864 3476 9916 3528
rect 10416 3476 10468 3528
rect 10692 3519 10744 3528
rect 10692 3485 10701 3519
rect 10701 3485 10735 3519
rect 10735 3485 10744 3519
rect 10692 3476 10744 3485
rect 11520 3544 11572 3596
rect 16856 3544 16908 3596
rect 18236 3680 18288 3732
rect 18052 3544 18104 3596
rect 1768 3383 1820 3392
rect 1768 3349 1777 3383
rect 1777 3349 1811 3383
rect 1811 3349 1820 3383
rect 1768 3340 1820 3349
rect 2504 3383 2556 3392
rect 2504 3349 2513 3383
rect 2513 3349 2547 3383
rect 2547 3349 2556 3383
rect 2504 3340 2556 3349
rect 2872 3340 2924 3392
rect 5908 3340 5960 3392
rect 8760 3340 8812 3392
rect 9496 3383 9548 3392
rect 9496 3349 9505 3383
rect 9505 3349 9539 3383
rect 9539 3349 9548 3383
rect 9496 3340 9548 3349
rect 10600 3340 10652 3392
rect 12992 3476 13044 3528
rect 14188 3519 14240 3528
rect 14188 3485 14197 3519
rect 14197 3485 14231 3519
rect 14231 3485 14240 3519
rect 14188 3476 14240 3485
rect 14372 3519 14424 3528
rect 14372 3485 14381 3519
rect 14381 3485 14415 3519
rect 14415 3485 14424 3519
rect 14372 3476 14424 3485
rect 14556 3476 14608 3528
rect 18328 3476 18380 3528
rect 15660 3408 15712 3460
rect 16948 3408 17000 3460
rect 14280 3383 14332 3392
rect 14280 3349 14289 3383
rect 14289 3349 14323 3383
rect 14323 3349 14332 3383
rect 14280 3340 14332 3349
rect 17224 3340 17276 3392
rect 17776 3340 17828 3392
rect 8214 3238 8266 3290
rect 8278 3238 8330 3290
rect 8342 3238 8394 3290
rect 8406 3238 8458 3290
rect 8470 3238 8522 3290
rect 16214 3238 16266 3290
rect 16278 3238 16330 3290
rect 16342 3238 16394 3290
rect 16406 3238 16458 3290
rect 16470 3238 16522 3290
rect 2228 3136 2280 3188
rect 2688 3179 2740 3188
rect 2688 3145 2697 3179
rect 2697 3145 2731 3179
rect 2731 3145 2740 3179
rect 2688 3136 2740 3145
rect 4068 3136 4120 3188
rect 4804 3179 4856 3188
rect 4804 3145 4813 3179
rect 4813 3145 4847 3179
rect 4847 3145 4856 3179
rect 4804 3136 4856 3145
rect 5816 3179 5868 3188
rect 5816 3145 5825 3179
rect 5825 3145 5859 3179
rect 5859 3145 5868 3179
rect 5816 3136 5868 3145
rect 7380 3136 7432 3188
rect 7748 3136 7800 3188
rect 8024 3179 8076 3188
rect 8024 3145 8033 3179
rect 8033 3145 8067 3179
rect 8067 3145 8076 3179
rect 8024 3136 8076 3145
rect 9220 3136 9272 3188
rect 1768 3043 1820 3052
rect 1768 3009 1777 3043
rect 1777 3009 1811 3043
rect 1811 3009 1820 3043
rect 1768 3000 1820 3009
rect 2136 3000 2188 3052
rect 4988 3043 5040 3052
rect 4988 3009 4997 3043
rect 4997 3009 5031 3043
rect 5031 3009 5040 3043
rect 4988 3000 5040 3009
rect 4160 2932 4212 2984
rect 5356 3043 5408 3052
rect 5356 3009 5365 3043
rect 5365 3009 5399 3043
rect 5399 3009 5408 3043
rect 5356 3000 5408 3009
rect 5908 3000 5960 3052
rect 8760 3068 8812 3120
rect 9496 3111 9548 3120
rect 9496 3077 9505 3111
rect 9505 3077 9539 3111
rect 9539 3077 9548 3111
rect 9496 3068 9548 3077
rect 11520 3068 11572 3120
rect 16120 3136 16172 3188
rect 17868 3179 17920 3188
rect 17868 3145 17877 3179
rect 17877 3145 17911 3179
rect 17911 3145 17920 3179
rect 17868 3136 17920 3145
rect 18052 3136 18104 3188
rect 5632 2932 5684 2984
rect 6736 3043 6788 3052
rect 6736 3009 6745 3043
rect 6745 3009 6779 3043
rect 6779 3009 6788 3043
rect 7656 3043 7708 3052
rect 6736 3000 6788 3009
rect 7656 3009 7665 3043
rect 7665 3009 7699 3043
rect 7699 3009 7708 3043
rect 7656 3000 7708 3009
rect 9772 3043 9824 3052
rect 9772 3009 9781 3043
rect 9781 3009 9815 3043
rect 9815 3009 9824 3043
rect 9772 3000 9824 3009
rect 10508 3000 10560 3052
rect 11612 3043 11664 3052
rect 11612 3009 11621 3043
rect 11621 3009 11655 3043
rect 11655 3009 11664 3043
rect 11612 3000 11664 3009
rect 11796 3043 11848 3052
rect 11796 3009 11805 3043
rect 11805 3009 11839 3043
rect 11839 3009 11848 3043
rect 11796 3000 11848 3009
rect 7104 2932 7156 2984
rect 2412 2864 2464 2916
rect 3332 2864 3384 2916
rect 5724 2864 5776 2916
rect 10232 2932 10284 2984
rect 11152 2975 11204 2984
rect 11152 2941 11161 2975
rect 11161 2941 11195 2975
rect 11195 2941 11204 2975
rect 11152 2932 11204 2941
rect 13820 3000 13872 3052
rect 17408 3068 17460 3120
rect 17224 3043 17276 3052
rect 17224 3009 17233 3043
rect 17233 3009 17267 3043
rect 17267 3009 17276 3043
rect 17224 3000 17276 3009
rect 14556 2975 14608 2984
rect 11060 2907 11112 2916
rect 11060 2873 11069 2907
rect 11069 2873 11103 2907
rect 11103 2873 11112 2907
rect 11060 2864 11112 2873
rect 8760 2796 8812 2848
rect 14556 2941 14565 2975
rect 14565 2941 14599 2975
rect 14599 2941 14608 2975
rect 14556 2932 14608 2941
rect 17500 2932 17552 2984
rect 17776 2975 17828 2984
rect 17776 2941 17785 2975
rect 17785 2941 17819 2975
rect 17819 2941 17828 2975
rect 17776 2932 17828 2941
rect 18236 2975 18288 2984
rect 18236 2941 18245 2975
rect 18245 2941 18279 2975
rect 18279 2941 18288 2975
rect 18236 2932 18288 2941
rect 12624 2864 12676 2916
rect 13360 2907 13412 2916
rect 13360 2873 13369 2907
rect 13369 2873 13403 2907
rect 13403 2873 13412 2907
rect 13360 2864 13412 2873
rect 11888 2796 11940 2848
rect 17040 2839 17092 2848
rect 17040 2805 17049 2839
rect 17049 2805 17083 2839
rect 17083 2805 17092 2839
rect 17040 2796 17092 2805
rect 4214 2694 4266 2746
rect 4278 2694 4330 2746
rect 4342 2694 4394 2746
rect 4406 2694 4458 2746
rect 4470 2694 4522 2746
rect 12214 2694 12266 2746
rect 12278 2694 12330 2746
rect 12342 2694 12394 2746
rect 12406 2694 12458 2746
rect 12470 2694 12522 2746
rect 2504 2635 2556 2644
rect 2504 2601 2513 2635
rect 2513 2601 2547 2635
rect 2547 2601 2556 2635
rect 2504 2592 2556 2601
rect 5356 2592 5408 2644
rect 3240 2567 3292 2576
rect 3240 2533 3249 2567
rect 3249 2533 3283 2567
rect 3283 2533 3292 2567
rect 3240 2524 3292 2533
rect 4620 2524 4672 2576
rect 2044 2388 2096 2440
rect 2872 2456 2924 2508
rect 5724 2499 5776 2508
rect 5724 2465 5733 2499
rect 5733 2465 5767 2499
rect 5767 2465 5776 2499
rect 5724 2456 5776 2465
rect 2780 2431 2832 2440
rect 2780 2397 2789 2431
rect 2789 2397 2823 2431
rect 2823 2397 2832 2431
rect 2780 2388 2832 2397
rect 3148 2388 3200 2440
rect 2872 2320 2924 2372
rect 3608 2252 3660 2304
rect 4160 2431 4212 2440
rect 4160 2397 4169 2431
rect 4169 2397 4203 2431
rect 4203 2397 4212 2431
rect 4160 2388 4212 2397
rect 5264 2431 5316 2440
rect 5264 2397 5273 2431
rect 5273 2397 5307 2431
rect 5307 2397 5316 2431
rect 5264 2388 5316 2397
rect 4988 2320 5040 2372
rect 4804 2252 4856 2304
rect 7564 2388 7616 2440
rect 10508 2592 10560 2644
rect 11796 2592 11848 2644
rect 11152 2524 11204 2576
rect 14188 2592 14240 2644
rect 17592 2567 17644 2576
rect 17592 2533 17601 2567
rect 17601 2533 17635 2567
rect 17635 2533 17644 2567
rect 17592 2524 17644 2533
rect 6000 2363 6052 2372
rect 6000 2329 6009 2363
rect 6009 2329 6043 2363
rect 6043 2329 6052 2363
rect 6000 2320 6052 2329
rect 6460 2320 6512 2372
rect 7748 2320 7800 2372
rect 8668 2388 8720 2440
rect 9220 2388 9272 2440
rect 10600 2456 10652 2508
rect 11612 2456 11664 2508
rect 14556 2456 14608 2508
rect 17040 2456 17092 2508
rect 17960 2456 18012 2508
rect 11060 2388 11112 2440
rect 13360 2388 13412 2440
rect 13912 2388 13964 2440
rect 11152 2320 11204 2372
rect 8576 2252 8628 2304
rect 9220 2295 9272 2304
rect 9220 2261 9229 2295
rect 9229 2261 9263 2295
rect 9263 2261 9272 2295
rect 9220 2252 9272 2261
rect 10232 2295 10284 2304
rect 10232 2261 10241 2295
rect 10241 2261 10275 2295
rect 10275 2261 10284 2295
rect 10232 2252 10284 2261
rect 11060 2252 11112 2304
rect 11980 2320 12032 2372
rect 14924 2252 14976 2304
rect 17776 2252 17828 2304
rect 17960 2320 18012 2372
rect 18328 2320 18380 2372
rect 8214 2150 8266 2202
rect 8278 2150 8330 2202
rect 8342 2150 8394 2202
rect 8406 2150 8458 2202
rect 8470 2150 8522 2202
rect 16214 2150 16266 2202
rect 16278 2150 16330 2202
rect 16342 2150 16394 2202
rect 16406 2150 16458 2202
rect 16470 2150 16522 2202
rect 2044 1980 2096 2032
rect 3148 2048 3200 2100
rect 4620 2048 4672 2100
rect 5264 2048 5316 2100
rect 6460 2048 6512 2100
rect 6644 2048 6696 2100
rect 8576 2048 8628 2100
rect 2596 1980 2648 2032
rect 3240 1980 3292 2032
rect 3608 2023 3660 2032
rect 3608 1989 3617 2023
rect 3617 1989 3651 2023
rect 3651 1989 3660 2023
rect 3608 1980 3660 1989
rect 5172 1980 5224 2032
rect 3332 1955 3384 1964
rect 3332 1921 3341 1955
rect 3341 1921 3375 1955
rect 3375 1921 3384 1955
rect 3332 1912 3384 1921
rect 5908 1912 5960 1964
rect 7380 1980 7432 2032
rect 9220 1980 9272 2032
rect 2780 1844 2832 1896
rect 4160 1844 4212 1896
rect 5356 1844 5408 1896
rect 6736 1912 6788 1964
rect 7564 1912 7616 1964
rect 11612 1980 11664 2032
rect 12624 1980 12676 2032
rect 4988 1776 5040 1828
rect 7748 1887 7800 1896
rect 7748 1853 7757 1887
rect 7757 1853 7791 1887
rect 7791 1853 7800 1887
rect 7748 1844 7800 1853
rect 9404 1844 9456 1896
rect 10692 1912 10744 1964
rect 11060 1955 11112 1964
rect 11060 1921 11069 1955
rect 11069 1921 11103 1955
rect 11103 1921 11112 1955
rect 11060 1912 11112 1921
rect 14556 2048 14608 2100
rect 14280 1980 14332 2032
rect 18236 2048 18288 2100
rect 15660 1912 15712 1964
rect 16948 1980 17000 2032
rect 16120 1955 16172 1964
rect 16120 1921 16129 1955
rect 16129 1921 16163 1955
rect 16163 1921 16172 1955
rect 16120 1912 16172 1921
rect 16764 1912 16816 1964
rect 11152 1887 11204 1896
rect 11152 1853 11161 1887
rect 11161 1853 11195 1887
rect 11195 1853 11204 1887
rect 11152 1844 11204 1853
rect 4804 1708 4856 1760
rect 9220 1708 9272 1760
rect 14924 1844 14976 1896
rect 16580 1844 16632 1896
rect 15936 1819 15988 1828
rect 15936 1785 15945 1819
rect 15945 1785 15979 1819
rect 15979 1785 15988 1819
rect 15936 1776 15988 1785
rect 10508 1708 10560 1760
rect 14832 1708 14884 1760
rect 4214 1606 4266 1658
rect 4278 1606 4330 1658
rect 4342 1606 4394 1658
rect 4406 1606 4458 1658
rect 4470 1606 4522 1658
rect 12214 1606 12266 1658
rect 12278 1606 12330 1658
rect 12342 1606 12394 1658
rect 12406 1606 12458 1658
rect 12470 1606 12522 1658
rect 2872 1504 2924 1556
rect 6000 1504 6052 1556
rect 11980 1504 12032 1556
rect 1492 1411 1544 1420
rect 1492 1377 1501 1411
rect 1501 1377 1535 1411
rect 1535 1377 1544 1411
rect 1492 1368 1544 1377
rect 4804 1368 4856 1420
rect 3332 1300 3384 1352
rect 4528 1275 4580 1284
rect 4528 1241 4537 1275
rect 4537 1241 4571 1275
rect 4571 1241 4580 1275
rect 4528 1232 4580 1241
rect 7748 1368 7800 1420
rect 9404 1411 9456 1420
rect 9404 1377 9413 1411
rect 9413 1377 9447 1411
rect 9447 1377 9456 1411
rect 9404 1368 9456 1377
rect 5172 1343 5224 1352
rect 5172 1309 5181 1343
rect 5181 1309 5215 1343
rect 5215 1309 5224 1343
rect 5172 1300 5224 1309
rect 5356 1343 5408 1352
rect 5356 1309 5365 1343
rect 5365 1309 5399 1343
rect 5399 1309 5408 1343
rect 5356 1300 5408 1309
rect 5908 1300 5960 1352
rect 8576 1300 8628 1352
rect 9220 1343 9272 1352
rect 7472 1275 7524 1284
rect 4620 1164 4672 1216
rect 6460 1207 6512 1216
rect 6460 1173 6469 1207
rect 6469 1173 6503 1207
rect 6503 1173 6512 1207
rect 6460 1164 6512 1173
rect 7472 1241 7481 1275
rect 7481 1241 7515 1275
rect 7515 1241 7524 1275
rect 7472 1232 7524 1241
rect 7564 1275 7616 1284
rect 7564 1241 7573 1275
rect 7573 1241 7607 1275
rect 7607 1241 7616 1275
rect 9220 1309 9229 1343
rect 9229 1309 9263 1343
rect 9263 1309 9272 1343
rect 9220 1300 9272 1309
rect 10232 1368 10284 1420
rect 11152 1411 11204 1420
rect 11152 1377 11161 1411
rect 11161 1377 11195 1411
rect 11195 1377 11204 1411
rect 11152 1368 11204 1377
rect 14556 1411 14608 1420
rect 14556 1377 14565 1411
rect 14565 1377 14599 1411
rect 14599 1377 14608 1411
rect 14556 1368 14608 1377
rect 14832 1411 14884 1420
rect 14832 1377 14841 1411
rect 14841 1377 14875 1411
rect 14875 1377 14884 1411
rect 14832 1368 14884 1377
rect 16120 1368 16172 1420
rect 9680 1300 9732 1352
rect 10508 1343 10560 1352
rect 10508 1309 10517 1343
rect 10517 1309 10551 1343
rect 10551 1309 10560 1343
rect 10508 1300 10560 1309
rect 11888 1300 11940 1352
rect 15936 1300 15988 1352
rect 16948 1343 17000 1352
rect 16948 1309 16957 1343
rect 16957 1309 16991 1343
rect 16991 1309 17000 1343
rect 16948 1300 17000 1309
rect 17592 1343 17644 1352
rect 17592 1309 17601 1343
rect 17601 1309 17635 1343
rect 17635 1309 17644 1343
rect 17592 1300 17644 1309
rect 18236 1300 18288 1352
rect 7564 1232 7616 1241
rect 11060 1232 11112 1284
rect 16580 1164 16632 1216
rect 16672 1164 16724 1216
rect 17500 1164 17552 1216
rect 18328 1207 18380 1216
rect 18328 1173 18337 1207
rect 18337 1173 18371 1207
rect 18371 1173 18380 1207
rect 18328 1164 18380 1173
rect 8214 1062 8266 1114
rect 8278 1062 8330 1114
rect 8342 1062 8394 1114
rect 8406 1062 8458 1114
rect 8470 1062 8522 1114
rect 16214 1062 16266 1114
rect 16278 1062 16330 1114
rect 16342 1062 16394 1114
rect 16406 1062 16458 1114
rect 16470 1062 16522 1114
rect 2780 960 2832 1012
rect 6460 960 6512 1012
rect 4528 892 4580 944
rect 5448 892 5500 944
rect 7564 892 7616 944
rect 18328 892 18380 944
<< metal2 >>
rect 1122 14362 1178 15000
rect 1122 14334 1348 14362
rect 1122 14200 1178 14334
rect 1320 13530 1348 14334
rect 2594 14200 2650 15000
rect 4066 14362 4122 15000
rect 3804 14334 4122 14362
rect 1308 13524 1360 13530
rect 1308 13466 1360 13472
rect 2228 13184 2280 13190
rect 2228 13126 2280 13132
rect 2320 13184 2372 13190
rect 2320 13126 2372 13132
rect 2240 12918 2268 13126
rect 2228 12912 2280 12918
rect 2228 12854 2280 12860
rect 1768 12640 1820 12646
rect 1768 12582 1820 12588
rect 1780 12306 1808 12582
rect 2240 12374 2268 12854
rect 2228 12368 2280 12374
rect 2228 12310 2280 12316
rect 1768 12300 1820 12306
rect 1768 12242 1820 12248
rect 2228 12164 2280 12170
rect 2228 12106 2280 12112
rect 1492 11688 1544 11694
rect 1492 11630 1544 11636
rect 1504 11150 1532 11630
rect 2240 11626 2268 12106
rect 2332 11830 2360 13126
rect 2320 11824 2372 11830
rect 2320 11766 2372 11772
rect 2228 11620 2280 11626
rect 2228 11562 2280 11568
rect 2240 11286 2268 11562
rect 2228 11280 2280 11286
rect 2228 11222 2280 11228
rect 1492 11144 1544 11150
rect 1492 11086 1544 11092
rect 1504 10742 1532 11086
rect 1492 10736 1544 10742
rect 1492 10678 1544 10684
rect 2044 10668 2096 10674
rect 2044 10610 2096 10616
rect 2056 10577 2084 10610
rect 2042 10568 2098 10577
rect 2042 10503 2098 10512
rect 1768 9920 1820 9926
rect 1768 9862 1820 9868
rect 1780 9489 1808 9862
rect 2240 9586 2268 11222
rect 2412 11008 2464 11014
rect 2412 10950 2464 10956
rect 2320 10600 2372 10606
rect 2320 10542 2372 10548
rect 2332 9926 2360 10542
rect 2424 10062 2452 10950
rect 2412 10056 2464 10062
rect 2412 9998 2464 10004
rect 2320 9920 2372 9926
rect 2320 9862 2372 9868
rect 2608 9722 2636 14200
rect 3422 13560 3478 13569
rect 3422 13495 3478 13504
rect 2964 13320 3016 13326
rect 2964 13262 3016 13268
rect 2688 13184 2740 13190
rect 2688 13126 2740 13132
rect 2700 12306 2728 13126
rect 2976 12850 3004 13262
rect 2964 12844 3016 12850
rect 2964 12786 3016 12792
rect 2778 12744 2834 12753
rect 2778 12679 2834 12688
rect 2688 12300 2740 12306
rect 2688 12242 2740 12248
rect 2792 10742 2820 12679
rect 2976 11898 3004 12786
rect 3148 12776 3200 12782
rect 3148 12718 3200 12724
rect 3160 12374 3188 12718
rect 3436 12442 3464 13495
rect 3424 12436 3476 12442
rect 3424 12378 3476 12384
rect 3148 12368 3200 12374
rect 3148 12310 3200 12316
rect 3436 12238 3464 12378
rect 3424 12232 3476 12238
rect 3424 12174 3476 12180
rect 3332 12096 3384 12102
rect 3332 12038 3384 12044
rect 2964 11892 3016 11898
rect 2964 11834 3016 11840
rect 2976 11150 3004 11834
rect 3344 11762 3372 12038
rect 3422 11928 3478 11937
rect 3422 11863 3478 11872
rect 3436 11830 3464 11863
rect 3424 11824 3476 11830
rect 3424 11766 3476 11772
rect 3332 11756 3384 11762
rect 3332 11698 3384 11704
rect 2964 11144 3016 11150
rect 2964 11086 3016 11092
rect 2780 10736 2832 10742
rect 2780 10678 2832 10684
rect 3148 10464 3200 10470
rect 3148 10406 3200 10412
rect 2780 10056 2832 10062
rect 2780 9998 2832 10004
rect 2596 9716 2648 9722
rect 2596 9658 2648 9664
rect 2792 9586 2820 9998
rect 3160 9654 3188 10406
rect 3344 9926 3372 11698
rect 3436 11354 3464 11766
rect 3424 11348 3476 11354
rect 3424 11290 3476 11296
rect 3424 10532 3476 10538
rect 3424 10474 3476 10480
rect 3332 9920 3384 9926
rect 3332 9862 3384 9868
rect 3436 9722 3464 10474
rect 3516 10464 3568 10470
rect 3804 10418 3832 14334
rect 4066 14200 4122 14334
rect 5538 14200 5594 15000
rect 7010 14200 7066 15000
rect 8482 14200 8538 15000
rect 9954 14200 10010 15000
rect 11426 14200 11482 15000
rect 12898 14200 12954 15000
rect 14370 14200 14426 15000
rect 15842 14200 15898 15000
rect 17314 14200 17370 15000
rect 18786 14200 18842 15000
rect 4214 13628 4522 13637
rect 4214 13626 4220 13628
rect 4276 13626 4300 13628
rect 4356 13626 4380 13628
rect 4436 13626 4460 13628
rect 4516 13626 4522 13628
rect 4276 13574 4278 13626
rect 4458 13574 4460 13626
rect 4214 13572 4220 13574
rect 4276 13572 4300 13574
rect 4356 13572 4380 13574
rect 4436 13572 4460 13574
rect 4516 13572 4522 13574
rect 4214 13563 4522 13572
rect 5552 13546 5580 14200
rect 5552 13518 5856 13546
rect 5540 13456 5592 13462
rect 5540 13398 5592 13404
rect 4436 13320 4488 13326
rect 4436 13262 4488 13268
rect 4528 13320 4580 13326
rect 4528 13262 4580 13268
rect 4344 13252 4396 13258
rect 4344 13194 4396 13200
rect 4356 12714 4384 13194
rect 4448 12918 4476 13262
rect 4436 12912 4488 12918
rect 4436 12854 4488 12860
rect 4540 12850 4568 13262
rect 5172 13184 5224 13190
rect 5172 13126 5224 13132
rect 4896 12912 4948 12918
rect 4896 12854 4948 12860
rect 4528 12844 4580 12850
rect 4580 12804 4660 12832
rect 4528 12786 4580 12792
rect 4344 12708 4396 12714
rect 4344 12650 4396 12656
rect 4214 12540 4522 12549
rect 4214 12538 4220 12540
rect 4276 12538 4300 12540
rect 4356 12538 4380 12540
rect 4436 12538 4460 12540
rect 4516 12538 4522 12540
rect 4276 12486 4278 12538
rect 4458 12486 4460 12538
rect 4214 12484 4220 12486
rect 4276 12484 4300 12486
rect 4356 12484 4380 12486
rect 4436 12484 4460 12486
rect 4516 12484 4522 12486
rect 4214 12475 4522 12484
rect 4632 12442 4660 12804
rect 4620 12436 4672 12442
rect 4620 12378 4672 12384
rect 4908 12374 4936 12854
rect 4896 12368 4948 12374
rect 4896 12310 4948 12316
rect 5184 11830 5212 13126
rect 5552 12306 5580 13398
rect 5632 13184 5684 13190
rect 5632 13126 5684 13132
rect 5644 12918 5672 13126
rect 5632 12912 5684 12918
rect 5632 12854 5684 12860
rect 5828 12434 5856 13518
rect 7024 13410 7052 14200
rect 8496 13530 8524 14200
rect 7104 13524 7156 13530
rect 7104 13466 7156 13472
rect 8484 13524 8536 13530
rect 8484 13466 8536 13472
rect 6552 13388 6604 13394
rect 6552 13330 6604 13336
rect 6840 13382 7052 13410
rect 6000 13252 6052 13258
rect 6000 13194 6052 13200
rect 5908 12844 5960 12850
rect 5908 12786 5960 12792
rect 5736 12406 5856 12434
rect 5540 12300 5592 12306
rect 5540 12242 5592 12248
rect 4068 11824 4120 11830
rect 4068 11766 4120 11772
rect 5172 11824 5224 11830
rect 5172 11766 5224 11772
rect 3884 11688 3936 11694
rect 3884 11630 3936 11636
rect 3896 11150 3924 11630
rect 3884 11144 3936 11150
rect 4080 11121 4108 11766
rect 5356 11688 5408 11694
rect 5356 11630 5408 11636
rect 5172 11620 5224 11626
rect 5172 11562 5224 11568
rect 4214 11452 4522 11461
rect 4214 11450 4220 11452
rect 4276 11450 4300 11452
rect 4356 11450 4380 11452
rect 4436 11450 4460 11452
rect 4516 11450 4522 11452
rect 4276 11398 4278 11450
rect 4458 11398 4460 11450
rect 4214 11396 4220 11398
rect 4276 11396 4300 11398
rect 4356 11396 4380 11398
rect 4436 11396 4460 11398
rect 4516 11396 4522 11398
rect 4214 11387 4522 11396
rect 5184 11286 5212 11562
rect 5172 11280 5224 11286
rect 5172 11222 5224 11228
rect 3884 11086 3936 11092
rect 4066 11112 4122 11121
rect 4066 11047 4122 11056
rect 3884 10736 3936 10742
rect 3884 10678 3936 10684
rect 3516 10406 3568 10412
rect 3528 10130 3556 10406
rect 3712 10390 3832 10418
rect 3516 10124 3568 10130
rect 3516 10066 3568 10072
rect 3712 9722 3740 10390
rect 3790 10296 3846 10305
rect 3790 10231 3846 10240
rect 3804 10130 3832 10231
rect 3896 10198 3924 10678
rect 4068 10668 4120 10674
rect 4068 10610 4120 10616
rect 3976 10600 4028 10606
rect 3976 10542 4028 10548
rect 3988 10266 4016 10542
rect 3976 10260 4028 10266
rect 3976 10202 4028 10208
rect 3884 10192 3936 10198
rect 3884 10134 3936 10140
rect 3792 10124 3844 10130
rect 3792 10066 3844 10072
rect 3424 9716 3476 9722
rect 3424 9658 3476 9664
rect 3700 9716 3752 9722
rect 3700 9658 3752 9664
rect 3148 9648 3200 9654
rect 3148 9590 3200 9596
rect 2228 9580 2280 9586
rect 2228 9522 2280 9528
rect 2780 9580 2832 9586
rect 2780 9522 2832 9528
rect 1766 9480 1822 9489
rect 1766 9415 1822 9424
rect 2044 9376 2096 9382
rect 2044 9318 2096 9324
rect 2056 8974 2084 9318
rect 2596 9036 2648 9042
rect 2596 8978 2648 8984
rect 2044 8968 2096 8974
rect 2044 8910 2096 8916
rect 1492 8900 1544 8906
rect 1492 8842 1544 8848
rect 1504 7886 1532 8842
rect 2608 8498 2636 8978
rect 2596 8492 2648 8498
rect 2596 8434 2648 8440
rect 1860 8288 1912 8294
rect 1860 8230 1912 8236
rect 1492 7880 1544 7886
rect 1492 7822 1544 7828
rect 1872 7410 1900 8230
rect 3160 7857 3188 9590
rect 3896 9450 3924 10134
rect 4080 10062 4108 10610
rect 4804 10600 4856 10606
rect 4804 10542 4856 10548
rect 4214 10364 4522 10373
rect 4214 10362 4220 10364
rect 4276 10362 4300 10364
rect 4356 10362 4380 10364
rect 4436 10362 4460 10364
rect 4516 10362 4522 10364
rect 4276 10310 4278 10362
rect 4458 10310 4460 10362
rect 4214 10308 4220 10310
rect 4276 10308 4300 10310
rect 4356 10308 4380 10310
rect 4436 10308 4460 10310
rect 4516 10308 4522 10310
rect 4214 10299 4522 10308
rect 4816 10062 4844 10542
rect 4068 10056 4120 10062
rect 4068 9998 4120 10004
rect 4804 10056 4856 10062
rect 4804 9998 4856 10004
rect 5264 10056 5316 10062
rect 5264 9998 5316 10004
rect 4252 9988 4304 9994
rect 4252 9930 4304 9936
rect 4264 9586 4292 9930
rect 4252 9580 4304 9586
rect 4252 9522 4304 9528
rect 5080 9580 5132 9586
rect 5080 9522 5132 9528
rect 3884 9444 3936 9450
rect 3884 9386 3936 9392
rect 4896 9376 4948 9382
rect 4896 9318 4948 9324
rect 4214 9276 4522 9285
rect 4214 9274 4220 9276
rect 4276 9274 4300 9276
rect 4356 9274 4380 9276
rect 4436 9274 4460 9276
rect 4516 9274 4522 9276
rect 4276 9222 4278 9274
rect 4458 9222 4460 9274
rect 4214 9220 4220 9222
rect 4276 9220 4300 9222
rect 4356 9220 4380 9222
rect 4436 9220 4460 9222
rect 4516 9220 4522 9222
rect 4214 9211 4522 9220
rect 4160 8900 4212 8906
rect 4160 8842 4212 8848
rect 3974 8664 4030 8673
rect 3974 8599 4030 8608
rect 3988 8430 4016 8599
rect 4172 8566 4200 8842
rect 4160 8560 4212 8566
rect 4160 8502 4212 8508
rect 4620 8492 4672 8498
rect 4620 8434 4672 8440
rect 3976 8424 4028 8430
rect 3976 8366 4028 8372
rect 4214 8188 4522 8197
rect 4214 8186 4220 8188
rect 4276 8186 4300 8188
rect 4356 8186 4380 8188
rect 4436 8186 4460 8188
rect 4516 8186 4522 8188
rect 4276 8134 4278 8186
rect 4458 8134 4460 8186
rect 4214 8132 4220 8134
rect 4276 8132 4300 8134
rect 4356 8132 4380 8134
rect 4436 8132 4460 8134
rect 4516 8132 4522 8134
rect 4214 8123 4522 8132
rect 4632 8022 4660 8434
rect 4620 8016 4672 8022
rect 4620 7958 4672 7964
rect 4908 7886 4936 9318
rect 5092 8566 5120 9522
rect 5276 9518 5304 9998
rect 5264 9512 5316 9518
rect 5264 9454 5316 9460
rect 5276 9110 5304 9454
rect 5264 9104 5316 9110
rect 5264 9046 5316 9052
rect 5080 8560 5132 8566
rect 5080 8502 5132 8508
rect 4988 8016 5040 8022
rect 4988 7958 5040 7964
rect 4896 7880 4948 7886
rect 3146 7848 3202 7857
rect 3056 7812 3108 7818
rect 4896 7822 4948 7828
rect 3146 7783 3202 7792
rect 3424 7812 3476 7818
rect 3056 7754 3108 7760
rect 3424 7754 3476 7760
rect 2596 7540 2648 7546
rect 2596 7482 2648 7488
rect 1860 7404 1912 7410
rect 1860 7346 1912 7352
rect 2044 7404 2096 7410
rect 2044 7346 2096 7352
rect 1872 6914 1900 7346
rect 2056 6934 2084 7346
rect 2412 7336 2464 7342
rect 2412 7278 2464 7284
rect 2044 6928 2096 6934
rect 1872 6886 1992 6914
rect 1676 6860 1728 6866
rect 1676 6802 1728 6808
rect 1584 6656 1636 6662
rect 1584 6598 1636 6604
rect 1596 6225 1624 6598
rect 1582 6216 1638 6225
rect 1582 6151 1638 6160
rect 1584 6112 1636 6118
rect 1584 6054 1636 6060
rect 1596 5409 1624 6054
rect 1582 5400 1638 5409
rect 1582 5335 1638 5344
rect 1688 4214 1716 6802
rect 1964 6798 1992 6886
rect 2044 6870 2096 6876
rect 2424 6798 2452 7278
rect 1952 6792 2004 6798
rect 1952 6734 2004 6740
rect 2412 6792 2464 6798
rect 2464 6752 2544 6780
rect 2412 6734 2464 6740
rect 1964 6322 1992 6734
rect 2412 6656 2464 6662
rect 2412 6598 2464 6604
rect 2424 6390 2452 6598
rect 2412 6384 2464 6390
rect 2412 6326 2464 6332
rect 1952 6316 2004 6322
rect 1952 6258 2004 6264
rect 2424 5914 2452 6326
rect 2516 5914 2544 6752
rect 2608 6322 2636 7482
rect 2780 7336 2832 7342
rect 2780 7278 2832 7284
rect 2792 7002 2820 7278
rect 2962 7032 3018 7041
rect 2780 6996 2832 7002
rect 2962 6967 3018 6976
rect 2780 6938 2832 6944
rect 2688 6928 2740 6934
rect 2688 6870 2740 6876
rect 2700 6458 2728 6870
rect 2792 6746 2820 6938
rect 2792 6718 2912 6746
rect 2780 6656 2832 6662
rect 2780 6598 2832 6604
rect 2688 6452 2740 6458
rect 2688 6394 2740 6400
rect 2792 6322 2820 6598
rect 2596 6316 2648 6322
rect 2596 6258 2648 6264
rect 2780 6316 2832 6322
rect 2780 6258 2832 6264
rect 2884 6254 2912 6718
rect 2872 6248 2924 6254
rect 2872 6190 2924 6196
rect 2596 6112 2648 6118
rect 2596 6054 2648 6060
rect 2412 5908 2464 5914
rect 2412 5850 2464 5856
rect 2504 5908 2556 5914
rect 2504 5850 2556 5856
rect 2608 5778 2636 6054
rect 2780 5840 2832 5846
rect 2780 5782 2832 5788
rect 2596 5772 2648 5778
rect 2596 5714 2648 5720
rect 2504 5704 2556 5710
rect 2504 5646 2556 5652
rect 2688 5704 2740 5710
rect 2792 5658 2820 5782
rect 2740 5652 2820 5658
rect 2688 5646 2820 5652
rect 2412 5024 2464 5030
rect 2412 4966 2464 4972
rect 1768 4684 1820 4690
rect 1768 4626 1820 4632
rect 1676 4208 1728 4214
rect 1676 4150 1728 4156
rect 1780 3777 1808 4626
rect 2136 4616 2188 4622
rect 2136 4558 2188 4564
rect 1860 4480 1912 4486
rect 1860 4422 1912 4428
rect 1872 4146 1900 4422
rect 1860 4140 1912 4146
rect 1860 4082 1912 4088
rect 1766 3768 1822 3777
rect 1766 3703 1822 3712
rect 1780 3534 1808 3703
rect 1872 3602 1900 4082
rect 1860 3596 1912 3602
rect 1860 3538 1912 3544
rect 1768 3528 1820 3534
rect 1768 3470 1820 3476
rect 1768 3392 1820 3398
rect 1768 3334 1820 3340
rect 1780 3058 1808 3334
rect 2148 3058 2176 4558
rect 2424 4146 2452 4966
rect 2516 4826 2544 5646
rect 2700 5630 2820 5646
rect 2780 5568 2832 5574
rect 2780 5510 2832 5516
rect 2792 5302 2820 5510
rect 2780 5296 2832 5302
rect 2780 5238 2832 5244
rect 2976 4826 3004 6967
rect 2504 4820 2556 4826
rect 2504 4762 2556 4768
rect 2964 4820 3016 4826
rect 2964 4762 3016 4768
rect 2596 4616 2648 4622
rect 2594 4584 2596 4593
rect 2648 4584 2650 4593
rect 2650 4542 2728 4570
rect 2594 4519 2650 4528
rect 2504 4276 2556 4282
rect 2504 4218 2556 4224
rect 2228 4140 2280 4146
rect 2228 4082 2280 4088
rect 2412 4140 2464 4146
rect 2412 4082 2464 4088
rect 2240 3602 2268 4082
rect 2228 3596 2280 3602
rect 2228 3538 2280 3544
rect 2240 3194 2268 3538
rect 2228 3188 2280 3194
rect 2228 3130 2280 3136
rect 1768 3052 1820 3058
rect 1768 2994 1820 3000
rect 2136 3052 2188 3058
rect 2136 2994 2188 3000
rect 2424 2922 2452 4082
rect 2516 3398 2544 4218
rect 2596 3460 2648 3466
rect 2596 3402 2648 3408
rect 2504 3392 2556 3398
rect 2504 3334 2556 3340
rect 2412 2916 2464 2922
rect 2412 2858 2464 2864
rect 2516 2650 2544 3334
rect 2504 2644 2556 2650
rect 2504 2586 2556 2592
rect 2044 2440 2096 2446
rect 2044 2382 2096 2388
rect 2056 2038 2084 2382
rect 2608 2038 2636 3402
rect 2700 3194 2728 4542
rect 2780 3460 2832 3466
rect 2780 3402 2832 3408
rect 2688 3188 2740 3194
rect 2688 3130 2740 3136
rect 2792 2961 2820 3402
rect 2872 3392 2924 3398
rect 2872 3334 2924 3340
rect 2778 2952 2834 2961
rect 2778 2887 2834 2896
rect 2792 2446 2820 2887
rect 2884 2514 2912 3334
rect 2872 2508 2924 2514
rect 2872 2450 2924 2456
rect 2780 2440 2832 2446
rect 2780 2382 2832 2388
rect 2044 2032 2096 2038
rect 2044 1974 2096 1980
rect 2596 2032 2648 2038
rect 2596 1974 2648 1980
rect 2792 1902 2820 2382
rect 2872 2372 2924 2378
rect 2872 2314 2924 2320
rect 2780 1896 2832 1902
rect 2780 1838 2832 1844
rect 1492 1420 1544 1426
rect 1492 1362 1544 1368
rect 1504 1329 1532 1362
rect 1490 1320 1546 1329
rect 1490 1255 1546 1264
rect 2792 1018 2820 1838
rect 2884 1562 2912 2314
rect 3068 2145 3096 7754
rect 3148 7404 3200 7410
rect 3148 7346 3200 7352
rect 3160 3738 3188 7346
rect 3436 7342 3464 7754
rect 4620 7744 4672 7750
rect 4620 7686 4672 7692
rect 4632 7410 4660 7686
rect 5000 7478 5028 7958
rect 5092 7546 5120 8502
rect 5368 8498 5396 11630
rect 5736 9586 5764 12406
rect 5920 12306 5948 12786
rect 5908 12300 5960 12306
rect 5908 12242 5960 12248
rect 6012 12238 6040 13194
rect 6092 13184 6144 13190
rect 6092 13126 6144 13132
rect 6184 13184 6236 13190
rect 6184 13126 6236 13132
rect 6104 12986 6132 13126
rect 6092 12980 6144 12986
rect 6092 12922 6144 12928
rect 6000 12232 6052 12238
rect 6000 12174 6052 12180
rect 5816 12096 5868 12102
rect 5816 12038 5868 12044
rect 5828 10742 5856 12038
rect 5908 11824 5960 11830
rect 5908 11766 5960 11772
rect 5920 11150 5948 11766
rect 5908 11144 5960 11150
rect 5908 11086 5960 11092
rect 5816 10736 5868 10742
rect 5816 10678 5868 10684
rect 5920 10674 5948 11086
rect 6012 11082 6040 12174
rect 6196 11898 6224 13126
rect 6276 12776 6328 12782
rect 6276 12718 6328 12724
rect 6288 12238 6316 12718
rect 6564 12714 6592 13330
rect 6840 12850 6868 13382
rect 7012 13320 7064 13326
rect 7012 13262 7064 13268
rect 6920 12980 6972 12986
rect 6920 12922 6972 12928
rect 6828 12844 6880 12850
rect 6748 12804 6828 12832
rect 6552 12708 6604 12714
rect 6552 12650 6604 12656
rect 6276 12232 6328 12238
rect 6276 12174 6328 12180
rect 6184 11892 6236 11898
rect 6184 11834 6236 11840
rect 6288 11830 6316 12174
rect 6276 11824 6328 11830
rect 6276 11766 6328 11772
rect 6092 11756 6144 11762
rect 6092 11698 6144 11704
rect 6104 11286 6132 11698
rect 6092 11280 6144 11286
rect 6092 11222 6144 11228
rect 6748 11218 6776 12804
rect 6828 12786 6880 12792
rect 6932 12782 6960 12922
rect 6920 12776 6972 12782
rect 6920 12718 6972 12724
rect 7024 11898 7052 13262
rect 7012 11892 7064 11898
rect 7012 11834 7064 11840
rect 6918 11792 6974 11801
rect 6918 11727 6974 11736
rect 7012 11756 7064 11762
rect 6826 11520 6882 11529
rect 6826 11455 6882 11464
rect 6736 11212 6788 11218
rect 6736 11154 6788 11160
rect 6840 11150 6868 11455
rect 6092 11144 6144 11150
rect 6092 11086 6144 11092
rect 6828 11144 6880 11150
rect 6828 11086 6880 11092
rect 6000 11076 6052 11082
rect 6000 11018 6052 11024
rect 6104 10674 6132 11086
rect 6736 10736 6788 10742
rect 6736 10678 6788 10684
rect 5908 10668 5960 10674
rect 5908 10610 5960 10616
rect 6092 10668 6144 10674
rect 6092 10610 6144 10616
rect 5908 10124 5960 10130
rect 5908 10066 5960 10072
rect 5920 9654 5948 10066
rect 6000 10056 6052 10062
rect 6052 10016 6132 10044
rect 6000 9998 6052 10004
rect 5908 9648 5960 9654
rect 5908 9590 5960 9596
rect 5724 9580 5776 9586
rect 5724 9522 5776 9528
rect 5736 9178 5764 9522
rect 5724 9172 5776 9178
rect 5724 9114 5776 9120
rect 5448 8900 5500 8906
rect 5448 8842 5500 8848
rect 5632 8900 5684 8906
rect 5632 8842 5684 8848
rect 5356 8492 5408 8498
rect 5356 8434 5408 8440
rect 5264 7880 5316 7886
rect 5368 7868 5396 8434
rect 5460 8090 5488 8842
rect 5644 8566 5672 8842
rect 5632 8560 5684 8566
rect 5632 8502 5684 8508
rect 5920 8430 5948 9590
rect 6104 9586 6132 10016
rect 6748 9994 6776 10678
rect 6932 10470 6960 11727
rect 7012 11698 7064 11704
rect 7024 11014 7052 11698
rect 7012 11008 7064 11014
rect 7012 10950 7064 10956
rect 7024 10713 7052 10950
rect 7116 10742 7144 13466
rect 8944 13388 8996 13394
rect 8944 13330 8996 13336
rect 7288 13252 7340 13258
rect 7288 13194 7340 13200
rect 7564 13252 7616 13258
rect 7564 13194 7616 13200
rect 7300 12832 7328 13194
rect 7380 12844 7432 12850
rect 7300 12804 7380 12832
rect 7380 12786 7432 12792
rect 7392 12306 7420 12786
rect 7576 12714 7604 13194
rect 8576 13184 8628 13190
rect 8576 13126 8628 13132
rect 8214 13084 8522 13093
rect 8214 13082 8220 13084
rect 8276 13082 8300 13084
rect 8356 13082 8380 13084
rect 8436 13082 8460 13084
rect 8516 13082 8522 13084
rect 8276 13030 8278 13082
rect 8458 13030 8460 13082
rect 8214 13028 8220 13030
rect 8276 13028 8300 13030
rect 8356 13028 8380 13030
rect 8436 13028 8460 13030
rect 8516 13028 8522 13030
rect 8214 13019 8522 13028
rect 7564 12708 7616 12714
rect 7564 12650 7616 12656
rect 7576 12374 7604 12650
rect 7748 12436 7800 12442
rect 7748 12378 7800 12384
rect 7564 12368 7616 12374
rect 7564 12310 7616 12316
rect 7380 12300 7432 12306
rect 7380 12242 7432 12248
rect 7760 12102 7788 12378
rect 8588 12306 8616 13126
rect 8956 12714 8984 13330
rect 9312 13320 9364 13326
rect 9312 13262 9364 13268
rect 9324 12850 9352 13262
rect 9588 13252 9640 13258
rect 9588 13194 9640 13200
rect 9772 13252 9824 13258
rect 9772 13194 9824 13200
rect 9600 12918 9628 13194
rect 9588 12912 9640 12918
rect 9588 12854 9640 12860
rect 9312 12844 9364 12850
rect 9312 12786 9364 12792
rect 8944 12708 8996 12714
rect 8944 12650 8996 12656
rect 8576 12300 8628 12306
rect 8576 12242 8628 12248
rect 8482 12200 8538 12209
rect 8482 12135 8484 12144
rect 8536 12135 8538 12144
rect 8850 12200 8906 12209
rect 8956 12170 8984 12650
rect 9140 12442 9260 12458
rect 9324 12442 9352 12786
rect 9128 12436 9260 12442
rect 9180 12430 9260 12436
rect 9128 12378 9180 12384
rect 9140 12347 9168 12378
rect 9128 12300 9180 12306
rect 9128 12242 9180 12248
rect 8850 12135 8906 12144
rect 8944 12164 8996 12170
rect 8484 12106 8536 12112
rect 7196 12096 7248 12102
rect 7196 12038 7248 12044
rect 7748 12096 7800 12102
rect 7748 12038 7800 12044
rect 7208 11082 7236 12038
rect 8214 11996 8522 12005
rect 8214 11994 8220 11996
rect 8276 11994 8300 11996
rect 8356 11994 8380 11996
rect 8436 11994 8460 11996
rect 8516 11994 8522 11996
rect 8276 11942 8278 11994
rect 8458 11942 8460 11994
rect 8214 11940 8220 11942
rect 8276 11940 8300 11942
rect 8356 11940 8380 11942
rect 8436 11940 8460 11942
rect 8516 11940 8522 11942
rect 8214 11931 8522 11940
rect 8208 11824 8260 11830
rect 8576 11824 8628 11830
rect 8260 11784 8576 11812
rect 8208 11766 8260 11772
rect 8576 11766 8628 11772
rect 8024 11756 8076 11762
rect 8024 11698 8076 11704
rect 7288 11280 7340 11286
rect 7288 11222 7340 11228
rect 7196 11076 7248 11082
rect 7196 11018 7248 11024
rect 7104 10736 7156 10742
rect 7010 10704 7066 10713
rect 7104 10678 7156 10684
rect 7010 10639 7066 10648
rect 6920 10464 6972 10470
rect 6920 10406 6972 10412
rect 7012 10464 7064 10470
rect 7012 10406 7064 10412
rect 7024 10062 7052 10406
rect 7012 10056 7064 10062
rect 7012 9998 7064 10004
rect 6736 9988 6788 9994
rect 6736 9930 6788 9936
rect 7208 9586 7236 11018
rect 7300 10674 7328 11222
rect 7840 11144 7892 11150
rect 7840 11086 7892 11092
rect 7472 11008 7524 11014
rect 7472 10950 7524 10956
rect 7484 10674 7512 10950
rect 7288 10668 7340 10674
rect 7288 10610 7340 10616
rect 7472 10668 7524 10674
rect 7472 10610 7524 10616
rect 7300 10130 7328 10610
rect 7852 10130 7880 11086
rect 7932 10668 7984 10674
rect 7932 10610 7984 10616
rect 7288 10124 7340 10130
rect 7288 10066 7340 10072
rect 7840 10124 7892 10130
rect 7840 10066 7892 10072
rect 7944 9926 7972 10610
rect 7932 9920 7984 9926
rect 7932 9862 7984 9868
rect 6092 9580 6144 9586
rect 6092 9522 6144 9528
rect 7196 9580 7248 9586
rect 7196 9522 7248 9528
rect 6000 8968 6052 8974
rect 5998 8936 6000 8945
rect 6052 8936 6054 8945
rect 5998 8871 6054 8880
rect 6104 8634 6132 9522
rect 7932 9512 7984 9518
rect 7932 9454 7984 9460
rect 7196 9444 7248 9450
rect 7248 9404 7328 9432
rect 7196 9386 7248 9392
rect 6920 9376 6972 9382
rect 6920 9318 6972 9324
rect 6932 9110 6960 9318
rect 7300 9178 7328 9404
rect 7288 9172 7340 9178
rect 7288 9114 7340 9120
rect 7944 9110 7972 9454
rect 6920 9104 6972 9110
rect 6642 9072 6698 9081
rect 6920 9046 6972 9052
rect 7932 9104 7984 9110
rect 7932 9046 7984 9052
rect 6642 9007 6698 9016
rect 6656 8634 6684 9007
rect 6828 8968 6880 8974
rect 6828 8910 6880 8916
rect 7196 8968 7248 8974
rect 7196 8910 7248 8916
rect 7656 8968 7708 8974
rect 7656 8910 7708 8916
rect 7748 8968 7800 8974
rect 7748 8910 7800 8916
rect 7838 8936 7894 8945
rect 6092 8628 6144 8634
rect 6092 8570 6144 8576
rect 6644 8628 6696 8634
rect 6644 8570 6696 8576
rect 6840 8566 6868 8910
rect 6828 8560 6880 8566
rect 6828 8502 6880 8508
rect 5540 8424 5592 8430
rect 5540 8366 5592 8372
rect 5908 8424 5960 8430
rect 5908 8366 5960 8372
rect 5448 8084 5500 8090
rect 5448 8026 5500 8032
rect 5316 7840 5396 7868
rect 5264 7822 5316 7828
rect 5552 7546 5580 8366
rect 5920 8090 5948 8366
rect 7208 8362 7236 8910
rect 7564 8832 7616 8838
rect 7564 8774 7616 8780
rect 7576 8498 7604 8774
rect 7668 8566 7696 8910
rect 7656 8560 7708 8566
rect 7656 8502 7708 8508
rect 7564 8492 7616 8498
rect 7564 8434 7616 8440
rect 7760 8430 7788 8910
rect 7838 8871 7894 8880
rect 7852 8838 7880 8871
rect 7840 8832 7892 8838
rect 7840 8774 7892 8780
rect 7748 8424 7800 8430
rect 7748 8366 7800 8372
rect 6644 8356 6696 8362
rect 6644 8298 6696 8304
rect 7196 8356 7248 8362
rect 7196 8298 7248 8304
rect 5908 8084 5960 8090
rect 5908 8026 5960 8032
rect 5920 7546 5948 8026
rect 6656 7886 6684 8298
rect 7852 8022 7880 8774
rect 7944 8634 7972 9046
rect 7932 8628 7984 8634
rect 7932 8570 7984 8576
rect 8036 8498 8064 11698
rect 8668 11688 8720 11694
rect 8220 11626 8340 11642
rect 8668 11630 8720 11636
rect 8208 11620 8340 11626
rect 8260 11614 8340 11620
rect 8208 11562 8260 11568
rect 8312 11257 8340 11614
rect 8576 11620 8628 11626
rect 8576 11562 8628 11568
rect 8298 11248 8354 11257
rect 8298 11183 8354 11192
rect 8116 11144 8168 11150
rect 8116 11086 8168 11092
rect 8128 10792 8156 11086
rect 8214 10908 8522 10917
rect 8214 10906 8220 10908
rect 8276 10906 8300 10908
rect 8356 10906 8380 10908
rect 8436 10906 8460 10908
rect 8516 10906 8522 10908
rect 8276 10854 8278 10906
rect 8458 10854 8460 10906
rect 8214 10852 8220 10854
rect 8276 10852 8300 10854
rect 8356 10852 8380 10854
rect 8436 10852 8460 10854
rect 8516 10852 8522 10854
rect 8214 10843 8522 10852
rect 8588 10810 8616 11562
rect 8680 11286 8708 11630
rect 8668 11280 8720 11286
rect 8668 11222 8720 11228
rect 8760 11144 8812 11150
rect 8666 11112 8722 11121
rect 8760 11086 8812 11092
rect 8666 11047 8722 11056
rect 8576 10804 8628 10810
rect 8128 10764 8524 10792
rect 8298 10704 8354 10713
rect 8496 10674 8524 10764
rect 8576 10746 8628 10752
rect 8298 10639 8300 10648
rect 8352 10639 8354 10648
rect 8484 10668 8536 10674
rect 8300 10610 8352 10616
rect 8484 10610 8536 10616
rect 8680 10554 8708 11047
rect 8208 10532 8260 10538
rect 8312 10526 8708 10554
rect 8312 10520 8340 10526
rect 8260 10492 8340 10520
rect 8208 10474 8260 10480
rect 8114 10432 8170 10441
rect 8114 10367 8170 10376
rect 8024 8492 8076 8498
rect 8024 8434 8076 8440
rect 7840 8016 7892 8022
rect 7840 7958 7892 7964
rect 7932 7948 7984 7954
rect 7932 7890 7984 7896
rect 6644 7880 6696 7886
rect 6644 7822 6696 7828
rect 7840 7880 7892 7886
rect 7840 7822 7892 7828
rect 7852 7546 7880 7822
rect 5080 7540 5132 7546
rect 5080 7482 5132 7488
rect 5540 7540 5592 7546
rect 5540 7482 5592 7488
rect 5908 7540 5960 7546
rect 5908 7482 5960 7488
rect 7840 7540 7892 7546
rect 7840 7482 7892 7488
rect 4988 7472 5040 7478
rect 4988 7414 5040 7420
rect 3608 7404 3660 7410
rect 3608 7346 3660 7352
rect 3976 7404 4028 7410
rect 3976 7346 4028 7352
rect 4620 7404 4672 7410
rect 4620 7346 4672 7352
rect 4712 7404 4764 7410
rect 4712 7346 4764 7352
rect 3424 7336 3476 7342
rect 3424 7278 3476 7284
rect 3240 6860 3292 6866
rect 3240 6802 3292 6808
rect 3252 5234 3280 6802
rect 3516 6316 3568 6322
rect 3516 6258 3568 6264
rect 3528 5914 3556 6258
rect 3620 6186 3648 7346
rect 3884 6792 3936 6798
rect 3884 6734 3936 6740
rect 3896 6662 3924 6734
rect 3884 6656 3936 6662
rect 3884 6598 3936 6604
rect 3700 6316 3752 6322
rect 3700 6258 3752 6264
rect 3608 6180 3660 6186
rect 3608 6122 3660 6128
rect 3516 5908 3568 5914
rect 3516 5850 3568 5856
rect 3712 5409 3740 6258
rect 3896 6254 3924 6598
rect 3988 6390 4016 7346
rect 4214 7100 4522 7109
rect 4214 7098 4220 7100
rect 4276 7098 4300 7100
rect 4356 7098 4380 7100
rect 4436 7098 4460 7100
rect 4516 7098 4522 7100
rect 4276 7046 4278 7098
rect 4458 7046 4460 7098
rect 4214 7044 4220 7046
rect 4276 7044 4300 7046
rect 4356 7044 4380 7046
rect 4436 7044 4460 7046
rect 4516 7044 4522 7046
rect 4214 7035 4522 7044
rect 4632 6934 4660 7346
rect 4620 6928 4672 6934
rect 4620 6870 4672 6876
rect 4724 6798 4752 7346
rect 4712 6792 4764 6798
rect 4712 6734 4764 6740
rect 3976 6384 4028 6390
rect 3976 6326 4028 6332
rect 4620 6384 4672 6390
rect 4620 6326 4672 6332
rect 4068 6316 4120 6322
rect 4068 6258 4120 6264
rect 3884 6248 3936 6254
rect 3884 6190 3936 6196
rect 4080 5914 4108 6258
rect 4214 6012 4522 6021
rect 4214 6010 4220 6012
rect 4276 6010 4300 6012
rect 4356 6010 4380 6012
rect 4436 6010 4460 6012
rect 4516 6010 4522 6012
rect 4276 5958 4278 6010
rect 4458 5958 4460 6010
rect 4214 5956 4220 5958
rect 4276 5956 4300 5958
rect 4356 5956 4380 5958
rect 4436 5956 4460 5958
rect 4516 5956 4522 5958
rect 4214 5947 4522 5956
rect 4068 5908 4120 5914
rect 4068 5850 4120 5856
rect 3884 5840 3936 5846
rect 3884 5782 3936 5788
rect 3698 5400 3754 5409
rect 3698 5335 3700 5344
rect 3752 5335 3754 5344
rect 3700 5306 3752 5312
rect 3712 5275 3740 5306
rect 3240 5228 3292 5234
rect 3240 5170 3292 5176
rect 3332 4480 3384 4486
rect 3332 4422 3384 4428
rect 3344 4078 3372 4422
rect 3332 4072 3384 4078
rect 3332 4014 3384 4020
rect 3148 3732 3200 3738
rect 3148 3674 3200 3680
rect 3896 3602 3924 5782
rect 4344 5636 4396 5642
rect 4344 5578 4396 5584
rect 4356 5234 4384 5578
rect 4632 5574 4660 6326
rect 4724 5846 4752 6734
rect 4896 6724 4948 6730
rect 4896 6666 4948 6672
rect 4908 6390 4936 6666
rect 4896 6384 4948 6390
rect 4896 6326 4948 6332
rect 5000 6118 5028 7414
rect 5920 7410 5948 7482
rect 7472 7472 7524 7478
rect 7472 7414 7524 7420
rect 5080 7404 5132 7410
rect 5080 7346 5132 7352
rect 5908 7404 5960 7410
rect 5908 7346 5960 7352
rect 5092 6798 5120 7346
rect 5356 7336 5408 7342
rect 5356 7278 5408 7284
rect 5080 6792 5132 6798
rect 5080 6734 5132 6740
rect 5368 6322 5396 7278
rect 6552 7200 6604 7206
rect 6552 7142 6604 7148
rect 5448 6384 5500 6390
rect 5448 6326 5500 6332
rect 5356 6316 5408 6322
rect 5356 6258 5408 6264
rect 4988 6112 5040 6118
rect 4988 6054 5040 6060
rect 5080 6112 5132 6118
rect 5080 6054 5132 6060
rect 4804 5908 4856 5914
rect 4804 5850 4856 5856
rect 4712 5840 4764 5846
rect 4712 5782 4764 5788
rect 4816 5642 4844 5850
rect 4804 5636 4856 5642
rect 4804 5578 4856 5584
rect 4620 5568 4672 5574
rect 4620 5510 4672 5516
rect 4712 5568 4764 5574
rect 4712 5510 4764 5516
rect 4632 5370 4660 5510
rect 4620 5364 4672 5370
rect 4620 5306 4672 5312
rect 4724 5250 4752 5510
rect 4632 5234 4752 5250
rect 4160 5228 4212 5234
rect 4160 5170 4212 5176
rect 4344 5228 4396 5234
rect 4344 5170 4396 5176
rect 4620 5228 4752 5234
rect 4672 5222 4752 5228
rect 4620 5170 4672 5176
rect 4172 5098 4200 5170
rect 4160 5092 4212 5098
rect 4160 5034 4212 5040
rect 4068 5024 4120 5030
rect 4068 4966 4120 4972
rect 4080 4690 4108 4966
rect 4214 4924 4522 4933
rect 4214 4922 4220 4924
rect 4276 4922 4300 4924
rect 4356 4922 4380 4924
rect 4436 4922 4460 4924
rect 4516 4922 4522 4924
rect 4276 4870 4278 4922
rect 4458 4870 4460 4922
rect 4214 4868 4220 4870
rect 4276 4868 4300 4870
rect 4356 4868 4380 4870
rect 4436 4868 4460 4870
rect 4516 4868 4522 4870
rect 4214 4859 4522 4868
rect 4068 4684 4120 4690
rect 4068 4626 4120 4632
rect 3884 3596 3936 3602
rect 3884 3538 3936 3544
rect 3240 3528 3292 3534
rect 3240 3470 3292 3476
rect 3252 2582 3280 3470
rect 4080 3194 4108 4626
rect 4252 4616 4304 4622
rect 4252 4558 4304 4564
rect 4264 4486 4292 4558
rect 4528 4548 4580 4554
rect 4528 4490 4580 4496
rect 4252 4480 4304 4486
rect 4252 4422 4304 4428
rect 4540 4010 4568 4490
rect 4528 4004 4580 4010
rect 4528 3946 4580 3952
rect 4214 3836 4522 3845
rect 4214 3834 4220 3836
rect 4276 3834 4300 3836
rect 4356 3834 4380 3836
rect 4436 3834 4460 3836
rect 4516 3834 4522 3836
rect 4276 3782 4278 3834
rect 4458 3782 4460 3834
rect 4214 3780 4220 3782
rect 4276 3780 4300 3782
rect 4356 3780 4380 3782
rect 4436 3780 4460 3782
rect 4516 3780 4522 3782
rect 4214 3771 4522 3780
rect 4632 3670 4660 5170
rect 4816 5098 4844 5578
rect 5092 5574 5120 6054
rect 5460 5642 5488 6326
rect 5540 5704 5592 5710
rect 5540 5646 5592 5652
rect 6368 5704 6420 5710
rect 6368 5646 6420 5652
rect 5264 5636 5316 5642
rect 5264 5578 5316 5584
rect 5448 5636 5500 5642
rect 5448 5578 5500 5584
rect 5080 5568 5132 5574
rect 5080 5510 5132 5516
rect 5276 5370 5304 5578
rect 5264 5364 5316 5370
rect 5264 5306 5316 5312
rect 5460 5302 5488 5578
rect 5448 5296 5500 5302
rect 5448 5238 5500 5244
rect 4896 5228 4948 5234
rect 4896 5170 4948 5176
rect 4712 5092 4764 5098
rect 4712 5034 4764 5040
rect 4804 5092 4856 5098
rect 4804 5034 4856 5040
rect 4724 4826 4752 5034
rect 4712 4820 4764 4826
rect 4712 4762 4764 4768
rect 4712 4480 4764 4486
rect 4712 4422 4764 4428
rect 4620 3664 4672 3670
rect 4620 3606 4672 3612
rect 4620 3528 4672 3534
rect 4620 3470 4672 3476
rect 4068 3188 4120 3194
rect 4068 3130 4120 3136
rect 4160 2984 4212 2990
rect 4080 2932 4160 2938
rect 4080 2926 4212 2932
rect 3332 2916 3384 2922
rect 3332 2858 3384 2864
rect 4080 2910 4200 2926
rect 3240 2576 3292 2582
rect 3240 2518 3292 2524
rect 3148 2440 3200 2446
rect 3148 2382 3200 2388
rect 3054 2136 3110 2145
rect 3160 2106 3188 2382
rect 3054 2071 3110 2080
rect 3148 2100 3200 2106
rect 3148 2042 3200 2048
rect 3252 2038 3280 2518
rect 3240 2032 3292 2038
rect 3240 1974 3292 1980
rect 3344 1970 3372 2858
rect 4080 2530 4108 2910
rect 4214 2748 4522 2757
rect 4214 2746 4220 2748
rect 4276 2746 4300 2748
rect 4356 2746 4380 2748
rect 4436 2746 4460 2748
rect 4516 2746 4522 2748
rect 4276 2694 4278 2746
rect 4458 2694 4460 2746
rect 4214 2692 4220 2694
rect 4276 2692 4300 2694
rect 4356 2692 4380 2694
rect 4436 2692 4460 2694
rect 4516 2692 4522 2694
rect 4214 2683 4522 2692
rect 4632 2582 4660 3470
rect 4620 2576 4672 2582
rect 4080 2502 4200 2530
rect 4620 2518 4672 2524
rect 4172 2446 4200 2502
rect 4160 2440 4212 2446
rect 4160 2382 4212 2388
rect 3608 2304 3660 2310
rect 3608 2246 3660 2252
rect 3620 2038 3648 2246
rect 3608 2032 3660 2038
rect 3608 1974 3660 1980
rect 3332 1964 3384 1970
rect 3332 1906 3384 1912
rect 2872 1556 2924 1562
rect 2872 1498 2924 1504
rect 3344 1358 3372 1906
rect 4172 1902 4200 2382
rect 4620 2100 4672 2106
rect 4620 2042 4672 2048
rect 4160 1896 4212 1902
rect 4160 1838 4212 1844
rect 4214 1660 4522 1669
rect 4214 1658 4220 1660
rect 4276 1658 4300 1660
rect 4356 1658 4380 1660
rect 4436 1658 4460 1660
rect 4516 1658 4522 1660
rect 4276 1606 4278 1658
rect 4458 1606 4460 1658
rect 4214 1604 4220 1606
rect 4276 1604 4300 1606
rect 4356 1604 4380 1606
rect 4436 1604 4460 1606
rect 4516 1604 4522 1606
rect 4214 1595 4522 1604
rect 3332 1352 3384 1358
rect 3332 1294 3384 1300
rect 4528 1284 4580 1290
rect 4528 1226 4580 1232
rect 2780 1012 2832 1018
rect 2780 954 2832 960
rect 4540 950 4568 1226
rect 4632 1222 4660 2042
rect 4620 1216 4672 1222
rect 4620 1158 4672 1164
rect 4528 944 4580 950
rect 4528 886 4580 892
rect 4724 762 4752 4422
rect 4816 3194 4844 5034
rect 4908 4622 4936 5170
rect 5080 5160 5132 5166
rect 5080 5102 5132 5108
rect 5092 4826 5120 5102
rect 5080 4820 5132 4826
rect 5080 4762 5132 4768
rect 5092 4622 5120 4762
rect 5552 4690 5580 5646
rect 6184 5160 6236 5166
rect 6184 5102 6236 5108
rect 5540 4684 5592 4690
rect 5540 4626 5592 4632
rect 6196 4622 6224 5102
rect 4896 4616 4948 4622
rect 4896 4558 4948 4564
rect 5080 4616 5132 4622
rect 5080 4558 5132 4564
rect 6000 4616 6052 4622
rect 6000 4558 6052 4564
rect 6184 4616 6236 4622
rect 6184 4558 6236 4564
rect 4908 4282 4936 4558
rect 4988 4480 5040 4486
rect 4988 4422 5040 4428
rect 4896 4276 4948 4282
rect 4896 4218 4948 4224
rect 5000 4214 5028 4422
rect 4988 4208 5040 4214
rect 4988 4150 5040 4156
rect 5092 4010 5120 4558
rect 5632 4140 5684 4146
rect 5632 4082 5684 4088
rect 5816 4140 5868 4146
rect 5816 4082 5868 4088
rect 5172 4072 5224 4078
rect 5172 4014 5224 4020
rect 5540 4072 5592 4078
rect 5540 4014 5592 4020
rect 5080 4004 5132 4010
rect 5080 3946 5132 3952
rect 5184 3602 5212 4014
rect 5172 3596 5224 3602
rect 5172 3538 5224 3544
rect 5448 3596 5500 3602
rect 5448 3538 5500 3544
rect 4804 3188 4856 3194
rect 4804 3130 4856 3136
rect 4988 3052 5040 3058
rect 4988 2994 5040 3000
rect 5356 3052 5408 3058
rect 5356 2994 5408 3000
rect 5000 2378 5028 2994
rect 5368 2650 5396 2994
rect 5356 2644 5408 2650
rect 5356 2586 5408 2592
rect 5264 2440 5316 2446
rect 5264 2382 5316 2388
rect 4988 2372 5040 2378
rect 4988 2314 5040 2320
rect 4804 2304 4856 2310
rect 4804 2246 4856 2252
rect 4816 1766 4844 2246
rect 5000 1834 5028 2314
rect 5276 2106 5304 2382
rect 5264 2100 5316 2106
rect 5264 2042 5316 2048
rect 5172 2032 5224 2038
rect 5172 1974 5224 1980
rect 4988 1828 5040 1834
rect 4988 1770 5040 1776
rect 4804 1760 4856 1766
rect 4804 1702 4856 1708
rect 4816 1426 4844 1702
rect 4804 1420 4856 1426
rect 4804 1362 4856 1368
rect 5184 1358 5212 1974
rect 5356 1896 5408 1902
rect 5356 1838 5408 1844
rect 5368 1358 5396 1838
rect 5172 1352 5224 1358
rect 5172 1294 5224 1300
rect 5356 1352 5408 1358
rect 5356 1294 5408 1300
rect 5460 950 5488 3538
rect 5552 3534 5580 4014
rect 5540 3528 5592 3534
rect 5540 3470 5592 3476
rect 5644 2990 5672 4082
rect 5724 4072 5776 4078
rect 5724 4014 5776 4020
rect 5632 2984 5684 2990
rect 5632 2926 5684 2932
rect 5736 2922 5764 4014
rect 5828 3194 5856 4082
rect 5908 3392 5960 3398
rect 5908 3334 5960 3340
rect 5816 3188 5868 3194
rect 5816 3130 5868 3136
rect 5920 3058 5948 3334
rect 5908 3052 5960 3058
rect 5908 2994 5960 3000
rect 5724 2916 5776 2922
rect 5724 2858 5776 2864
rect 5736 2514 5764 2858
rect 6012 2530 6040 4558
rect 6196 4078 6224 4558
rect 6184 4072 6236 4078
rect 6184 4014 6236 4020
rect 6380 3738 6408 5646
rect 6460 5024 6512 5030
rect 6460 4966 6512 4972
rect 6472 4690 6500 4966
rect 6564 4826 6592 7142
rect 7484 6866 7512 7414
rect 7944 7410 7972 7890
rect 8036 7410 8064 8434
rect 8128 8430 8156 10367
rect 8220 10062 8248 10474
rect 8392 10464 8444 10470
rect 8772 10441 8800 11086
rect 8864 10554 8892 12135
rect 8944 12106 8996 12112
rect 9036 11076 9088 11082
rect 9036 11018 9088 11024
rect 9048 10577 9076 11018
rect 9034 10568 9090 10577
rect 8864 10526 8984 10554
rect 8852 10464 8904 10470
rect 8392 10406 8444 10412
rect 8758 10432 8814 10441
rect 8404 10146 8432 10406
rect 8852 10406 8904 10412
rect 8758 10367 8814 10376
rect 8312 10130 8432 10146
rect 8300 10124 8432 10130
rect 8352 10118 8432 10124
rect 8668 10124 8720 10130
rect 8300 10066 8352 10072
rect 8668 10066 8720 10072
rect 8208 10056 8260 10062
rect 8208 9998 8260 10004
rect 8576 9988 8628 9994
rect 8576 9930 8628 9936
rect 8214 9820 8522 9829
rect 8214 9818 8220 9820
rect 8276 9818 8300 9820
rect 8356 9818 8380 9820
rect 8436 9818 8460 9820
rect 8516 9818 8522 9820
rect 8276 9766 8278 9818
rect 8458 9766 8460 9818
rect 8214 9764 8220 9766
rect 8276 9764 8300 9766
rect 8356 9764 8380 9766
rect 8436 9764 8460 9766
rect 8516 9764 8522 9766
rect 8214 9755 8522 9764
rect 8300 9580 8352 9586
rect 8300 9522 8352 9528
rect 8484 9580 8536 9586
rect 8588 9568 8616 9930
rect 8680 9654 8708 10066
rect 8760 10056 8812 10062
rect 8760 9998 8812 10004
rect 8668 9648 8720 9654
rect 8668 9590 8720 9596
rect 8536 9540 8616 9568
rect 8484 9522 8536 9528
rect 8312 8922 8340 9522
rect 8680 9518 8708 9590
rect 8668 9512 8720 9518
rect 8668 9454 8720 9460
rect 8576 9376 8628 9382
rect 8576 9318 8628 9324
rect 8588 9110 8616 9318
rect 8576 9104 8628 9110
rect 8576 9046 8628 9052
rect 8680 9042 8708 9454
rect 8668 9036 8720 9042
rect 8668 8978 8720 8984
rect 8772 8922 8800 9998
rect 8312 8894 8800 8922
rect 8680 8838 8708 8894
rect 8576 8832 8628 8838
rect 8576 8774 8628 8780
rect 8668 8832 8720 8838
rect 8668 8774 8720 8780
rect 8214 8732 8522 8741
rect 8214 8730 8220 8732
rect 8276 8730 8300 8732
rect 8356 8730 8380 8732
rect 8436 8730 8460 8732
rect 8516 8730 8522 8732
rect 8276 8678 8278 8730
rect 8458 8678 8460 8730
rect 8214 8676 8220 8678
rect 8276 8676 8300 8678
rect 8356 8676 8380 8678
rect 8436 8676 8460 8678
rect 8516 8676 8522 8678
rect 8214 8667 8522 8676
rect 8116 8424 8168 8430
rect 8116 8366 8168 8372
rect 8128 7546 8156 8366
rect 8588 7886 8616 8774
rect 8680 8566 8708 8774
rect 8668 8560 8720 8566
rect 8668 8502 8720 8508
rect 8864 8498 8892 10406
rect 8956 9586 8984 10526
rect 9034 10503 9036 10512
rect 9088 10503 9090 10512
rect 9036 10474 9088 10480
rect 9048 10443 9076 10474
rect 9140 9654 9168 12242
rect 9232 12170 9260 12430
rect 9312 12436 9364 12442
rect 9312 12378 9364 12384
rect 9496 12436 9548 12442
rect 9496 12378 9548 12384
rect 9404 12232 9456 12238
rect 9404 12174 9456 12180
rect 9220 12164 9272 12170
rect 9220 12106 9272 12112
rect 9232 12073 9260 12106
rect 9218 12064 9274 12073
rect 9218 11999 9274 12008
rect 9416 11898 9444 12174
rect 9404 11892 9456 11898
rect 9404 11834 9456 11840
rect 9508 11762 9536 12378
rect 9586 12200 9642 12209
rect 9586 12135 9642 12144
rect 9600 12102 9628 12135
rect 9588 12096 9640 12102
rect 9588 12038 9640 12044
rect 9680 12096 9732 12102
rect 9680 12038 9732 12044
rect 9784 12084 9812 13194
rect 9864 12096 9916 12102
rect 9784 12056 9864 12084
rect 9692 11898 9720 12038
rect 9680 11892 9732 11898
rect 9680 11834 9732 11840
rect 9784 11801 9812 12056
rect 9864 12038 9916 12044
rect 9968 11830 9996 14200
rect 10140 13320 10192 13326
rect 10140 13262 10192 13268
rect 10152 12850 10180 13262
rect 11336 13252 11388 13258
rect 11336 13194 11388 13200
rect 10600 13184 10652 13190
rect 10600 13126 10652 13132
rect 10784 13184 10836 13190
rect 10784 13126 10836 13132
rect 11060 13184 11112 13190
rect 11060 13126 11112 13132
rect 10612 12986 10640 13126
rect 10600 12980 10652 12986
rect 10600 12922 10652 12928
rect 10796 12850 10824 13126
rect 11072 12918 11100 13126
rect 11060 12912 11112 12918
rect 11060 12854 11112 12860
rect 10140 12844 10192 12850
rect 10140 12786 10192 12792
rect 10784 12844 10836 12850
rect 10784 12786 10836 12792
rect 10322 12744 10378 12753
rect 10322 12679 10378 12688
rect 10046 12336 10102 12345
rect 10046 12271 10102 12280
rect 9956 11824 10008 11830
rect 9770 11792 9826 11801
rect 9496 11756 9548 11762
rect 9956 11766 10008 11772
rect 9770 11727 9826 11736
rect 9864 11756 9916 11762
rect 9496 11698 9548 11704
rect 9864 11698 9916 11704
rect 9876 11665 9904 11698
rect 9956 11688 10008 11694
rect 9862 11656 9918 11665
rect 9496 11620 9548 11626
rect 9956 11630 10008 11636
rect 9862 11591 9918 11600
rect 9496 11562 9548 11568
rect 9508 11150 9536 11562
rect 9968 11218 9996 11630
rect 10060 11286 10088 12271
rect 10336 12170 10364 12679
rect 11348 12442 11376 13194
rect 11336 12436 11388 12442
rect 11336 12378 11388 12384
rect 10414 12336 10470 12345
rect 10414 12271 10470 12280
rect 10508 12300 10560 12306
rect 10428 12238 10456 12271
rect 10508 12242 10560 12248
rect 10416 12232 10468 12238
rect 10416 12174 10468 12180
rect 10324 12164 10376 12170
rect 10324 12106 10376 12112
rect 10520 11898 10548 12242
rect 10600 12232 10652 12238
rect 10600 12174 10652 12180
rect 11152 12232 11204 12238
rect 11152 12174 11204 12180
rect 11244 12232 11296 12238
rect 11244 12174 11296 12180
rect 10612 11937 10640 12174
rect 10968 12164 11020 12170
rect 11020 12124 11100 12152
rect 10968 12106 11020 12112
rect 10598 11928 10654 11937
rect 10508 11892 10560 11898
rect 11072 11898 11100 12124
rect 10598 11863 10600 11872
rect 10508 11834 10560 11840
rect 10652 11863 10654 11872
rect 11060 11892 11112 11898
rect 10600 11834 10652 11840
rect 11060 11834 11112 11840
rect 10140 11824 10192 11830
rect 10612 11803 10640 11834
rect 10140 11766 10192 11772
rect 10782 11792 10838 11801
rect 10048 11280 10100 11286
rect 10048 11222 10100 11228
rect 9956 11212 10008 11218
rect 9956 11154 10008 11160
rect 9496 11144 9548 11150
rect 9218 11112 9274 11121
rect 9496 11086 9548 11092
rect 9218 11047 9274 11056
rect 9128 9648 9180 9654
rect 9128 9590 9180 9596
rect 8944 9580 8996 9586
rect 8944 9522 8996 9528
rect 8852 8492 8904 8498
rect 8852 8434 8904 8440
rect 8944 8492 8996 8498
rect 8944 8434 8996 8440
rect 8956 8090 8984 8434
rect 9232 8294 9260 11047
rect 9600 10764 9996 10792
rect 9494 10568 9550 10577
rect 9600 10538 9628 10764
rect 9968 10674 9996 10764
rect 10152 10713 10180 11766
rect 10232 11756 10284 11762
rect 10782 11727 10838 11736
rect 10232 11698 10284 11704
rect 10244 11014 10272 11698
rect 10508 11688 10560 11694
rect 10506 11656 10508 11665
rect 10560 11656 10562 11665
rect 10506 11591 10562 11600
rect 10414 11384 10470 11393
rect 10414 11319 10470 11328
rect 10428 11150 10456 11319
rect 10520 11286 10548 11591
rect 10508 11280 10560 11286
rect 10508 11222 10560 11228
rect 10796 11234 10824 11727
rect 10874 11656 10930 11665
rect 10874 11591 10930 11600
rect 10888 11558 10916 11591
rect 10876 11552 10928 11558
rect 10968 11552 11020 11558
rect 10876 11494 10928 11500
rect 10966 11520 10968 11529
rect 11020 11520 11022 11529
rect 10966 11455 11022 11464
rect 10968 11348 11020 11354
rect 10968 11290 11020 11296
rect 10980 11257 11008 11290
rect 10966 11248 11022 11257
rect 10796 11218 10916 11234
rect 10796 11212 10928 11218
rect 10796 11206 10876 11212
rect 10966 11183 11022 11192
rect 10876 11154 10928 11160
rect 10416 11144 10468 11150
rect 10416 11086 10468 11092
rect 10784 11144 10836 11150
rect 10784 11086 10836 11092
rect 10968 11144 11020 11150
rect 10968 11086 11020 11092
rect 10232 11008 10284 11014
rect 10232 10950 10284 10956
rect 10244 10742 10272 10950
rect 10232 10736 10284 10742
rect 10138 10704 10194 10713
rect 9864 10668 9916 10674
rect 9864 10610 9916 10616
rect 9956 10668 10008 10674
rect 10284 10713 10364 10724
rect 10284 10704 10378 10713
rect 10284 10696 10322 10704
rect 10232 10678 10284 10684
rect 10138 10639 10194 10648
rect 10322 10639 10378 10648
rect 9956 10610 10008 10616
rect 9494 10503 9550 10512
rect 9588 10532 9640 10538
rect 9508 10470 9536 10503
rect 9772 10532 9824 10538
rect 9588 10474 9640 10480
rect 9692 10492 9772 10520
rect 9496 10464 9548 10470
rect 9496 10406 9548 10412
rect 9692 9926 9720 10492
rect 9772 10474 9824 10480
rect 9876 10470 9904 10610
rect 10232 10600 10284 10606
rect 10232 10542 10284 10548
rect 9864 10464 9916 10470
rect 9864 10406 9916 10412
rect 10046 10160 10102 10169
rect 9772 10124 9824 10130
rect 10046 10095 10048 10104
rect 9772 10066 9824 10072
rect 10100 10095 10102 10104
rect 10048 10066 10100 10072
rect 9784 10033 9812 10066
rect 9864 10056 9916 10062
rect 9770 10024 9826 10033
rect 9864 9998 9916 10004
rect 9770 9959 9826 9968
rect 9496 9920 9548 9926
rect 9496 9862 9548 9868
rect 9680 9920 9732 9926
rect 9680 9862 9732 9868
rect 9508 8974 9536 9862
rect 9692 9586 9720 9862
rect 9588 9580 9640 9586
rect 9588 9522 9640 9528
rect 9680 9580 9732 9586
rect 9680 9522 9732 9528
rect 9600 9110 9628 9522
rect 9588 9104 9640 9110
rect 9588 9046 9640 9052
rect 9404 8968 9456 8974
rect 9404 8910 9456 8916
rect 9496 8968 9548 8974
rect 9496 8910 9548 8916
rect 9416 8634 9444 8910
rect 9588 8832 9640 8838
rect 9588 8774 9640 8780
rect 9404 8628 9456 8634
rect 9404 8570 9456 8576
rect 9494 8528 9550 8537
rect 9494 8463 9550 8472
rect 9508 8430 9536 8463
rect 9496 8424 9548 8430
rect 9496 8366 9548 8372
rect 9600 8294 9628 8774
rect 9692 8566 9720 9522
rect 9876 9178 9904 9998
rect 10060 9654 10088 10066
rect 10140 9988 10192 9994
rect 10140 9930 10192 9936
rect 10152 9654 10180 9930
rect 10048 9648 10100 9654
rect 10048 9590 10100 9596
rect 10140 9648 10192 9654
rect 10140 9590 10192 9596
rect 9956 9376 10008 9382
rect 9956 9318 10008 9324
rect 9864 9172 9916 9178
rect 9864 9114 9916 9120
rect 9772 9104 9824 9110
rect 9772 9046 9824 9052
rect 9784 8906 9812 9046
rect 9772 8900 9824 8906
rect 9772 8842 9824 8848
rect 9680 8560 9732 8566
rect 9680 8502 9732 8508
rect 9772 8492 9824 8498
rect 9772 8434 9824 8440
rect 9220 8288 9272 8294
rect 9220 8230 9272 8236
rect 9588 8288 9640 8294
rect 9588 8230 9640 8236
rect 8944 8084 8996 8090
rect 8944 8026 8996 8032
rect 8576 7880 8628 7886
rect 8576 7822 8628 7828
rect 8668 7744 8720 7750
rect 8668 7686 8720 7692
rect 8214 7644 8522 7653
rect 8214 7642 8220 7644
rect 8276 7642 8300 7644
rect 8356 7642 8380 7644
rect 8436 7642 8460 7644
rect 8516 7642 8522 7644
rect 8276 7590 8278 7642
rect 8458 7590 8460 7642
rect 8214 7588 8220 7590
rect 8276 7588 8300 7590
rect 8356 7588 8380 7590
rect 8436 7588 8460 7590
rect 8516 7588 8522 7590
rect 8214 7579 8522 7588
rect 8116 7540 8168 7546
rect 8116 7482 8168 7488
rect 8680 7478 8708 7686
rect 8668 7472 8720 7478
rect 8668 7414 8720 7420
rect 8956 7410 8984 8026
rect 9784 7936 9812 8434
rect 9876 8430 9904 9114
rect 9968 8566 9996 9318
rect 10140 8628 10192 8634
rect 10140 8570 10192 8576
rect 9956 8560 10008 8566
rect 9956 8502 10008 8508
rect 9864 8424 9916 8430
rect 9864 8366 9916 8372
rect 10152 8362 10180 8570
rect 10244 8430 10272 10542
rect 10428 10470 10456 11086
rect 10692 11076 10744 11082
rect 10692 11018 10744 11024
rect 10508 10668 10560 10674
rect 10508 10610 10560 10616
rect 10416 10464 10468 10470
rect 10416 10406 10468 10412
rect 10416 10124 10468 10130
rect 10416 10066 10468 10072
rect 10322 8800 10378 8809
rect 10322 8735 10378 8744
rect 10336 8498 10364 8735
rect 10428 8498 10456 10066
rect 10520 9586 10548 10610
rect 10704 9926 10732 11018
rect 10796 10849 10824 11086
rect 10980 10985 11008 11086
rect 10966 10976 11022 10985
rect 10966 10911 11022 10920
rect 10782 10840 10838 10849
rect 10782 10775 10838 10784
rect 10876 10464 10928 10470
rect 10876 10406 10928 10412
rect 10888 10062 10916 10406
rect 10784 10056 10836 10062
rect 10784 9998 10836 10004
rect 10876 10056 10928 10062
rect 10876 9998 10928 10004
rect 10692 9920 10744 9926
rect 10692 9862 10744 9868
rect 10796 9586 10824 9998
rect 10980 9674 11008 10911
rect 11072 10742 11100 11834
rect 11164 11286 11192 12174
rect 11256 11830 11284 12174
rect 11244 11824 11296 11830
rect 11244 11766 11296 11772
rect 11152 11280 11204 11286
rect 11152 11222 11204 11228
rect 11060 10736 11112 10742
rect 11060 10678 11112 10684
rect 11072 10418 11100 10678
rect 11164 10538 11192 11222
rect 11440 10674 11468 14200
rect 12716 13728 12768 13734
rect 12716 13670 12768 13676
rect 12214 13628 12522 13637
rect 12214 13626 12220 13628
rect 12276 13626 12300 13628
rect 12356 13626 12380 13628
rect 12436 13626 12460 13628
rect 12516 13626 12522 13628
rect 12276 13574 12278 13626
rect 12458 13574 12460 13626
rect 12214 13572 12220 13574
rect 12276 13572 12300 13574
rect 12356 13572 12380 13574
rect 12436 13572 12460 13574
rect 12516 13572 12522 13574
rect 12214 13563 12522 13572
rect 11612 13320 11664 13326
rect 11612 13262 11664 13268
rect 12624 13320 12676 13326
rect 12624 13262 12676 13268
rect 11624 12986 11652 13262
rect 12256 13252 12308 13258
rect 12256 13194 12308 13200
rect 11612 12980 11664 12986
rect 11612 12922 11664 12928
rect 11624 12850 11652 12922
rect 11612 12844 11664 12850
rect 11612 12786 11664 12792
rect 11624 12753 11652 12786
rect 12072 12776 12124 12782
rect 11610 12744 11666 12753
rect 12072 12718 12124 12724
rect 11610 12679 11666 12688
rect 12084 12442 12112 12718
rect 12268 12646 12296 13194
rect 12256 12640 12308 12646
rect 12256 12582 12308 12588
rect 12214 12540 12522 12549
rect 12214 12538 12220 12540
rect 12276 12538 12300 12540
rect 12356 12538 12380 12540
rect 12436 12538 12460 12540
rect 12516 12538 12522 12540
rect 12276 12486 12278 12538
rect 12458 12486 12460 12538
rect 12214 12484 12220 12486
rect 12276 12484 12300 12486
rect 12356 12484 12380 12486
rect 12436 12484 12460 12486
rect 12516 12484 12522 12486
rect 12214 12475 12522 12484
rect 12072 12436 12124 12442
rect 12072 12378 12124 12384
rect 11796 12368 11848 12374
rect 11796 12310 11848 12316
rect 11888 12368 11940 12374
rect 11888 12310 11940 12316
rect 11808 12209 11836 12310
rect 11794 12200 11850 12209
rect 11794 12135 11850 12144
rect 11796 12096 11848 12102
rect 11796 12038 11848 12044
rect 11704 11824 11756 11830
rect 11704 11766 11756 11772
rect 11520 11756 11572 11762
rect 11520 11698 11572 11704
rect 11532 11218 11560 11698
rect 11612 11620 11664 11626
rect 11612 11562 11664 11568
rect 11520 11212 11572 11218
rect 11520 11154 11572 11160
rect 11520 11008 11572 11014
rect 11520 10950 11572 10956
rect 11428 10668 11480 10674
rect 11428 10610 11480 10616
rect 11152 10532 11204 10538
rect 11152 10474 11204 10480
rect 11072 10390 11192 10418
rect 11060 9988 11112 9994
rect 11060 9930 11112 9936
rect 11072 9722 11100 9930
rect 10888 9646 11008 9674
rect 11060 9716 11112 9722
rect 11060 9658 11112 9664
rect 10508 9580 10560 9586
rect 10508 9522 10560 9528
rect 10784 9580 10836 9586
rect 10784 9522 10836 9528
rect 10508 9376 10560 9382
rect 10508 9318 10560 9324
rect 10520 9178 10548 9318
rect 10796 9178 10824 9522
rect 10508 9172 10560 9178
rect 10508 9114 10560 9120
rect 10784 9172 10836 9178
rect 10784 9114 10836 9120
rect 10692 9104 10744 9110
rect 10692 9046 10744 9052
rect 10600 8968 10652 8974
rect 10598 8936 10600 8945
rect 10652 8936 10654 8945
rect 10508 8900 10560 8906
rect 10598 8871 10654 8880
rect 10508 8842 10560 8848
rect 10520 8537 10548 8842
rect 10506 8528 10562 8537
rect 10324 8492 10376 8498
rect 10324 8434 10376 8440
rect 10416 8492 10468 8498
rect 10506 8463 10562 8472
rect 10416 8434 10468 8440
rect 10232 8424 10284 8430
rect 10232 8366 10284 8372
rect 10140 8356 10192 8362
rect 10140 8298 10192 8304
rect 10416 8356 10468 8362
rect 10416 8298 10468 8304
rect 9508 7908 9812 7936
rect 9508 7818 9536 7908
rect 9864 7880 9916 7886
rect 9864 7822 9916 7828
rect 9496 7812 9548 7818
rect 9496 7754 9548 7760
rect 9128 7744 9180 7750
rect 9128 7686 9180 7692
rect 9140 7410 9168 7686
rect 7932 7404 7984 7410
rect 7932 7346 7984 7352
rect 8024 7404 8076 7410
rect 8024 7346 8076 7352
rect 8944 7404 8996 7410
rect 8944 7346 8996 7352
rect 9128 7404 9180 7410
rect 9128 7346 9180 7352
rect 7472 6860 7524 6866
rect 7472 6802 7524 6808
rect 6920 6792 6972 6798
rect 6920 6734 6972 6740
rect 8116 6792 8168 6798
rect 8116 6734 8168 6740
rect 6932 6390 6960 6734
rect 7012 6724 7064 6730
rect 7012 6666 7064 6672
rect 6920 6384 6972 6390
rect 6920 6326 6972 6332
rect 7024 6322 7052 6666
rect 7472 6384 7524 6390
rect 7472 6326 7524 6332
rect 7012 6316 7064 6322
rect 7012 6258 7064 6264
rect 6920 5840 6972 5846
rect 6920 5782 6972 5788
rect 6736 5568 6788 5574
rect 6736 5510 6788 5516
rect 6552 4820 6604 4826
rect 6552 4762 6604 4768
rect 6460 4684 6512 4690
rect 6460 4626 6512 4632
rect 6748 4078 6776 5510
rect 6932 5234 6960 5782
rect 7024 5574 7052 6258
rect 7288 6112 7340 6118
rect 7288 6054 7340 6060
rect 7012 5568 7064 5574
rect 7012 5510 7064 5516
rect 7300 5302 7328 6054
rect 7484 5710 7512 6326
rect 8128 5778 8156 6734
rect 8576 6724 8628 6730
rect 8576 6666 8628 6672
rect 8214 6556 8522 6565
rect 8214 6554 8220 6556
rect 8276 6554 8300 6556
rect 8356 6554 8380 6556
rect 8436 6554 8460 6556
rect 8516 6554 8522 6556
rect 8276 6502 8278 6554
rect 8458 6502 8460 6554
rect 8214 6500 8220 6502
rect 8276 6500 8300 6502
rect 8356 6500 8380 6502
rect 8436 6500 8460 6502
rect 8516 6500 8522 6502
rect 8214 6491 8522 6500
rect 8588 6458 8616 6666
rect 8576 6452 8628 6458
rect 8576 6394 8628 6400
rect 8956 6254 8984 7346
rect 9508 7002 9536 7754
rect 9678 7440 9734 7449
rect 9678 7375 9680 7384
rect 9732 7375 9734 7384
rect 9680 7346 9732 7352
rect 9876 7342 9904 7822
rect 10428 7410 10456 8298
rect 10704 7750 10732 9046
rect 10888 8537 10916 9646
rect 10968 9580 11020 9586
rect 10968 9522 11020 9528
rect 10980 9110 11008 9522
rect 10968 9104 11020 9110
rect 10968 9046 11020 9052
rect 10874 8528 10930 8537
rect 10874 8463 10930 8472
rect 11164 8362 11192 10390
rect 11428 10192 11480 10198
rect 11428 10134 11480 10140
rect 11440 9625 11468 10134
rect 11532 9926 11560 10950
rect 11624 10606 11652 11562
rect 11716 11150 11744 11766
rect 11704 11144 11756 11150
rect 11704 11086 11756 11092
rect 11702 10704 11758 10713
rect 11702 10639 11758 10648
rect 11716 10606 11744 10639
rect 11612 10600 11664 10606
rect 11612 10542 11664 10548
rect 11704 10600 11756 10606
rect 11704 10542 11756 10548
rect 11704 9988 11756 9994
rect 11704 9930 11756 9936
rect 11520 9920 11572 9926
rect 11520 9862 11572 9868
rect 11426 9616 11482 9625
rect 11716 9586 11744 9930
rect 11808 9654 11836 12038
rect 11900 10674 11928 12310
rect 12360 12294 12572 12322
rect 11980 12096 12032 12102
rect 11980 12038 12032 12044
rect 11992 11762 12020 12038
rect 12162 11928 12218 11937
rect 12162 11863 12164 11872
rect 12216 11863 12218 11872
rect 12164 11834 12216 11840
rect 12360 11830 12388 12294
rect 12544 12238 12572 12294
rect 12440 12232 12492 12238
rect 12440 12174 12492 12180
rect 12532 12232 12584 12238
rect 12532 12174 12584 12180
rect 12348 11824 12400 11830
rect 12254 11792 12310 11801
rect 11980 11756 12032 11762
rect 12348 11766 12400 11772
rect 12254 11727 12310 11736
rect 11980 11698 12032 11704
rect 12072 11688 12124 11694
rect 12268 11676 12296 11727
rect 12452 11676 12480 12174
rect 12636 11676 12664 13262
rect 12728 13258 12756 13670
rect 12716 13252 12768 13258
rect 12716 13194 12768 13200
rect 12728 12714 12756 13194
rect 12716 12708 12768 12714
rect 12716 12650 12768 12656
rect 12808 12436 12860 12442
rect 12808 12378 12860 12384
rect 12716 12368 12768 12374
rect 12716 12310 12768 12316
rect 12728 11744 12756 12310
rect 12820 12102 12848 12378
rect 12912 12374 12940 14200
rect 13820 13456 13872 13462
rect 13820 13398 13872 13404
rect 13084 13320 13136 13326
rect 13084 13262 13136 13268
rect 13096 12850 13124 13262
rect 13728 13184 13780 13190
rect 13728 13126 13780 13132
rect 13084 12844 13136 12850
rect 13084 12786 13136 12792
rect 13096 12442 13124 12786
rect 13740 12442 13768 13126
rect 13832 12918 13860 13398
rect 14188 13320 14240 13326
rect 14188 13262 14240 13268
rect 13820 12912 13872 12918
rect 13820 12854 13872 12860
rect 13912 12844 13964 12850
rect 13912 12786 13964 12792
rect 14004 12844 14056 12850
rect 14004 12786 14056 12792
rect 13084 12436 13136 12442
rect 13084 12378 13136 12384
rect 13728 12436 13780 12442
rect 13728 12378 13780 12384
rect 12900 12368 12952 12374
rect 12900 12310 12952 12316
rect 12912 12238 12940 12310
rect 12992 12300 13044 12306
rect 12992 12242 13044 12248
rect 12900 12232 12952 12238
rect 13004 12209 13032 12242
rect 13084 12232 13136 12238
rect 12900 12174 12952 12180
rect 12990 12200 13046 12209
rect 13084 12174 13136 12180
rect 13636 12232 13688 12238
rect 13636 12174 13688 12180
rect 12990 12135 13046 12144
rect 12808 12096 12860 12102
rect 12808 12038 12860 12044
rect 12728 11716 12848 11744
rect 12268 11648 12388 11676
rect 12452 11648 12756 11676
rect 12072 11630 12124 11636
rect 12084 11393 12112 11630
rect 12360 11540 12388 11648
rect 12624 11552 12676 11558
rect 12360 11512 12624 11540
rect 12624 11494 12676 11500
rect 12214 11452 12522 11461
rect 12214 11450 12220 11452
rect 12276 11450 12300 11452
rect 12356 11450 12380 11452
rect 12436 11450 12460 11452
rect 12516 11450 12522 11452
rect 12276 11398 12278 11450
rect 12458 11398 12460 11450
rect 12214 11396 12220 11398
rect 12276 11396 12300 11398
rect 12356 11396 12380 11398
rect 12436 11396 12460 11398
rect 12516 11396 12522 11398
rect 12070 11384 12126 11393
rect 12214 11387 12522 11396
rect 12070 11319 12126 11328
rect 12636 11286 12664 11494
rect 12624 11280 12676 11286
rect 12624 11222 12676 11228
rect 12440 11144 12492 11150
rect 12492 11104 12664 11132
rect 12440 11086 12492 11092
rect 12348 11008 12400 11014
rect 12348 10950 12400 10956
rect 12162 10840 12218 10849
rect 12162 10775 12218 10784
rect 12256 10804 12308 10810
rect 12176 10674 12204 10775
rect 12256 10746 12308 10752
rect 12268 10713 12296 10746
rect 12360 10742 12388 10950
rect 12348 10736 12400 10742
rect 12254 10704 12310 10713
rect 11888 10668 11940 10674
rect 12164 10668 12216 10674
rect 11888 10610 11940 10616
rect 11992 10628 12164 10656
rect 11992 10266 12020 10628
rect 12348 10678 12400 10684
rect 12532 10736 12584 10742
rect 12532 10678 12584 10684
rect 12254 10639 12310 10648
rect 12164 10610 12216 10616
rect 12544 10577 12572 10678
rect 12636 10674 12664 11104
rect 12624 10668 12676 10674
rect 12624 10610 12676 10616
rect 12530 10568 12586 10577
rect 12636 10538 12664 10610
rect 12530 10503 12586 10512
rect 12624 10532 12676 10538
rect 12624 10474 12676 10480
rect 12214 10364 12522 10373
rect 12214 10362 12220 10364
rect 12276 10362 12300 10364
rect 12356 10362 12380 10364
rect 12436 10362 12460 10364
rect 12516 10362 12522 10364
rect 12276 10310 12278 10362
rect 12458 10310 12460 10362
rect 12214 10308 12220 10310
rect 12276 10308 12300 10310
rect 12356 10308 12380 10310
rect 12436 10308 12460 10310
rect 12516 10308 12522 10310
rect 12214 10299 12522 10308
rect 11980 10260 12032 10266
rect 11980 10202 12032 10208
rect 11886 10024 11942 10033
rect 11886 9959 11942 9968
rect 11796 9648 11848 9654
rect 11796 9590 11848 9596
rect 11426 9551 11482 9560
rect 11704 9580 11756 9586
rect 11704 9522 11756 9528
rect 11716 8974 11744 9522
rect 11900 9518 11928 9959
rect 12072 9920 12124 9926
rect 12072 9862 12124 9868
rect 12624 9920 12676 9926
rect 12624 9862 12676 9868
rect 11888 9512 11940 9518
rect 11940 9472 12020 9500
rect 11888 9454 11940 9460
rect 11704 8968 11756 8974
rect 11704 8910 11756 8916
rect 11888 8900 11940 8906
rect 11888 8842 11940 8848
rect 11900 8809 11928 8842
rect 11886 8800 11942 8809
rect 11886 8735 11942 8744
rect 11702 8664 11758 8673
rect 11702 8599 11758 8608
rect 11426 8392 11482 8401
rect 11152 8356 11204 8362
rect 11716 8362 11744 8599
rect 11426 8327 11482 8336
rect 11704 8356 11756 8362
rect 11152 8298 11204 8304
rect 11440 7954 11468 8327
rect 11704 8298 11756 8304
rect 11992 8294 12020 9472
rect 12084 9160 12112 9862
rect 12636 9586 12664 9862
rect 12532 9580 12584 9586
rect 12532 9522 12584 9528
rect 12624 9580 12676 9586
rect 12624 9522 12676 9528
rect 12544 9466 12572 9522
rect 12544 9438 12664 9466
rect 12728 9450 12756 11648
rect 12820 11558 12848 11716
rect 12898 11656 12954 11665
rect 12898 11591 12954 11600
rect 12808 11552 12860 11558
rect 12808 11494 12860 11500
rect 12912 11218 12940 11591
rect 12992 11348 13044 11354
rect 12992 11290 13044 11296
rect 12900 11212 12952 11218
rect 12900 11154 12952 11160
rect 13004 10554 13032 11290
rect 13096 10674 13124 12174
rect 13360 11552 13412 11558
rect 13360 11494 13412 11500
rect 13544 11552 13596 11558
rect 13544 11494 13596 11500
rect 13268 11212 13320 11218
rect 13268 11154 13320 11160
rect 13176 11144 13228 11150
rect 13280 11121 13308 11154
rect 13176 11086 13228 11092
rect 13266 11112 13322 11121
rect 13188 10742 13216 11086
rect 13266 11047 13322 11056
rect 13176 10736 13228 10742
rect 13176 10678 13228 10684
rect 13280 10674 13308 11047
rect 13372 10742 13400 11494
rect 13452 11144 13504 11150
rect 13452 11086 13504 11092
rect 13464 10985 13492 11086
rect 13450 10976 13506 10985
rect 13450 10911 13506 10920
rect 13360 10736 13412 10742
rect 13360 10678 13412 10684
rect 13084 10668 13136 10674
rect 13084 10610 13136 10616
rect 13268 10668 13320 10674
rect 13268 10610 13320 10616
rect 12912 10538 13032 10554
rect 12900 10532 13032 10538
rect 12952 10526 13032 10532
rect 13096 10554 13124 10610
rect 13096 10526 13400 10554
rect 12900 10474 12952 10480
rect 12808 10464 12860 10470
rect 12808 10406 12860 10412
rect 12820 10198 12848 10406
rect 12808 10192 12860 10198
rect 12808 10134 12860 10140
rect 12820 10062 12848 10134
rect 12808 10056 12860 10062
rect 12808 9998 12860 10004
rect 12636 9330 12664 9438
rect 12716 9444 12768 9450
rect 12716 9386 12768 9392
rect 12808 9444 12860 9450
rect 12808 9386 12860 9392
rect 12820 9330 12848 9386
rect 12636 9302 12848 9330
rect 12214 9276 12522 9285
rect 12214 9274 12220 9276
rect 12276 9274 12300 9276
rect 12356 9274 12380 9276
rect 12436 9274 12460 9276
rect 12516 9274 12522 9276
rect 12276 9222 12278 9274
rect 12458 9222 12460 9274
rect 12214 9220 12220 9222
rect 12276 9220 12300 9222
rect 12356 9220 12380 9222
rect 12436 9220 12460 9222
rect 12516 9220 12522 9222
rect 12214 9211 12522 9220
rect 12440 9172 12492 9178
rect 12084 9132 12204 9160
rect 12176 8974 12204 9132
rect 12440 9114 12492 9120
rect 12452 9042 12480 9114
rect 12532 9104 12584 9110
rect 12532 9046 12584 9052
rect 12440 9036 12492 9042
rect 12440 8978 12492 8984
rect 12164 8968 12216 8974
rect 12164 8910 12216 8916
rect 12176 8430 12204 8910
rect 12256 8560 12308 8566
rect 12254 8528 12256 8537
rect 12308 8528 12310 8537
rect 12544 8514 12572 9046
rect 12808 8968 12860 8974
rect 12912 8945 12940 10474
rect 13268 10192 13320 10198
rect 13268 10134 13320 10140
rect 13280 10062 13308 10134
rect 13268 10056 13320 10062
rect 13268 9998 13320 10004
rect 13084 9920 13136 9926
rect 13084 9862 13136 9868
rect 13176 9920 13228 9926
rect 13176 9862 13228 9868
rect 13096 9518 13124 9862
rect 13188 9586 13216 9862
rect 13176 9580 13228 9586
rect 13176 9522 13228 9528
rect 13084 9512 13136 9518
rect 13084 9454 13136 9460
rect 13096 9110 13124 9454
rect 13084 9104 13136 9110
rect 13084 9046 13136 9052
rect 12992 9036 13044 9042
rect 12992 8978 13044 8984
rect 12808 8910 12860 8916
rect 12898 8936 12954 8945
rect 12716 8832 12768 8838
rect 12716 8774 12768 8780
rect 12452 8498 12572 8514
rect 12254 8463 12310 8472
rect 12440 8492 12572 8498
rect 12492 8486 12572 8492
rect 12440 8434 12492 8440
rect 12164 8424 12216 8430
rect 12164 8366 12216 8372
rect 11520 8288 11572 8294
rect 11520 8230 11572 8236
rect 11980 8288 12032 8294
rect 11980 8230 12032 8236
rect 11532 7993 11560 8230
rect 11518 7984 11574 7993
rect 11428 7948 11480 7954
rect 11518 7919 11574 7928
rect 11428 7890 11480 7896
rect 10508 7744 10560 7750
rect 10508 7686 10560 7692
rect 10692 7744 10744 7750
rect 10692 7686 10744 7692
rect 10520 7449 10548 7686
rect 10506 7440 10562 7449
rect 9956 7404 10008 7410
rect 9956 7346 10008 7352
rect 10416 7404 10468 7410
rect 10506 7375 10508 7384
rect 10416 7346 10468 7352
rect 10560 7375 10562 7384
rect 10508 7346 10560 7352
rect 9588 7336 9640 7342
rect 9588 7278 9640 7284
rect 9864 7336 9916 7342
rect 9864 7278 9916 7284
rect 9496 6996 9548 7002
rect 9496 6938 9548 6944
rect 9128 6724 9180 6730
rect 9128 6666 9180 6672
rect 9140 6458 9168 6666
rect 9128 6452 9180 6458
rect 9128 6394 9180 6400
rect 8484 6248 8536 6254
rect 8484 6190 8536 6196
rect 8944 6248 8996 6254
rect 8944 6190 8996 6196
rect 8496 5914 8524 6190
rect 8484 5908 8536 5914
rect 8484 5850 8536 5856
rect 8760 5908 8812 5914
rect 8760 5850 8812 5856
rect 8116 5772 8168 5778
rect 8116 5714 8168 5720
rect 7472 5704 7524 5710
rect 7472 5646 7524 5652
rect 8024 5704 8076 5710
rect 8024 5646 8076 5652
rect 7932 5568 7984 5574
rect 7932 5510 7984 5516
rect 7288 5296 7340 5302
rect 7288 5238 7340 5244
rect 6920 5228 6972 5234
rect 6920 5170 6972 5176
rect 7944 4826 7972 5510
rect 7932 4820 7984 4826
rect 7932 4762 7984 4768
rect 7840 4684 7892 4690
rect 7840 4626 7892 4632
rect 7472 4208 7524 4214
rect 7472 4150 7524 4156
rect 6736 4072 6788 4078
rect 6736 4014 6788 4020
rect 6460 3936 6512 3942
rect 6460 3878 6512 3884
rect 6736 3936 6788 3942
rect 6736 3878 6788 3884
rect 6472 3738 6500 3878
rect 6368 3732 6420 3738
rect 6368 3674 6420 3680
rect 6460 3732 6512 3738
rect 6460 3674 6512 3680
rect 6644 3528 6696 3534
rect 6644 3470 6696 3476
rect 5724 2508 5776 2514
rect 5724 2450 5776 2456
rect 5920 2502 6040 2530
rect 5920 1970 5948 2502
rect 6000 2372 6052 2378
rect 6000 2314 6052 2320
rect 6460 2372 6512 2378
rect 6460 2314 6512 2320
rect 5908 1964 5960 1970
rect 5908 1906 5960 1912
rect 5920 1358 5948 1906
rect 6012 1562 6040 2314
rect 6472 2106 6500 2314
rect 6656 2106 6684 3470
rect 6748 3058 6776 3878
rect 7484 3602 7512 4150
rect 7748 4072 7800 4078
rect 7748 4014 7800 4020
rect 7472 3596 7524 3602
rect 7472 3538 7524 3544
rect 7104 3528 7156 3534
rect 7104 3470 7156 3476
rect 7656 3528 7708 3534
rect 7656 3470 7708 3476
rect 6736 3052 6788 3058
rect 6736 2994 6788 3000
rect 6460 2100 6512 2106
rect 6460 2042 6512 2048
rect 6644 2100 6696 2106
rect 6644 2042 6696 2048
rect 6748 1970 6776 2994
rect 7116 2990 7144 3470
rect 7380 3188 7432 3194
rect 7380 3130 7432 3136
rect 7104 2984 7156 2990
rect 7104 2926 7156 2932
rect 7392 2038 7420 3130
rect 7668 3058 7696 3470
rect 7760 3194 7788 4014
rect 7852 3534 7880 4626
rect 7840 3528 7892 3534
rect 7840 3470 7892 3476
rect 8036 3466 8064 5646
rect 8214 5468 8522 5477
rect 8214 5466 8220 5468
rect 8276 5466 8300 5468
rect 8356 5466 8380 5468
rect 8436 5466 8460 5468
rect 8516 5466 8522 5468
rect 8276 5414 8278 5466
rect 8458 5414 8460 5466
rect 8214 5412 8220 5414
rect 8276 5412 8300 5414
rect 8356 5412 8380 5414
rect 8436 5412 8460 5414
rect 8516 5412 8522 5414
rect 8214 5403 8522 5412
rect 8772 5370 8800 5850
rect 9508 5778 9536 6938
rect 9600 5914 9628 7278
rect 9680 7200 9732 7206
rect 9680 7142 9732 7148
rect 9864 7200 9916 7206
rect 9864 7142 9916 7148
rect 9692 6798 9720 7142
rect 9876 7002 9904 7142
rect 9864 6996 9916 7002
rect 9864 6938 9916 6944
rect 9680 6792 9732 6798
rect 9680 6734 9732 6740
rect 9968 6186 9996 7346
rect 9956 6180 10008 6186
rect 9956 6122 10008 6128
rect 9680 6112 9732 6118
rect 9680 6054 9732 6060
rect 9588 5908 9640 5914
rect 9588 5850 9640 5856
rect 9496 5772 9548 5778
rect 9496 5714 9548 5720
rect 9600 5710 9628 5850
rect 9588 5704 9640 5710
rect 9588 5646 9640 5652
rect 9404 5636 9456 5642
rect 9404 5578 9456 5584
rect 8760 5364 8812 5370
rect 8760 5306 8812 5312
rect 9128 5296 9180 5302
rect 9128 5238 9180 5244
rect 9140 4690 9168 5238
rect 9128 4684 9180 4690
rect 9128 4626 9180 4632
rect 9312 4616 9364 4622
rect 9312 4558 9364 4564
rect 8576 4480 8628 4486
rect 8576 4422 8628 4428
rect 8214 4380 8522 4389
rect 8214 4378 8220 4380
rect 8276 4378 8300 4380
rect 8356 4378 8380 4380
rect 8436 4378 8460 4380
rect 8516 4378 8522 4380
rect 8276 4326 8278 4378
rect 8458 4326 8460 4378
rect 8214 4324 8220 4326
rect 8276 4324 8300 4326
rect 8356 4324 8380 4326
rect 8436 4324 8460 4326
rect 8516 4324 8522 4326
rect 8214 4315 8522 4324
rect 8588 4146 8616 4422
rect 9324 4214 9352 4558
rect 9312 4208 9364 4214
rect 9312 4150 9364 4156
rect 8576 4140 8628 4146
rect 8576 4082 8628 4088
rect 8484 4004 8536 4010
rect 8484 3946 8536 3952
rect 8496 3534 8524 3946
rect 8588 3602 8616 4082
rect 9324 4010 9352 4150
rect 9312 4004 9364 4010
rect 9312 3946 9364 3952
rect 9220 3936 9272 3942
rect 9220 3878 9272 3884
rect 8576 3596 8628 3602
rect 8576 3538 8628 3544
rect 8484 3528 8536 3534
rect 8484 3470 8536 3476
rect 8668 3528 8720 3534
rect 8668 3470 8720 3476
rect 8024 3460 8076 3466
rect 8024 3402 8076 3408
rect 8036 3194 8064 3402
rect 8214 3292 8522 3301
rect 8214 3290 8220 3292
rect 8276 3290 8300 3292
rect 8356 3290 8380 3292
rect 8436 3290 8460 3292
rect 8516 3290 8522 3292
rect 8276 3238 8278 3290
rect 8458 3238 8460 3290
rect 8214 3236 8220 3238
rect 8276 3236 8300 3238
rect 8356 3236 8380 3238
rect 8436 3236 8460 3238
rect 8516 3236 8522 3238
rect 8214 3227 8522 3236
rect 7748 3188 7800 3194
rect 7748 3130 7800 3136
rect 8024 3188 8076 3194
rect 8024 3130 8076 3136
rect 7656 3052 7708 3058
rect 7656 2994 7708 3000
rect 8680 2802 8708 3470
rect 8760 3392 8812 3398
rect 8760 3334 8812 3340
rect 8772 3126 8800 3334
rect 9232 3194 9260 3878
rect 9416 3670 9444 5578
rect 9692 5302 9720 6054
rect 9968 5710 9996 6122
rect 9956 5704 10008 5710
rect 9956 5646 10008 5652
rect 10428 5370 10456 7346
rect 10704 7290 10732 7686
rect 11888 7540 11940 7546
rect 11888 7482 11940 7488
rect 11060 7404 11112 7410
rect 11060 7346 11112 7352
rect 10508 7268 10560 7274
rect 10508 7210 10560 7216
rect 10612 7262 10732 7290
rect 10876 7336 10928 7342
rect 10876 7278 10928 7284
rect 10520 6322 10548 7210
rect 10508 6316 10560 6322
rect 10508 6258 10560 6264
rect 10612 5778 10640 7262
rect 10692 7200 10744 7206
rect 10692 7142 10744 7148
rect 10704 6866 10732 7142
rect 10692 6860 10744 6866
rect 10692 6802 10744 6808
rect 10704 6322 10732 6802
rect 10888 6798 10916 7278
rect 11072 6798 11100 7346
rect 11900 6798 11928 7482
rect 11992 7410 12020 8230
rect 12214 8188 12522 8197
rect 12214 8186 12220 8188
rect 12276 8186 12300 8188
rect 12356 8186 12380 8188
rect 12436 8186 12460 8188
rect 12516 8186 12522 8188
rect 12276 8134 12278 8186
rect 12458 8134 12460 8186
rect 12214 8132 12220 8134
rect 12276 8132 12300 8134
rect 12356 8132 12380 8134
rect 12436 8132 12460 8134
rect 12516 8132 12522 8134
rect 12214 8123 12522 8132
rect 12728 7886 12756 8774
rect 12716 7880 12768 7886
rect 12716 7822 12768 7828
rect 12256 7812 12308 7818
rect 12256 7754 12308 7760
rect 12164 7744 12216 7750
rect 12164 7686 12216 7692
rect 12176 7546 12204 7686
rect 12164 7540 12216 7546
rect 12164 7482 12216 7488
rect 12268 7478 12296 7754
rect 12256 7472 12308 7478
rect 12256 7414 12308 7420
rect 11980 7404 12032 7410
rect 11980 7346 12032 7352
rect 12728 7342 12756 7822
rect 12716 7336 12768 7342
rect 12716 7278 12768 7284
rect 12214 7100 12522 7109
rect 12214 7098 12220 7100
rect 12276 7098 12300 7100
rect 12356 7098 12380 7100
rect 12436 7098 12460 7100
rect 12516 7098 12522 7100
rect 12276 7046 12278 7098
rect 12458 7046 12460 7098
rect 12214 7044 12220 7046
rect 12276 7044 12300 7046
rect 12356 7044 12380 7046
rect 12436 7044 12460 7046
rect 12516 7044 12522 7046
rect 12214 7035 12522 7044
rect 10876 6792 10928 6798
rect 10876 6734 10928 6740
rect 11060 6792 11112 6798
rect 11060 6734 11112 6740
rect 11888 6792 11940 6798
rect 11888 6734 11940 6740
rect 12256 6792 12308 6798
rect 12256 6734 12308 6740
rect 11072 6390 11100 6734
rect 12164 6656 12216 6662
rect 12164 6598 12216 6604
rect 12176 6458 12204 6598
rect 12164 6452 12216 6458
rect 12164 6394 12216 6400
rect 12268 6390 12296 6734
rect 12716 6656 12768 6662
rect 12716 6598 12768 6604
rect 11060 6384 11112 6390
rect 11060 6326 11112 6332
rect 12256 6384 12308 6390
rect 12256 6326 12308 6332
rect 10692 6316 10744 6322
rect 10692 6258 10744 6264
rect 11520 6112 11572 6118
rect 11520 6054 11572 6060
rect 10600 5772 10652 5778
rect 10600 5714 10652 5720
rect 11532 5710 11560 6054
rect 12214 6012 12522 6021
rect 12214 6010 12220 6012
rect 12276 6010 12300 6012
rect 12356 6010 12380 6012
rect 12436 6010 12460 6012
rect 12516 6010 12522 6012
rect 12276 5958 12278 6010
rect 12458 5958 12460 6010
rect 12214 5956 12220 5958
rect 12276 5956 12300 5958
rect 12356 5956 12380 5958
rect 12436 5956 12460 5958
rect 12516 5956 12522 5958
rect 12214 5947 12522 5956
rect 11520 5704 11572 5710
rect 11520 5646 11572 5652
rect 11336 5568 11388 5574
rect 11336 5510 11388 5516
rect 10416 5364 10468 5370
rect 10416 5306 10468 5312
rect 11348 5302 11376 5510
rect 9680 5296 9732 5302
rect 9680 5238 9732 5244
rect 10140 5296 10192 5302
rect 10140 5238 10192 5244
rect 11336 5296 11388 5302
rect 11336 5238 11388 5244
rect 12624 5296 12676 5302
rect 12624 5238 12676 5244
rect 9772 5160 9824 5166
rect 9772 5102 9824 5108
rect 9680 4072 9732 4078
rect 9680 4014 9732 4020
rect 9404 3664 9456 3670
rect 9404 3606 9456 3612
rect 9416 3534 9444 3606
rect 9404 3528 9456 3534
rect 9404 3470 9456 3476
rect 9496 3392 9548 3398
rect 9496 3334 9548 3340
rect 9220 3188 9272 3194
rect 9220 3130 9272 3136
rect 8760 3120 8812 3126
rect 8760 3062 8812 3068
rect 8760 2848 8812 2854
rect 8680 2796 8760 2802
rect 8680 2790 8812 2796
rect 8680 2774 8800 2790
rect 8680 2446 8708 2774
rect 9232 2446 9260 3130
rect 9508 3126 9536 3334
rect 9496 3120 9548 3126
rect 9496 3062 9548 3068
rect 7564 2440 7616 2446
rect 7564 2382 7616 2388
rect 8668 2440 8720 2446
rect 8668 2382 8720 2388
rect 9220 2440 9272 2446
rect 9220 2382 9272 2388
rect 7380 2032 7432 2038
rect 7380 1974 7432 1980
rect 7576 1970 7604 2382
rect 7748 2372 7800 2378
rect 7748 2314 7800 2320
rect 6736 1964 6788 1970
rect 7564 1964 7616 1970
rect 6736 1906 6788 1912
rect 7484 1924 7564 1952
rect 6000 1556 6052 1562
rect 6000 1498 6052 1504
rect 5908 1352 5960 1358
rect 5908 1294 5960 1300
rect 7484 1290 7512 1924
rect 7564 1906 7616 1912
rect 7760 1902 7788 2314
rect 8576 2304 8628 2310
rect 8576 2246 8628 2252
rect 9220 2304 9272 2310
rect 9220 2246 9272 2252
rect 8214 2204 8522 2213
rect 8214 2202 8220 2204
rect 8276 2202 8300 2204
rect 8356 2202 8380 2204
rect 8436 2202 8460 2204
rect 8516 2202 8522 2204
rect 8276 2150 8278 2202
rect 8458 2150 8460 2202
rect 8214 2148 8220 2150
rect 8276 2148 8300 2150
rect 8356 2148 8380 2150
rect 8436 2148 8460 2150
rect 8516 2148 8522 2150
rect 8214 2139 8522 2148
rect 8588 2106 8616 2246
rect 8576 2100 8628 2106
rect 8576 2042 8628 2048
rect 7748 1896 7800 1902
rect 7748 1838 7800 1844
rect 7760 1426 7788 1838
rect 7748 1420 7800 1426
rect 7748 1362 7800 1368
rect 8588 1358 8616 2042
rect 9232 2038 9260 2246
rect 9220 2032 9272 2038
rect 9220 1974 9272 1980
rect 9404 1896 9456 1902
rect 9404 1838 9456 1844
rect 9220 1760 9272 1766
rect 9220 1702 9272 1708
rect 9232 1358 9260 1702
rect 9416 1426 9444 1838
rect 9404 1420 9456 1426
rect 9404 1362 9456 1368
rect 9692 1358 9720 4014
rect 9784 3058 9812 5102
rect 10152 4758 10180 5238
rect 11980 5160 12032 5166
rect 11980 5102 12032 5108
rect 10140 4752 10192 4758
rect 10140 4694 10192 4700
rect 11992 4690 12020 5102
rect 12214 4924 12522 4933
rect 12214 4922 12220 4924
rect 12276 4922 12300 4924
rect 12356 4922 12380 4924
rect 12436 4922 12460 4924
rect 12516 4922 12522 4924
rect 12276 4870 12278 4922
rect 12458 4870 12460 4922
rect 12214 4868 12220 4870
rect 12276 4868 12300 4870
rect 12356 4868 12380 4870
rect 12436 4868 12460 4870
rect 12516 4868 12522 4870
rect 12214 4859 12522 4868
rect 11980 4684 12032 4690
rect 11980 4626 12032 4632
rect 10876 4548 10928 4554
rect 10876 4490 10928 4496
rect 11980 4548 12032 4554
rect 11980 4490 12032 4496
rect 9864 4140 9916 4146
rect 9864 4082 9916 4088
rect 10416 4140 10468 4146
rect 10416 4082 10468 4088
rect 10600 4140 10652 4146
rect 10600 4082 10652 4088
rect 9876 3534 9904 4082
rect 10428 3942 10456 4082
rect 10416 3936 10468 3942
rect 10416 3878 10468 3884
rect 10428 3534 10456 3878
rect 9864 3528 9916 3534
rect 9864 3470 9916 3476
rect 10416 3528 10468 3534
rect 10416 3470 10468 3476
rect 10612 3398 10640 4082
rect 10888 4078 10916 4490
rect 11992 4282 12020 4490
rect 12636 4282 12664 5238
rect 12728 4554 12756 6598
rect 12820 6254 12848 8910
rect 12898 8871 12954 8880
rect 12900 8356 12952 8362
rect 12900 8298 12952 8304
rect 12912 8090 12940 8298
rect 12900 8084 12952 8090
rect 12900 8026 12952 8032
rect 13004 7886 13032 8978
rect 13084 8968 13136 8974
rect 13084 8910 13136 8916
rect 13096 8022 13124 8910
rect 13188 8498 13216 9522
rect 13176 8492 13228 8498
rect 13176 8434 13228 8440
rect 13280 8378 13308 9998
rect 13188 8350 13308 8378
rect 13372 9602 13400 10526
rect 13464 9722 13492 10911
rect 13556 10266 13584 11494
rect 13648 11354 13676 12174
rect 13820 11892 13872 11898
rect 13820 11834 13872 11840
rect 13832 11354 13860 11834
rect 13924 11830 13952 12786
rect 14016 12646 14044 12786
rect 14004 12640 14056 12646
rect 14004 12582 14056 12588
rect 13912 11824 13964 11830
rect 13912 11766 13964 11772
rect 13636 11348 13688 11354
rect 13636 11290 13688 11296
rect 13820 11348 13872 11354
rect 13820 11290 13872 11296
rect 13832 11234 13860 11290
rect 13832 11206 13952 11234
rect 13728 11144 13780 11150
rect 13728 11086 13780 11092
rect 13636 11008 13688 11014
rect 13636 10950 13688 10956
rect 13648 10742 13676 10950
rect 13636 10736 13688 10742
rect 13636 10678 13688 10684
rect 13544 10260 13596 10266
rect 13544 10202 13596 10208
rect 13452 9716 13504 9722
rect 13452 9658 13504 9664
rect 13372 9586 13492 9602
rect 13372 9580 13504 9586
rect 13372 9574 13452 9580
rect 13084 8016 13136 8022
rect 13084 7958 13136 7964
rect 12992 7880 13044 7886
rect 12992 7822 13044 7828
rect 13188 7478 13216 8350
rect 13268 8016 13320 8022
rect 13268 7958 13320 7964
rect 13176 7472 13228 7478
rect 13176 7414 13228 7420
rect 13084 7200 13136 7206
rect 13084 7142 13136 7148
rect 13096 6662 13124 7142
rect 13280 6934 13308 7958
rect 13372 7834 13400 9574
rect 13452 9522 13504 9528
rect 13556 9466 13584 10202
rect 13740 10062 13768 11086
rect 13820 11076 13872 11082
rect 13820 11018 13872 11024
rect 13832 10742 13860 11018
rect 13820 10736 13872 10742
rect 13820 10678 13872 10684
rect 13924 10470 13952 11206
rect 14016 10713 14044 12582
rect 14200 12238 14228 13262
rect 14280 12436 14332 12442
rect 14280 12378 14332 12384
rect 14188 12232 14240 12238
rect 14188 12174 14240 12180
rect 14094 12064 14150 12073
rect 14094 11999 14150 12008
rect 14108 11898 14136 11999
rect 14096 11892 14148 11898
rect 14096 11834 14148 11840
rect 14096 11756 14148 11762
rect 14096 11698 14148 11704
rect 14002 10704 14058 10713
rect 14002 10639 14058 10648
rect 13912 10464 13964 10470
rect 13912 10406 13964 10412
rect 13728 10056 13780 10062
rect 13728 9998 13780 10004
rect 13740 9586 13768 9998
rect 14004 9648 14056 9654
rect 14004 9590 14056 9596
rect 13728 9580 13780 9586
rect 13728 9522 13780 9528
rect 14016 9489 14044 9590
rect 13464 9438 13584 9466
rect 14002 9480 14058 9489
rect 13464 8974 13492 9438
rect 14002 9415 14058 9424
rect 13544 9376 13596 9382
rect 13544 9318 13596 9324
rect 13636 9376 13688 9382
rect 13636 9318 13688 9324
rect 13820 9376 13872 9382
rect 13820 9318 13872 9324
rect 13556 9178 13584 9318
rect 13544 9172 13596 9178
rect 13544 9114 13596 9120
rect 13452 8968 13504 8974
rect 13452 8910 13504 8916
rect 13648 8906 13676 9318
rect 13832 8956 13860 9318
rect 13910 9072 13966 9081
rect 13910 9007 13966 9016
rect 13740 8928 13860 8956
rect 13636 8900 13688 8906
rect 13636 8842 13688 8848
rect 13450 8392 13506 8401
rect 13450 8327 13452 8336
rect 13504 8327 13506 8336
rect 13544 8356 13596 8362
rect 13452 8298 13504 8304
rect 13544 8298 13596 8304
rect 13372 7806 13492 7834
rect 13464 7342 13492 7806
rect 13452 7336 13504 7342
rect 13452 7278 13504 7284
rect 13268 6928 13320 6934
rect 13268 6870 13320 6876
rect 13084 6656 13136 6662
rect 13084 6598 13136 6604
rect 13280 6254 13308 6870
rect 13464 6780 13492 7278
rect 13556 7274 13584 8298
rect 13648 8294 13676 8842
rect 13740 8537 13768 8928
rect 13820 8832 13872 8838
rect 13820 8774 13872 8780
rect 13726 8528 13782 8537
rect 13832 8498 13860 8774
rect 13924 8566 13952 9007
rect 14108 8974 14136 11698
rect 14200 10266 14228 12174
rect 14292 11830 14320 12378
rect 14280 11824 14332 11830
rect 14280 11766 14332 11772
rect 14384 11762 14412 14200
rect 15198 13560 15254 13569
rect 15198 13495 15254 13504
rect 14648 13252 14700 13258
rect 14648 13194 14700 13200
rect 14660 12918 14688 13194
rect 14648 12912 14700 12918
rect 14648 12854 14700 12860
rect 15212 12306 15240 13495
rect 15384 13320 15436 13326
rect 15384 13262 15436 13268
rect 15396 12646 15424 13262
rect 15752 13184 15804 13190
rect 15752 13126 15804 13132
rect 15476 12912 15528 12918
rect 15476 12854 15528 12860
rect 15384 12640 15436 12646
rect 15384 12582 15436 12588
rect 15200 12300 15252 12306
rect 15200 12242 15252 12248
rect 15396 12238 15424 12582
rect 15488 12374 15516 12854
rect 15764 12850 15792 13126
rect 15752 12844 15804 12850
rect 15752 12786 15804 12792
rect 15856 12434 15884 14200
rect 17328 13734 17356 14200
rect 17316 13728 17368 13734
rect 17316 13670 17368 13676
rect 17224 13388 17276 13394
rect 17224 13330 17276 13336
rect 16764 13320 16816 13326
rect 16764 13262 16816 13268
rect 16028 13252 16080 13258
rect 16028 13194 16080 13200
rect 16040 12714 16068 13194
rect 16214 13084 16522 13093
rect 16214 13082 16220 13084
rect 16276 13082 16300 13084
rect 16356 13082 16380 13084
rect 16436 13082 16460 13084
rect 16516 13082 16522 13084
rect 16276 13030 16278 13082
rect 16458 13030 16460 13082
rect 16214 13028 16220 13030
rect 16276 13028 16300 13030
rect 16356 13028 16380 13030
rect 16436 13028 16460 13030
rect 16516 13028 16522 13030
rect 16214 13019 16522 13028
rect 16776 12986 16804 13262
rect 16764 12980 16816 12986
rect 16764 12922 16816 12928
rect 17040 12844 17092 12850
rect 17040 12786 17092 12792
rect 16028 12708 16080 12714
rect 16028 12650 16080 12656
rect 15764 12406 15884 12434
rect 15476 12368 15528 12374
rect 15476 12310 15528 12316
rect 15384 12232 15436 12238
rect 15384 12174 15436 12180
rect 15292 12164 15344 12170
rect 15292 12106 15344 12112
rect 14832 12096 14884 12102
rect 14832 12038 14884 12044
rect 14372 11756 14424 11762
rect 14372 11698 14424 11704
rect 14280 11008 14332 11014
rect 14280 10950 14332 10956
rect 14292 10606 14320 10950
rect 14280 10600 14332 10606
rect 14280 10542 14332 10548
rect 14188 10260 14240 10266
rect 14188 10202 14240 10208
rect 14188 10124 14240 10130
rect 14188 10066 14240 10072
rect 14004 8968 14056 8974
rect 14004 8910 14056 8916
rect 14096 8968 14148 8974
rect 14096 8910 14148 8916
rect 14016 8616 14044 8910
rect 14108 8838 14136 8910
rect 14096 8832 14148 8838
rect 14096 8774 14148 8780
rect 14016 8588 14136 8616
rect 13912 8560 13964 8566
rect 13964 8520 14044 8548
rect 13912 8502 13964 8508
rect 13726 8463 13782 8472
rect 13820 8492 13872 8498
rect 13820 8434 13872 8440
rect 13636 8288 13688 8294
rect 13636 8230 13688 8236
rect 13832 7410 13860 8434
rect 13820 7404 13872 7410
rect 13820 7346 13872 7352
rect 13544 7268 13596 7274
rect 13544 7210 13596 7216
rect 13728 7200 13780 7206
rect 13728 7142 13780 7148
rect 13740 6798 13768 7142
rect 13544 6792 13596 6798
rect 13464 6752 13544 6780
rect 13544 6734 13596 6740
rect 13728 6792 13780 6798
rect 13728 6734 13780 6740
rect 12808 6248 12860 6254
rect 12808 6190 12860 6196
rect 13268 6248 13320 6254
rect 13268 6190 13320 6196
rect 12820 5370 12848 6190
rect 12808 5364 12860 5370
rect 12808 5306 12860 5312
rect 13556 4826 13584 6734
rect 14016 6202 14044 8520
rect 14108 8498 14136 8588
rect 14096 8492 14148 8498
rect 14096 8434 14148 8440
rect 14200 8022 14228 10066
rect 14280 9580 14332 9586
rect 14280 9522 14332 9528
rect 14292 9110 14320 9522
rect 14280 9104 14332 9110
rect 14280 9046 14332 9052
rect 14384 8090 14412 11698
rect 14648 11552 14700 11558
rect 14648 11494 14700 11500
rect 14660 11218 14688 11494
rect 14648 11212 14700 11218
rect 14648 11154 14700 11160
rect 14844 11150 14872 12038
rect 14924 11824 14976 11830
rect 14924 11766 14976 11772
rect 15016 11824 15068 11830
rect 15016 11766 15068 11772
rect 14936 11626 14964 11766
rect 14924 11620 14976 11626
rect 14924 11562 14976 11568
rect 14832 11144 14884 11150
rect 14832 11086 14884 11092
rect 14924 10804 14976 10810
rect 14924 10746 14976 10752
rect 14464 10736 14516 10742
rect 14464 10678 14516 10684
rect 14476 9450 14504 10678
rect 14556 10600 14608 10606
rect 14556 10542 14608 10548
rect 14568 9976 14596 10542
rect 14936 10198 14964 10746
rect 15028 10470 15056 11766
rect 15304 11354 15332 12106
rect 15384 11892 15436 11898
rect 15384 11834 15436 11840
rect 15292 11348 15344 11354
rect 15292 11290 15344 11296
rect 15200 11280 15252 11286
rect 15200 11222 15252 11228
rect 15212 10810 15240 11222
rect 15200 10804 15252 10810
rect 15200 10746 15252 10752
rect 15292 10668 15344 10674
rect 15292 10610 15344 10616
rect 15016 10464 15068 10470
rect 15016 10406 15068 10412
rect 14924 10192 14976 10198
rect 14924 10134 14976 10140
rect 15028 10130 15056 10406
rect 15106 10160 15162 10169
rect 15016 10124 15068 10130
rect 15106 10095 15162 10104
rect 15016 10066 15068 10072
rect 15120 10062 15148 10095
rect 14740 10056 14792 10062
rect 14740 9998 14792 10004
rect 14832 10056 14884 10062
rect 14832 9998 14884 10004
rect 15108 10056 15160 10062
rect 15108 9998 15160 10004
rect 14648 9988 14700 9994
rect 14568 9948 14648 9976
rect 14568 9586 14596 9948
rect 14648 9930 14700 9936
rect 14752 9722 14780 9998
rect 14740 9716 14792 9722
rect 14740 9658 14792 9664
rect 14556 9580 14608 9586
rect 14556 9522 14608 9528
rect 14752 9450 14780 9658
rect 14464 9444 14516 9450
rect 14464 9386 14516 9392
rect 14740 9444 14792 9450
rect 14740 9386 14792 9392
rect 14476 9110 14504 9386
rect 14464 9104 14516 9110
rect 14464 9046 14516 9052
rect 14556 8968 14608 8974
rect 14554 8936 14556 8945
rect 14608 8936 14610 8945
rect 14554 8871 14610 8880
rect 14568 8362 14596 8871
rect 14844 8566 14872 9998
rect 15120 9674 15148 9998
rect 15120 9646 15240 9674
rect 15304 9654 15332 10610
rect 15396 10130 15424 11834
rect 15764 11762 15792 12406
rect 16040 12238 16068 12650
rect 17052 12442 17080 12786
rect 17040 12436 17092 12442
rect 17040 12378 17092 12384
rect 16028 12232 16080 12238
rect 16028 12174 16080 12180
rect 16948 12232 17000 12238
rect 16948 12174 17000 12180
rect 16028 12096 16080 12102
rect 16028 12038 16080 12044
rect 16120 12096 16172 12102
rect 16120 12038 16172 12044
rect 16764 12096 16816 12102
rect 16764 12038 16816 12044
rect 15752 11756 15804 11762
rect 15752 11698 15804 11704
rect 15476 11688 15528 11694
rect 15476 11630 15528 11636
rect 15568 11688 15620 11694
rect 15568 11630 15620 11636
rect 15488 10810 15516 11630
rect 15580 11286 15608 11630
rect 15568 11280 15620 11286
rect 15568 11222 15620 11228
rect 15568 11076 15620 11082
rect 15568 11018 15620 11024
rect 15476 10804 15528 10810
rect 15476 10746 15528 10752
rect 15476 10668 15528 10674
rect 15476 10610 15528 10616
rect 15384 10124 15436 10130
rect 15384 10066 15436 10072
rect 15212 9586 15240 9646
rect 15292 9648 15344 9654
rect 15292 9590 15344 9596
rect 15200 9580 15252 9586
rect 15200 9522 15252 9528
rect 15384 9580 15436 9586
rect 15384 9522 15436 9528
rect 15212 9058 15240 9522
rect 15396 9450 15424 9522
rect 15384 9444 15436 9450
rect 15384 9386 15436 9392
rect 15212 9030 15332 9058
rect 15198 8936 15254 8945
rect 15198 8871 15254 8880
rect 15016 8832 15068 8838
rect 15212 8786 15240 8871
rect 15016 8774 15068 8780
rect 15028 8673 15056 8774
rect 15120 8758 15240 8786
rect 15014 8664 15070 8673
rect 15120 8634 15148 8758
rect 15014 8599 15070 8608
rect 15108 8628 15160 8634
rect 15108 8570 15160 8576
rect 15200 8628 15252 8634
rect 15200 8570 15252 8576
rect 14832 8560 14884 8566
rect 15212 8514 15240 8570
rect 14832 8502 14884 8508
rect 15120 8498 15240 8514
rect 15304 8498 15332 9030
rect 15108 8492 15240 8498
rect 15160 8486 15240 8492
rect 15292 8492 15344 8498
rect 15108 8434 15160 8440
rect 15292 8434 15344 8440
rect 14556 8356 14608 8362
rect 14556 8298 14608 8304
rect 14832 8288 14884 8294
rect 14832 8230 14884 8236
rect 14372 8084 14424 8090
rect 14372 8026 14424 8032
rect 14188 8016 14240 8022
rect 14844 7993 14872 8230
rect 14188 7958 14240 7964
rect 14830 7984 14886 7993
rect 14830 7919 14886 7928
rect 14844 7886 14872 7919
rect 14832 7880 14884 7886
rect 14832 7822 14884 7828
rect 15304 7546 15332 8434
rect 15396 8294 15424 9386
rect 15488 8945 15516 10610
rect 15580 9450 15608 11018
rect 15660 10056 15712 10062
rect 15660 9998 15712 10004
rect 15672 9586 15700 9998
rect 15660 9580 15712 9586
rect 15660 9522 15712 9528
rect 15672 9489 15700 9522
rect 15658 9480 15714 9489
rect 15568 9444 15620 9450
rect 15658 9415 15714 9424
rect 15568 9386 15620 9392
rect 15568 8968 15620 8974
rect 15474 8936 15530 8945
rect 15568 8910 15620 8916
rect 15474 8871 15530 8880
rect 15476 8832 15528 8838
rect 15476 8774 15528 8780
rect 15488 8566 15516 8774
rect 15476 8560 15528 8566
rect 15476 8502 15528 8508
rect 15384 8288 15436 8294
rect 15384 8230 15436 8236
rect 15292 7540 15344 7546
rect 15292 7482 15344 7488
rect 14096 7404 14148 7410
rect 14096 7346 14148 7352
rect 15200 7404 15252 7410
rect 15200 7346 15252 7352
rect 14108 7206 14136 7346
rect 15016 7268 15068 7274
rect 15016 7210 15068 7216
rect 14096 7200 14148 7206
rect 14096 7142 14148 7148
rect 14108 6866 14136 7142
rect 14096 6860 14148 6866
rect 14096 6802 14148 6808
rect 14108 6254 14136 6802
rect 14832 6384 14884 6390
rect 14832 6326 14884 6332
rect 13924 6174 14044 6202
rect 14096 6248 14148 6254
rect 14096 6190 14148 6196
rect 13924 5710 13952 6174
rect 14004 6112 14056 6118
rect 14004 6054 14056 6060
rect 13912 5704 13964 5710
rect 13912 5646 13964 5652
rect 13728 5636 13780 5642
rect 13728 5578 13780 5584
rect 13544 4820 13596 4826
rect 13544 4762 13596 4768
rect 13740 4622 13768 5578
rect 13820 4820 13872 4826
rect 13820 4762 13872 4768
rect 13728 4616 13780 4622
rect 13728 4558 13780 4564
rect 12716 4548 12768 4554
rect 12716 4490 12768 4496
rect 11980 4276 12032 4282
rect 11980 4218 12032 4224
rect 12624 4276 12676 4282
rect 12624 4218 12676 4224
rect 13740 4214 13768 4558
rect 13728 4208 13780 4214
rect 13728 4150 13780 4156
rect 13832 4146 13860 4762
rect 13924 4622 13952 5646
rect 14016 5302 14044 6054
rect 14188 5704 14240 5710
rect 14188 5646 14240 5652
rect 14740 5704 14792 5710
rect 14740 5646 14792 5652
rect 14004 5296 14056 5302
rect 14004 5238 14056 5244
rect 13912 4616 13964 4622
rect 13912 4558 13964 4564
rect 12440 4140 12492 4146
rect 12440 4082 12492 4088
rect 13820 4140 13872 4146
rect 13820 4082 13872 4088
rect 10784 4072 10836 4078
rect 10784 4014 10836 4020
rect 10876 4072 10928 4078
rect 10876 4014 10928 4020
rect 10796 3738 10824 4014
rect 12452 3942 12480 4082
rect 12992 4072 13044 4078
rect 12992 4014 13044 4020
rect 12440 3936 12492 3942
rect 12440 3878 12492 3884
rect 12214 3836 12522 3845
rect 12214 3834 12220 3836
rect 12276 3834 12300 3836
rect 12356 3834 12380 3836
rect 12436 3834 12460 3836
rect 12516 3834 12522 3836
rect 12276 3782 12278 3834
rect 12458 3782 12460 3834
rect 12214 3780 12220 3782
rect 12276 3780 12300 3782
rect 12356 3780 12380 3782
rect 12436 3780 12460 3782
rect 12516 3780 12522 3782
rect 12214 3771 12522 3780
rect 10784 3732 10836 3738
rect 10784 3674 10836 3680
rect 11520 3596 11572 3602
rect 11520 3538 11572 3544
rect 10692 3528 10744 3534
rect 10692 3470 10744 3476
rect 10600 3392 10652 3398
rect 10600 3334 10652 3340
rect 9772 3052 9824 3058
rect 9772 2994 9824 3000
rect 10508 3052 10560 3058
rect 10508 2994 10560 3000
rect 10232 2984 10284 2990
rect 10232 2926 10284 2932
rect 10244 2310 10272 2926
rect 10520 2650 10548 2994
rect 10508 2644 10560 2650
rect 10508 2586 10560 2592
rect 10232 2304 10284 2310
rect 10232 2246 10284 2252
rect 10244 1426 10272 2246
rect 10520 1766 10548 2586
rect 10612 2514 10640 3334
rect 10704 3097 10732 3470
rect 11532 3126 11560 3538
rect 13004 3534 13032 4014
rect 12992 3528 13044 3534
rect 12992 3470 13044 3476
rect 11520 3120 11572 3126
rect 10690 3088 10746 3097
rect 11520 3062 11572 3068
rect 11610 3088 11666 3097
rect 10690 3023 10746 3032
rect 10600 2508 10652 2514
rect 10600 2450 10652 2456
rect 10704 1970 10732 3023
rect 11152 2984 11204 2990
rect 11152 2926 11204 2932
rect 11060 2916 11112 2922
rect 11060 2858 11112 2864
rect 11072 2446 11100 2858
rect 11164 2582 11192 2926
rect 11532 2774 11560 3062
rect 13832 3058 13860 4082
rect 11610 3023 11612 3032
rect 11664 3023 11666 3032
rect 11796 3052 11848 3058
rect 11612 2994 11664 3000
rect 11796 2994 11848 3000
rect 13820 3052 13872 3058
rect 13820 2994 13872 3000
rect 11532 2746 11652 2774
rect 11152 2576 11204 2582
rect 11152 2518 11204 2524
rect 11060 2440 11112 2446
rect 11060 2382 11112 2388
rect 11164 2378 11192 2518
rect 11624 2514 11652 2746
rect 11808 2650 11836 2994
rect 12624 2916 12676 2922
rect 12624 2858 12676 2864
rect 13360 2916 13412 2922
rect 13360 2858 13412 2864
rect 11888 2848 11940 2854
rect 11888 2790 11940 2796
rect 11796 2644 11848 2650
rect 11796 2586 11848 2592
rect 11612 2508 11664 2514
rect 11612 2450 11664 2456
rect 11152 2372 11204 2378
rect 11152 2314 11204 2320
rect 11060 2304 11112 2310
rect 11060 2246 11112 2252
rect 11072 1970 11100 2246
rect 11624 2038 11652 2450
rect 11612 2032 11664 2038
rect 11612 1974 11664 1980
rect 10692 1964 10744 1970
rect 10692 1906 10744 1912
rect 11060 1964 11112 1970
rect 11060 1906 11112 1912
rect 10508 1760 10560 1766
rect 10508 1702 10560 1708
rect 10232 1420 10284 1426
rect 10232 1362 10284 1368
rect 10520 1358 10548 1702
rect 8576 1352 8628 1358
rect 8576 1294 8628 1300
rect 9220 1352 9272 1358
rect 9220 1294 9272 1300
rect 9680 1352 9732 1358
rect 9680 1294 9732 1300
rect 10508 1352 10560 1358
rect 10508 1294 10560 1300
rect 11072 1290 11100 1906
rect 11152 1896 11204 1902
rect 11152 1838 11204 1844
rect 11164 1426 11192 1838
rect 11152 1420 11204 1426
rect 11152 1362 11204 1368
rect 11900 1358 11928 2790
rect 12214 2748 12522 2757
rect 12214 2746 12220 2748
rect 12276 2746 12300 2748
rect 12356 2746 12380 2748
rect 12436 2746 12460 2748
rect 12516 2746 12522 2748
rect 12276 2694 12278 2746
rect 12458 2694 12460 2746
rect 12214 2692 12220 2694
rect 12276 2692 12300 2694
rect 12356 2692 12380 2694
rect 12436 2692 12460 2694
rect 12516 2692 12522 2694
rect 12214 2683 12522 2692
rect 11980 2372 12032 2378
rect 11980 2314 12032 2320
rect 11992 1562 12020 2314
rect 12636 2038 12664 2858
rect 13372 2446 13400 2858
rect 13924 2446 13952 4558
rect 14096 4140 14148 4146
rect 14200 4128 14228 5646
rect 14464 5296 14516 5302
rect 14464 5238 14516 5244
rect 14476 4758 14504 5238
rect 14752 5166 14780 5646
rect 14844 5370 14872 6326
rect 15028 6322 15056 7210
rect 15212 6866 15240 7346
rect 15200 6860 15252 6866
rect 15200 6802 15252 6808
rect 15304 6798 15332 7482
rect 15476 7336 15528 7342
rect 15476 7278 15528 7284
rect 15488 6798 15516 7278
rect 15292 6792 15344 6798
rect 15292 6734 15344 6740
rect 15476 6792 15528 6798
rect 15476 6734 15528 6740
rect 15016 6316 15068 6322
rect 15016 6258 15068 6264
rect 15304 6254 15332 6734
rect 15292 6248 15344 6254
rect 15292 6190 15344 6196
rect 15292 6112 15344 6118
rect 15292 6054 15344 6060
rect 14832 5364 14884 5370
rect 14832 5306 14884 5312
rect 14740 5160 14792 5166
rect 14740 5102 14792 5108
rect 14464 4752 14516 4758
rect 14464 4694 14516 4700
rect 14752 4690 14780 5102
rect 14740 4684 14792 4690
rect 14740 4626 14792 4632
rect 15304 4554 15332 6054
rect 15292 4548 15344 4554
rect 15292 4490 15344 4496
rect 15476 4548 15528 4554
rect 15476 4490 15528 4496
rect 15488 4282 15516 4490
rect 15476 4276 15528 4282
rect 15476 4218 15528 4224
rect 14148 4100 14228 4128
rect 14096 4082 14148 4088
rect 14200 3942 14228 4100
rect 14372 4072 14424 4078
rect 14372 4014 14424 4020
rect 14556 4072 14608 4078
rect 14556 4014 14608 4020
rect 14188 3936 14240 3942
rect 14188 3878 14240 3884
rect 14200 3534 14228 3878
rect 14384 3534 14412 4014
rect 14568 3534 14596 4014
rect 14188 3528 14240 3534
rect 14188 3470 14240 3476
rect 14372 3528 14424 3534
rect 14372 3470 14424 3476
rect 14556 3528 14608 3534
rect 14556 3470 14608 3476
rect 14200 2650 14228 3470
rect 14280 3392 14332 3398
rect 14280 3334 14332 3340
rect 14188 2644 14240 2650
rect 14188 2586 14240 2592
rect 13360 2440 13412 2446
rect 13360 2382 13412 2388
rect 13912 2440 13964 2446
rect 13912 2382 13964 2388
rect 14292 2038 14320 3334
rect 14568 2990 14596 3470
rect 14556 2984 14608 2990
rect 14556 2926 14608 2932
rect 14568 2514 14596 2926
rect 14556 2508 14608 2514
rect 14556 2450 14608 2456
rect 14568 2106 14596 2450
rect 14924 2304 14976 2310
rect 14924 2246 14976 2252
rect 14556 2100 14608 2106
rect 14556 2042 14608 2048
rect 12624 2032 12676 2038
rect 12624 1974 12676 1980
rect 14280 2032 14332 2038
rect 14280 1974 14332 1980
rect 12214 1660 12522 1669
rect 12214 1658 12220 1660
rect 12276 1658 12300 1660
rect 12356 1658 12380 1660
rect 12436 1658 12460 1660
rect 12516 1658 12522 1660
rect 12276 1606 12278 1658
rect 12458 1606 12460 1658
rect 12214 1604 12220 1606
rect 12276 1604 12300 1606
rect 12356 1604 12380 1606
rect 12436 1604 12460 1606
rect 12516 1604 12522 1606
rect 12214 1595 12522 1604
rect 11980 1556 12032 1562
rect 11980 1498 12032 1504
rect 14568 1426 14596 2042
rect 14936 1902 14964 2246
rect 14924 1896 14976 1902
rect 14924 1838 14976 1844
rect 14832 1760 14884 1766
rect 14832 1702 14884 1708
rect 14844 1426 14872 1702
rect 14556 1420 14608 1426
rect 14556 1362 14608 1368
rect 14832 1420 14884 1426
rect 14832 1362 14884 1368
rect 11888 1352 11940 1358
rect 11888 1294 11940 1300
rect 7472 1284 7524 1290
rect 7472 1226 7524 1232
rect 7564 1284 7616 1290
rect 7564 1226 7616 1232
rect 11060 1284 11112 1290
rect 11060 1226 11112 1232
rect 6460 1216 6512 1222
rect 6460 1158 6512 1164
rect 6472 1018 6500 1158
rect 6460 1012 6512 1018
rect 6460 954 6512 960
rect 7576 950 7604 1226
rect 8214 1116 8522 1125
rect 8214 1114 8220 1116
rect 8276 1114 8300 1116
rect 8356 1114 8380 1116
rect 8436 1114 8460 1116
rect 8516 1114 8522 1116
rect 8276 1062 8278 1114
rect 8458 1062 8460 1114
rect 8214 1060 8220 1062
rect 8276 1060 8300 1062
rect 8356 1060 8380 1062
rect 8436 1060 8460 1062
rect 8516 1060 8522 1062
rect 8214 1051 8522 1060
rect 5448 944 5500 950
rect 4908 870 5028 898
rect 5448 886 5500 892
rect 7564 944 7616 950
rect 7564 886 7616 892
rect 4908 762 4936 870
rect 5000 800 5028 870
rect 14936 800 14964 1838
rect 15580 1329 15608 8910
rect 15660 7744 15712 7750
rect 15660 7686 15712 7692
rect 15672 5778 15700 7686
rect 15660 5772 15712 5778
rect 15660 5714 15712 5720
rect 15764 5370 15792 11698
rect 15934 11248 15990 11257
rect 15934 11183 15990 11192
rect 15844 11144 15896 11150
rect 15844 11086 15896 11092
rect 15856 10742 15884 11086
rect 15844 10736 15896 10742
rect 15844 10678 15896 10684
rect 15842 9616 15898 9625
rect 15842 9551 15898 9560
rect 15856 6390 15884 9551
rect 15948 7954 15976 11183
rect 16040 11121 16068 12038
rect 16132 11762 16160 12038
rect 16214 11996 16522 12005
rect 16214 11994 16220 11996
rect 16276 11994 16300 11996
rect 16356 11994 16380 11996
rect 16436 11994 16460 11996
rect 16516 11994 16522 11996
rect 16276 11942 16278 11994
rect 16458 11942 16460 11994
rect 16214 11940 16220 11942
rect 16276 11940 16300 11942
rect 16356 11940 16380 11942
rect 16436 11940 16460 11942
rect 16516 11940 16522 11942
rect 16214 11931 16522 11940
rect 16120 11756 16172 11762
rect 16120 11698 16172 11704
rect 16776 11626 16804 12038
rect 16764 11620 16816 11626
rect 16764 11562 16816 11568
rect 16856 11620 16908 11626
rect 16856 11562 16908 11568
rect 16672 11144 16724 11150
rect 16026 11112 16082 11121
rect 16672 11086 16724 11092
rect 16026 11047 16082 11056
rect 16040 9382 16068 11047
rect 16214 10908 16522 10917
rect 16214 10906 16220 10908
rect 16276 10906 16300 10908
rect 16356 10906 16380 10908
rect 16436 10906 16460 10908
rect 16516 10906 16522 10908
rect 16276 10854 16278 10906
rect 16458 10854 16460 10906
rect 16214 10852 16220 10854
rect 16276 10852 16300 10854
rect 16356 10852 16380 10854
rect 16436 10852 16460 10854
rect 16516 10852 16522 10854
rect 16214 10843 16522 10852
rect 16684 10810 16712 11086
rect 16868 11082 16896 11562
rect 16856 11076 16908 11082
rect 16856 11018 16908 11024
rect 16672 10804 16724 10810
rect 16672 10746 16724 10752
rect 16764 10600 16816 10606
rect 16764 10542 16816 10548
rect 16776 10062 16804 10542
rect 16764 10056 16816 10062
rect 16764 9998 16816 10004
rect 16672 9988 16724 9994
rect 16672 9930 16724 9936
rect 16214 9820 16522 9829
rect 16214 9818 16220 9820
rect 16276 9818 16300 9820
rect 16356 9818 16380 9820
rect 16436 9818 16460 9820
rect 16516 9818 16522 9820
rect 16276 9766 16278 9818
rect 16458 9766 16460 9818
rect 16214 9764 16220 9766
rect 16276 9764 16300 9766
rect 16356 9764 16380 9766
rect 16436 9764 16460 9766
rect 16516 9764 16522 9766
rect 16214 9755 16522 9764
rect 16684 9654 16712 9930
rect 16776 9654 16804 9998
rect 16672 9648 16724 9654
rect 16672 9590 16724 9596
rect 16764 9648 16816 9654
rect 16764 9590 16816 9596
rect 16672 9512 16724 9518
rect 16672 9454 16724 9460
rect 16028 9376 16080 9382
rect 16028 9318 16080 9324
rect 16120 9104 16172 9110
rect 16120 9046 16172 9052
rect 16028 8492 16080 8498
rect 16028 8434 16080 8440
rect 15936 7948 15988 7954
rect 15936 7890 15988 7896
rect 15936 6656 15988 6662
rect 15936 6598 15988 6604
rect 15844 6384 15896 6390
rect 15844 6326 15896 6332
rect 15856 5778 15884 6326
rect 15948 6322 15976 6598
rect 15936 6316 15988 6322
rect 15936 6258 15988 6264
rect 15844 5772 15896 5778
rect 15844 5714 15896 5720
rect 16040 5574 16068 8434
rect 16132 6798 16160 9046
rect 16684 8974 16712 9454
rect 16672 8968 16724 8974
rect 16672 8910 16724 8916
rect 16960 8906 16988 12174
rect 17236 12102 17264 13330
rect 17776 13184 17828 13190
rect 17776 13126 17828 13132
rect 17788 12850 17816 13126
rect 17776 12844 17828 12850
rect 17776 12786 17828 12792
rect 17788 12374 17816 12786
rect 18236 12640 18288 12646
rect 18236 12582 18288 12588
rect 17776 12368 17828 12374
rect 17776 12310 17828 12316
rect 18248 12306 18276 12582
rect 18800 12345 18828 14200
rect 18786 12336 18842 12345
rect 18236 12300 18288 12306
rect 18786 12271 18842 12280
rect 18236 12242 18288 12248
rect 17224 12096 17276 12102
rect 17224 12038 17276 12044
rect 17132 11552 17184 11558
rect 17132 11494 17184 11500
rect 17144 11218 17172 11494
rect 17132 11212 17184 11218
rect 17132 11154 17184 11160
rect 17236 9654 17264 12038
rect 17684 11756 17736 11762
rect 17684 11698 17736 11704
rect 17500 11280 17552 11286
rect 17500 11222 17552 11228
rect 17512 10742 17540 11222
rect 17500 10736 17552 10742
rect 17500 10678 17552 10684
rect 17696 10606 17724 11698
rect 18144 11620 18196 11626
rect 18144 11562 18196 11568
rect 18052 11144 18104 11150
rect 18052 11086 18104 11092
rect 17684 10600 17736 10606
rect 17684 10542 17736 10548
rect 17408 10532 17460 10538
rect 17408 10474 17460 10480
rect 17420 9994 17448 10474
rect 18064 10266 18092 11086
rect 18156 10742 18184 11562
rect 18144 10736 18196 10742
rect 18144 10678 18196 10684
rect 18052 10260 18104 10266
rect 18052 10202 18104 10208
rect 18156 10062 18184 10678
rect 17684 10056 17736 10062
rect 17684 9998 17736 10004
rect 18144 10056 18196 10062
rect 18144 9998 18196 10004
rect 17408 9988 17460 9994
rect 17408 9930 17460 9936
rect 17224 9648 17276 9654
rect 17224 9590 17276 9596
rect 16948 8900 17000 8906
rect 16948 8842 17000 8848
rect 16214 8732 16522 8741
rect 16214 8730 16220 8732
rect 16276 8730 16300 8732
rect 16356 8730 16380 8732
rect 16436 8730 16460 8732
rect 16516 8730 16522 8732
rect 16276 8678 16278 8730
rect 16458 8678 16460 8730
rect 16214 8676 16220 8678
rect 16276 8676 16300 8678
rect 16356 8676 16380 8678
rect 16436 8676 16460 8678
rect 16516 8676 16522 8678
rect 16214 8667 16522 8676
rect 17236 8514 17264 9590
rect 17696 8974 17724 9998
rect 17776 9580 17828 9586
rect 17776 9522 17828 9528
rect 17684 8968 17736 8974
rect 17684 8910 17736 8916
rect 17052 8486 17264 8514
rect 16672 8356 16724 8362
rect 16672 8298 16724 8304
rect 16580 7812 16632 7818
rect 16580 7754 16632 7760
rect 16214 7644 16522 7653
rect 16214 7642 16220 7644
rect 16276 7642 16300 7644
rect 16356 7642 16380 7644
rect 16436 7642 16460 7644
rect 16516 7642 16522 7644
rect 16276 7590 16278 7642
rect 16458 7590 16460 7642
rect 16214 7588 16220 7590
rect 16276 7588 16300 7590
rect 16356 7588 16380 7590
rect 16436 7588 16460 7590
rect 16516 7588 16522 7590
rect 16214 7579 16522 7588
rect 16592 7546 16620 7754
rect 16580 7540 16632 7546
rect 16580 7482 16632 7488
rect 16684 7410 16712 8298
rect 16212 7404 16264 7410
rect 16212 7346 16264 7352
rect 16672 7404 16724 7410
rect 16672 7346 16724 7352
rect 16120 6792 16172 6798
rect 16120 6734 16172 6740
rect 16224 6644 16252 7346
rect 16132 6616 16252 6644
rect 16028 5568 16080 5574
rect 16028 5510 16080 5516
rect 15752 5364 15804 5370
rect 15752 5306 15804 5312
rect 16132 4826 16160 6616
rect 16214 6556 16522 6565
rect 16214 6554 16220 6556
rect 16276 6554 16300 6556
rect 16356 6554 16380 6556
rect 16436 6554 16460 6556
rect 16516 6554 16522 6556
rect 16276 6502 16278 6554
rect 16458 6502 16460 6554
rect 16214 6500 16220 6502
rect 16276 6500 16300 6502
rect 16356 6500 16380 6502
rect 16436 6500 16460 6502
rect 16516 6500 16522 6502
rect 16214 6491 16522 6500
rect 17052 6458 17080 8486
rect 17224 8356 17276 8362
rect 17224 8298 17276 8304
rect 17236 7478 17264 8298
rect 17408 7744 17460 7750
rect 17408 7686 17460 7692
rect 17224 7472 17276 7478
rect 17224 7414 17276 7420
rect 17316 6860 17368 6866
rect 17316 6802 17368 6808
rect 16580 6452 16632 6458
rect 16580 6394 16632 6400
rect 17040 6452 17092 6458
rect 17040 6394 17092 6400
rect 16592 5914 16620 6394
rect 17132 6384 17184 6390
rect 17132 6326 17184 6332
rect 16580 5908 16632 5914
rect 16580 5850 16632 5856
rect 16214 5468 16522 5477
rect 16214 5466 16220 5468
rect 16276 5466 16300 5468
rect 16356 5466 16380 5468
rect 16436 5466 16460 5468
rect 16516 5466 16522 5468
rect 16276 5414 16278 5466
rect 16458 5414 16460 5466
rect 16214 5412 16220 5414
rect 16276 5412 16300 5414
rect 16356 5412 16380 5414
rect 16436 5412 16460 5414
rect 16516 5412 16522 5414
rect 16214 5403 16522 5412
rect 16592 5370 16620 5850
rect 16580 5364 16632 5370
rect 16580 5306 16632 5312
rect 16120 4820 16172 4826
rect 16120 4762 16172 4768
rect 16856 4684 16908 4690
rect 16856 4626 16908 4632
rect 16028 4480 16080 4486
rect 16028 4422 16080 4428
rect 15660 3460 15712 3466
rect 15660 3402 15712 3408
rect 15672 1970 15700 3402
rect 16040 2774 16068 4422
rect 16214 4380 16522 4389
rect 16214 4378 16220 4380
rect 16276 4378 16300 4380
rect 16356 4378 16380 4380
rect 16436 4378 16460 4380
rect 16516 4378 16522 4380
rect 16276 4326 16278 4378
rect 16458 4326 16460 4378
rect 16214 4324 16220 4326
rect 16276 4324 16300 4326
rect 16356 4324 16380 4326
rect 16436 4324 16460 4326
rect 16516 4324 16522 4326
rect 16214 4315 16522 4324
rect 16672 4208 16724 4214
rect 16672 4150 16724 4156
rect 16580 4072 16632 4078
rect 16580 4014 16632 4020
rect 16120 4004 16172 4010
rect 16120 3946 16172 3952
rect 16132 3194 16160 3946
rect 16214 3292 16522 3301
rect 16214 3290 16220 3292
rect 16276 3290 16300 3292
rect 16356 3290 16380 3292
rect 16436 3290 16460 3292
rect 16516 3290 16522 3292
rect 16276 3238 16278 3290
rect 16458 3238 16460 3290
rect 16214 3236 16220 3238
rect 16276 3236 16300 3238
rect 16356 3236 16380 3238
rect 16436 3236 16460 3238
rect 16516 3236 16522 3238
rect 16214 3227 16522 3236
rect 16120 3188 16172 3194
rect 16120 3130 16172 3136
rect 16040 2746 16160 2774
rect 16132 1970 16160 2746
rect 16214 2204 16522 2213
rect 16214 2202 16220 2204
rect 16276 2202 16300 2204
rect 16356 2202 16380 2204
rect 16436 2202 16460 2204
rect 16516 2202 16522 2204
rect 16276 2150 16278 2202
rect 16458 2150 16460 2202
rect 16214 2148 16220 2150
rect 16276 2148 16300 2150
rect 16356 2148 16380 2150
rect 16436 2148 16460 2150
rect 16516 2148 16522 2150
rect 16214 2139 16522 2148
rect 15660 1964 15712 1970
rect 15660 1906 15712 1912
rect 16120 1964 16172 1970
rect 16120 1906 16172 1912
rect 15936 1828 15988 1834
rect 15936 1770 15988 1776
rect 15948 1358 15976 1770
rect 16132 1426 16160 1906
rect 16592 1902 16620 4014
rect 16580 1896 16632 1902
rect 16580 1838 16632 1844
rect 16120 1420 16172 1426
rect 16120 1362 16172 1368
rect 15936 1352 15988 1358
rect 15566 1320 15622 1329
rect 15936 1294 15988 1300
rect 15566 1255 15622 1264
rect 16592 1222 16620 1838
rect 16684 1222 16712 4150
rect 16764 3936 16816 3942
rect 16764 3878 16816 3884
rect 16776 1970 16804 3878
rect 16868 3602 16896 4626
rect 17144 4622 17172 6326
rect 17328 5370 17356 6802
rect 17316 5364 17368 5370
rect 17316 5306 17368 5312
rect 17224 5296 17276 5302
rect 17224 5238 17276 5244
rect 17236 4622 17264 5238
rect 17132 4616 17184 4622
rect 17132 4558 17184 4564
rect 17224 4616 17276 4622
rect 17224 4558 17276 4564
rect 16948 4548 17000 4554
rect 16948 4490 17000 4496
rect 17040 4548 17092 4554
rect 17040 4490 17092 4496
rect 16856 3596 16908 3602
rect 16856 3538 16908 3544
rect 16960 3466 16988 4490
rect 17052 4282 17080 4490
rect 17040 4276 17092 4282
rect 17040 4218 17092 4224
rect 16948 3460 17000 3466
rect 16948 3402 17000 3408
rect 17052 3097 17080 4218
rect 17144 4214 17172 4558
rect 17236 4282 17264 4558
rect 17224 4276 17276 4282
rect 17224 4218 17276 4224
rect 17132 4208 17184 4214
rect 17132 4150 17184 4156
rect 17144 4010 17172 4150
rect 17132 4004 17184 4010
rect 17132 3946 17184 3952
rect 17224 3392 17276 3398
rect 17224 3334 17276 3340
rect 17038 3088 17094 3097
rect 17236 3058 17264 3334
rect 17420 3126 17448 7686
rect 17500 6928 17552 6934
rect 17500 6870 17552 6876
rect 17512 6186 17540 6870
rect 17788 6225 17816 9522
rect 18052 9444 18104 9450
rect 18052 9386 18104 9392
rect 18064 9110 18092 9386
rect 18052 9104 18104 9110
rect 18052 9046 18104 9052
rect 18064 8566 18092 9046
rect 18052 8560 18104 8566
rect 18052 8502 18104 8508
rect 17960 8424 18012 8430
rect 17960 8366 18012 8372
rect 17868 8288 17920 8294
rect 17868 8230 17920 8236
rect 17880 7886 17908 8230
rect 17868 7880 17920 7886
rect 17868 7822 17920 7828
rect 17880 7478 17908 7822
rect 17972 7546 18000 8366
rect 18420 8356 18472 8362
rect 18420 8298 18472 8304
rect 18052 8016 18104 8022
rect 18052 7958 18104 7964
rect 17960 7540 18012 7546
rect 17960 7482 18012 7488
rect 17868 7472 17920 7478
rect 17868 7414 17920 7420
rect 18064 6730 18092 7958
rect 18052 6724 18104 6730
rect 18052 6666 18104 6672
rect 18144 6724 18196 6730
rect 18144 6666 18196 6672
rect 18064 6322 18092 6666
rect 18052 6316 18104 6322
rect 18052 6258 18104 6264
rect 17774 6216 17830 6225
rect 17500 6180 17552 6186
rect 17774 6151 17830 6160
rect 17500 6122 17552 6128
rect 17512 5846 17540 6122
rect 17788 5846 17816 6151
rect 17500 5840 17552 5846
rect 17500 5782 17552 5788
rect 17776 5840 17828 5846
rect 17776 5782 17828 5788
rect 17512 3942 17540 5782
rect 18064 5710 18092 6258
rect 18156 5914 18184 6666
rect 18144 5908 18196 5914
rect 18144 5850 18196 5856
rect 18052 5704 18104 5710
rect 18052 5646 18104 5652
rect 17592 5636 17644 5642
rect 17592 5578 17644 5584
rect 17604 5302 17632 5578
rect 17592 5296 17644 5302
rect 17592 5238 17644 5244
rect 17684 5160 17736 5166
rect 17684 5102 17736 5108
rect 17696 4146 17724 5102
rect 18052 4616 18104 4622
rect 18052 4558 18104 4564
rect 17960 4208 18012 4214
rect 17960 4150 18012 4156
rect 17684 4140 17736 4146
rect 17684 4082 17736 4088
rect 17500 3936 17552 3942
rect 17500 3878 17552 3884
rect 17776 3392 17828 3398
rect 17776 3334 17828 3340
rect 17408 3120 17460 3126
rect 17408 3062 17460 3068
rect 17038 3023 17094 3032
rect 17224 3052 17276 3058
rect 17224 2994 17276 3000
rect 17788 2990 17816 3334
rect 17868 3188 17920 3194
rect 17868 3130 17920 3136
rect 17500 2984 17552 2990
rect 17500 2926 17552 2932
rect 17776 2984 17828 2990
rect 17776 2926 17828 2932
rect 17040 2848 17092 2854
rect 17040 2790 17092 2796
rect 17052 2514 17080 2790
rect 17040 2508 17092 2514
rect 17040 2450 17092 2456
rect 16948 2032 17000 2038
rect 16948 1974 17000 1980
rect 16764 1964 16816 1970
rect 16764 1906 16816 1912
rect 16960 1358 16988 1974
rect 16948 1352 17000 1358
rect 16948 1294 17000 1300
rect 17512 1222 17540 2926
rect 17592 2576 17644 2582
rect 17592 2518 17644 2524
rect 17604 1358 17632 2518
rect 17788 2310 17816 2926
rect 17880 2394 17908 3130
rect 17972 2514 18000 4150
rect 18064 3602 18092 4558
rect 18236 4140 18288 4146
rect 18236 4082 18288 4088
rect 18248 3738 18276 4082
rect 18328 4072 18380 4078
rect 18328 4014 18380 4020
rect 18236 3732 18288 3738
rect 18236 3674 18288 3680
rect 18052 3596 18104 3602
rect 18052 3538 18104 3544
rect 18064 3194 18092 3538
rect 18340 3534 18368 4014
rect 18432 3777 18460 8298
rect 18418 3768 18474 3777
rect 18418 3703 18474 3712
rect 18328 3528 18380 3534
rect 18328 3470 18380 3476
rect 18052 3188 18104 3194
rect 18052 3130 18104 3136
rect 18236 2984 18288 2990
rect 18236 2926 18288 2932
rect 17960 2508 18012 2514
rect 17960 2450 18012 2456
rect 17880 2378 18000 2394
rect 17880 2372 18012 2378
rect 17880 2366 17960 2372
rect 17960 2314 18012 2320
rect 17776 2304 17828 2310
rect 17776 2246 17828 2252
rect 18248 2106 18276 2926
rect 18340 2378 18368 3470
rect 18328 2372 18380 2378
rect 18328 2314 18380 2320
rect 18236 2100 18288 2106
rect 18236 2042 18288 2048
rect 18248 1358 18276 2042
rect 17592 1352 17644 1358
rect 17592 1294 17644 1300
rect 18236 1352 18288 1358
rect 18236 1294 18288 1300
rect 18340 1222 18368 2314
rect 16580 1216 16632 1222
rect 16580 1158 16632 1164
rect 16672 1216 16724 1222
rect 16672 1158 16724 1164
rect 17500 1216 17552 1222
rect 17500 1158 17552 1164
rect 18328 1216 18380 1222
rect 18328 1158 18380 1164
rect 16214 1116 16522 1125
rect 16214 1114 16220 1116
rect 16276 1114 16300 1116
rect 16356 1114 16380 1116
rect 16436 1114 16460 1116
rect 16516 1114 16522 1116
rect 16276 1062 16278 1114
rect 16458 1062 16460 1114
rect 16214 1060 16220 1062
rect 16276 1060 16300 1062
rect 16356 1060 16380 1062
rect 16436 1060 16460 1062
rect 16516 1060 16522 1062
rect 16214 1051 16522 1060
rect 18340 950 18368 1158
rect 18328 944 18380 950
rect 18328 886 18380 892
rect 4724 734 4936 762
rect 4986 0 5042 800
rect 14922 0 14978 800
<< via2 >>
rect 2042 10512 2098 10568
rect 3422 13504 3478 13560
rect 2778 12688 2834 12744
rect 3422 11872 3478 11928
rect 4220 13626 4276 13628
rect 4300 13626 4356 13628
rect 4380 13626 4436 13628
rect 4460 13626 4516 13628
rect 4220 13574 4266 13626
rect 4266 13574 4276 13626
rect 4300 13574 4330 13626
rect 4330 13574 4342 13626
rect 4342 13574 4356 13626
rect 4380 13574 4394 13626
rect 4394 13574 4406 13626
rect 4406 13574 4436 13626
rect 4460 13574 4470 13626
rect 4470 13574 4516 13626
rect 4220 13572 4276 13574
rect 4300 13572 4356 13574
rect 4380 13572 4436 13574
rect 4460 13572 4516 13574
rect 4220 12538 4276 12540
rect 4300 12538 4356 12540
rect 4380 12538 4436 12540
rect 4460 12538 4516 12540
rect 4220 12486 4266 12538
rect 4266 12486 4276 12538
rect 4300 12486 4330 12538
rect 4330 12486 4342 12538
rect 4342 12486 4356 12538
rect 4380 12486 4394 12538
rect 4394 12486 4406 12538
rect 4406 12486 4436 12538
rect 4460 12486 4470 12538
rect 4470 12486 4516 12538
rect 4220 12484 4276 12486
rect 4300 12484 4356 12486
rect 4380 12484 4436 12486
rect 4460 12484 4516 12486
rect 4220 11450 4276 11452
rect 4300 11450 4356 11452
rect 4380 11450 4436 11452
rect 4460 11450 4516 11452
rect 4220 11398 4266 11450
rect 4266 11398 4276 11450
rect 4300 11398 4330 11450
rect 4330 11398 4342 11450
rect 4342 11398 4356 11450
rect 4380 11398 4394 11450
rect 4394 11398 4406 11450
rect 4406 11398 4436 11450
rect 4460 11398 4470 11450
rect 4470 11398 4516 11450
rect 4220 11396 4276 11398
rect 4300 11396 4356 11398
rect 4380 11396 4436 11398
rect 4460 11396 4516 11398
rect 4066 11056 4122 11112
rect 3790 10240 3846 10296
rect 1766 9424 1822 9480
rect 4220 10362 4276 10364
rect 4300 10362 4356 10364
rect 4380 10362 4436 10364
rect 4460 10362 4516 10364
rect 4220 10310 4266 10362
rect 4266 10310 4276 10362
rect 4300 10310 4330 10362
rect 4330 10310 4342 10362
rect 4342 10310 4356 10362
rect 4380 10310 4394 10362
rect 4394 10310 4406 10362
rect 4406 10310 4436 10362
rect 4460 10310 4470 10362
rect 4470 10310 4516 10362
rect 4220 10308 4276 10310
rect 4300 10308 4356 10310
rect 4380 10308 4436 10310
rect 4460 10308 4516 10310
rect 4220 9274 4276 9276
rect 4300 9274 4356 9276
rect 4380 9274 4436 9276
rect 4460 9274 4516 9276
rect 4220 9222 4266 9274
rect 4266 9222 4276 9274
rect 4300 9222 4330 9274
rect 4330 9222 4342 9274
rect 4342 9222 4356 9274
rect 4380 9222 4394 9274
rect 4394 9222 4406 9274
rect 4406 9222 4436 9274
rect 4460 9222 4470 9274
rect 4470 9222 4516 9274
rect 4220 9220 4276 9222
rect 4300 9220 4356 9222
rect 4380 9220 4436 9222
rect 4460 9220 4516 9222
rect 3974 8608 4030 8664
rect 4220 8186 4276 8188
rect 4300 8186 4356 8188
rect 4380 8186 4436 8188
rect 4460 8186 4516 8188
rect 4220 8134 4266 8186
rect 4266 8134 4276 8186
rect 4300 8134 4330 8186
rect 4330 8134 4342 8186
rect 4342 8134 4356 8186
rect 4380 8134 4394 8186
rect 4394 8134 4406 8186
rect 4406 8134 4436 8186
rect 4460 8134 4470 8186
rect 4470 8134 4516 8186
rect 4220 8132 4276 8134
rect 4300 8132 4356 8134
rect 4380 8132 4436 8134
rect 4460 8132 4516 8134
rect 3146 7792 3202 7848
rect 1582 6160 1638 6216
rect 1582 5344 1638 5400
rect 2962 6976 3018 7032
rect 1766 3712 1822 3768
rect 2594 4564 2596 4584
rect 2596 4564 2648 4584
rect 2648 4564 2650 4584
rect 2594 4528 2650 4564
rect 2778 2896 2834 2952
rect 1490 1264 1546 1320
rect 6918 11736 6974 11792
rect 6826 11464 6882 11520
rect 8220 13082 8276 13084
rect 8300 13082 8356 13084
rect 8380 13082 8436 13084
rect 8460 13082 8516 13084
rect 8220 13030 8266 13082
rect 8266 13030 8276 13082
rect 8300 13030 8330 13082
rect 8330 13030 8342 13082
rect 8342 13030 8356 13082
rect 8380 13030 8394 13082
rect 8394 13030 8406 13082
rect 8406 13030 8436 13082
rect 8460 13030 8470 13082
rect 8470 13030 8516 13082
rect 8220 13028 8276 13030
rect 8300 13028 8356 13030
rect 8380 13028 8436 13030
rect 8460 13028 8516 13030
rect 8482 12164 8538 12200
rect 8482 12144 8484 12164
rect 8484 12144 8536 12164
rect 8536 12144 8538 12164
rect 8850 12144 8906 12200
rect 8220 11994 8276 11996
rect 8300 11994 8356 11996
rect 8380 11994 8436 11996
rect 8460 11994 8516 11996
rect 8220 11942 8266 11994
rect 8266 11942 8276 11994
rect 8300 11942 8330 11994
rect 8330 11942 8342 11994
rect 8342 11942 8356 11994
rect 8380 11942 8394 11994
rect 8394 11942 8406 11994
rect 8406 11942 8436 11994
rect 8460 11942 8470 11994
rect 8470 11942 8516 11994
rect 8220 11940 8276 11942
rect 8300 11940 8356 11942
rect 8380 11940 8436 11942
rect 8460 11940 8516 11942
rect 7010 10648 7066 10704
rect 5998 8916 6000 8936
rect 6000 8916 6052 8936
rect 6052 8916 6054 8936
rect 5998 8880 6054 8916
rect 6642 9016 6698 9072
rect 7838 8880 7894 8936
rect 8298 11192 8354 11248
rect 8220 10906 8276 10908
rect 8300 10906 8356 10908
rect 8380 10906 8436 10908
rect 8460 10906 8516 10908
rect 8220 10854 8266 10906
rect 8266 10854 8276 10906
rect 8300 10854 8330 10906
rect 8330 10854 8342 10906
rect 8342 10854 8356 10906
rect 8380 10854 8394 10906
rect 8394 10854 8406 10906
rect 8406 10854 8436 10906
rect 8460 10854 8470 10906
rect 8470 10854 8516 10906
rect 8220 10852 8276 10854
rect 8300 10852 8356 10854
rect 8380 10852 8436 10854
rect 8460 10852 8516 10854
rect 8666 11056 8722 11112
rect 8298 10668 8354 10704
rect 8298 10648 8300 10668
rect 8300 10648 8352 10668
rect 8352 10648 8354 10668
rect 8114 10376 8170 10432
rect 4220 7098 4276 7100
rect 4300 7098 4356 7100
rect 4380 7098 4436 7100
rect 4460 7098 4516 7100
rect 4220 7046 4266 7098
rect 4266 7046 4276 7098
rect 4300 7046 4330 7098
rect 4330 7046 4342 7098
rect 4342 7046 4356 7098
rect 4380 7046 4394 7098
rect 4394 7046 4406 7098
rect 4406 7046 4436 7098
rect 4460 7046 4470 7098
rect 4470 7046 4516 7098
rect 4220 7044 4276 7046
rect 4300 7044 4356 7046
rect 4380 7044 4436 7046
rect 4460 7044 4516 7046
rect 4220 6010 4276 6012
rect 4300 6010 4356 6012
rect 4380 6010 4436 6012
rect 4460 6010 4516 6012
rect 4220 5958 4266 6010
rect 4266 5958 4276 6010
rect 4300 5958 4330 6010
rect 4330 5958 4342 6010
rect 4342 5958 4356 6010
rect 4380 5958 4394 6010
rect 4394 5958 4406 6010
rect 4406 5958 4436 6010
rect 4460 5958 4470 6010
rect 4470 5958 4516 6010
rect 4220 5956 4276 5958
rect 4300 5956 4356 5958
rect 4380 5956 4436 5958
rect 4460 5956 4516 5958
rect 3698 5364 3754 5400
rect 3698 5344 3700 5364
rect 3700 5344 3752 5364
rect 3752 5344 3754 5364
rect 4220 4922 4276 4924
rect 4300 4922 4356 4924
rect 4380 4922 4436 4924
rect 4460 4922 4516 4924
rect 4220 4870 4266 4922
rect 4266 4870 4276 4922
rect 4300 4870 4330 4922
rect 4330 4870 4342 4922
rect 4342 4870 4356 4922
rect 4380 4870 4394 4922
rect 4394 4870 4406 4922
rect 4406 4870 4436 4922
rect 4460 4870 4470 4922
rect 4470 4870 4516 4922
rect 4220 4868 4276 4870
rect 4300 4868 4356 4870
rect 4380 4868 4436 4870
rect 4460 4868 4516 4870
rect 4220 3834 4276 3836
rect 4300 3834 4356 3836
rect 4380 3834 4436 3836
rect 4460 3834 4516 3836
rect 4220 3782 4266 3834
rect 4266 3782 4276 3834
rect 4300 3782 4330 3834
rect 4330 3782 4342 3834
rect 4342 3782 4356 3834
rect 4380 3782 4394 3834
rect 4394 3782 4406 3834
rect 4406 3782 4436 3834
rect 4460 3782 4470 3834
rect 4470 3782 4516 3834
rect 4220 3780 4276 3782
rect 4300 3780 4356 3782
rect 4380 3780 4436 3782
rect 4460 3780 4516 3782
rect 3054 2080 3110 2136
rect 4220 2746 4276 2748
rect 4300 2746 4356 2748
rect 4380 2746 4436 2748
rect 4460 2746 4516 2748
rect 4220 2694 4266 2746
rect 4266 2694 4276 2746
rect 4300 2694 4330 2746
rect 4330 2694 4342 2746
rect 4342 2694 4356 2746
rect 4380 2694 4394 2746
rect 4394 2694 4406 2746
rect 4406 2694 4436 2746
rect 4460 2694 4470 2746
rect 4470 2694 4516 2746
rect 4220 2692 4276 2694
rect 4300 2692 4356 2694
rect 4380 2692 4436 2694
rect 4460 2692 4516 2694
rect 4220 1658 4276 1660
rect 4300 1658 4356 1660
rect 4380 1658 4436 1660
rect 4460 1658 4516 1660
rect 4220 1606 4266 1658
rect 4266 1606 4276 1658
rect 4300 1606 4330 1658
rect 4330 1606 4342 1658
rect 4342 1606 4356 1658
rect 4380 1606 4394 1658
rect 4394 1606 4406 1658
rect 4406 1606 4436 1658
rect 4460 1606 4470 1658
rect 4470 1606 4516 1658
rect 4220 1604 4276 1606
rect 4300 1604 4356 1606
rect 4380 1604 4436 1606
rect 4460 1604 4516 1606
rect 8758 10376 8814 10432
rect 8220 9818 8276 9820
rect 8300 9818 8356 9820
rect 8380 9818 8436 9820
rect 8460 9818 8516 9820
rect 8220 9766 8266 9818
rect 8266 9766 8276 9818
rect 8300 9766 8330 9818
rect 8330 9766 8342 9818
rect 8342 9766 8356 9818
rect 8380 9766 8394 9818
rect 8394 9766 8406 9818
rect 8406 9766 8436 9818
rect 8460 9766 8470 9818
rect 8470 9766 8516 9818
rect 8220 9764 8276 9766
rect 8300 9764 8356 9766
rect 8380 9764 8436 9766
rect 8460 9764 8516 9766
rect 8220 8730 8276 8732
rect 8300 8730 8356 8732
rect 8380 8730 8436 8732
rect 8460 8730 8516 8732
rect 8220 8678 8266 8730
rect 8266 8678 8276 8730
rect 8300 8678 8330 8730
rect 8330 8678 8342 8730
rect 8342 8678 8356 8730
rect 8380 8678 8394 8730
rect 8394 8678 8406 8730
rect 8406 8678 8436 8730
rect 8460 8678 8470 8730
rect 8470 8678 8516 8730
rect 8220 8676 8276 8678
rect 8300 8676 8356 8678
rect 8380 8676 8436 8678
rect 8460 8676 8516 8678
rect 9034 10532 9090 10568
rect 9034 10512 9036 10532
rect 9036 10512 9088 10532
rect 9088 10512 9090 10532
rect 9218 12008 9274 12064
rect 9586 12144 9642 12200
rect 10322 12688 10378 12744
rect 10046 12280 10102 12336
rect 9770 11736 9826 11792
rect 9862 11600 9918 11656
rect 10414 12280 10470 12336
rect 10598 11892 10654 11928
rect 10598 11872 10600 11892
rect 10600 11872 10652 11892
rect 10652 11872 10654 11892
rect 9218 11056 9274 11112
rect 9494 10512 9550 10568
rect 10782 11736 10838 11792
rect 10506 11636 10508 11656
rect 10508 11636 10560 11656
rect 10560 11636 10562 11656
rect 10506 11600 10562 11636
rect 10414 11328 10470 11384
rect 10874 11600 10930 11656
rect 10966 11500 10968 11520
rect 10968 11500 11020 11520
rect 11020 11500 11022 11520
rect 10966 11464 11022 11500
rect 10966 11192 11022 11248
rect 10138 10648 10194 10704
rect 10322 10648 10378 10704
rect 10046 10124 10102 10160
rect 10046 10104 10048 10124
rect 10048 10104 10100 10124
rect 10100 10104 10102 10124
rect 9770 9968 9826 10024
rect 9494 8472 9550 8528
rect 8220 7642 8276 7644
rect 8300 7642 8356 7644
rect 8380 7642 8436 7644
rect 8460 7642 8516 7644
rect 8220 7590 8266 7642
rect 8266 7590 8276 7642
rect 8300 7590 8330 7642
rect 8330 7590 8342 7642
rect 8342 7590 8356 7642
rect 8380 7590 8394 7642
rect 8394 7590 8406 7642
rect 8406 7590 8436 7642
rect 8460 7590 8470 7642
rect 8470 7590 8516 7642
rect 8220 7588 8276 7590
rect 8300 7588 8356 7590
rect 8380 7588 8436 7590
rect 8460 7588 8516 7590
rect 10322 8744 10378 8800
rect 10966 10920 11022 10976
rect 10782 10784 10838 10840
rect 12220 13626 12276 13628
rect 12300 13626 12356 13628
rect 12380 13626 12436 13628
rect 12460 13626 12516 13628
rect 12220 13574 12266 13626
rect 12266 13574 12276 13626
rect 12300 13574 12330 13626
rect 12330 13574 12342 13626
rect 12342 13574 12356 13626
rect 12380 13574 12394 13626
rect 12394 13574 12406 13626
rect 12406 13574 12436 13626
rect 12460 13574 12470 13626
rect 12470 13574 12516 13626
rect 12220 13572 12276 13574
rect 12300 13572 12356 13574
rect 12380 13572 12436 13574
rect 12460 13572 12516 13574
rect 11610 12688 11666 12744
rect 12220 12538 12276 12540
rect 12300 12538 12356 12540
rect 12380 12538 12436 12540
rect 12460 12538 12516 12540
rect 12220 12486 12266 12538
rect 12266 12486 12276 12538
rect 12300 12486 12330 12538
rect 12330 12486 12342 12538
rect 12342 12486 12356 12538
rect 12380 12486 12394 12538
rect 12394 12486 12406 12538
rect 12406 12486 12436 12538
rect 12460 12486 12470 12538
rect 12470 12486 12516 12538
rect 12220 12484 12276 12486
rect 12300 12484 12356 12486
rect 12380 12484 12436 12486
rect 12460 12484 12516 12486
rect 11794 12144 11850 12200
rect 10598 8916 10600 8936
rect 10600 8916 10652 8936
rect 10652 8916 10654 8936
rect 10598 8880 10654 8916
rect 10506 8472 10562 8528
rect 8220 6554 8276 6556
rect 8300 6554 8356 6556
rect 8380 6554 8436 6556
rect 8460 6554 8516 6556
rect 8220 6502 8266 6554
rect 8266 6502 8276 6554
rect 8300 6502 8330 6554
rect 8330 6502 8342 6554
rect 8342 6502 8356 6554
rect 8380 6502 8394 6554
rect 8394 6502 8406 6554
rect 8406 6502 8436 6554
rect 8460 6502 8470 6554
rect 8470 6502 8516 6554
rect 8220 6500 8276 6502
rect 8300 6500 8356 6502
rect 8380 6500 8436 6502
rect 8460 6500 8516 6502
rect 9678 7404 9734 7440
rect 9678 7384 9680 7404
rect 9680 7384 9732 7404
rect 9732 7384 9734 7404
rect 10874 8472 10930 8528
rect 11702 10648 11758 10704
rect 11426 9560 11482 9616
rect 12162 11892 12218 11928
rect 12162 11872 12164 11892
rect 12164 11872 12216 11892
rect 12216 11872 12218 11892
rect 12254 11736 12310 11792
rect 12990 12144 13046 12200
rect 12220 11450 12276 11452
rect 12300 11450 12356 11452
rect 12380 11450 12436 11452
rect 12460 11450 12516 11452
rect 12220 11398 12266 11450
rect 12266 11398 12276 11450
rect 12300 11398 12330 11450
rect 12330 11398 12342 11450
rect 12342 11398 12356 11450
rect 12380 11398 12394 11450
rect 12394 11398 12406 11450
rect 12406 11398 12436 11450
rect 12460 11398 12470 11450
rect 12470 11398 12516 11450
rect 12220 11396 12276 11398
rect 12300 11396 12356 11398
rect 12380 11396 12436 11398
rect 12460 11396 12516 11398
rect 12070 11328 12126 11384
rect 12162 10784 12218 10840
rect 12254 10648 12310 10704
rect 12530 10512 12586 10568
rect 12220 10362 12276 10364
rect 12300 10362 12356 10364
rect 12380 10362 12436 10364
rect 12460 10362 12516 10364
rect 12220 10310 12266 10362
rect 12266 10310 12276 10362
rect 12300 10310 12330 10362
rect 12330 10310 12342 10362
rect 12342 10310 12356 10362
rect 12380 10310 12394 10362
rect 12394 10310 12406 10362
rect 12406 10310 12436 10362
rect 12460 10310 12470 10362
rect 12470 10310 12516 10362
rect 12220 10308 12276 10310
rect 12300 10308 12356 10310
rect 12380 10308 12436 10310
rect 12460 10308 12516 10310
rect 11886 9968 11942 10024
rect 11886 8744 11942 8800
rect 11702 8608 11758 8664
rect 11426 8336 11482 8392
rect 12898 11600 12954 11656
rect 13266 11056 13322 11112
rect 13450 10920 13506 10976
rect 12220 9274 12276 9276
rect 12300 9274 12356 9276
rect 12380 9274 12436 9276
rect 12460 9274 12516 9276
rect 12220 9222 12266 9274
rect 12266 9222 12276 9274
rect 12300 9222 12330 9274
rect 12330 9222 12342 9274
rect 12342 9222 12356 9274
rect 12380 9222 12394 9274
rect 12394 9222 12406 9274
rect 12406 9222 12436 9274
rect 12460 9222 12470 9274
rect 12470 9222 12516 9274
rect 12220 9220 12276 9222
rect 12300 9220 12356 9222
rect 12380 9220 12436 9222
rect 12460 9220 12516 9222
rect 12254 8508 12256 8528
rect 12256 8508 12308 8528
rect 12308 8508 12310 8528
rect 12254 8472 12310 8508
rect 11518 7928 11574 7984
rect 10506 7404 10562 7440
rect 10506 7384 10508 7404
rect 10508 7384 10560 7404
rect 10560 7384 10562 7404
rect 8220 5466 8276 5468
rect 8300 5466 8356 5468
rect 8380 5466 8436 5468
rect 8460 5466 8516 5468
rect 8220 5414 8266 5466
rect 8266 5414 8276 5466
rect 8300 5414 8330 5466
rect 8330 5414 8342 5466
rect 8342 5414 8356 5466
rect 8380 5414 8394 5466
rect 8394 5414 8406 5466
rect 8406 5414 8436 5466
rect 8460 5414 8470 5466
rect 8470 5414 8516 5466
rect 8220 5412 8276 5414
rect 8300 5412 8356 5414
rect 8380 5412 8436 5414
rect 8460 5412 8516 5414
rect 8220 4378 8276 4380
rect 8300 4378 8356 4380
rect 8380 4378 8436 4380
rect 8460 4378 8516 4380
rect 8220 4326 8266 4378
rect 8266 4326 8276 4378
rect 8300 4326 8330 4378
rect 8330 4326 8342 4378
rect 8342 4326 8356 4378
rect 8380 4326 8394 4378
rect 8394 4326 8406 4378
rect 8406 4326 8436 4378
rect 8460 4326 8470 4378
rect 8470 4326 8516 4378
rect 8220 4324 8276 4326
rect 8300 4324 8356 4326
rect 8380 4324 8436 4326
rect 8460 4324 8516 4326
rect 8220 3290 8276 3292
rect 8300 3290 8356 3292
rect 8380 3290 8436 3292
rect 8460 3290 8516 3292
rect 8220 3238 8266 3290
rect 8266 3238 8276 3290
rect 8300 3238 8330 3290
rect 8330 3238 8342 3290
rect 8342 3238 8356 3290
rect 8380 3238 8394 3290
rect 8394 3238 8406 3290
rect 8406 3238 8436 3290
rect 8460 3238 8470 3290
rect 8470 3238 8516 3290
rect 8220 3236 8276 3238
rect 8300 3236 8356 3238
rect 8380 3236 8436 3238
rect 8460 3236 8516 3238
rect 12220 8186 12276 8188
rect 12300 8186 12356 8188
rect 12380 8186 12436 8188
rect 12460 8186 12516 8188
rect 12220 8134 12266 8186
rect 12266 8134 12276 8186
rect 12300 8134 12330 8186
rect 12330 8134 12342 8186
rect 12342 8134 12356 8186
rect 12380 8134 12394 8186
rect 12394 8134 12406 8186
rect 12406 8134 12436 8186
rect 12460 8134 12470 8186
rect 12470 8134 12516 8186
rect 12220 8132 12276 8134
rect 12300 8132 12356 8134
rect 12380 8132 12436 8134
rect 12460 8132 12516 8134
rect 12220 7098 12276 7100
rect 12300 7098 12356 7100
rect 12380 7098 12436 7100
rect 12460 7098 12516 7100
rect 12220 7046 12266 7098
rect 12266 7046 12276 7098
rect 12300 7046 12330 7098
rect 12330 7046 12342 7098
rect 12342 7046 12356 7098
rect 12380 7046 12394 7098
rect 12394 7046 12406 7098
rect 12406 7046 12436 7098
rect 12460 7046 12470 7098
rect 12470 7046 12516 7098
rect 12220 7044 12276 7046
rect 12300 7044 12356 7046
rect 12380 7044 12436 7046
rect 12460 7044 12516 7046
rect 12220 6010 12276 6012
rect 12300 6010 12356 6012
rect 12380 6010 12436 6012
rect 12460 6010 12516 6012
rect 12220 5958 12266 6010
rect 12266 5958 12276 6010
rect 12300 5958 12330 6010
rect 12330 5958 12342 6010
rect 12342 5958 12356 6010
rect 12380 5958 12394 6010
rect 12394 5958 12406 6010
rect 12406 5958 12436 6010
rect 12460 5958 12470 6010
rect 12470 5958 12516 6010
rect 12220 5956 12276 5958
rect 12300 5956 12356 5958
rect 12380 5956 12436 5958
rect 12460 5956 12516 5958
rect 8220 2202 8276 2204
rect 8300 2202 8356 2204
rect 8380 2202 8436 2204
rect 8460 2202 8516 2204
rect 8220 2150 8266 2202
rect 8266 2150 8276 2202
rect 8300 2150 8330 2202
rect 8330 2150 8342 2202
rect 8342 2150 8356 2202
rect 8380 2150 8394 2202
rect 8394 2150 8406 2202
rect 8406 2150 8436 2202
rect 8460 2150 8470 2202
rect 8470 2150 8516 2202
rect 8220 2148 8276 2150
rect 8300 2148 8356 2150
rect 8380 2148 8436 2150
rect 8460 2148 8516 2150
rect 12220 4922 12276 4924
rect 12300 4922 12356 4924
rect 12380 4922 12436 4924
rect 12460 4922 12516 4924
rect 12220 4870 12266 4922
rect 12266 4870 12276 4922
rect 12300 4870 12330 4922
rect 12330 4870 12342 4922
rect 12342 4870 12356 4922
rect 12380 4870 12394 4922
rect 12394 4870 12406 4922
rect 12406 4870 12436 4922
rect 12460 4870 12470 4922
rect 12470 4870 12516 4922
rect 12220 4868 12276 4870
rect 12300 4868 12356 4870
rect 12380 4868 12436 4870
rect 12460 4868 12516 4870
rect 12898 8880 12954 8936
rect 14094 12008 14150 12064
rect 14002 10648 14058 10704
rect 14002 9424 14058 9480
rect 13910 9016 13966 9072
rect 13450 8356 13506 8392
rect 13450 8336 13452 8356
rect 13452 8336 13504 8356
rect 13504 8336 13506 8356
rect 13726 8472 13782 8528
rect 15198 13504 15254 13560
rect 16220 13082 16276 13084
rect 16300 13082 16356 13084
rect 16380 13082 16436 13084
rect 16460 13082 16516 13084
rect 16220 13030 16266 13082
rect 16266 13030 16276 13082
rect 16300 13030 16330 13082
rect 16330 13030 16342 13082
rect 16342 13030 16356 13082
rect 16380 13030 16394 13082
rect 16394 13030 16406 13082
rect 16406 13030 16436 13082
rect 16460 13030 16470 13082
rect 16470 13030 16516 13082
rect 16220 13028 16276 13030
rect 16300 13028 16356 13030
rect 16380 13028 16436 13030
rect 16460 13028 16516 13030
rect 15106 10104 15162 10160
rect 14554 8916 14556 8936
rect 14556 8916 14608 8936
rect 14608 8916 14610 8936
rect 14554 8880 14610 8916
rect 15198 8880 15254 8936
rect 15014 8608 15070 8664
rect 14830 7928 14886 7984
rect 15658 9424 15714 9480
rect 15474 8880 15530 8936
rect 12220 3834 12276 3836
rect 12300 3834 12356 3836
rect 12380 3834 12436 3836
rect 12460 3834 12516 3836
rect 12220 3782 12266 3834
rect 12266 3782 12276 3834
rect 12300 3782 12330 3834
rect 12330 3782 12342 3834
rect 12342 3782 12356 3834
rect 12380 3782 12394 3834
rect 12394 3782 12406 3834
rect 12406 3782 12436 3834
rect 12460 3782 12470 3834
rect 12470 3782 12516 3834
rect 12220 3780 12276 3782
rect 12300 3780 12356 3782
rect 12380 3780 12436 3782
rect 12460 3780 12516 3782
rect 10690 3032 10746 3088
rect 11610 3052 11666 3088
rect 11610 3032 11612 3052
rect 11612 3032 11664 3052
rect 11664 3032 11666 3052
rect 12220 2746 12276 2748
rect 12300 2746 12356 2748
rect 12380 2746 12436 2748
rect 12460 2746 12516 2748
rect 12220 2694 12266 2746
rect 12266 2694 12276 2746
rect 12300 2694 12330 2746
rect 12330 2694 12342 2746
rect 12342 2694 12356 2746
rect 12380 2694 12394 2746
rect 12394 2694 12406 2746
rect 12406 2694 12436 2746
rect 12460 2694 12470 2746
rect 12470 2694 12516 2746
rect 12220 2692 12276 2694
rect 12300 2692 12356 2694
rect 12380 2692 12436 2694
rect 12460 2692 12516 2694
rect 12220 1658 12276 1660
rect 12300 1658 12356 1660
rect 12380 1658 12436 1660
rect 12460 1658 12516 1660
rect 12220 1606 12266 1658
rect 12266 1606 12276 1658
rect 12300 1606 12330 1658
rect 12330 1606 12342 1658
rect 12342 1606 12356 1658
rect 12380 1606 12394 1658
rect 12394 1606 12406 1658
rect 12406 1606 12436 1658
rect 12460 1606 12470 1658
rect 12470 1606 12516 1658
rect 12220 1604 12276 1606
rect 12300 1604 12356 1606
rect 12380 1604 12436 1606
rect 12460 1604 12516 1606
rect 8220 1114 8276 1116
rect 8300 1114 8356 1116
rect 8380 1114 8436 1116
rect 8460 1114 8516 1116
rect 8220 1062 8266 1114
rect 8266 1062 8276 1114
rect 8300 1062 8330 1114
rect 8330 1062 8342 1114
rect 8342 1062 8356 1114
rect 8380 1062 8394 1114
rect 8394 1062 8406 1114
rect 8406 1062 8436 1114
rect 8460 1062 8470 1114
rect 8470 1062 8516 1114
rect 8220 1060 8276 1062
rect 8300 1060 8356 1062
rect 8380 1060 8436 1062
rect 8460 1060 8516 1062
rect 15934 11192 15990 11248
rect 15842 9560 15898 9616
rect 16220 11994 16276 11996
rect 16300 11994 16356 11996
rect 16380 11994 16436 11996
rect 16460 11994 16516 11996
rect 16220 11942 16266 11994
rect 16266 11942 16276 11994
rect 16300 11942 16330 11994
rect 16330 11942 16342 11994
rect 16342 11942 16356 11994
rect 16380 11942 16394 11994
rect 16394 11942 16406 11994
rect 16406 11942 16436 11994
rect 16460 11942 16470 11994
rect 16470 11942 16516 11994
rect 16220 11940 16276 11942
rect 16300 11940 16356 11942
rect 16380 11940 16436 11942
rect 16460 11940 16516 11942
rect 16026 11056 16082 11112
rect 16220 10906 16276 10908
rect 16300 10906 16356 10908
rect 16380 10906 16436 10908
rect 16460 10906 16516 10908
rect 16220 10854 16266 10906
rect 16266 10854 16276 10906
rect 16300 10854 16330 10906
rect 16330 10854 16342 10906
rect 16342 10854 16356 10906
rect 16380 10854 16394 10906
rect 16394 10854 16406 10906
rect 16406 10854 16436 10906
rect 16460 10854 16470 10906
rect 16470 10854 16516 10906
rect 16220 10852 16276 10854
rect 16300 10852 16356 10854
rect 16380 10852 16436 10854
rect 16460 10852 16516 10854
rect 16220 9818 16276 9820
rect 16300 9818 16356 9820
rect 16380 9818 16436 9820
rect 16460 9818 16516 9820
rect 16220 9766 16266 9818
rect 16266 9766 16276 9818
rect 16300 9766 16330 9818
rect 16330 9766 16342 9818
rect 16342 9766 16356 9818
rect 16380 9766 16394 9818
rect 16394 9766 16406 9818
rect 16406 9766 16436 9818
rect 16460 9766 16470 9818
rect 16470 9766 16516 9818
rect 16220 9764 16276 9766
rect 16300 9764 16356 9766
rect 16380 9764 16436 9766
rect 16460 9764 16516 9766
rect 18786 12280 18842 12336
rect 16220 8730 16276 8732
rect 16300 8730 16356 8732
rect 16380 8730 16436 8732
rect 16460 8730 16516 8732
rect 16220 8678 16266 8730
rect 16266 8678 16276 8730
rect 16300 8678 16330 8730
rect 16330 8678 16342 8730
rect 16342 8678 16356 8730
rect 16380 8678 16394 8730
rect 16394 8678 16406 8730
rect 16406 8678 16436 8730
rect 16460 8678 16470 8730
rect 16470 8678 16516 8730
rect 16220 8676 16276 8678
rect 16300 8676 16356 8678
rect 16380 8676 16436 8678
rect 16460 8676 16516 8678
rect 16220 7642 16276 7644
rect 16300 7642 16356 7644
rect 16380 7642 16436 7644
rect 16460 7642 16516 7644
rect 16220 7590 16266 7642
rect 16266 7590 16276 7642
rect 16300 7590 16330 7642
rect 16330 7590 16342 7642
rect 16342 7590 16356 7642
rect 16380 7590 16394 7642
rect 16394 7590 16406 7642
rect 16406 7590 16436 7642
rect 16460 7590 16470 7642
rect 16470 7590 16516 7642
rect 16220 7588 16276 7590
rect 16300 7588 16356 7590
rect 16380 7588 16436 7590
rect 16460 7588 16516 7590
rect 16220 6554 16276 6556
rect 16300 6554 16356 6556
rect 16380 6554 16436 6556
rect 16460 6554 16516 6556
rect 16220 6502 16266 6554
rect 16266 6502 16276 6554
rect 16300 6502 16330 6554
rect 16330 6502 16342 6554
rect 16342 6502 16356 6554
rect 16380 6502 16394 6554
rect 16394 6502 16406 6554
rect 16406 6502 16436 6554
rect 16460 6502 16470 6554
rect 16470 6502 16516 6554
rect 16220 6500 16276 6502
rect 16300 6500 16356 6502
rect 16380 6500 16436 6502
rect 16460 6500 16516 6502
rect 16220 5466 16276 5468
rect 16300 5466 16356 5468
rect 16380 5466 16436 5468
rect 16460 5466 16516 5468
rect 16220 5414 16266 5466
rect 16266 5414 16276 5466
rect 16300 5414 16330 5466
rect 16330 5414 16342 5466
rect 16342 5414 16356 5466
rect 16380 5414 16394 5466
rect 16394 5414 16406 5466
rect 16406 5414 16436 5466
rect 16460 5414 16470 5466
rect 16470 5414 16516 5466
rect 16220 5412 16276 5414
rect 16300 5412 16356 5414
rect 16380 5412 16436 5414
rect 16460 5412 16516 5414
rect 16220 4378 16276 4380
rect 16300 4378 16356 4380
rect 16380 4378 16436 4380
rect 16460 4378 16516 4380
rect 16220 4326 16266 4378
rect 16266 4326 16276 4378
rect 16300 4326 16330 4378
rect 16330 4326 16342 4378
rect 16342 4326 16356 4378
rect 16380 4326 16394 4378
rect 16394 4326 16406 4378
rect 16406 4326 16436 4378
rect 16460 4326 16470 4378
rect 16470 4326 16516 4378
rect 16220 4324 16276 4326
rect 16300 4324 16356 4326
rect 16380 4324 16436 4326
rect 16460 4324 16516 4326
rect 16220 3290 16276 3292
rect 16300 3290 16356 3292
rect 16380 3290 16436 3292
rect 16460 3290 16516 3292
rect 16220 3238 16266 3290
rect 16266 3238 16276 3290
rect 16300 3238 16330 3290
rect 16330 3238 16342 3290
rect 16342 3238 16356 3290
rect 16380 3238 16394 3290
rect 16394 3238 16406 3290
rect 16406 3238 16436 3290
rect 16460 3238 16470 3290
rect 16470 3238 16516 3290
rect 16220 3236 16276 3238
rect 16300 3236 16356 3238
rect 16380 3236 16436 3238
rect 16460 3236 16516 3238
rect 16220 2202 16276 2204
rect 16300 2202 16356 2204
rect 16380 2202 16436 2204
rect 16460 2202 16516 2204
rect 16220 2150 16266 2202
rect 16266 2150 16276 2202
rect 16300 2150 16330 2202
rect 16330 2150 16342 2202
rect 16342 2150 16356 2202
rect 16380 2150 16394 2202
rect 16394 2150 16406 2202
rect 16406 2150 16436 2202
rect 16460 2150 16470 2202
rect 16470 2150 16516 2202
rect 16220 2148 16276 2150
rect 16300 2148 16356 2150
rect 16380 2148 16436 2150
rect 16460 2148 16516 2150
rect 15566 1264 15622 1320
rect 17038 3032 17094 3088
rect 17774 6160 17830 6216
rect 18418 3712 18474 3768
rect 16220 1114 16276 1116
rect 16300 1114 16356 1116
rect 16380 1114 16436 1116
rect 16460 1114 16516 1116
rect 16220 1062 16266 1114
rect 16266 1062 16276 1114
rect 16300 1062 16330 1114
rect 16330 1062 16342 1114
rect 16342 1062 16356 1114
rect 16380 1062 16394 1114
rect 16394 1062 16406 1114
rect 16406 1062 16436 1114
rect 16460 1062 16470 1114
rect 16470 1062 16516 1114
rect 16220 1060 16276 1062
rect 16300 1060 16356 1062
rect 16380 1060 16436 1062
rect 16460 1060 16516 1062
<< metal3 >>
rect 4210 13632 4526 13633
rect 0 13562 800 13592
rect 4210 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4526 13632
rect 4210 13567 4526 13568
rect 12210 13632 12526 13633
rect 12210 13568 12216 13632
rect 12280 13568 12296 13632
rect 12360 13568 12376 13632
rect 12440 13568 12456 13632
rect 12520 13568 12526 13632
rect 12210 13567 12526 13568
rect 3417 13562 3483 13565
rect 0 13560 3483 13562
rect 0 13504 3422 13560
rect 3478 13504 3483 13560
rect 0 13502 3483 13504
rect 0 13472 800 13502
rect 3417 13499 3483 13502
rect 15193 13562 15259 13565
rect 19200 13562 20000 13592
rect 15193 13560 20000 13562
rect 15193 13504 15198 13560
rect 15254 13504 20000 13560
rect 15193 13502 20000 13504
rect 15193 13499 15259 13502
rect 19200 13472 20000 13502
rect 8210 13088 8526 13089
rect 8210 13024 8216 13088
rect 8280 13024 8296 13088
rect 8360 13024 8376 13088
rect 8440 13024 8456 13088
rect 8520 13024 8526 13088
rect 8210 13023 8526 13024
rect 16210 13088 16526 13089
rect 16210 13024 16216 13088
rect 16280 13024 16296 13088
rect 16360 13024 16376 13088
rect 16440 13024 16456 13088
rect 16520 13024 16526 13088
rect 16210 13023 16526 13024
rect 0 12746 800 12776
rect 2773 12746 2839 12749
rect 0 12744 2839 12746
rect 0 12688 2778 12744
rect 2834 12688 2839 12744
rect 0 12686 2839 12688
rect 0 12656 800 12686
rect 2773 12683 2839 12686
rect 10317 12746 10383 12749
rect 11605 12746 11671 12749
rect 10317 12744 11671 12746
rect 10317 12688 10322 12744
rect 10378 12688 11610 12744
rect 11666 12688 11671 12744
rect 10317 12686 11671 12688
rect 10317 12683 10383 12686
rect 11605 12683 11671 12686
rect 4210 12544 4526 12545
rect 4210 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4526 12544
rect 4210 12479 4526 12480
rect 12210 12544 12526 12545
rect 12210 12480 12216 12544
rect 12280 12480 12296 12544
rect 12360 12480 12376 12544
rect 12440 12480 12456 12544
rect 12520 12480 12526 12544
rect 12210 12479 12526 12480
rect 10041 12338 10107 12341
rect 10409 12338 10475 12341
rect 18781 12338 18847 12341
rect 10041 12336 18847 12338
rect 10041 12280 10046 12336
rect 10102 12280 10414 12336
rect 10470 12280 18786 12336
rect 18842 12280 18847 12336
rect 10041 12278 18847 12280
rect 10041 12275 10107 12278
rect 10409 12275 10475 12278
rect 18781 12275 18847 12278
rect 8477 12202 8543 12205
rect 8845 12202 8911 12205
rect 9581 12202 9647 12205
rect 8477 12200 9647 12202
rect 8477 12144 8482 12200
rect 8538 12144 8850 12200
rect 8906 12144 9586 12200
rect 9642 12144 9647 12200
rect 8477 12142 9647 12144
rect 8477 12139 8543 12142
rect 8845 12139 8911 12142
rect 9581 12139 9647 12142
rect 11789 12202 11855 12205
rect 12985 12202 13051 12205
rect 11789 12200 13051 12202
rect 11789 12144 11794 12200
rect 11850 12144 12990 12200
rect 13046 12144 13051 12200
rect 11789 12142 13051 12144
rect 11789 12139 11855 12142
rect 12985 12139 13051 12142
rect 9213 12066 9279 12069
rect 14089 12066 14155 12069
rect 9213 12064 14155 12066
rect 9213 12008 9218 12064
rect 9274 12008 14094 12064
rect 14150 12008 14155 12064
rect 9213 12006 14155 12008
rect 9213 12003 9279 12006
rect 14089 12003 14155 12006
rect 8210 12000 8526 12001
rect 0 11930 800 11960
rect 8210 11936 8216 12000
rect 8280 11936 8296 12000
rect 8360 11936 8376 12000
rect 8440 11936 8456 12000
rect 8520 11936 8526 12000
rect 8210 11935 8526 11936
rect 16210 12000 16526 12001
rect 16210 11936 16216 12000
rect 16280 11936 16296 12000
rect 16360 11936 16376 12000
rect 16440 11936 16456 12000
rect 16520 11936 16526 12000
rect 16210 11935 16526 11936
rect 3417 11930 3483 11933
rect 0 11928 3483 11930
rect 0 11872 3422 11928
rect 3478 11872 3483 11928
rect 0 11870 3483 11872
rect 0 11840 800 11870
rect 3417 11867 3483 11870
rect 10593 11930 10659 11933
rect 12157 11930 12223 11933
rect 10593 11928 12223 11930
rect 10593 11872 10598 11928
rect 10654 11872 12162 11928
rect 12218 11872 12223 11928
rect 10593 11870 12223 11872
rect 10593 11867 10659 11870
rect 12157 11867 12223 11870
rect 6913 11794 6979 11797
rect 9765 11794 9831 11797
rect 6913 11792 9831 11794
rect 6913 11736 6918 11792
rect 6974 11736 9770 11792
rect 9826 11736 9831 11792
rect 6913 11734 9831 11736
rect 6913 11731 6979 11734
rect 9765 11731 9831 11734
rect 10777 11794 10843 11797
rect 12249 11794 12315 11797
rect 10777 11792 12315 11794
rect 10777 11736 10782 11792
rect 10838 11736 12254 11792
rect 12310 11736 12315 11792
rect 10777 11734 12315 11736
rect 10777 11731 10843 11734
rect 12249 11731 12315 11734
rect 9857 11658 9923 11661
rect 10501 11658 10567 11661
rect 9857 11656 10567 11658
rect 9857 11600 9862 11656
rect 9918 11600 10506 11656
rect 10562 11600 10567 11656
rect 9857 11598 10567 11600
rect 9857 11595 9923 11598
rect 10501 11595 10567 11598
rect 10869 11658 10935 11661
rect 12893 11658 12959 11661
rect 10869 11656 12959 11658
rect 10869 11600 10874 11656
rect 10930 11600 12898 11656
rect 12954 11600 12959 11656
rect 10869 11598 12959 11600
rect 10869 11595 10935 11598
rect 12893 11595 12959 11598
rect 6821 11522 6887 11525
rect 10961 11522 11027 11525
rect 6821 11520 11027 11522
rect 6821 11464 6826 11520
rect 6882 11464 10966 11520
rect 11022 11464 11027 11520
rect 6821 11462 11027 11464
rect 6821 11459 6887 11462
rect 10961 11459 11027 11462
rect 4210 11456 4526 11457
rect 4210 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4526 11456
rect 4210 11391 4526 11392
rect 12210 11456 12526 11457
rect 12210 11392 12216 11456
rect 12280 11392 12296 11456
rect 12360 11392 12376 11456
rect 12440 11392 12456 11456
rect 12520 11392 12526 11456
rect 12210 11391 12526 11392
rect 10409 11386 10475 11389
rect 12065 11386 12131 11389
rect 10409 11384 12131 11386
rect 10409 11328 10414 11384
rect 10470 11328 12070 11384
rect 12126 11328 12131 11384
rect 10409 11326 12131 11328
rect 10409 11323 10475 11326
rect 12065 11323 12131 11326
rect 8293 11250 8359 11253
rect 10961 11250 11027 11253
rect 15929 11250 15995 11253
rect 8293 11248 8402 11250
rect 8293 11192 8298 11248
rect 8354 11192 8402 11248
rect 8293 11187 8402 11192
rect 10961 11248 15995 11250
rect 10961 11192 10966 11248
rect 11022 11192 15934 11248
rect 15990 11192 15995 11248
rect 10961 11190 15995 11192
rect 10961 11187 11027 11190
rect 15929 11187 15995 11190
rect 0 11114 800 11144
rect 4061 11114 4127 11117
rect 0 11112 4127 11114
rect 0 11056 4066 11112
rect 4122 11056 4127 11112
rect 0 11054 4127 11056
rect 8342 11114 8402 11187
rect 8661 11114 8727 11117
rect 9213 11114 9279 11117
rect 13261 11114 13327 11117
rect 8342 11112 13327 11114
rect 8342 11056 8666 11112
rect 8722 11056 9218 11112
rect 9274 11056 13266 11112
rect 13322 11056 13327 11112
rect 8342 11054 13327 11056
rect 0 11024 800 11054
rect 4061 11051 4127 11054
rect 8661 11051 8727 11054
rect 9213 11051 9279 11054
rect 13261 11051 13327 11054
rect 16021 11114 16087 11117
rect 19200 11114 20000 11144
rect 16021 11112 20000 11114
rect 16021 11056 16026 11112
rect 16082 11056 20000 11112
rect 16021 11054 20000 11056
rect 16021 11051 16087 11054
rect 19200 11024 20000 11054
rect 10961 10978 11027 10981
rect 13445 10978 13511 10981
rect 10961 10976 13511 10978
rect 10961 10920 10966 10976
rect 11022 10920 13450 10976
rect 13506 10920 13511 10976
rect 10961 10918 13511 10920
rect 10961 10915 11027 10918
rect 13445 10915 13511 10918
rect 8210 10912 8526 10913
rect 8210 10848 8216 10912
rect 8280 10848 8296 10912
rect 8360 10848 8376 10912
rect 8440 10848 8456 10912
rect 8520 10848 8526 10912
rect 8210 10847 8526 10848
rect 16210 10912 16526 10913
rect 16210 10848 16216 10912
rect 16280 10848 16296 10912
rect 16360 10848 16376 10912
rect 16440 10848 16456 10912
rect 16520 10848 16526 10912
rect 16210 10847 16526 10848
rect 10777 10842 10843 10845
rect 12157 10842 12223 10845
rect 10777 10840 12223 10842
rect 10777 10784 10782 10840
rect 10838 10784 12162 10840
rect 12218 10784 12223 10840
rect 10777 10782 12223 10784
rect 10777 10779 10843 10782
rect 12157 10779 12223 10782
rect 7005 10706 7071 10709
rect 8293 10706 8359 10709
rect 10133 10706 10199 10709
rect 7005 10704 10199 10706
rect 7005 10648 7010 10704
rect 7066 10648 8298 10704
rect 8354 10648 10138 10704
rect 10194 10648 10199 10704
rect 7005 10646 10199 10648
rect 7005 10643 7071 10646
rect 8293 10643 8359 10646
rect 10133 10643 10199 10646
rect 10317 10706 10383 10709
rect 11697 10706 11763 10709
rect 10317 10704 11763 10706
rect 10317 10648 10322 10704
rect 10378 10648 11702 10704
rect 11758 10648 11763 10704
rect 10317 10646 11763 10648
rect 10317 10643 10383 10646
rect 11697 10643 11763 10646
rect 12249 10706 12315 10709
rect 13997 10706 14063 10709
rect 12249 10704 14063 10706
rect 12249 10648 12254 10704
rect 12310 10648 14002 10704
rect 14058 10648 14063 10704
rect 12249 10646 14063 10648
rect 12249 10643 12315 10646
rect 13997 10643 14063 10646
rect 2037 10570 2103 10573
rect 9029 10570 9095 10573
rect 2037 10568 9095 10570
rect 2037 10512 2042 10568
rect 2098 10512 9034 10568
rect 9090 10512 9095 10568
rect 2037 10510 9095 10512
rect 2037 10507 2103 10510
rect 9029 10507 9095 10510
rect 9489 10570 9555 10573
rect 12525 10570 12591 10573
rect 9489 10568 12591 10570
rect 9489 10512 9494 10568
rect 9550 10512 12530 10568
rect 12586 10512 12591 10568
rect 9489 10510 12591 10512
rect 9489 10507 9555 10510
rect 12525 10507 12591 10510
rect 8109 10434 8175 10437
rect 8753 10434 8819 10437
rect 8109 10432 8819 10434
rect 8109 10376 8114 10432
rect 8170 10376 8758 10432
rect 8814 10376 8819 10432
rect 8109 10374 8819 10376
rect 8109 10371 8175 10374
rect 8753 10371 8819 10374
rect 4210 10368 4526 10369
rect 0 10298 800 10328
rect 4210 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4526 10368
rect 4210 10303 4526 10304
rect 12210 10368 12526 10369
rect 12210 10304 12216 10368
rect 12280 10304 12296 10368
rect 12360 10304 12376 10368
rect 12440 10304 12456 10368
rect 12520 10304 12526 10368
rect 12210 10303 12526 10304
rect 3785 10298 3851 10301
rect 0 10296 3851 10298
rect 0 10240 3790 10296
rect 3846 10240 3851 10296
rect 0 10238 3851 10240
rect 0 10208 800 10238
rect 3785 10235 3851 10238
rect 10041 10162 10107 10165
rect 15101 10162 15167 10165
rect 10041 10160 15167 10162
rect 10041 10104 10046 10160
rect 10102 10104 15106 10160
rect 15162 10104 15167 10160
rect 10041 10102 15167 10104
rect 10041 10099 10107 10102
rect 15101 10099 15167 10102
rect 9765 10026 9831 10029
rect 11881 10026 11947 10029
rect 9765 10024 11947 10026
rect 9765 9968 9770 10024
rect 9826 9968 11886 10024
rect 11942 9968 11947 10024
rect 9765 9966 11947 9968
rect 9765 9963 9831 9966
rect 11881 9963 11947 9966
rect 8210 9824 8526 9825
rect 8210 9760 8216 9824
rect 8280 9760 8296 9824
rect 8360 9760 8376 9824
rect 8440 9760 8456 9824
rect 8520 9760 8526 9824
rect 8210 9759 8526 9760
rect 16210 9824 16526 9825
rect 16210 9760 16216 9824
rect 16280 9760 16296 9824
rect 16360 9760 16376 9824
rect 16440 9760 16456 9824
rect 16520 9760 16526 9824
rect 16210 9759 16526 9760
rect 11421 9618 11487 9621
rect 15837 9618 15903 9621
rect 11421 9616 15903 9618
rect 11421 9560 11426 9616
rect 11482 9560 15842 9616
rect 15898 9560 15903 9616
rect 11421 9558 15903 9560
rect 11421 9555 11487 9558
rect 15837 9555 15903 9558
rect 0 9482 800 9512
rect 1761 9482 1827 9485
rect 0 9480 1827 9482
rect 0 9424 1766 9480
rect 1822 9424 1827 9480
rect 0 9422 1827 9424
rect 0 9392 800 9422
rect 1761 9419 1827 9422
rect 13997 9482 14063 9485
rect 15653 9482 15719 9485
rect 13997 9480 15719 9482
rect 13997 9424 14002 9480
rect 14058 9424 15658 9480
rect 15714 9424 15719 9480
rect 13997 9422 15719 9424
rect 13997 9419 14063 9422
rect 15653 9419 15719 9422
rect 4210 9280 4526 9281
rect 4210 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4526 9280
rect 4210 9215 4526 9216
rect 12210 9280 12526 9281
rect 12210 9216 12216 9280
rect 12280 9216 12296 9280
rect 12360 9216 12376 9280
rect 12440 9216 12456 9280
rect 12520 9216 12526 9280
rect 12210 9215 12526 9216
rect 6637 9074 6703 9077
rect 13905 9074 13971 9077
rect 6637 9072 13971 9074
rect 6637 9016 6642 9072
rect 6698 9016 13910 9072
rect 13966 9016 13971 9072
rect 6637 9014 13971 9016
rect 6637 9011 6703 9014
rect 13905 9011 13971 9014
rect 5993 8938 6059 8941
rect 7833 8938 7899 8941
rect 5993 8936 7899 8938
rect 5993 8880 5998 8936
rect 6054 8880 7838 8936
rect 7894 8880 7899 8936
rect 5993 8878 7899 8880
rect 5993 8875 6059 8878
rect 7833 8875 7899 8878
rect 10593 8938 10659 8941
rect 12893 8938 12959 8941
rect 14549 8938 14615 8941
rect 10593 8936 14615 8938
rect 10593 8880 10598 8936
rect 10654 8880 12898 8936
rect 12954 8880 14554 8936
rect 14610 8880 14615 8936
rect 10593 8878 14615 8880
rect 10593 8875 10659 8878
rect 12893 8875 12959 8878
rect 14549 8875 14615 8878
rect 15193 8938 15259 8941
rect 15469 8938 15535 8941
rect 15193 8936 16682 8938
rect 15193 8880 15198 8936
rect 15254 8880 15474 8936
rect 15530 8880 16682 8936
rect 15193 8878 16682 8880
rect 15193 8875 15259 8878
rect 15469 8875 15535 8878
rect 10317 8802 10383 8805
rect 11881 8802 11947 8805
rect 10317 8800 11947 8802
rect 10317 8744 10322 8800
rect 10378 8744 11886 8800
rect 11942 8744 11947 8800
rect 10317 8742 11947 8744
rect 10317 8739 10383 8742
rect 11881 8739 11947 8742
rect 8210 8736 8526 8737
rect 0 8666 800 8696
rect 8210 8672 8216 8736
rect 8280 8672 8296 8736
rect 8360 8672 8376 8736
rect 8440 8672 8456 8736
rect 8520 8672 8526 8736
rect 8210 8671 8526 8672
rect 16210 8736 16526 8737
rect 16210 8672 16216 8736
rect 16280 8672 16296 8736
rect 16360 8672 16376 8736
rect 16440 8672 16456 8736
rect 16520 8672 16526 8736
rect 16210 8671 16526 8672
rect 3969 8666 4035 8669
rect 0 8664 4035 8666
rect 0 8608 3974 8664
rect 4030 8608 4035 8664
rect 0 8606 4035 8608
rect 0 8576 800 8606
rect 3969 8603 4035 8606
rect 11697 8666 11763 8669
rect 15009 8666 15075 8669
rect 11697 8664 15075 8666
rect 11697 8608 11702 8664
rect 11758 8608 15014 8664
rect 15070 8608 15075 8664
rect 11697 8606 15075 8608
rect 16622 8666 16682 8878
rect 19200 8666 20000 8696
rect 16622 8606 20000 8666
rect 11697 8603 11763 8606
rect 15009 8603 15075 8606
rect 19200 8576 20000 8606
rect 9489 8530 9555 8533
rect 10501 8530 10567 8533
rect 10869 8530 10935 8533
rect 9489 8528 10935 8530
rect 9489 8472 9494 8528
rect 9550 8472 10506 8528
rect 10562 8472 10874 8528
rect 10930 8472 10935 8528
rect 9489 8470 10935 8472
rect 9489 8467 9555 8470
rect 10501 8467 10567 8470
rect 10869 8467 10935 8470
rect 12249 8530 12315 8533
rect 13721 8530 13787 8533
rect 12249 8528 13787 8530
rect 12249 8472 12254 8528
rect 12310 8472 13726 8528
rect 13782 8472 13787 8528
rect 12249 8470 13787 8472
rect 12249 8467 12315 8470
rect 13721 8467 13787 8470
rect 11421 8394 11487 8397
rect 13445 8394 13511 8397
rect 11421 8392 13511 8394
rect 11421 8336 11426 8392
rect 11482 8336 13450 8392
rect 13506 8336 13511 8392
rect 11421 8334 13511 8336
rect 11421 8331 11487 8334
rect 13445 8331 13511 8334
rect 4210 8192 4526 8193
rect 4210 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4526 8192
rect 4210 8127 4526 8128
rect 12210 8192 12526 8193
rect 12210 8128 12216 8192
rect 12280 8128 12296 8192
rect 12360 8128 12376 8192
rect 12440 8128 12456 8192
rect 12520 8128 12526 8192
rect 12210 8127 12526 8128
rect 11513 7986 11579 7989
rect 14825 7986 14891 7989
rect 11513 7984 14891 7986
rect 11513 7928 11518 7984
rect 11574 7928 14830 7984
rect 14886 7928 14891 7984
rect 11513 7926 14891 7928
rect 11513 7923 11579 7926
rect 14825 7923 14891 7926
rect 0 7850 800 7880
rect 3141 7850 3207 7853
rect 0 7848 3207 7850
rect 0 7792 3146 7848
rect 3202 7792 3207 7848
rect 0 7790 3207 7792
rect 0 7760 800 7790
rect 3141 7787 3207 7790
rect 8210 7648 8526 7649
rect 8210 7584 8216 7648
rect 8280 7584 8296 7648
rect 8360 7584 8376 7648
rect 8440 7584 8456 7648
rect 8520 7584 8526 7648
rect 8210 7583 8526 7584
rect 16210 7648 16526 7649
rect 16210 7584 16216 7648
rect 16280 7584 16296 7648
rect 16360 7584 16376 7648
rect 16440 7584 16456 7648
rect 16520 7584 16526 7648
rect 16210 7583 16526 7584
rect 9673 7442 9739 7445
rect 10501 7442 10567 7445
rect 9673 7440 10567 7442
rect 9673 7384 9678 7440
rect 9734 7384 10506 7440
rect 10562 7384 10567 7440
rect 9673 7382 10567 7384
rect 9673 7379 9739 7382
rect 10501 7379 10567 7382
rect 4210 7104 4526 7105
rect 0 7034 800 7064
rect 4210 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4526 7104
rect 4210 7039 4526 7040
rect 12210 7104 12526 7105
rect 12210 7040 12216 7104
rect 12280 7040 12296 7104
rect 12360 7040 12376 7104
rect 12440 7040 12456 7104
rect 12520 7040 12526 7104
rect 12210 7039 12526 7040
rect 2957 7034 3023 7037
rect 0 7032 3023 7034
rect 0 6976 2962 7032
rect 3018 6976 3023 7032
rect 0 6974 3023 6976
rect 0 6944 800 6974
rect 2957 6971 3023 6974
rect 8210 6560 8526 6561
rect 8210 6496 8216 6560
rect 8280 6496 8296 6560
rect 8360 6496 8376 6560
rect 8440 6496 8456 6560
rect 8520 6496 8526 6560
rect 8210 6495 8526 6496
rect 16210 6560 16526 6561
rect 16210 6496 16216 6560
rect 16280 6496 16296 6560
rect 16360 6496 16376 6560
rect 16440 6496 16456 6560
rect 16520 6496 16526 6560
rect 16210 6495 16526 6496
rect 0 6218 800 6248
rect 1577 6218 1643 6221
rect 0 6216 1643 6218
rect 0 6160 1582 6216
rect 1638 6160 1643 6216
rect 0 6158 1643 6160
rect 0 6128 800 6158
rect 1577 6155 1643 6158
rect 17769 6218 17835 6221
rect 19200 6218 20000 6248
rect 17769 6216 20000 6218
rect 17769 6160 17774 6216
rect 17830 6160 20000 6216
rect 17769 6158 20000 6160
rect 17769 6155 17835 6158
rect 19200 6128 20000 6158
rect 4210 6016 4526 6017
rect 4210 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4526 6016
rect 4210 5951 4526 5952
rect 12210 6016 12526 6017
rect 12210 5952 12216 6016
rect 12280 5952 12296 6016
rect 12360 5952 12376 6016
rect 12440 5952 12456 6016
rect 12520 5952 12526 6016
rect 12210 5951 12526 5952
rect 8210 5472 8526 5473
rect 0 5402 800 5432
rect 8210 5408 8216 5472
rect 8280 5408 8296 5472
rect 8360 5408 8376 5472
rect 8440 5408 8456 5472
rect 8520 5408 8526 5472
rect 8210 5407 8526 5408
rect 16210 5472 16526 5473
rect 16210 5408 16216 5472
rect 16280 5408 16296 5472
rect 16360 5408 16376 5472
rect 16440 5408 16456 5472
rect 16520 5408 16526 5472
rect 16210 5407 16526 5408
rect 1577 5402 1643 5405
rect 3693 5402 3759 5405
rect 0 5400 3759 5402
rect 0 5344 1582 5400
rect 1638 5344 3698 5400
rect 3754 5344 3759 5400
rect 0 5342 3759 5344
rect 0 5312 800 5342
rect 1577 5339 1643 5342
rect 3693 5339 3759 5342
rect 4210 4928 4526 4929
rect 4210 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4526 4928
rect 4210 4863 4526 4864
rect 12210 4928 12526 4929
rect 12210 4864 12216 4928
rect 12280 4864 12296 4928
rect 12360 4864 12376 4928
rect 12440 4864 12456 4928
rect 12520 4864 12526 4928
rect 12210 4863 12526 4864
rect 0 4586 800 4616
rect 2589 4586 2655 4589
rect 0 4584 2655 4586
rect 0 4528 2594 4584
rect 2650 4528 2655 4584
rect 0 4526 2655 4528
rect 0 4496 800 4526
rect 2589 4523 2655 4526
rect 8210 4384 8526 4385
rect 8210 4320 8216 4384
rect 8280 4320 8296 4384
rect 8360 4320 8376 4384
rect 8440 4320 8456 4384
rect 8520 4320 8526 4384
rect 8210 4319 8526 4320
rect 16210 4384 16526 4385
rect 16210 4320 16216 4384
rect 16280 4320 16296 4384
rect 16360 4320 16376 4384
rect 16440 4320 16456 4384
rect 16520 4320 16526 4384
rect 16210 4319 16526 4320
rect 4210 3840 4526 3841
rect 0 3770 800 3800
rect 4210 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4526 3840
rect 4210 3775 4526 3776
rect 12210 3840 12526 3841
rect 12210 3776 12216 3840
rect 12280 3776 12296 3840
rect 12360 3776 12376 3840
rect 12440 3776 12456 3840
rect 12520 3776 12526 3840
rect 12210 3775 12526 3776
rect 1761 3770 1827 3773
rect 0 3768 1827 3770
rect 0 3712 1766 3768
rect 1822 3712 1827 3768
rect 0 3710 1827 3712
rect 0 3680 800 3710
rect 1761 3707 1827 3710
rect 18413 3770 18479 3773
rect 19200 3770 20000 3800
rect 18413 3768 20000 3770
rect 18413 3712 18418 3768
rect 18474 3712 20000 3768
rect 18413 3710 20000 3712
rect 18413 3707 18479 3710
rect 19200 3680 20000 3710
rect 8210 3296 8526 3297
rect 8210 3232 8216 3296
rect 8280 3232 8296 3296
rect 8360 3232 8376 3296
rect 8440 3232 8456 3296
rect 8520 3232 8526 3296
rect 8210 3231 8526 3232
rect 16210 3296 16526 3297
rect 16210 3232 16216 3296
rect 16280 3232 16296 3296
rect 16360 3232 16376 3296
rect 16440 3232 16456 3296
rect 16520 3232 16526 3296
rect 16210 3231 16526 3232
rect 10685 3090 10751 3093
rect 11605 3090 11671 3093
rect 17033 3090 17099 3093
rect 10685 3088 17099 3090
rect 10685 3032 10690 3088
rect 10746 3032 11610 3088
rect 11666 3032 17038 3088
rect 17094 3032 17099 3088
rect 10685 3030 17099 3032
rect 10685 3027 10751 3030
rect 11605 3027 11671 3030
rect 17033 3027 17099 3030
rect 0 2954 800 2984
rect 2773 2954 2839 2957
rect 0 2952 2839 2954
rect 0 2896 2778 2952
rect 2834 2896 2839 2952
rect 0 2894 2839 2896
rect 0 2864 800 2894
rect 2773 2891 2839 2894
rect 4210 2752 4526 2753
rect 4210 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4526 2752
rect 4210 2687 4526 2688
rect 12210 2752 12526 2753
rect 12210 2688 12216 2752
rect 12280 2688 12296 2752
rect 12360 2688 12376 2752
rect 12440 2688 12456 2752
rect 12520 2688 12526 2752
rect 12210 2687 12526 2688
rect 8210 2208 8526 2209
rect 0 2138 800 2168
rect 8210 2144 8216 2208
rect 8280 2144 8296 2208
rect 8360 2144 8376 2208
rect 8440 2144 8456 2208
rect 8520 2144 8526 2208
rect 8210 2143 8526 2144
rect 16210 2208 16526 2209
rect 16210 2144 16216 2208
rect 16280 2144 16296 2208
rect 16360 2144 16376 2208
rect 16440 2144 16456 2208
rect 16520 2144 16526 2208
rect 16210 2143 16526 2144
rect 3049 2138 3115 2141
rect 0 2136 3115 2138
rect 0 2080 3054 2136
rect 3110 2080 3115 2136
rect 0 2078 3115 2080
rect 0 2048 800 2078
rect 3049 2075 3115 2078
rect 4210 1664 4526 1665
rect 4210 1600 4216 1664
rect 4280 1600 4296 1664
rect 4360 1600 4376 1664
rect 4440 1600 4456 1664
rect 4520 1600 4526 1664
rect 4210 1599 4526 1600
rect 12210 1664 12526 1665
rect 12210 1600 12216 1664
rect 12280 1600 12296 1664
rect 12360 1600 12376 1664
rect 12440 1600 12456 1664
rect 12520 1600 12526 1664
rect 12210 1599 12526 1600
rect 0 1322 800 1352
rect 1485 1322 1551 1325
rect 0 1320 1551 1322
rect 0 1264 1490 1320
rect 1546 1264 1551 1320
rect 0 1262 1551 1264
rect 0 1232 800 1262
rect 1485 1259 1551 1262
rect 15561 1322 15627 1325
rect 19200 1322 20000 1352
rect 15561 1320 20000 1322
rect 15561 1264 15566 1320
rect 15622 1264 20000 1320
rect 15561 1262 20000 1264
rect 15561 1259 15627 1262
rect 19200 1232 20000 1262
rect 8210 1120 8526 1121
rect 8210 1056 8216 1120
rect 8280 1056 8296 1120
rect 8360 1056 8376 1120
rect 8440 1056 8456 1120
rect 8520 1056 8526 1120
rect 8210 1055 8526 1056
rect 16210 1120 16526 1121
rect 16210 1056 16216 1120
rect 16280 1056 16296 1120
rect 16360 1056 16376 1120
rect 16440 1056 16456 1120
rect 16520 1056 16526 1120
rect 16210 1055 16526 1056
<< via3 >>
rect 4216 13628 4280 13632
rect 4216 13572 4220 13628
rect 4220 13572 4276 13628
rect 4276 13572 4280 13628
rect 4216 13568 4280 13572
rect 4296 13628 4360 13632
rect 4296 13572 4300 13628
rect 4300 13572 4356 13628
rect 4356 13572 4360 13628
rect 4296 13568 4360 13572
rect 4376 13628 4440 13632
rect 4376 13572 4380 13628
rect 4380 13572 4436 13628
rect 4436 13572 4440 13628
rect 4376 13568 4440 13572
rect 4456 13628 4520 13632
rect 4456 13572 4460 13628
rect 4460 13572 4516 13628
rect 4516 13572 4520 13628
rect 4456 13568 4520 13572
rect 12216 13628 12280 13632
rect 12216 13572 12220 13628
rect 12220 13572 12276 13628
rect 12276 13572 12280 13628
rect 12216 13568 12280 13572
rect 12296 13628 12360 13632
rect 12296 13572 12300 13628
rect 12300 13572 12356 13628
rect 12356 13572 12360 13628
rect 12296 13568 12360 13572
rect 12376 13628 12440 13632
rect 12376 13572 12380 13628
rect 12380 13572 12436 13628
rect 12436 13572 12440 13628
rect 12376 13568 12440 13572
rect 12456 13628 12520 13632
rect 12456 13572 12460 13628
rect 12460 13572 12516 13628
rect 12516 13572 12520 13628
rect 12456 13568 12520 13572
rect 8216 13084 8280 13088
rect 8216 13028 8220 13084
rect 8220 13028 8276 13084
rect 8276 13028 8280 13084
rect 8216 13024 8280 13028
rect 8296 13084 8360 13088
rect 8296 13028 8300 13084
rect 8300 13028 8356 13084
rect 8356 13028 8360 13084
rect 8296 13024 8360 13028
rect 8376 13084 8440 13088
rect 8376 13028 8380 13084
rect 8380 13028 8436 13084
rect 8436 13028 8440 13084
rect 8376 13024 8440 13028
rect 8456 13084 8520 13088
rect 8456 13028 8460 13084
rect 8460 13028 8516 13084
rect 8516 13028 8520 13084
rect 8456 13024 8520 13028
rect 16216 13084 16280 13088
rect 16216 13028 16220 13084
rect 16220 13028 16276 13084
rect 16276 13028 16280 13084
rect 16216 13024 16280 13028
rect 16296 13084 16360 13088
rect 16296 13028 16300 13084
rect 16300 13028 16356 13084
rect 16356 13028 16360 13084
rect 16296 13024 16360 13028
rect 16376 13084 16440 13088
rect 16376 13028 16380 13084
rect 16380 13028 16436 13084
rect 16436 13028 16440 13084
rect 16376 13024 16440 13028
rect 16456 13084 16520 13088
rect 16456 13028 16460 13084
rect 16460 13028 16516 13084
rect 16516 13028 16520 13084
rect 16456 13024 16520 13028
rect 4216 12540 4280 12544
rect 4216 12484 4220 12540
rect 4220 12484 4276 12540
rect 4276 12484 4280 12540
rect 4216 12480 4280 12484
rect 4296 12540 4360 12544
rect 4296 12484 4300 12540
rect 4300 12484 4356 12540
rect 4356 12484 4360 12540
rect 4296 12480 4360 12484
rect 4376 12540 4440 12544
rect 4376 12484 4380 12540
rect 4380 12484 4436 12540
rect 4436 12484 4440 12540
rect 4376 12480 4440 12484
rect 4456 12540 4520 12544
rect 4456 12484 4460 12540
rect 4460 12484 4516 12540
rect 4516 12484 4520 12540
rect 4456 12480 4520 12484
rect 12216 12540 12280 12544
rect 12216 12484 12220 12540
rect 12220 12484 12276 12540
rect 12276 12484 12280 12540
rect 12216 12480 12280 12484
rect 12296 12540 12360 12544
rect 12296 12484 12300 12540
rect 12300 12484 12356 12540
rect 12356 12484 12360 12540
rect 12296 12480 12360 12484
rect 12376 12540 12440 12544
rect 12376 12484 12380 12540
rect 12380 12484 12436 12540
rect 12436 12484 12440 12540
rect 12376 12480 12440 12484
rect 12456 12540 12520 12544
rect 12456 12484 12460 12540
rect 12460 12484 12516 12540
rect 12516 12484 12520 12540
rect 12456 12480 12520 12484
rect 8216 11996 8280 12000
rect 8216 11940 8220 11996
rect 8220 11940 8276 11996
rect 8276 11940 8280 11996
rect 8216 11936 8280 11940
rect 8296 11996 8360 12000
rect 8296 11940 8300 11996
rect 8300 11940 8356 11996
rect 8356 11940 8360 11996
rect 8296 11936 8360 11940
rect 8376 11996 8440 12000
rect 8376 11940 8380 11996
rect 8380 11940 8436 11996
rect 8436 11940 8440 11996
rect 8376 11936 8440 11940
rect 8456 11996 8520 12000
rect 8456 11940 8460 11996
rect 8460 11940 8516 11996
rect 8516 11940 8520 11996
rect 8456 11936 8520 11940
rect 16216 11996 16280 12000
rect 16216 11940 16220 11996
rect 16220 11940 16276 11996
rect 16276 11940 16280 11996
rect 16216 11936 16280 11940
rect 16296 11996 16360 12000
rect 16296 11940 16300 11996
rect 16300 11940 16356 11996
rect 16356 11940 16360 11996
rect 16296 11936 16360 11940
rect 16376 11996 16440 12000
rect 16376 11940 16380 11996
rect 16380 11940 16436 11996
rect 16436 11940 16440 11996
rect 16376 11936 16440 11940
rect 16456 11996 16520 12000
rect 16456 11940 16460 11996
rect 16460 11940 16516 11996
rect 16516 11940 16520 11996
rect 16456 11936 16520 11940
rect 4216 11452 4280 11456
rect 4216 11396 4220 11452
rect 4220 11396 4276 11452
rect 4276 11396 4280 11452
rect 4216 11392 4280 11396
rect 4296 11452 4360 11456
rect 4296 11396 4300 11452
rect 4300 11396 4356 11452
rect 4356 11396 4360 11452
rect 4296 11392 4360 11396
rect 4376 11452 4440 11456
rect 4376 11396 4380 11452
rect 4380 11396 4436 11452
rect 4436 11396 4440 11452
rect 4376 11392 4440 11396
rect 4456 11452 4520 11456
rect 4456 11396 4460 11452
rect 4460 11396 4516 11452
rect 4516 11396 4520 11452
rect 4456 11392 4520 11396
rect 12216 11452 12280 11456
rect 12216 11396 12220 11452
rect 12220 11396 12276 11452
rect 12276 11396 12280 11452
rect 12216 11392 12280 11396
rect 12296 11452 12360 11456
rect 12296 11396 12300 11452
rect 12300 11396 12356 11452
rect 12356 11396 12360 11452
rect 12296 11392 12360 11396
rect 12376 11452 12440 11456
rect 12376 11396 12380 11452
rect 12380 11396 12436 11452
rect 12436 11396 12440 11452
rect 12376 11392 12440 11396
rect 12456 11452 12520 11456
rect 12456 11396 12460 11452
rect 12460 11396 12516 11452
rect 12516 11396 12520 11452
rect 12456 11392 12520 11396
rect 8216 10908 8280 10912
rect 8216 10852 8220 10908
rect 8220 10852 8276 10908
rect 8276 10852 8280 10908
rect 8216 10848 8280 10852
rect 8296 10908 8360 10912
rect 8296 10852 8300 10908
rect 8300 10852 8356 10908
rect 8356 10852 8360 10908
rect 8296 10848 8360 10852
rect 8376 10908 8440 10912
rect 8376 10852 8380 10908
rect 8380 10852 8436 10908
rect 8436 10852 8440 10908
rect 8376 10848 8440 10852
rect 8456 10908 8520 10912
rect 8456 10852 8460 10908
rect 8460 10852 8516 10908
rect 8516 10852 8520 10908
rect 8456 10848 8520 10852
rect 16216 10908 16280 10912
rect 16216 10852 16220 10908
rect 16220 10852 16276 10908
rect 16276 10852 16280 10908
rect 16216 10848 16280 10852
rect 16296 10908 16360 10912
rect 16296 10852 16300 10908
rect 16300 10852 16356 10908
rect 16356 10852 16360 10908
rect 16296 10848 16360 10852
rect 16376 10908 16440 10912
rect 16376 10852 16380 10908
rect 16380 10852 16436 10908
rect 16436 10852 16440 10908
rect 16376 10848 16440 10852
rect 16456 10908 16520 10912
rect 16456 10852 16460 10908
rect 16460 10852 16516 10908
rect 16516 10852 16520 10908
rect 16456 10848 16520 10852
rect 4216 10364 4280 10368
rect 4216 10308 4220 10364
rect 4220 10308 4276 10364
rect 4276 10308 4280 10364
rect 4216 10304 4280 10308
rect 4296 10364 4360 10368
rect 4296 10308 4300 10364
rect 4300 10308 4356 10364
rect 4356 10308 4360 10364
rect 4296 10304 4360 10308
rect 4376 10364 4440 10368
rect 4376 10308 4380 10364
rect 4380 10308 4436 10364
rect 4436 10308 4440 10364
rect 4376 10304 4440 10308
rect 4456 10364 4520 10368
rect 4456 10308 4460 10364
rect 4460 10308 4516 10364
rect 4516 10308 4520 10364
rect 4456 10304 4520 10308
rect 12216 10364 12280 10368
rect 12216 10308 12220 10364
rect 12220 10308 12276 10364
rect 12276 10308 12280 10364
rect 12216 10304 12280 10308
rect 12296 10364 12360 10368
rect 12296 10308 12300 10364
rect 12300 10308 12356 10364
rect 12356 10308 12360 10364
rect 12296 10304 12360 10308
rect 12376 10364 12440 10368
rect 12376 10308 12380 10364
rect 12380 10308 12436 10364
rect 12436 10308 12440 10364
rect 12376 10304 12440 10308
rect 12456 10364 12520 10368
rect 12456 10308 12460 10364
rect 12460 10308 12516 10364
rect 12516 10308 12520 10364
rect 12456 10304 12520 10308
rect 8216 9820 8280 9824
rect 8216 9764 8220 9820
rect 8220 9764 8276 9820
rect 8276 9764 8280 9820
rect 8216 9760 8280 9764
rect 8296 9820 8360 9824
rect 8296 9764 8300 9820
rect 8300 9764 8356 9820
rect 8356 9764 8360 9820
rect 8296 9760 8360 9764
rect 8376 9820 8440 9824
rect 8376 9764 8380 9820
rect 8380 9764 8436 9820
rect 8436 9764 8440 9820
rect 8376 9760 8440 9764
rect 8456 9820 8520 9824
rect 8456 9764 8460 9820
rect 8460 9764 8516 9820
rect 8516 9764 8520 9820
rect 8456 9760 8520 9764
rect 16216 9820 16280 9824
rect 16216 9764 16220 9820
rect 16220 9764 16276 9820
rect 16276 9764 16280 9820
rect 16216 9760 16280 9764
rect 16296 9820 16360 9824
rect 16296 9764 16300 9820
rect 16300 9764 16356 9820
rect 16356 9764 16360 9820
rect 16296 9760 16360 9764
rect 16376 9820 16440 9824
rect 16376 9764 16380 9820
rect 16380 9764 16436 9820
rect 16436 9764 16440 9820
rect 16376 9760 16440 9764
rect 16456 9820 16520 9824
rect 16456 9764 16460 9820
rect 16460 9764 16516 9820
rect 16516 9764 16520 9820
rect 16456 9760 16520 9764
rect 4216 9276 4280 9280
rect 4216 9220 4220 9276
rect 4220 9220 4276 9276
rect 4276 9220 4280 9276
rect 4216 9216 4280 9220
rect 4296 9276 4360 9280
rect 4296 9220 4300 9276
rect 4300 9220 4356 9276
rect 4356 9220 4360 9276
rect 4296 9216 4360 9220
rect 4376 9276 4440 9280
rect 4376 9220 4380 9276
rect 4380 9220 4436 9276
rect 4436 9220 4440 9276
rect 4376 9216 4440 9220
rect 4456 9276 4520 9280
rect 4456 9220 4460 9276
rect 4460 9220 4516 9276
rect 4516 9220 4520 9276
rect 4456 9216 4520 9220
rect 12216 9276 12280 9280
rect 12216 9220 12220 9276
rect 12220 9220 12276 9276
rect 12276 9220 12280 9276
rect 12216 9216 12280 9220
rect 12296 9276 12360 9280
rect 12296 9220 12300 9276
rect 12300 9220 12356 9276
rect 12356 9220 12360 9276
rect 12296 9216 12360 9220
rect 12376 9276 12440 9280
rect 12376 9220 12380 9276
rect 12380 9220 12436 9276
rect 12436 9220 12440 9276
rect 12376 9216 12440 9220
rect 12456 9276 12520 9280
rect 12456 9220 12460 9276
rect 12460 9220 12516 9276
rect 12516 9220 12520 9276
rect 12456 9216 12520 9220
rect 8216 8732 8280 8736
rect 8216 8676 8220 8732
rect 8220 8676 8276 8732
rect 8276 8676 8280 8732
rect 8216 8672 8280 8676
rect 8296 8732 8360 8736
rect 8296 8676 8300 8732
rect 8300 8676 8356 8732
rect 8356 8676 8360 8732
rect 8296 8672 8360 8676
rect 8376 8732 8440 8736
rect 8376 8676 8380 8732
rect 8380 8676 8436 8732
rect 8436 8676 8440 8732
rect 8376 8672 8440 8676
rect 8456 8732 8520 8736
rect 8456 8676 8460 8732
rect 8460 8676 8516 8732
rect 8516 8676 8520 8732
rect 8456 8672 8520 8676
rect 16216 8732 16280 8736
rect 16216 8676 16220 8732
rect 16220 8676 16276 8732
rect 16276 8676 16280 8732
rect 16216 8672 16280 8676
rect 16296 8732 16360 8736
rect 16296 8676 16300 8732
rect 16300 8676 16356 8732
rect 16356 8676 16360 8732
rect 16296 8672 16360 8676
rect 16376 8732 16440 8736
rect 16376 8676 16380 8732
rect 16380 8676 16436 8732
rect 16436 8676 16440 8732
rect 16376 8672 16440 8676
rect 16456 8732 16520 8736
rect 16456 8676 16460 8732
rect 16460 8676 16516 8732
rect 16516 8676 16520 8732
rect 16456 8672 16520 8676
rect 4216 8188 4280 8192
rect 4216 8132 4220 8188
rect 4220 8132 4276 8188
rect 4276 8132 4280 8188
rect 4216 8128 4280 8132
rect 4296 8188 4360 8192
rect 4296 8132 4300 8188
rect 4300 8132 4356 8188
rect 4356 8132 4360 8188
rect 4296 8128 4360 8132
rect 4376 8188 4440 8192
rect 4376 8132 4380 8188
rect 4380 8132 4436 8188
rect 4436 8132 4440 8188
rect 4376 8128 4440 8132
rect 4456 8188 4520 8192
rect 4456 8132 4460 8188
rect 4460 8132 4516 8188
rect 4516 8132 4520 8188
rect 4456 8128 4520 8132
rect 12216 8188 12280 8192
rect 12216 8132 12220 8188
rect 12220 8132 12276 8188
rect 12276 8132 12280 8188
rect 12216 8128 12280 8132
rect 12296 8188 12360 8192
rect 12296 8132 12300 8188
rect 12300 8132 12356 8188
rect 12356 8132 12360 8188
rect 12296 8128 12360 8132
rect 12376 8188 12440 8192
rect 12376 8132 12380 8188
rect 12380 8132 12436 8188
rect 12436 8132 12440 8188
rect 12376 8128 12440 8132
rect 12456 8188 12520 8192
rect 12456 8132 12460 8188
rect 12460 8132 12516 8188
rect 12516 8132 12520 8188
rect 12456 8128 12520 8132
rect 8216 7644 8280 7648
rect 8216 7588 8220 7644
rect 8220 7588 8276 7644
rect 8276 7588 8280 7644
rect 8216 7584 8280 7588
rect 8296 7644 8360 7648
rect 8296 7588 8300 7644
rect 8300 7588 8356 7644
rect 8356 7588 8360 7644
rect 8296 7584 8360 7588
rect 8376 7644 8440 7648
rect 8376 7588 8380 7644
rect 8380 7588 8436 7644
rect 8436 7588 8440 7644
rect 8376 7584 8440 7588
rect 8456 7644 8520 7648
rect 8456 7588 8460 7644
rect 8460 7588 8516 7644
rect 8516 7588 8520 7644
rect 8456 7584 8520 7588
rect 16216 7644 16280 7648
rect 16216 7588 16220 7644
rect 16220 7588 16276 7644
rect 16276 7588 16280 7644
rect 16216 7584 16280 7588
rect 16296 7644 16360 7648
rect 16296 7588 16300 7644
rect 16300 7588 16356 7644
rect 16356 7588 16360 7644
rect 16296 7584 16360 7588
rect 16376 7644 16440 7648
rect 16376 7588 16380 7644
rect 16380 7588 16436 7644
rect 16436 7588 16440 7644
rect 16376 7584 16440 7588
rect 16456 7644 16520 7648
rect 16456 7588 16460 7644
rect 16460 7588 16516 7644
rect 16516 7588 16520 7644
rect 16456 7584 16520 7588
rect 4216 7100 4280 7104
rect 4216 7044 4220 7100
rect 4220 7044 4276 7100
rect 4276 7044 4280 7100
rect 4216 7040 4280 7044
rect 4296 7100 4360 7104
rect 4296 7044 4300 7100
rect 4300 7044 4356 7100
rect 4356 7044 4360 7100
rect 4296 7040 4360 7044
rect 4376 7100 4440 7104
rect 4376 7044 4380 7100
rect 4380 7044 4436 7100
rect 4436 7044 4440 7100
rect 4376 7040 4440 7044
rect 4456 7100 4520 7104
rect 4456 7044 4460 7100
rect 4460 7044 4516 7100
rect 4516 7044 4520 7100
rect 4456 7040 4520 7044
rect 12216 7100 12280 7104
rect 12216 7044 12220 7100
rect 12220 7044 12276 7100
rect 12276 7044 12280 7100
rect 12216 7040 12280 7044
rect 12296 7100 12360 7104
rect 12296 7044 12300 7100
rect 12300 7044 12356 7100
rect 12356 7044 12360 7100
rect 12296 7040 12360 7044
rect 12376 7100 12440 7104
rect 12376 7044 12380 7100
rect 12380 7044 12436 7100
rect 12436 7044 12440 7100
rect 12376 7040 12440 7044
rect 12456 7100 12520 7104
rect 12456 7044 12460 7100
rect 12460 7044 12516 7100
rect 12516 7044 12520 7100
rect 12456 7040 12520 7044
rect 8216 6556 8280 6560
rect 8216 6500 8220 6556
rect 8220 6500 8276 6556
rect 8276 6500 8280 6556
rect 8216 6496 8280 6500
rect 8296 6556 8360 6560
rect 8296 6500 8300 6556
rect 8300 6500 8356 6556
rect 8356 6500 8360 6556
rect 8296 6496 8360 6500
rect 8376 6556 8440 6560
rect 8376 6500 8380 6556
rect 8380 6500 8436 6556
rect 8436 6500 8440 6556
rect 8376 6496 8440 6500
rect 8456 6556 8520 6560
rect 8456 6500 8460 6556
rect 8460 6500 8516 6556
rect 8516 6500 8520 6556
rect 8456 6496 8520 6500
rect 16216 6556 16280 6560
rect 16216 6500 16220 6556
rect 16220 6500 16276 6556
rect 16276 6500 16280 6556
rect 16216 6496 16280 6500
rect 16296 6556 16360 6560
rect 16296 6500 16300 6556
rect 16300 6500 16356 6556
rect 16356 6500 16360 6556
rect 16296 6496 16360 6500
rect 16376 6556 16440 6560
rect 16376 6500 16380 6556
rect 16380 6500 16436 6556
rect 16436 6500 16440 6556
rect 16376 6496 16440 6500
rect 16456 6556 16520 6560
rect 16456 6500 16460 6556
rect 16460 6500 16516 6556
rect 16516 6500 16520 6556
rect 16456 6496 16520 6500
rect 4216 6012 4280 6016
rect 4216 5956 4220 6012
rect 4220 5956 4276 6012
rect 4276 5956 4280 6012
rect 4216 5952 4280 5956
rect 4296 6012 4360 6016
rect 4296 5956 4300 6012
rect 4300 5956 4356 6012
rect 4356 5956 4360 6012
rect 4296 5952 4360 5956
rect 4376 6012 4440 6016
rect 4376 5956 4380 6012
rect 4380 5956 4436 6012
rect 4436 5956 4440 6012
rect 4376 5952 4440 5956
rect 4456 6012 4520 6016
rect 4456 5956 4460 6012
rect 4460 5956 4516 6012
rect 4516 5956 4520 6012
rect 4456 5952 4520 5956
rect 12216 6012 12280 6016
rect 12216 5956 12220 6012
rect 12220 5956 12276 6012
rect 12276 5956 12280 6012
rect 12216 5952 12280 5956
rect 12296 6012 12360 6016
rect 12296 5956 12300 6012
rect 12300 5956 12356 6012
rect 12356 5956 12360 6012
rect 12296 5952 12360 5956
rect 12376 6012 12440 6016
rect 12376 5956 12380 6012
rect 12380 5956 12436 6012
rect 12436 5956 12440 6012
rect 12376 5952 12440 5956
rect 12456 6012 12520 6016
rect 12456 5956 12460 6012
rect 12460 5956 12516 6012
rect 12516 5956 12520 6012
rect 12456 5952 12520 5956
rect 8216 5468 8280 5472
rect 8216 5412 8220 5468
rect 8220 5412 8276 5468
rect 8276 5412 8280 5468
rect 8216 5408 8280 5412
rect 8296 5468 8360 5472
rect 8296 5412 8300 5468
rect 8300 5412 8356 5468
rect 8356 5412 8360 5468
rect 8296 5408 8360 5412
rect 8376 5468 8440 5472
rect 8376 5412 8380 5468
rect 8380 5412 8436 5468
rect 8436 5412 8440 5468
rect 8376 5408 8440 5412
rect 8456 5468 8520 5472
rect 8456 5412 8460 5468
rect 8460 5412 8516 5468
rect 8516 5412 8520 5468
rect 8456 5408 8520 5412
rect 16216 5468 16280 5472
rect 16216 5412 16220 5468
rect 16220 5412 16276 5468
rect 16276 5412 16280 5468
rect 16216 5408 16280 5412
rect 16296 5468 16360 5472
rect 16296 5412 16300 5468
rect 16300 5412 16356 5468
rect 16356 5412 16360 5468
rect 16296 5408 16360 5412
rect 16376 5468 16440 5472
rect 16376 5412 16380 5468
rect 16380 5412 16436 5468
rect 16436 5412 16440 5468
rect 16376 5408 16440 5412
rect 16456 5468 16520 5472
rect 16456 5412 16460 5468
rect 16460 5412 16516 5468
rect 16516 5412 16520 5468
rect 16456 5408 16520 5412
rect 4216 4924 4280 4928
rect 4216 4868 4220 4924
rect 4220 4868 4276 4924
rect 4276 4868 4280 4924
rect 4216 4864 4280 4868
rect 4296 4924 4360 4928
rect 4296 4868 4300 4924
rect 4300 4868 4356 4924
rect 4356 4868 4360 4924
rect 4296 4864 4360 4868
rect 4376 4924 4440 4928
rect 4376 4868 4380 4924
rect 4380 4868 4436 4924
rect 4436 4868 4440 4924
rect 4376 4864 4440 4868
rect 4456 4924 4520 4928
rect 4456 4868 4460 4924
rect 4460 4868 4516 4924
rect 4516 4868 4520 4924
rect 4456 4864 4520 4868
rect 12216 4924 12280 4928
rect 12216 4868 12220 4924
rect 12220 4868 12276 4924
rect 12276 4868 12280 4924
rect 12216 4864 12280 4868
rect 12296 4924 12360 4928
rect 12296 4868 12300 4924
rect 12300 4868 12356 4924
rect 12356 4868 12360 4924
rect 12296 4864 12360 4868
rect 12376 4924 12440 4928
rect 12376 4868 12380 4924
rect 12380 4868 12436 4924
rect 12436 4868 12440 4924
rect 12376 4864 12440 4868
rect 12456 4924 12520 4928
rect 12456 4868 12460 4924
rect 12460 4868 12516 4924
rect 12516 4868 12520 4924
rect 12456 4864 12520 4868
rect 8216 4380 8280 4384
rect 8216 4324 8220 4380
rect 8220 4324 8276 4380
rect 8276 4324 8280 4380
rect 8216 4320 8280 4324
rect 8296 4380 8360 4384
rect 8296 4324 8300 4380
rect 8300 4324 8356 4380
rect 8356 4324 8360 4380
rect 8296 4320 8360 4324
rect 8376 4380 8440 4384
rect 8376 4324 8380 4380
rect 8380 4324 8436 4380
rect 8436 4324 8440 4380
rect 8376 4320 8440 4324
rect 8456 4380 8520 4384
rect 8456 4324 8460 4380
rect 8460 4324 8516 4380
rect 8516 4324 8520 4380
rect 8456 4320 8520 4324
rect 16216 4380 16280 4384
rect 16216 4324 16220 4380
rect 16220 4324 16276 4380
rect 16276 4324 16280 4380
rect 16216 4320 16280 4324
rect 16296 4380 16360 4384
rect 16296 4324 16300 4380
rect 16300 4324 16356 4380
rect 16356 4324 16360 4380
rect 16296 4320 16360 4324
rect 16376 4380 16440 4384
rect 16376 4324 16380 4380
rect 16380 4324 16436 4380
rect 16436 4324 16440 4380
rect 16376 4320 16440 4324
rect 16456 4380 16520 4384
rect 16456 4324 16460 4380
rect 16460 4324 16516 4380
rect 16516 4324 16520 4380
rect 16456 4320 16520 4324
rect 4216 3836 4280 3840
rect 4216 3780 4220 3836
rect 4220 3780 4276 3836
rect 4276 3780 4280 3836
rect 4216 3776 4280 3780
rect 4296 3836 4360 3840
rect 4296 3780 4300 3836
rect 4300 3780 4356 3836
rect 4356 3780 4360 3836
rect 4296 3776 4360 3780
rect 4376 3836 4440 3840
rect 4376 3780 4380 3836
rect 4380 3780 4436 3836
rect 4436 3780 4440 3836
rect 4376 3776 4440 3780
rect 4456 3836 4520 3840
rect 4456 3780 4460 3836
rect 4460 3780 4516 3836
rect 4516 3780 4520 3836
rect 4456 3776 4520 3780
rect 12216 3836 12280 3840
rect 12216 3780 12220 3836
rect 12220 3780 12276 3836
rect 12276 3780 12280 3836
rect 12216 3776 12280 3780
rect 12296 3836 12360 3840
rect 12296 3780 12300 3836
rect 12300 3780 12356 3836
rect 12356 3780 12360 3836
rect 12296 3776 12360 3780
rect 12376 3836 12440 3840
rect 12376 3780 12380 3836
rect 12380 3780 12436 3836
rect 12436 3780 12440 3836
rect 12376 3776 12440 3780
rect 12456 3836 12520 3840
rect 12456 3780 12460 3836
rect 12460 3780 12516 3836
rect 12516 3780 12520 3836
rect 12456 3776 12520 3780
rect 8216 3292 8280 3296
rect 8216 3236 8220 3292
rect 8220 3236 8276 3292
rect 8276 3236 8280 3292
rect 8216 3232 8280 3236
rect 8296 3292 8360 3296
rect 8296 3236 8300 3292
rect 8300 3236 8356 3292
rect 8356 3236 8360 3292
rect 8296 3232 8360 3236
rect 8376 3292 8440 3296
rect 8376 3236 8380 3292
rect 8380 3236 8436 3292
rect 8436 3236 8440 3292
rect 8376 3232 8440 3236
rect 8456 3292 8520 3296
rect 8456 3236 8460 3292
rect 8460 3236 8516 3292
rect 8516 3236 8520 3292
rect 8456 3232 8520 3236
rect 16216 3292 16280 3296
rect 16216 3236 16220 3292
rect 16220 3236 16276 3292
rect 16276 3236 16280 3292
rect 16216 3232 16280 3236
rect 16296 3292 16360 3296
rect 16296 3236 16300 3292
rect 16300 3236 16356 3292
rect 16356 3236 16360 3292
rect 16296 3232 16360 3236
rect 16376 3292 16440 3296
rect 16376 3236 16380 3292
rect 16380 3236 16436 3292
rect 16436 3236 16440 3292
rect 16376 3232 16440 3236
rect 16456 3292 16520 3296
rect 16456 3236 16460 3292
rect 16460 3236 16516 3292
rect 16516 3236 16520 3292
rect 16456 3232 16520 3236
rect 4216 2748 4280 2752
rect 4216 2692 4220 2748
rect 4220 2692 4276 2748
rect 4276 2692 4280 2748
rect 4216 2688 4280 2692
rect 4296 2748 4360 2752
rect 4296 2692 4300 2748
rect 4300 2692 4356 2748
rect 4356 2692 4360 2748
rect 4296 2688 4360 2692
rect 4376 2748 4440 2752
rect 4376 2692 4380 2748
rect 4380 2692 4436 2748
rect 4436 2692 4440 2748
rect 4376 2688 4440 2692
rect 4456 2748 4520 2752
rect 4456 2692 4460 2748
rect 4460 2692 4516 2748
rect 4516 2692 4520 2748
rect 4456 2688 4520 2692
rect 12216 2748 12280 2752
rect 12216 2692 12220 2748
rect 12220 2692 12276 2748
rect 12276 2692 12280 2748
rect 12216 2688 12280 2692
rect 12296 2748 12360 2752
rect 12296 2692 12300 2748
rect 12300 2692 12356 2748
rect 12356 2692 12360 2748
rect 12296 2688 12360 2692
rect 12376 2748 12440 2752
rect 12376 2692 12380 2748
rect 12380 2692 12436 2748
rect 12436 2692 12440 2748
rect 12376 2688 12440 2692
rect 12456 2748 12520 2752
rect 12456 2692 12460 2748
rect 12460 2692 12516 2748
rect 12516 2692 12520 2748
rect 12456 2688 12520 2692
rect 8216 2204 8280 2208
rect 8216 2148 8220 2204
rect 8220 2148 8276 2204
rect 8276 2148 8280 2204
rect 8216 2144 8280 2148
rect 8296 2204 8360 2208
rect 8296 2148 8300 2204
rect 8300 2148 8356 2204
rect 8356 2148 8360 2204
rect 8296 2144 8360 2148
rect 8376 2204 8440 2208
rect 8376 2148 8380 2204
rect 8380 2148 8436 2204
rect 8436 2148 8440 2204
rect 8376 2144 8440 2148
rect 8456 2204 8520 2208
rect 8456 2148 8460 2204
rect 8460 2148 8516 2204
rect 8516 2148 8520 2204
rect 8456 2144 8520 2148
rect 16216 2204 16280 2208
rect 16216 2148 16220 2204
rect 16220 2148 16276 2204
rect 16276 2148 16280 2204
rect 16216 2144 16280 2148
rect 16296 2204 16360 2208
rect 16296 2148 16300 2204
rect 16300 2148 16356 2204
rect 16356 2148 16360 2204
rect 16296 2144 16360 2148
rect 16376 2204 16440 2208
rect 16376 2148 16380 2204
rect 16380 2148 16436 2204
rect 16436 2148 16440 2204
rect 16376 2144 16440 2148
rect 16456 2204 16520 2208
rect 16456 2148 16460 2204
rect 16460 2148 16516 2204
rect 16516 2148 16520 2204
rect 16456 2144 16520 2148
rect 4216 1660 4280 1664
rect 4216 1604 4220 1660
rect 4220 1604 4276 1660
rect 4276 1604 4280 1660
rect 4216 1600 4280 1604
rect 4296 1660 4360 1664
rect 4296 1604 4300 1660
rect 4300 1604 4356 1660
rect 4356 1604 4360 1660
rect 4296 1600 4360 1604
rect 4376 1660 4440 1664
rect 4376 1604 4380 1660
rect 4380 1604 4436 1660
rect 4436 1604 4440 1660
rect 4376 1600 4440 1604
rect 4456 1660 4520 1664
rect 4456 1604 4460 1660
rect 4460 1604 4516 1660
rect 4516 1604 4520 1660
rect 4456 1600 4520 1604
rect 12216 1660 12280 1664
rect 12216 1604 12220 1660
rect 12220 1604 12276 1660
rect 12276 1604 12280 1660
rect 12216 1600 12280 1604
rect 12296 1660 12360 1664
rect 12296 1604 12300 1660
rect 12300 1604 12356 1660
rect 12356 1604 12360 1660
rect 12296 1600 12360 1604
rect 12376 1660 12440 1664
rect 12376 1604 12380 1660
rect 12380 1604 12436 1660
rect 12436 1604 12440 1660
rect 12376 1600 12440 1604
rect 12456 1660 12520 1664
rect 12456 1604 12460 1660
rect 12460 1604 12516 1660
rect 12516 1604 12520 1660
rect 12456 1600 12520 1604
rect 8216 1116 8280 1120
rect 8216 1060 8220 1116
rect 8220 1060 8276 1116
rect 8276 1060 8280 1116
rect 8216 1056 8280 1060
rect 8296 1116 8360 1120
rect 8296 1060 8300 1116
rect 8300 1060 8356 1116
rect 8356 1060 8360 1116
rect 8296 1056 8360 1060
rect 8376 1116 8440 1120
rect 8376 1060 8380 1116
rect 8380 1060 8436 1116
rect 8436 1060 8440 1116
rect 8376 1056 8440 1060
rect 8456 1116 8520 1120
rect 8456 1060 8460 1116
rect 8460 1060 8516 1116
rect 8516 1060 8520 1116
rect 8456 1056 8520 1060
rect 16216 1116 16280 1120
rect 16216 1060 16220 1116
rect 16220 1060 16276 1116
rect 16276 1060 16280 1116
rect 16216 1056 16280 1060
rect 16296 1116 16360 1120
rect 16296 1060 16300 1116
rect 16300 1060 16356 1116
rect 16356 1060 16360 1116
rect 16296 1056 16360 1060
rect 16376 1116 16440 1120
rect 16376 1060 16380 1116
rect 16380 1060 16436 1116
rect 16436 1060 16440 1116
rect 16376 1056 16440 1060
rect 16456 1116 16520 1120
rect 16456 1060 16460 1116
rect 16460 1060 16516 1116
rect 16516 1060 16520 1116
rect 16456 1056 16520 1060
<< metal4 >>
rect 4208 13632 4528 13648
rect 4208 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4528 13632
rect 4208 12544 4528 13568
rect 4208 12480 4216 12544
rect 4280 12488 4296 12544
rect 4360 12488 4376 12544
rect 4440 12488 4456 12544
rect 4520 12480 4528 12544
rect 4208 12252 4250 12480
rect 4486 12252 4528 12480
rect 4208 11456 4528 12252
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 4208 10368 4528 11392
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 4208 9280 4528 10304
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 8192 4528 9216
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 7104 4528 8128
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 6016 4528 7040
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 4928 4528 5952
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 4488 4528 4864
rect 4208 4252 4250 4488
rect 4486 4252 4528 4488
rect 4208 3840 4528 4252
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 2752 4528 3776
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 1664 4528 2688
rect 4208 1600 4216 1664
rect 4280 1600 4296 1664
rect 4360 1600 4376 1664
rect 4440 1600 4456 1664
rect 4520 1600 4528 1664
rect 4208 1040 4528 1600
rect 8208 13088 8528 13648
rect 8208 13024 8216 13088
rect 8280 13024 8296 13088
rect 8360 13024 8376 13088
rect 8440 13024 8456 13088
rect 8520 13024 8528 13088
rect 8208 12000 8528 13024
rect 8208 11936 8216 12000
rect 8280 11936 8296 12000
rect 8360 11936 8376 12000
rect 8440 11936 8456 12000
rect 8520 11936 8528 12000
rect 8208 10912 8528 11936
rect 8208 10848 8216 10912
rect 8280 10848 8296 10912
rect 8360 10848 8376 10912
rect 8440 10848 8456 10912
rect 8520 10848 8528 10912
rect 8208 9824 8528 10848
rect 8208 9760 8216 9824
rect 8280 9760 8296 9824
rect 8360 9760 8376 9824
rect 8440 9760 8456 9824
rect 8520 9760 8528 9824
rect 8208 8736 8528 9760
rect 8208 8672 8216 8736
rect 8280 8672 8296 8736
rect 8360 8672 8376 8736
rect 8440 8672 8456 8736
rect 8520 8672 8528 8736
rect 8208 8488 8528 8672
rect 8208 8252 8250 8488
rect 8486 8252 8528 8488
rect 8208 7648 8528 8252
rect 8208 7584 8216 7648
rect 8280 7584 8296 7648
rect 8360 7584 8376 7648
rect 8440 7584 8456 7648
rect 8520 7584 8528 7648
rect 8208 6560 8528 7584
rect 8208 6496 8216 6560
rect 8280 6496 8296 6560
rect 8360 6496 8376 6560
rect 8440 6496 8456 6560
rect 8520 6496 8528 6560
rect 8208 5472 8528 6496
rect 8208 5408 8216 5472
rect 8280 5408 8296 5472
rect 8360 5408 8376 5472
rect 8440 5408 8456 5472
rect 8520 5408 8528 5472
rect 8208 4384 8528 5408
rect 8208 4320 8216 4384
rect 8280 4320 8296 4384
rect 8360 4320 8376 4384
rect 8440 4320 8456 4384
rect 8520 4320 8528 4384
rect 8208 3296 8528 4320
rect 8208 3232 8216 3296
rect 8280 3232 8296 3296
rect 8360 3232 8376 3296
rect 8440 3232 8456 3296
rect 8520 3232 8528 3296
rect 8208 2208 8528 3232
rect 8208 2144 8216 2208
rect 8280 2144 8296 2208
rect 8360 2144 8376 2208
rect 8440 2144 8456 2208
rect 8520 2144 8528 2208
rect 8208 1120 8528 2144
rect 8208 1056 8216 1120
rect 8280 1056 8296 1120
rect 8360 1056 8376 1120
rect 8440 1056 8456 1120
rect 8520 1056 8528 1120
rect 8208 1040 8528 1056
rect 12208 13632 12528 13648
rect 12208 13568 12216 13632
rect 12280 13568 12296 13632
rect 12360 13568 12376 13632
rect 12440 13568 12456 13632
rect 12520 13568 12528 13632
rect 12208 12544 12528 13568
rect 12208 12480 12216 12544
rect 12280 12488 12296 12544
rect 12360 12488 12376 12544
rect 12440 12488 12456 12544
rect 12520 12480 12528 12544
rect 12208 12252 12250 12480
rect 12486 12252 12528 12480
rect 12208 11456 12528 12252
rect 12208 11392 12216 11456
rect 12280 11392 12296 11456
rect 12360 11392 12376 11456
rect 12440 11392 12456 11456
rect 12520 11392 12528 11456
rect 12208 10368 12528 11392
rect 12208 10304 12216 10368
rect 12280 10304 12296 10368
rect 12360 10304 12376 10368
rect 12440 10304 12456 10368
rect 12520 10304 12528 10368
rect 12208 9280 12528 10304
rect 12208 9216 12216 9280
rect 12280 9216 12296 9280
rect 12360 9216 12376 9280
rect 12440 9216 12456 9280
rect 12520 9216 12528 9280
rect 12208 8192 12528 9216
rect 12208 8128 12216 8192
rect 12280 8128 12296 8192
rect 12360 8128 12376 8192
rect 12440 8128 12456 8192
rect 12520 8128 12528 8192
rect 12208 7104 12528 8128
rect 12208 7040 12216 7104
rect 12280 7040 12296 7104
rect 12360 7040 12376 7104
rect 12440 7040 12456 7104
rect 12520 7040 12528 7104
rect 12208 6016 12528 7040
rect 12208 5952 12216 6016
rect 12280 5952 12296 6016
rect 12360 5952 12376 6016
rect 12440 5952 12456 6016
rect 12520 5952 12528 6016
rect 12208 4928 12528 5952
rect 12208 4864 12216 4928
rect 12280 4864 12296 4928
rect 12360 4864 12376 4928
rect 12440 4864 12456 4928
rect 12520 4864 12528 4928
rect 12208 4488 12528 4864
rect 12208 4252 12250 4488
rect 12486 4252 12528 4488
rect 12208 3840 12528 4252
rect 12208 3776 12216 3840
rect 12280 3776 12296 3840
rect 12360 3776 12376 3840
rect 12440 3776 12456 3840
rect 12520 3776 12528 3840
rect 12208 2752 12528 3776
rect 12208 2688 12216 2752
rect 12280 2688 12296 2752
rect 12360 2688 12376 2752
rect 12440 2688 12456 2752
rect 12520 2688 12528 2752
rect 12208 1664 12528 2688
rect 12208 1600 12216 1664
rect 12280 1600 12296 1664
rect 12360 1600 12376 1664
rect 12440 1600 12456 1664
rect 12520 1600 12528 1664
rect 12208 1040 12528 1600
rect 16208 13088 16528 13648
rect 16208 13024 16216 13088
rect 16280 13024 16296 13088
rect 16360 13024 16376 13088
rect 16440 13024 16456 13088
rect 16520 13024 16528 13088
rect 16208 12000 16528 13024
rect 16208 11936 16216 12000
rect 16280 11936 16296 12000
rect 16360 11936 16376 12000
rect 16440 11936 16456 12000
rect 16520 11936 16528 12000
rect 16208 10912 16528 11936
rect 16208 10848 16216 10912
rect 16280 10848 16296 10912
rect 16360 10848 16376 10912
rect 16440 10848 16456 10912
rect 16520 10848 16528 10912
rect 16208 9824 16528 10848
rect 16208 9760 16216 9824
rect 16280 9760 16296 9824
rect 16360 9760 16376 9824
rect 16440 9760 16456 9824
rect 16520 9760 16528 9824
rect 16208 8736 16528 9760
rect 16208 8672 16216 8736
rect 16280 8672 16296 8736
rect 16360 8672 16376 8736
rect 16440 8672 16456 8736
rect 16520 8672 16528 8736
rect 16208 8488 16528 8672
rect 16208 8252 16250 8488
rect 16486 8252 16528 8488
rect 16208 7648 16528 8252
rect 16208 7584 16216 7648
rect 16280 7584 16296 7648
rect 16360 7584 16376 7648
rect 16440 7584 16456 7648
rect 16520 7584 16528 7648
rect 16208 6560 16528 7584
rect 16208 6496 16216 6560
rect 16280 6496 16296 6560
rect 16360 6496 16376 6560
rect 16440 6496 16456 6560
rect 16520 6496 16528 6560
rect 16208 5472 16528 6496
rect 16208 5408 16216 5472
rect 16280 5408 16296 5472
rect 16360 5408 16376 5472
rect 16440 5408 16456 5472
rect 16520 5408 16528 5472
rect 16208 4384 16528 5408
rect 16208 4320 16216 4384
rect 16280 4320 16296 4384
rect 16360 4320 16376 4384
rect 16440 4320 16456 4384
rect 16520 4320 16528 4384
rect 16208 3296 16528 4320
rect 16208 3232 16216 3296
rect 16280 3232 16296 3296
rect 16360 3232 16376 3296
rect 16440 3232 16456 3296
rect 16520 3232 16528 3296
rect 16208 2208 16528 3232
rect 16208 2144 16216 2208
rect 16280 2144 16296 2208
rect 16360 2144 16376 2208
rect 16440 2144 16456 2208
rect 16520 2144 16528 2208
rect 16208 1120 16528 2144
rect 16208 1056 16216 1120
rect 16280 1056 16296 1120
rect 16360 1056 16376 1120
rect 16440 1056 16456 1120
rect 16520 1056 16528 1120
rect 16208 1040 16528 1056
<< via4 >>
rect 4250 12480 4280 12488
rect 4280 12480 4296 12488
rect 4296 12480 4360 12488
rect 4360 12480 4376 12488
rect 4376 12480 4440 12488
rect 4440 12480 4456 12488
rect 4456 12480 4486 12488
rect 4250 12252 4486 12480
rect 4250 4252 4486 4488
rect 8250 8252 8486 8488
rect 12250 12480 12280 12488
rect 12280 12480 12296 12488
rect 12296 12480 12360 12488
rect 12360 12480 12376 12488
rect 12376 12480 12440 12488
rect 12440 12480 12456 12488
rect 12456 12480 12486 12488
rect 12250 12252 12486 12480
rect 12250 4252 12486 4488
rect 16250 8252 16486 8488
<< metal5 >>
rect 1056 12488 18908 12530
rect 1056 12252 4250 12488
rect 4486 12252 12250 12488
rect 12486 12252 18908 12488
rect 1056 12210 18908 12252
rect 1056 8488 18908 8530
rect 1056 8252 8250 8488
rect 8486 8252 16250 8488
rect 16486 8252 18908 8488
rect 1056 8210 18908 8252
rect 1056 4488 18908 4530
rect 1056 4252 4250 4488
rect 4486 4252 12250 4488
rect 12486 4252 18908 4488
rect 1056 4210 18908 4252
use sky130_fd_sc_hd__diode_2  ANTENNA__243__A $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform -1 0 1932 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__244__A
timestamp 1665323087
transform -1 0 2760 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__252__A
timestamp 1665323087
transform -1 0 4508 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__257__A_N
timestamp 1665323087
transform -1 0 5428 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__258__A
timestamp 1665323087
transform -1 0 6164 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__260__A1
timestamp 1665323087
transform 1 0 1564 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__266__A
timestamp 1665323087
transform 1 0 1564 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__267__A1
timestamp 1665323087
transform 1 0 1472 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__270__A1
timestamp 1665323087
transform 1 0 4048 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__287__B1
timestamp 1665323087
transform -1 0 6624 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__289__A1
timestamp 1665323087
transform -1 0 3588 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__348__A
timestamp 1665323087
transform 1 0 5796 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__349__A
timestamp 1665323087
transform 1 0 7728 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__350__A
timestamp 1665323087
transform -1 0 5704 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__358__A
timestamp 1665323087
transform -1 0 3312 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__360__A2
timestamp 1665323087
transform -1 0 1932 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__361__B
timestamp 1665323087
transform -1 0 13892 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__363__A2
timestamp 1665323087
transform -1 0 14352 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__364__A2
timestamp 1665323087
transform -1 0 5244 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__369__A2
timestamp 1665323087
transform -1 0 3496 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__373__A2
timestamp 1665323087
transform -1 0 2760 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__374__B1
timestamp 1665323087
transform 1 0 8740 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__375__A2
timestamp 1665323087
transform 1 0 3404 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__378__A2
timestamp 1665323087
transform 1 0 3864 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__379__A
timestamp 1665323087
transform 1 0 11132 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__380__A2
timestamp 1665323087
transform 1 0 10948 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__383__A2
timestamp 1665323087
transform -1 0 12144 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__384__A_N
timestamp 1665323087
transform -1 0 3588 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__387__B1
timestamp 1665323087
transform -1 0 6164 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__389__A2
timestamp 1665323087
transform -1 0 6808 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__392__A1
timestamp 1665323087
transform -1 0 6624 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__392__A2
timestamp 1665323087
transform -1 0 7820 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__396__A2
timestamp 1665323087
transform -1 0 12972 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__399__A2
timestamp 1665323087
transform -1 0 18492 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__404__A1
timestamp 1665323087
transform 1 0 15824 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__404__A2
timestamp 1665323087
transform -1 0 13892 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__409__B1
timestamp 1665323087
transform -1 0 16008 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__410__A1
timestamp 1665323087
transform -1 0 18216 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__410__A2
timestamp 1665323087
transform -1 0 6164 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__411__A2
timestamp 1665323087
transform -1 0 10120 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__417__B1
timestamp 1665323087
transform -1 0 9200 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__419__A1
timestamp 1665323087
transform 1 0 16744 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__419__A2
timestamp 1665323087
transform -1 0 10948 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__421__B1
timestamp 1665323087
transform -1 0 12880 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__422__A1
timestamp 1665323087
transform 1 0 15640 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__422__A2
timestamp 1665323087
transform -1 0 18492 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__423__A2
timestamp 1665323087
transform 1 0 18308 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__424__A2
timestamp 1665323087
transform -1 0 16192 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__425__A
timestamp 1665323087
transform 1 0 2852 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__425__B
timestamp 1665323087
transform -1 0 4048 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__427__A
timestamp 1665323087
transform 1 0 16284 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__428__A
timestamp 1665323087
transform -1 0 18492 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__447__A
timestamp 1665323087
transform -1 0 6164 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__470__D
timestamp 1665323087
transform -1 0 14904 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ringosc.dstage\[0\].id.delaybuf0_A
timestamp 1665323087
transform -1 0 4324 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ringosc.ibufp00_A
timestamp 1665323087
transform -1 0 1656 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform 1 0 1380 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform 1 0 3312 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29
timestamp 1665323087
transform 1 0 3772 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_39
timestamp 1665323087
transform 1 0 4692 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43
timestamp 1665323087
transform 1 0 5060 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_49 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform 1 0 5612 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55
timestamp 1665323087
transform 1 0 6164 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57
timestamp 1665323087
transform 1 0 6348 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_60 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform 1 0 6624 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_72 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform 1 0 7728 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_78
timestamp 1665323087
transform 1 0 8280 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_83
timestamp 1665323087
transform 1 0 8740 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_85
timestamp 1665323087
transform 1 0 8924 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_94
timestamp 1665323087
transform 1 0 9752 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_111
timestamp 1665323087
transform 1 0 11316 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_113
timestamp 1665323087
transform 1 0 11500 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_117
timestamp 1665323087
transform 1 0 11868 0 1 1088
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_122 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform 1 0 12328 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_134
timestamp 1665323087
transform 1 0 13432 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_141
timestamp 1665323087
transform 1 0 14076 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_145
timestamp 1665323087
transform 1 0 14444 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_167
timestamp 1665323087
transform 1 0 16468 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_169
timestamp 1665323087
transform 1 0 16652 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_175
timestamp 1665323087
transform 1 0 17204 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_183
timestamp 1665323087
transform 1 0 17940 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_189
timestamp 1665323087
transform 1 0 18492 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_1_3
timestamp 1665323087
transform 1 0 1380 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_11
timestamp 1665323087
transform 1 0 2116 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_20
timestamp 1665323087
transform 1 0 2944 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_45
timestamp 1665323087
transform 1 0 5244 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_49
timestamp 1665323087
transform 1 0 5612 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_55
timestamp 1665323087
transform 1 0 6164 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_57
timestamp 1665323087
transform 1 0 6348 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_61
timestamp 1665323087
transform 1 0 6716 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_76
timestamp 1665323087
transform 1 0 8096 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_1_99
timestamp 1665323087
transform 1 0 10212 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_1_111
timestamp 1665323087
transform 1 0 11316 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_113
timestamp 1665323087
transform 1 0 11500 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_135
timestamp 1665323087
transform 1 0 13524 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_158
timestamp 1665323087
transform 1 0 15640 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_1_165
timestamp 1665323087
transform 1 0 16284 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_169
timestamp 1665323087
transform 1 0 16652 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_186
timestamp 1665323087
transform 1 0 18216 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_3
timestamp 1665323087
transform 1 0 1380 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_9
timestamp 1665323087
transform 1 0 1932 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_20
timestamp 1665323087
transform 1 0 2944 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_2_27
timestamp 1665323087
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_29
timestamp 1665323087
transform 1 0 3772 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_38
timestamp 1665323087
transform 1 0 4600 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_48
timestamp 1665323087
transform 1 0 5520 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_71
timestamp 1665323087
transform 1 0 7636 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_79
timestamp 1665323087
transform 1 0 8372 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_83
timestamp 1665323087
transform 1 0 8740 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_85
timestamp 1665323087
transform 1 0 8924 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_92
timestamp 1665323087
transform 1 0 9568 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_96
timestamp 1665323087
transform 1 0 9936 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_103
timestamp 1665323087
transform 1 0 10580 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_2_112
timestamp 1665323087
transform 1 0 11408 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_139
timestamp 1665323087
transform 1 0 13892 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_141
timestamp 1665323087
transform 1 0 14076 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_146
timestamp 1665323087
transform 1 0 14536 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_150
timestamp 1665323087
transform 1 0 14904 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_173
timestamp 1665323087
transform 1 0 17020 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_177
timestamp 1665323087
transform 1 0 17388 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_2_187
timestamp 1665323087
transform 1 0 18308 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_3
timestamp 1665323087
transform 1 0 1380 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_14
timestamp 1665323087
transform 1 0 2392 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_18
timestamp 1665323087
transform 1 0 2760 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_33
timestamp 1665323087
transform 1 0 4140 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_37
timestamp 1665323087
transform 1 0 4508 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_3_47
timestamp 1665323087
transform 1 0 5428 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_3_55
timestamp 1665323087
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_3_57
timestamp 1665323087
transform 1 0 6348 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_64
timestamp 1665323087
transform 1 0 6992 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_72
timestamp 1665323087
transform 1 0 7728 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_3_95 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform 1 0 9844 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_110
timestamp 1665323087
transform 1 0 11224 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_3_113
timestamp 1665323087
transform 1 0 11500 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_120
timestamp 1665323087
transform 1 0 12144 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_127
timestamp 1665323087
transform 1 0 12788 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_131
timestamp 1665323087
transform 1 0 13156 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_137
timestamp 1665323087
transform 1 0 13708 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_144
timestamp 1665323087
transform 1 0 14352 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_3_167
timestamp 1665323087
transform 1 0 16468 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_3_169
timestamp 1665323087
transform 1 0 16652 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_176
timestamp 1665323087
transform 1 0 17296 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_3_187
timestamp 1665323087
transform 1 0 18308 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_3
timestamp 1665323087
transform 1 0 1380 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_9
timestamp 1665323087
transform 1 0 1932 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_20
timestamp 1665323087
transform 1 0 2944 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_4_25
timestamp 1665323087
transform 1 0 3404 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_4_29
timestamp 1665323087
transform 1 0 3772 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_43
timestamp 1665323087
transform 1 0 5060 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_47
timestamp 1665323087
transform 1 0 5428 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_58
timestamp 1665323087
transform 1 0 6440 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_67
timestamp 1665323087
transform 1 0 7268 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_74
timestamp 1665323087
transform 1 0 7912 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_83
timestamp 1665323087
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_85
timestamp 1665323087
transform 1 0 8924 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_93
timestamp 1665323087
transform 1 0 9660 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_102
timestamp 1665323087
transform 1 0 10488 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_112
timestamp 1665323087
transform 1 0 11408 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_135
timestamp 1665323087
transform 1 0 13524 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_139
timestamp 1665323087
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_141
timestamp 1665323087
transform 1 0 14076 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_147
timestamp 1665323087
transform 1 0 14628 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_151
timestamp 1665323087
transform 1 0 14996 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_4_173
timestamp 1665323087
transform 1 0 17020 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_185
timestamp 1665323087
transform 1 0 18124 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_4_189
timestamp 1665323087
transform 1 0 18492 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_3
timestamp 1665323087
transform 1 0 1380 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_12
timestamp 1665323087
transform 1 0 2208 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_35
timestamp 1665323087
transform 1 0 4324 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_46
timestamp 1665323087
transform 1 0 5336 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_5_53
timestamp 1665323087
transform 1 0 5980 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_5_57
timestamp 1665323087
transform 1 0 6348 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_79
timestamp 1665323087
transform 1 0 8372 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_85
timestamp 1665323087
transform 1 0 8924 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_91
timestamp 1665323087
transform 1 0 9476 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_98
timestamp 1665323087
transform 1 0 10120 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_5_106
timestamp 1665323087
transform 1 0 10856 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_5_113
timestamp 1665323087
transform 1 0 11500 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_120
timestamp 1665323087
transform 1 0 12144 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_127
timestamp 1665323087
transform 1 0 12788 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_134
timestamp 1665323087
transform 1 0 13432 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_138
timestamp 1665323087
transform 1 0 13800 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_144
timestamp 1665323087
transform 1 0 14352 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_5_167
timestamp 1665323087
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_5_169
timestamp 1665323087
transform 1 0 16652 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_174
timestamp 1665323087
transform 1 0 17112 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_181
timestamp 1665323087
transform 1 0 17756 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_188
timestamp 1665323087
transform 1 0 18400 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_6_3
timestamp 1665323087
transform 1 0 1380 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_12
timestamp 1665323087
transform 1 0 2208 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_17
timestamp 1665323087
transform 1 0 2668 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_21
timestamp 1665323087
transform 1 0 3036 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp 1665323087
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_29
timestamp 1665323087
transform 1 0 3772 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_32
timestamp 1665323087
transform 1 0 4048 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_39
timestamp 1665323087
transform 1 0 4692 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_46
timestamp 1665323087
transform 1 0 5336 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_53
timestamp 1665323087
transform 1 0 5980 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_76
timestamp 1665323087
transform 1 0 8096 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_6_83
timestamp 1665323087
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_6_85
timestamp 1665323087
transform 1 0 8924 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_93
timestamp 1665323087
transform 1 0 9660 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_6_100
timestamp 1665323087
transform 1 0 10304 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_108
timestamp 1665323087
transform 1 0 11040 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_130
timestamp 1665323087
transform 1 0 13064 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_139
timestamp 1665323087
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_141
timestamp 1665323087
transform 1 0 14076 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_146
timestamp 1665323087
transform 1 0 14536 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_6_169
timestamp 1665323087
transform 1 0 16652 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_177
timestamp 1665323087
transform 1 0 17388 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_186
timestamp 1665323087
transform 1 0 18216 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_3
timestamp 1665323087
transform 1 0 1380 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_17
timestamp 1665323087
transform 1 0 2668 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_23
timestamp 1665323087
transform 1 0 3220 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_27
timestamp 1665323087
transform 1 0 3588 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_34
timestamp 1665323087
transform 1 0 4232 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_43
timestamp 1665323087
transform 1 0 5060 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_51
timestamp 1665323087
transform 1 0 5796 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_7_55
timestamp 1665323087
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_57
timestamp 1665323087
transform 1 0 6348 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_62
timestamp 1665323087
transform 1 0 6808 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_85
timestamp 1665323087
transform 1 0 8924 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_108
timestamp 1665323087
transform 1 0 11040 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_113
timestamp 1665323087
transform 1 0 11500 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_135
timestamp 1665323087
transform 1 0 13524 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_158
timestamp 1665323087
transform 1 0 15640 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_7_162
timestamp 1665323087
transform 1 0 16008 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_7_167
timestamp 1665323087
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_169
timestamp 1665323087
transform 1 0 16652 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_172
timestamp 1665323087
transform 1 0 16928 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_179
timestamp 1665323087
transform 1 0 17572 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_186
timestamp 1665323087
transform 1 0 18216 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_3
timestamp 1665323087
transform 1 0 1380 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_6
timestamp 1665323087
transform 1 0 1656 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_13
timestamp 1665323087
transform 1 0 2300 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_24
timestamp 1665323087
transform 1 0 3312 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_29
timestamp 1665323087
transform 1 0 3772 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_37
timestamp 1665323087
transform 1 0 4508 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_46
timestamp 1665323087
transform 1 0 5336 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_55
timestamp 1665323087
transform 1 0 6164 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_61
timestamp 1665323087
transform 1 0 6716 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_74
timestamp 1665323087
transform 1 0 7912 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_8_81
timestamp 1665323087
transform 1 0 8556 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_8_85
timestamp 1665323087
transform 1 0 8924 0 1 5440
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_8_98
timestamp 1665323087
transform 1 0 10120 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_114
timestamp 1665323087
transform 1 0 11592 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_126
timestamp 1665323087
transform 1 0 12696 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_130
timestamp 1665323087
transform 1 0 13064 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_135
timestamp 1665323087
transform 1 0 13524 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_139
timestamp 1665323087
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_8_141
timestamp 1665323087
transform 1 0 14076 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_8_147
timestamp 1665323087
transform 1 0 14628 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_171
timestamp 1665323087
transform 1 0 16836 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_180
timestamp 1665323087
transform 1 0 17664 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_185
timestamp 1665323087
transform 1 0 18124 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_8_189
timestamp 1665323087
transform 1 0 18492 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_3
timestamp 1665323087
transform 1 0 1380 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_7
timestamp 1665323087
transform 1 0 1748 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_12
timestamp 1665323087
transform 1 0 2208 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_22
timestamp 1665323087
transform 1 0 3128 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_32
timestamp 1665323087
transform 1 0 4048 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_39
timestamp 1665323087
transform 1 0 4692 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_49
timestamp 1665323087
transform 1 0 5612 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_54
timestamp 1665323087
transform 1 0 6072 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_9_57
timestamp 1665323087
transform 1 0 6348 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_63
timestamp 1665323087
transform 1 0 6900 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_67
timestamp 1665323087
transform 1 0 7268 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_72
timestamp 1665323087
transform 1 0 7728 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_83
timestamp 1665323087
transform 1 0 8740 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_94
timestamp 1665323087
transform 1 0 9752 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_100
timestamp 1665323087
transform 1 0 10304 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_107
timestamp 1665323087
transform 1 0 10948 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_111
timestamp 1665323087
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_9_113
timestamp 1665323087
transform 1 0 11500 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_123
timestamp 1665323087
transform 1 0 12420 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_138
timestamp 1665323087
transform 1 0 13800 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_9_145
timestamp 1665323087
transform 1 0 14444 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_156
timestamp 1665323087
transform 1 0 15456 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_160
timestamp 1665323087
transform 1 0 15824 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_9_167
timestamp 1665323087
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_169
timestamp 1665323087
transform 1 0 16652 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_9_189
timestamp 1665323087
transform 1 0 18492 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_3
timestamp 1665323087
transform 1 0 1380 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_7
timestamp 1665323087
transform 1 0 1748 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_19
timestamp 1665323087
transform 1 0 2852 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_10_27
timestamp 1665323087
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_10_29
timestamp 1665323087
transform 1 0 3772 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_34
timestamp 1665323087
transform 1 0 4232 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_49
timestamp 1665323087
transform 1 0 5612 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_64
timestamp 1665323087
transform 1 0 6992 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_79
timestamp 1665323087
transform 1 0 8372 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_83
timestamp 1665323087
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_85
timestamp 1665323087
transform 1 0 8924 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_99
timestamp 1665323087
transform 1 0 10212 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_110
timestamp 1665323087
transform 1 0 11224 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_125
timestamp 1665323087
transform 1 0 12604 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_136
timestamp 1665323087
transform 1 0 13616 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_141
timestamp 1665323087
transform 1 0 14076 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_155
timestamp 1665323087
transform 1 0 15364 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_10_163
timestamp 1665323087
transform 1 0 16100 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_177
timestamp 1665323087
transform 1 0 17388 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_186
timestamp 1665323087
transform 1 0 18216 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_3
timestamp 1665323087
transform 1 0 1380 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_6
timestamp 1665323087
transform 1 0 1656 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_16
timestamp 1665323087
transform 1 0 2576 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_30
timestamp 1665323087
transform 1 0 3864 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_38
timestamp 1665323087
transform 1 0 4600 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_45
timestamp 1665323087
transform 1 0 5244 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_50
timestamp 1665323087
transform 1 0 5704 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_11_55
timestamp 1665323087
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_11_57
timestamp 1665323087
transform 1 0 6348 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_62
timestamp 1665323087
transform 1 0 6808 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_70
timestamp 1665323087
transform 1 0 7544 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_81
timestamp 1665323087
transform 1 0 8556 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_90
timestamp 1665323087
transform 1 0 9384 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_98
timestamp 1665323087
transform 1 0 10120 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_11_106
timestamp 1665323087
transform 1 0 10856 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_113
timestamp 1665323087
transform 1 0 11500 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_123
timestamp 1665323087
transform 1 0 12420 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_127
timestamp 1665323087
transform 1 0 12788 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_137
timestamp 1665323087
transform 1 0 13708 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_143
timestamp 1665323087
transform 1 0 14260 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_154
timestamp 1665323087
transform 1 0 15272 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_160
timestamp 1665323087
transform 1 0 15824 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_167
timestamp 1665323087
transform 1 0 16468 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_11_169
timestamp 1665323087
transform 1 0 16652 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_181
timestamp 1665323087
transform 1 0 17756 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_186
timestamp 1665323087
transform 1 0 18216 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_3
timestamp 1665323087
transform 1 0 1380 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_24
timestamp 1665323087
transform 1 0 3312 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_29
timestamp 1665323087
transform 1 0 3772 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_35
timestamp 1665323087
transform 1 0 4324 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_44
timestamp 1665323087
transform 1 0 5152 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_49
timestamp 1665323087
transform 1 0 5612 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_53
timestamp 1665323087
transform 1 0 5980 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_68
timestamp 1665323087
transform 1 0 7360 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_12_83
timestamp 1665323087
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_85
timestamp 1665323087
transform 1 0 8924 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_93
timestamp 1665323087
transform 1 0 9660 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_99
timestamp 1665323087
transform 1 0 10212 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_12_107
timestamp 1665323087
transform 1 0 10948 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_118
timestamp 1665323087
transform 1 0 11960 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_133
timestamp 1665323087
transform 1 0 13340 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_139
timestamp 1665323087
transform 1 0 13892 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_141
timestamp 1665323087
transform 1 0 14076 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_144
timestamp 1665323087
transform 1 0 14352 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_12_159
timestamp 1665323087
transform 1 0 15732 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_169
timestamp 1665323087
transform 1 0 16652 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_12_189
timestamp 1665323087
transform 1 0 18492 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_3
timestamp 1665323087
transform 1 0 1380 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_13_9
timestamp 1665323087
transform 1 0 1932 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_15
timestamp 1665323087
transform 1 0 2484 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_34
timestamp 1665323087
transform 1 0 4232 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_13_47
timestamp 1665323087
transform 1 0 5428 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_13_55
timestamp 1665323087
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_57
timestamp 1665323087
transform 1 0 6348 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_13_62
timestamp 1665323087
transform 1 0 6808 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_70
timestamp 1665323087
transform 1 0 7544 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_74
timestamp 1665323087
transform 1 0 7912 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_81
timestamp 1665323087
transform 1 0 8556 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_90
timestamp 1665323087
transform 1 0 9384 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_13_102
timestamp 1665323087
transform 1 0 10488 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_107
timestamp 1665323087
transform 1 0 10948 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_13_111
timestamp 1665323087
transform 1 0 11316 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_113
timestamp 1665323087
transform 1 0 11500 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_118
timestamp 1665323087
transform 1 0 11960 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_13_123
timestamp 1665323087
transform 1 0 12420 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_128
timestamp 1665323087
transform 1 0 12880 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_138
timestamp 1665323087
transform 1 0 13800 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_145
timestamp 1665323087
transform 1 0 14444 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_151
timestamp 1665323087
transform 1 0 14996 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_161
timestamp 1665323087
transform 1 0 15916 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_166
timestamp 1665323087
transform 1 0 16376 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_13_169
timestamp 1665323087
transform 1 0 16652 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_177
timestamp 1665323087
transform 1 0 17388 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_185
timestamp 1665323087
transform 1 0 18124 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_13_189
timestamp 1665323087
transform 1 0 18492 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_3
timestamp 1665323087
transform 1 0 1380 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_14_17
timestamp 1665323087
transform 1 0 2668 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_27
timestamp 1665323087
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_29
timestamp 1665323087
transform 1 0 3772 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_38
timestamp 1665323087
transform 1 0 4600 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_44
timestamp 1665323087
transform 1 0 5152 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_48
timestamp 1665323087
transform 1 0 5520 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_14_56
timestamp 1665323087
transform 1 0 6256 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_63
timestamp 1665323087
transform 1 0 6900 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_70
timestamp 1665323087
transform 1 0 7544 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_14_77
timestamp 1665323087
transform 1 0 8188 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_14_83
timestamp 1665323087
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_85
timestamp 1665323087
transform 1 0 8924 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_89
timestamp 1665323087
transform 1 0 9292 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_97
timestamp 1665323087
transform 1 0 10028 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_109
timestamp 1665323087
transform 1 0 11132 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_113
timestamp 1665323087
transform 1 0 11500 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_117
timestamp 1665323087
transform 1 0 11868 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_124
timestamp 1665323087
transform 1 0 12512 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_128
timestamp 1665323087
transform 1 0 12880 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_14_137
timestamp 1665323087
transform 1 0 13708 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_14_141
timestamp 1665323087
transform 1 0 14076 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_150
timestamp 1665323087
transform 1 0 14904 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_160
timestamp 1665323087
transform 1 0 15824 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_164
timestamp 1665323087
transform 1 0 16192 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_168
timestamp 1665323087
transform 1 0 16560 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_14_187
timestamp 1665323087
transform 1 0 18308 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_15_3
timestamp 1665323087
transform 1 0 1380 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_15_13
timestamp 1665323087
transform 1 0 2300 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_17
timestamp 1665323087
transform 1 0 2668 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_36
timestamp 1665323087
transform 1 0 4416 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_40
timestamp 1665323087
transform 1 0 4784 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_44
timestamp 1665323087
transform 1 0 5152 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_55
timestamp 1665323087
transform 1 0 6164 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_15_57
timestamp 1665323087
transform 1 0 6348 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_62
timestamp 1665323087
transform 1 0 6808 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_72
timestamp 1665323087
transform 1 0 7728 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_81
timestamp 1665323087
transform 1 0 8556 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_85
timestamp 1665323087
transform 1 0 8924 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_92
timestamp 1665323087
transform 1 0 9568 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_15_102
timestamp 1665323087
transform 1 0 10488 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_15_111
timestamp 1665323087
transform 1 0 11316 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_15_113
timestamp 1665323087
transform 1 0 11500 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_119
timestamp 1665323087
transform 1 0 12052 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_127
timestamp 1665323087
transform 1 0 12788 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_134
timestamp 1665323087
transform 1 0 13432 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_15_139
timestamp 1665323087
transform 1 0 13892 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_151
timestamp 1665323087
transform 1 0 14996 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_15_161
timestamp 1665323087
transform 1 0 15916 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_15_167
timestamp 1665323087
transform 1 0 16468 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_15_169
timestamp 1665323087
transform 1 0 16652 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_177
timestamp 1665323087
transform 1 0 17388 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_186
timestamp 1665323087
transform 1 0 18216 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_3
timestamp 1665323087
transform 1 0 1380 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_9
timestamp 1665323087
transform 1 0 1932 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_18
timestamp 1665323087
transform 1 0 2760 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_16_27
timestamp 1665323087
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_29
timestamp 1665323087
transform 1 0 3772 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_41
timestamp 1665323087
transform 1 0 4876 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_46
timestamp 1665323087
transform 1 0 5336 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_52
timestamp 1665323087
transform 1 0 5888 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_59
timestamp 1665323087
transform 1 0 6532 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_68
timestamp 1665323087
transform 1 0 7360 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_72
timestamp 1665323087
transform 1 0 7728 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_16_81
timestamp 1665323087
transform 1 0 8556 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_16_85
timestamp 1665323087
transform 1 0 8924 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_91
timestamp 1665323087
transform 1 0 9476 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_100
timestamp 1665323087
transform 1 0 10304 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_107
timestamp 1665323087
transform 1 0 10948 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_114
timestamp 1665323087
transform 1 0 11592 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_122
timestamp 1665323087
transform 1 0 12328 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_16_127
timestamp 1665323087
transform 1 0 12788 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_135
timestamp 1665323087
transform 1 0 13524 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_16_139
timestamp 1665323087
transform 1 0 13892 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_141
timestamp 1665323087
transform 1 0 14076 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_150
timestamp 1665323087
transform 1 0 14904 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_160
timestamp 1665323087
transform 1 0 15824 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_166
timestamp 1665323087
transform 1 0 16376 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_181
timestamp 1665323087
transform 1 0 17756 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_16_187
timestamp 1665323087
transform 1 0 18308 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_17_3
timestamp 1665323087
transform 1 0 1380 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_14
timestamp 1665323087
transform 1 0 2392 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_18
timestamp 1665323087
transform 1 0 2760 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_24
timestamp 1665323087
transform 1 0 3312 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_29
timestamp 1665323087
transform 1 0 3772 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_38
timestamp 1665323087
transform 1 0 4600 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_44
timestamp 1665323087
transform 1 0 5152 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_55
timestamp 1665323087
transform 1 0 6164 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_17_57
timestamp 1665323087
transform 1 0 6348 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_62
timestamp 1665323087
transform 1 0 6808 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_71
timestamp 1665323087
transform 1 0 7636 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_17_82
timestamp 1665323087
transform 1 0 8648 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_90
timestamp 1665323087
transform 1 0 9384 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_17_99
timestamp 1665323087
transform 1 0 10212 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_110
timestamp 1665323087
transform 1 0 11224 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_113
timestamp 1665323087
transform 1 0 11500 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_122
timestamp 1665323087
transform 1 0 12328 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_129
timestamp 1665323087
transform 1 0 12972 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_138
timestamp 1665323087
transform 1 0 13800 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_142
timestamp 1665323087
transform 1 0 14168 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_17_149
timestamp 1665323087
transform 1 0 14812 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_17_161
timestamp 1665323087
transform 1 0 15916 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_17_167
timestamp 1665323087
transform 1 0 16468 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_17_169
timestamp 1665323087
transform 1 0 16652 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_179
timestamp 1665323087
transform 1 0 17572 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_188
timestamp 1665323087
transform 1 0 18400 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_18_3
timestamp 1665323087
transform 1 0 1380 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_22
timestamp 1665323087
transform 1 0 3128 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_26
timestamp 1665323087
transform 1 0 3496 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_18_29
timestamp 1665323087
transform 1 0 3772 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_48
timestamp 1665323087
transform 1 0 5520 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_61
timestamp 1665323087
transform 1 0 6716 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_18_72
timestamp 1665323087
transform 1 0 7728 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_18_83
timestamp 1665323087
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_18_85
timestamp 1665323087
transform 1 0 8924 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_94
timestamp 1665323087
transform 1 0 9752 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_98
timestamp 1665323087
transform 1 0 10120 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_105
timestamp 1665323087
transform 1 0 10764 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_115
timestamp 1665323087
transform 1 0 11684 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_125
timestamp 1665323087
transform 1 0 12604 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_129
timestamp 1665323087
transform 1 0 12972 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_18_139
timestamp 1665323087
transform 1 0 13892 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_18_141
timestamp 1665323087
transform 1 0 14076 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_151
timestamp 1665323087
transform 1 0 14996 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_18_158
timestamp 1665323087
transform 1 0 15640 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_172
timestamp 1665323087
transform 1 0 16928 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_181
timestamp 1665323087
transform 1 0 17756 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_186
timestamp 1665323087
transform 1 0 18216 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_3
timestamp 1665323087
transform 1 0 1380 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_14
timestamp 1665323087
transform 1 0 2392 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_18
timestamp 1665323087
transform 1 0 2760 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_23
timestamp 1665323087
transform 1 0 3220 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_32
timestamp 1665323087
transform 1 0 4048 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_41
timestamp 1665323087
transform 1 0 4876 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_46
timestamp 1665323087
transform 1 0 5336 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_19_55
timestamp 1665323087
transform 1 0 6164 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_19_57
timestamp 1665323087
transform 1 0 6348 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_60
timestamp 1665323087
transform 1 0 6624 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_69
timestamp 1665323087
transform 1 0 7452 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_73
timestamp 1665323087
transform 1 0 7820 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_82
timestamp 1665323087
transform 1 0 8648 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_88
timestamp 1665323087
transform 1 0 9200 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_100
timestamp 1665323087
transform 1 0 10304 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_108
timestamp 1665323087
transform 1 0 11040 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_113
timestamp 1665323087
transform 1 0 11500 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_122
timestamp 1665323087
transform 1 0 12328 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_19_127
timestamp 1665323087
transform 1 0 12788 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_136
timestamp 1665323087
transform 1 0 13616 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_145
timestamp 1665323087
transform 1 0 14444 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_158
timestamp 1665323087
transform 1 0 15640 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_162
timestamp 1665323087
transform 1 0 16008 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_19_167
timestamp 1665323087
transform 1 0 16468 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_169
timestamp 1665323087
transform 1 0 16652 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_19_189
timestamp 1665323087
transform 1 0 18492 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_3
timestamp 1665323087
transform 1 0 1380 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_14
timestamp 1665323087
transform 1 0 2392 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_18
timestamp 1665323087
transform 1 0 2760 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_23
timestamp 1665323087
transform 1 0 3220 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_20_27
timestamp 1665323087
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_20_29
timestamp 1665323087
transform 1 0 3772 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_20_37
timestamp 1665323087
transform 1 0 4508 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_20_47
timestamp 1665323087
transform 1 0 5428 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_54
timestamp 1665323087
transform 1 0 6072 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_74
timestamp 1665323087
transform 1 0 7912 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_20_83
timestamp 1665323087
transform 1 0 8740 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_20_85
timestamp 1665323087
transform 1 0 8924 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_20_95
timestamp 1665323087
transform 1 0 9844 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_106
timestamp 1665323087
transform 1 0 10856 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_116
timestamp 1665323087
transform 1 0 11776 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_20_120
timestamp 1665323087
transform 1 0 12144 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_131
timestamp 1665323087
transform 1 0 13156 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_138
timestamp 1665323087
transform 1 0 13800 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_20_141
timestamp 1665323087
transform 1 0 14076 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_20_160
timestamp 1665323087
transform 1 0 15824 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_167
timestamp 1665323087
transform 1 0 16468 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_176
timestamp 1665323087
transform 1 0 17296 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_185
timestamp 1665323087
transform 1 0 18124 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_20_189
timestamp 1665323087
transform 1 0 18492 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_21_3
timestamp 1665323087
transform 1 0 1380 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_21_17
timestamp 1665323087
transform 1 0 2668 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_38
timestamp 1665323087
transform 1 0 4600 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_51
timestamp 1665323087
transform 1 0 5796 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_21_55
timestamp 1665323087
transform 1 0 6164 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_21_57
timestamp 1665323087
transform 1 0 6348 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_67
timestamp 1665323087
transform 1 0 7268 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_87
timestamp 1665323087
transform 1 0 9108 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_100
timestamp 1665323087
transform 1 0 10304 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_111
timestamp 1665323087
transform 1 0 11316 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_21_113
timestamp 1665323087
transform 1 0 11500 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_125
timestamp 1665323087
transform 1 0 12604 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_129
timestamp 1665323087
transform 1 0 12972 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_141
timestamp 1665323087
transform 1 0 14076 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_147
timestamp 1665323087
transform 1 0 14628 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_21_167
timestamp 1665323087
transform 1 0 16468 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_169
timestamp 1665323087
transform 1 0 16652 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_184
timestamp 1665323087
transform 1 0 18032 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_21_189
timestamp 1665323087
transform 1 0 18492 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_3
timestamp 1665323087
transform 1 0 1380 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_11
timestamp 1665323087
transform 1 0 2116 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_15
timestamp 1665323087
transform 1 0 2484 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_20
timestamp 1665323087
transform 1 0 2944 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_27
timestamp 1665323087
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_22_29
timestamp 1665323087
transform 1 0 3772 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_32
timestamp 1665323087
transform 1 0 4048 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_41
timestamp 1665323087
transform 1 0 4876 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_45
timestamp 1665323087
transform 1 0 5244 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_51
timestamp 1665323087
transform 1 0 5796 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_22_55
timestamp 1665323087
transform 1 0 6164 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_22_57
timestamp 1665323087
transform 1 0 6348 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_65
timestamp 1665323087
transform 1 0 7084 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_71
timestamp 1665323087
transform 1 0 7636 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_76
timestamp 1665323087
transform 1 0 8096 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_83
timestamp 1665323087
transform 1 0 8740 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_85
timestamp 1665323087
transform 1 0 8924 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_94
timestamp 1665323087
transform 1 0 9752 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_22_99
timestamp 1665323087
transform 1 0 10212 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_22_105
timestamp 1665323087
transform 1 0 10764 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_22_109
timestamp 1665323087
transform 1 0 11132 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_22_113
timestamp 1665323087
transform 1 0 11500 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_22_117
timestamp 1665323087
transform 1 0 11868 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_22_127
timestamp 1665323087
transform 1 0 12788 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_131
timestamp 1665323087
transform 1 0 13156 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_22_139
timestamp 1665323087
transform 1 0 13892 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_22_141
timestamp 1665323087
transform 1 0 14076 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_149
timestamp 1665323087
transform 1 0 14812 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_22_154
timestamp 1665323087
transform 1 0 15272 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_22_161
timestamp 1665323087
transform 1 0 15916 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_166
timestamp 1665323087
transform 1 0 16376 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_22_169
timestamp 1665323087
transform 1 0 16652 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_177
timestamp 1665323087
transform 1 0 17388 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_182
timestamp 1665323087
transform 1 0 17848 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_186
timestamp 1665323087
transform 1 0 18216 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1665323087
transform 1 0 1104 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1665323087
transform -1 0 18860 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1665323087
transform 1 0 1104 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1665323087
transform -1 0 18860 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1665323087
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1665323087
transform -1 0 18860 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1665323087
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1665323087
transform -1 0 18860 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1665323087
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1665323087
transform -1 0 18860 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1665323087
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1665323087
transform -1 0 18860 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1665323087
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1665323087
transform -1 0 18860 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1665323087
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1665323087
transform -1 0 18860 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1665323087
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1665323087
transform -1 0 18860 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1665323087
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1665323087
transform -1 0 18860 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1665323087
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1665323087
transform -1 0 18860 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1665323087
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1665323087
transform -1 0 18860 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1665323087
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1665323087
transform -1 0 18860 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1665323087
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1665323087
transform -1 0 18860 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1665323087
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1665323087
transform -1 0 18860 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1665323087
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1665323087
transform -1 0 18860 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1665323087
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1665323087
transform -1 0 18860 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1665323087
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1665323087
transform -1 0 18860 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1665323087
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1665323087
transform -1 0 18860 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1665323087
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1665323087
transform -1 0 18860 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1665323087
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1665323087
transform -1 0 18860 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1665323087
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1665323087
transform -1 0 18860 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1665323087
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1665323087
transform -1 0 18860 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_46 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform 1 0 3680 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_47
timestamp 1665323087
transform 1 0 6256 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_48
timestamp 1665323087
transform 1 0 8832 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_49
timestamp 1665323087
transform 1 0 11408 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_50
timestamp 1665323087
transform 1 0 13984 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_51
timestamp 1665323087
transform 1 0 16560 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_52
timestamp 1665323087
transform 1 0 6256 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_53
timestamp 1665323087
transform 1 0 11408 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_54
timestamp 1665323087
transform 1 0 16560 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_55
timestamp 1665323087
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_56
timestamp 1665323087
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_57
timestamp 1665323087
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_58
timestamp 1665323087
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_59
timestamp 1665323087
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_60
timestamp 1665323087
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_61
timestamp 1665323087
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_62
timestamp 1665323087
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_63
timestamp 1665323087
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_64
timestamp 1665323087
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_65
timestamp 1665323087
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_66
timestamp 1665323087
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_67
timestamp 1665323087
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_68
timestamp 1665323087
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_69
timestamp 1665323087
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_70
timestamp 1665323087
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_71
timestamp 1665323087
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_72
timestamp 1665323087
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_73
timestamp 1665323087
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_74
timestamp 1665323087
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_75
timestamp 1665323087
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_76
timestamp 1665323087
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_77
timestamp 1665323087
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_78
timestamp 1665323087
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_79
timestamp 1665323087
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_80
timestamp 1665323087
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_81
timestamp 1665323087
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_82
timestamp 1665323087
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_83
timestamp 1665323087
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_84
timestamp 1665323087
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_85
timestamp 1665323087
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_86
timestamp 1665323087
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_87
timestamp 1665323087
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_88
timestamp 1665323087
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_89
timestamp 1665323087
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_90
timestamp 1665323087
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_91
timestamp 1665323087
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_92
timestamp 1665323087
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_93
timestamp 1665323087
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_94
timestamp 1665323087
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_95
timestamp 1665323087
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_96
timestamp 1665323087
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_97
timestamp 1665323087
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_98
timestamp 1665323087
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_99
timestamp 1665323087
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_100
timestamp 1665323087
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_101
timestamp 1665323087
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_102
timestamp 1665323087
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_103
timestamp 1665323087
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_104
timestamp 1665323087
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_105
timestamp 1665323087
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_106
timestamp 1665323087
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_107
timestamp 1665323087
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_108
timestamp 1665323087
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_109
timestamp 1665323087
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_110
timestamp 1665323087
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_111
timestamp 1665323087
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_112
timestamp 1665323087
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_113
timestamp 1665323087
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_114
timestamp 1665323087
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_115
timestamp 1665323087
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_116
timestamp 1665323087
transform 1 0 6256 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_117
timestamp 1665323087
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_118
timestamp 1665323087
transform 1 0 11408 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_119
timestamp 1665323087
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_120
timestamp 1665323087
transform 1 0 16560 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__xnor2_2  _214_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform 1 0 17020 0 -1 2176
box -38 -48 1234 592
use sky130_fd_sc_hd__buf_2  _215_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform 1 0 18124 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _216_
timestamp 1665323087
transform -1 0 17112 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_2  _217_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform 1 0 7084 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _218_
timestamp 1665323087
transform -1 0 6808 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_2  _219_
timestamp 1665323087
transform 1 0 4508 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _220_
timestamp 1665323087
transform -1 0 3588 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_2  _221_
timestamp 1665323087
transform -1 0 6440 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _222_
timestamp 1665323087
transform 1 0 6348 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_2  _223_
timestamp 1665323087
transform 1 0 6900 0 1 1088
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _224_
timestamp 1665323087
transform -1 0 6164 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _225_
timestamp 1665323087
transform 1 0 8372 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_2  _226_
timestamp 1665323087
transform 1 0 3864 0 1 1088
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _227_
timestamp 1665323087
transform -1 0 1932 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _228_
timestamp 1665323087
transform -1 0 15824 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _229_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform -1 0 11868 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _230_
timestamp 1665323087
transform 1 0 6440 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__nand2b_2  _231_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform -1 0 7268 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__and2_2  _232_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform -1 0 5520 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_2  _233_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform -1 0 8096 0 -1 2176
box -38 -48 1234 592
use sky130_fd_sc_hd__and2_2  _234_
timestamp 1665323087
transform -1 0 6992 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__and2_2  _235_
timestamp 1665323087
transform -1 0 8372 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__a211o_2  _236_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform 1 0 4692 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_2  _237_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform -1 0 4232 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _238_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform 1 0 4876 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_2  _239_
timestamp 1665323087
transform -1 0 6164 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__and3_2  _240_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform -1 0 4508 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_2  _241_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform -1 0 5060 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_2  _242_
timestamp 1665323087
transform 1 0 4232 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _243_
timestamp 1665323087
transform 1 0 1932 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _244_
timestamp 1665323087
transform -1 0 2668 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_2  _245_
timestamp 1665323087
transform 1 0 3956 0 1 2176
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_2  _246_
timestamp 1665323087
transform -1 0 6164 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _247_
timestamp 1665323087
transform -1 0 5980 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_2  _248_
timestamp 1665323087
transform -1 0 5060 0 1 3264
box -38 -48 1234 592
use sky130_fd_sc_hd__o32a_2  _249_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform -1 0 3312 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_2  _250_
timestamp 1665323087
transform -1 0 2300 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_2  _251_
timestamp 1665323087
transform -1 0 4140 0 -1 3264
box -38 -48 1234 592
use sky130_fd_sc_hd__inv_2  _252_
timestamp 1665323087
transform 1 0 1656 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__nand2b_2  _253_
timestamp 1665323087
transform -1 0 2392 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_2  _254_
timestamp 1665323087
transform -1 0 2116 0 -1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _255_
timestamp 1665323087
transform -1 0 3588 0 1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _256_
timestamp 1665323087
transform -1 0 3404 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__nand3b_2  _257_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform -1 0 2944 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__and2_2  _258_
timestamp 1665323087
transform 1 0 1656 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_2  _259_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform 1 0 1564 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__o2111a_2  _260_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform -1 0 2852 0 1 6528
box -38 -48 958 592
use sky130_fd_sc_hd__xor2_2  _261_
timestamp 1665323087
transform -1 0 6992 0 1 6528
box -38 -48 1234 592
use sky130_fd_sc_hd__inv_2  _262_
timestamp 1665323087
transform 1 0 5796 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__and2_2  _263_
timestamp 1665323087
transform -1 0 5796 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_2  _264_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform 1 0 4692 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_2  _265_
timestamp 1665323087
transform -1 0 5612 0 1 6528
box -38 -48 1234 592
use sky130_fd_sc_hd__and2_2  _266_
timestamp 1665323087
transform -1 0 3588 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_2  _267_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform -1 0 2576 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_2  _268_
timestamp 1665323087
transform 1 0 4784 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _269_
timestamp 1665323087
transform -1 0 6900 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_2  _270_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform -1 0 5612 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__o31a_2  _271_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform -1 0 3128 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _272_
timestamp 1665323087
transform 1 0 7176 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _273_
timestamp 1665323087
transform 1 0 9844 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__and2_2  _274_
timestamp 1665323087
transform 1 0 9568 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _275_
timestamp 1665323087
transform -1 0 16376 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _276_
timestamp 1665323087
transform 1 0 13616 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _277_
timestamp 1665323087
transform -1 0 7544 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__nand4_2  _278_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform 1 0 9568 0 -1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__nand2_2  _279_
timestamp 1665323087
transform 1 0 7084 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _280_
timestamp 1665323087
transform -1 0 12788 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _281_
timestamp 1665323087
transform -1 0 12512 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _282_
timestamp 1665323087
transform -1 0 12052 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _283_
timestamp 1665323087
transform 1 0 7728 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _284_
timestamp 1665323087
transform 1 0 9660 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__and3_2  _285_
timestamp 1665323087
transform 1 0 10396 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__and4b_2  _286_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform -1 0 18308 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__o21ai_2  _287_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform -1 0 2944 0 -1 2176
box -38 -48 682 592
use sky130_fd_sc_hd__and4b_2  _288_
timestamp 1665323087
transform 1 0 2116 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__o211a_2  _289_
timestamp 1665323087
transform 1 0 3312 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__nand4b_2  _290_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform 1 0 2760 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__and3b_2  _291_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform 1 0 11224 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__o31a_2  _292_
timestamp 1665323087
transform -1 0 13708 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _293_
timestamp 1665323087
transform 1 0 13892 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_2  _294_
timestamp 1665323087
transform -1 0 13340 0 1 7616
box -38 -48 1234 592
use sky130_fd_sc_hd__nor2_2  _295_
timestamp 1665323087
transform 1 0 8924 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__and2_2  _296_
timestamp 1665323087
transform 1 0 10304 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_2  _297_
timestamp 1665323087
transform 1 0 10488 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _298_
timestamp 1665323087
transform -1 0 6900 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _299_
timestamp 1665323087
transform -1 0 14996 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_2  _300_
timestamp 1665323087
transform -1 0 12972 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _301_
timestamp 1665323087
transform -1 0 8556 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_2  _302_
timestamp 1665323087
transform 1 0 6164 0 1 7616
box -38 -48 1234 592
use sky130_fd_sc_hd__inv_2  _303_
timestamp 1665323087
transform 1 0 8464 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_2  _304_
timestamp 1665323087
transform -1 0 9660 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__a32o_2  _305_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform -1 0 8556 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _306_
timestamp 1665323087
transform -1 0 12420 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_2  _307_
timestamp 1665323087
transform -1 0 12420 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__xnor2_2  _308_
timestamp 1665323087
transform 1 0 14168 0 1 6528
box -38 -48 1234 592
use sky130_fd_sc_hd__and2_2  _309_
timestamp 1665323087
transform 1 0 15548 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_2  _310_
timestamp 1665323087
transform -1 0 15272 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_2  _311_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform -1 0 15456 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_2  _312_
timestamp 1665323087
transform -1 0 11224 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_2  _313_
timestamp 1665323087
transform 1 0 11408 0 1 6528
box -38 -48 1234 592
use sky130_fd_sc_hd__mux2_2  _314_
timestamp 1665323087
transform 1 0 11592 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _315_
timestamp 1665323087
transform -1 0 11592 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__xor2_2  _316_
timestamp 1665323087
transform -1 0 10212 0 1 6528
box -38 -48 1234 592
use sky130_fd_sc_hd__mux2_2  _317_
timestamp 1665323087
transform -1 0 9752 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _318_
timestamp 1665323087
transform 1 0 9936 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_2  _319_
timestamp 1665323087
transform -1 0 13708 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__o211a_2  _320_
timestamp 1665323087
transform -1 0 13800 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_2  _321_
timestamp 1665323087
transform 1 0 14536 0 1 7616
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_2  _322_
timestamp 1665323087
transform 1 0 7544 0 1 7616
box -38 -48 1234 592
use sky130_fd_sc_hd__o2bb2a_2  _323_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform 1 0 12788 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_2  _324_
timestamp 1665323087
transform -1 0 8556 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_2  _325_
timestamp 1665323087
transform 1 0 7176 0 1 6528
box -38 -48 1234 592
use sky130_fd_sc_hd__mux2_2  _326_
timestamp 1665323087
transform 1 0 7912 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _327_
timestamp 1665323087
transform -1 0 7728 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_2  _328_
timestamp 1665323087
transform -1 0 14444 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_2  _329_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform -1 0 13800 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__and3_2  _330_
timestamp 1665323087
transform 1 0 10028 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__and2_2  _331_
timestamp 1665323087
transform -1 0 10856 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_2  _332_
timestamp 1665323087
transform -1 0 9660 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__nand2b_2  _333_
timestamp 1665323087
transform 1 0 9844 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_2  _334_
timestamp 1665323087
transform 1 0 10672 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_2  _335_
timestamp 1665323087
transform 1 0 10580 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_2  _336_
timestamp 1665323087
transform -1 0 10120 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_2  _337_
timestamp 1665323087
transform 1 0 10764 0 1 2176
box -38 -48 682 592
use sky130_fd_sc_hd__and2_2  _338_
timestamp 1665323087
transform 1 0 11592 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _339_
timestamp 1665323087
transform 1 0 11960 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_2  _340_
timestamp 1665323087
transform 1 0 10120 0 1 1088
box -38 -48 1234 592
use sky130_fd_sc_hd__a21boi_2  _341_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform 1 0 10488 0 -1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__nand3_2  _342_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform 1 0 9016 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_2  _343_
timestamp 1665323087
transform 1 0 17480 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _344_
timestamp 1665323087
transform 1 0 17572 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_2  _345_
timestamp 1665323087
transform 1 0 17296 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _346_
timestamp 1665323087
transform -1 0 17296 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__nand2b_2  _347_
timestamp 1665323087
transform -1 0 18216 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _348_
timestamp 1665323087
transform 1 0 6440 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _349_
timestamp 1665323087
transform 1 0 6440 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_2  _350_
timestamp 1665323087
transform -1 0 6164 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_2  _351_
timestamp 1665323087
transform -1 0 6256 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _352_
timestamp 1665323087
transform -1 0 5888 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_2  _353_
timestamp 1665323087
transform -1 0 10948 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__and2b_2  _354_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform -1 0 10212 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__and3_2  _355_
timestamp 1665323087
transform -1 0 12328 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_2  _356_
timestamp 1665323087
transform 1 0 10304 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _357_
timestamp 1665323087
transform -1 0 9476 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _358_
timestamp 1665323087
transform 1 0 6072 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__and2_2  _359_
timestamp 1665323087
transform 1 0 10488 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_2  _360_
timestamp 1665323087
transform -1 0 2760 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_2  _361_
timestamp 1665323087
transform 1 0 12972 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _362_
timestamp 1665323087
transform 1 0 13984 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__a211o_2  _363_
timestamp 1665323087
transform 1 0 14168 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_2  _364_
timestamp 1665323087
transform -1 0 6164 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _365_
timestamp 1665323087
transform 1 0 12512 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__and2_2  _366_
timestamp 1665323087
transform 1 0 10764 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_2  _367_
timestamp 1665323087
transform -1 0 11592 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_2  _368_
timestamp 1665323087
transform 1 0 11868 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_2  _369_
timestamp 1665323087
transform -1 0 4048 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_2  _370_
timestamp 1665323087
transform -1 0 13800 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _371_
timestamp 1665323087
transform -1 0 12328 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_2  _372_
timestamp 1665323087
transform -1 0 9752 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_2  _373_
timestamp 1665323087
transform 1 0 1748 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_2  _374_
timestamp 1665323087
transform -1 0 8556 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_2  _375_
timestamp 1665323087
transform -1 0 4508 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_2  _376_
timestamp 1665323087
transform -1 0 9384 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_2  _377_
timestamp 1665323087
transform 1 0 6808 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_2  _378_
timestamp 1665323087
transform -1 0 7084 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _379_
timestamp 1665323087
transform -1 0 11960 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_2  _380_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform 1 0 11040 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _381_
timestamp 1665323087
transform 1 0 16008 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_2  _382_
timestamp 1665323087
transform -1 0 11684 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _383_
timestamp 1665323087
transform 1 0 11592 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__nand2b_2  _384_
timestamp 1665323087
transform 1 0 5520 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__o31a_2  _385_
timestamp 1665323087
transform -1 0 7728 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_2  _386_
timestamp 1665323087
transform -1 0 9384 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_2  _387_
timestamp 1665323087
transform 1 0 6900 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__o21a_2  _388_
timestamp 1665323087
transform 1 0 6992 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_2  _389_
timestamp 1665323087
transform -1 0 7360 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _390_
timestamp 1665323087
transform 1 0 13156 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_2  _391_
timestamp 1665323087
transform -1 0 8648 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_2  _392_
timestamp 1665323087
transform 1 0 8004 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_2  _393_
timestamp 1665323087
transform 1 0 10396 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_2  _394_
timestamp 1665323087
transform 1 0 9660 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_2  _395_
timestamp 1665323087
transform 1 0 9752 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _396_
timestamp 1665323087
transform 1 0 10488 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_2  _397_
timestamp 1665323087
transform 1 0 15180 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__and2_2  _398_
timestamp 1665323087
transform 1 0 12236 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_2  _399_
timestamp 1665323087
transform 1 0 12420 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__nand2b_2  _400_
timestamp 1665323087
transform 1 0 13156 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_2  _401_
timestamp 1665323087
transform 1 0 13064 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__o22a_2  _402_
timestamp 1665323087
transform -1 0 13892 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__and3_2  _403_
timestamp 1665323087
transform 1 0 13064 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_2  _404_
timestamp 1665323087
transform 1 0 13800 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__nand3_2  _405_
timestamp 1665323087
transform 1 0 15088 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__nand3b_2  _406_
timestamp 1665323087
transform 1 0 14168 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__and3_2  _407_
timestamp 1665323087
transform 1 0 14260 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_2  _408_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform 1 0 14168 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__a32o_2  _409_
timestamp 1665323087
transform 1 0 14812 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_2  _410_
timestamp 1665323087
transform 1 0 12144 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_2  _411_
timestamp 1665323087
transform -1 0 10856 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__o22a_2  _412_
timestamp 1665323087
transform 1 0 7820 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_2  _413_
timestamp 1665323087
transform 1 0 8004 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__o2111a_2  _414_
timestamp 1665323087
transform 1 0 9384 0 -1 11968
box -38 -48 958 592
use sky130_fd_sc_hd__o21ai_2  _415_
timestamp 1665323087
transform 1 0 9384 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_2  _416_
timestamp 1665323087
transform -1 0 9568 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_2  _417_
timestamp 1665323087
transform 1 0 9016 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__o31a_2  _418_
timestamp 1665323087
transform -1 0 14904 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_2  _419_
timestamp 1665323087
transform -1 0 17296 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__nand3_2  _420_
timestamp 1665323087
transform 1 0 15180 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__a32o_2  _421_
timestamp 1665323087
transform -1 0 15916 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_2  _422_
timestamp 1665323087
transform 1 0 16744 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_2  _423_
timestamp 1665323087
transform 1 0 15180 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _424_
timestamp 1665323087
transform 1 0 15088 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_2  _425_
timestamp 1665323087
transform 1 0 4232 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _426_
timestamp 1665323087
transform 1 0 8556 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_2  _427_
timestamp 1665323087
transform -1 0 17388 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _428_
timestamp 1665323087
transform -1 0 18400 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _429_
timestamp 1665323087
transform 1 0 14168 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_2  _430_
timestamp 1665323087
transform 1 0 13892 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _431_
timestamp 1665323087
transform 1 0 9108 0 1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _432_
timestamp 1665323087
transform -1 0 12788 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _433_
timestamp 1665323087
transform -1 0 13708 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _434_
timestamp 1665323087
transform 1 0 9108 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_2  _435_
timestamp 1665323087
transform -1 0 13432 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _436_
timestamp 1665323087
transform -1 0 8740 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _437_
timestamp 1665323087
transform 1 0 13432 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _438_
timestamp 1665323087
transform 1 0 14168 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_2  _439_
timestamp 1665323087
transform -1 0 9660 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _440_
timestamp 1665323087
transform -1 0 12144 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _441_
timestamp 1665323087
transform 1 0 14168 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _442_
timestamp 1665323087
transform 1 0 9844 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _443_
timestamp 1665323087
transform -1 0 7728 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_2  _444_
timestamp 1665323087
transform 1 0 12328 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _445_
timestamp 1665323087
transform 1 0 13892 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _446_
timestamp 1665323087
transform 1 0 14168 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _447_
timestamp 1665323087
transform -1 0 6808 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_2  _448_
timestamp 1665323087
transform -1 0 16284 0 -1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _449_
timestamp 1665323087
transform 1 0 16744 0 1 1088
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _450_
timestamp 1665323087
transform -1 0 5612 0 1 1088
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _451_
timestamp 1665323087
transform 1 0 5704 0 -1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _452_
timestamp 1665323087
transform -1 0 7912 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _453_
timestamp 1665323087
transform -1 0 5980 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _454_
timestamp 1665323087
transform -1 0 8740 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__dfrtp_2  _455_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform 1 0 15088 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _456_
timestamp 1665323087
transform 1 0 15088 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _457_
timestamp 1665323087
transform 1 0 14536 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _458_
timestamp 1665323087
transform -1 0 10212 0 -1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _459_
timestamp 1665323087
transform -1 0 13524 0 -1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _460_
timestamp 1665323087
transform 1 0 11960 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _461_
timestamp 1665323087
transform 1 0 11592 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _462_
timestamp 1665323087
transform -1 0 9844 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _463_
timestamp 1665323087
transform 1 0 13708 0 -1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _464_
timestamp 1665323087
transform 1 0 6992 0 -1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _465_
timestamp 1665323087
transform -1 0 13064 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _466_
timestamp 1665323087
transform 1 0 14904 0 1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _467_
timestamp 1665323087
transform 1 0 9108 0 -1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _468_
timestamp 1665323087
transform 1 0 11592 0 -1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _469_
timestamp 1665323087
transform 1 0 14720 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _470_
timestamp 1665323087
transform -1 0 15640 0 -1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _471_
timestamp 1665323087
transform 1 0 14536 0 1 1088
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _472_
timestamp 1665323087
transform 1 0 14536 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _473_
timestamp 1665323087
transform 1 0 3312 0 -1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _474_
timestamp 1665323087
transform 1 0 5704 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _475_
timestamp 1665323087
transform 1 0 6440 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _476_
timestamp 1665323087
transform 1 0 2392 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _477_
timestamp 1665323087
transform 1 0 6164 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__clkbuf_16  clockp_buffer_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform -1 0 3312 0 1 1088
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clockp_buffer_1
timestamp 1665323087
transform 1 0 1472 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[0\].id.delaybuf0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform -1 0 4600 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[0\].id.delaybuf1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform 1 0 4876 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[0\].id.delayen0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform 1 0 3956 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[0\].id.delayen1
timestamp 1665323087
transform -1 0 5152 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__einvn_8  ringosc.dstage\[0\].id.delayenb0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform 1 0 2576 0 -1 8704
box -38 -48 1694 592
use sky130_fd_sc_hd__einvn_4  ringosc.dstage\[0\].id.delayenb1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform -1 0 5428 0 -1 8704
box -38 -48 1050 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[0\].id.delayint0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform 1 0 5336 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[1\].id.delaybuf0
timestamp 1665323087
transform 1 0 4784 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[1\].id.delaybuf1
timestamp 1665323087
transform 1 0 5060 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[1\].id.delayen0
timestamp 1665323087
transform 1 0 2944 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[1\].id.delayen1
timestamp 1665323087
transform -1 0 4600 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__einvn_8  ringosc.dstage\[1\].id.delayenb0
timestamp 1665323087
transform 1 0 2760 0 -1 9792
box -38 -48 1694 592
use sky130_fd_sc_hd__einvn_4  ringosc.dstage\[1\].id.delayenb1
timestamp 1665323087
transform -1 0 4876 0 1 9792
box -38 -48 1050 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[1\].id.delayint0
timestamp 1665323087
transform -1 0 3772 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[2\].id.delaybuf0
timestamp 1665323087
transform 1 0 4784 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[2\].id.delaybuf1
timestamp 1665323087
transform 1 0 14996 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[2\].id.delayen0
timestamp 1665323087
transform 1 0 14168 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[2\].id.delayen1
timestamp 1665323087
transform 1 0 13248 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__einvn_8  ringosc.dstage\[2\].id.delayenb0
timestamp 1665323087
transform 1 0 14168 0 1 11968
box -38 -48 1694 592
use sky130_fd_sc_hd__einvn_4  ringosc.dstage\[2\].id.delayenb1
timestamp 1665323087
transform 1 0 13064 0 -1 13056
box -38 -48 1050 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[2\].id.delayint0
timestamp 1665323087
transform 1 0 16100 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[3\].id.delaybuf0
timestamp 1665323087
transform -1 0 14628 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[3\].id.delaybuf1
timestamp 1665323087
transform 1 0 11592 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[3\].id.delayen0
timestamp 1665323087
transform 1 0 6624 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[3\].id.delayen1
timestamp 1665323087
transform -1 0 11316 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__einvn_8  ringosc.dstage\[3\].id.delayenb0
timestamp 1665323087
transform 1 0 6256 0 1 11968
box -38 -48 1694 592
use sky130_fd_sc_hd__einvn_4  ringosc.dstage\[3\].id.delayenb1
timestamp 1665323087
transform -1 0 12604 0 -1 13056
box -38 -48 1050 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[3\].id.delayint0
timestamp 1665323087
transform -1 0 10764 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[4\].id.delaybuf0
timestamp 1665323087
transform -1 0 7636 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[4\].id.delaybuf1
timestamp 1665323087
transform 1 0 5796 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[4\].id.delayen0
timestamp 1665323087
transform 1 0 4232 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[4\].id.delayen1
timestamp 1665323087
transform -1 0 6164 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__einvn_8  ringosc.dstage\[4\].id.delayenb0
timestamp 1665323087
transform 1 0 3864 0 1 10880
box -38 -48 1694 592
use sky130_fd_sc_hd__einvn_4  ringosc.dstage\[4\].id.delayenb1
timestamp 1665323087
transform -1 0 6716 0 1 10880
box -38 -48 1050 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[4\].id.delayint0
timestamp 1665323087
transform -1 0 5336 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[5\].id.delaybuf0
timestamp 1665323087
transform -1 0 3220 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[5\].id.delaybuf1
timestamp 1665323087
transform 1 0 2668 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[5\].id.delayen0
timestamp 1665323087
transform 1 0 1748 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[5\].id.delayen1
timestamp 1665323087
transform 1 0 1748 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__einvn_8  ringosc.dstage\[5\].id.delayenb0
timestamp 1665323087
transform 1 0 1472 0 1 10880
box -38 -48 1694 592
use sky130_fd_sc_hd__einvn_4  ringosc.dstage\[5\].id.delayenb1
timestamp 1665323087
transform 1 0 1656 0 -1 13056
box -38 -48 1050 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[5\].id.delayint0
timestamp 1665323087
transform 1 0 2208 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[6\].id.delaybuf0
timestamp 1665323087
transform 1 0 2852 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[6\].id.delaybuf1
timestamp 1665323087
transform 1 0 7820 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[6\].id.delayen0
timestamp 1665323087
transform -1 0 4876 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[6\].id.delayen1
timestamp 1665323087
transform -1 0 5428 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__einvn_8  ringosc.dstage\[6\].id.delayenb0
timestamp 1665323087
transform -1 0 4600 0 -1 13056
box -38 -48 1694 592
use sky130_fd_sc_hd__einvn_4  ringosc.dstage\[6\].id.delayenb1
timestamp 1665323087
transform -1 0 5796 0 -1 13056
box -38 -48 1050 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[6\].id.delayint0
timestamp 1665323087
transform -1 0 3588 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[7\].id.delaybuf0
timestamp 1665323087
transform 1 0 5428 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[7\].id.delaybuf1
timestamp 1665323087
transform 1 0 9936 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[7\].id.delayen0
timestamp 1665323087
transform 1 0 8096 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[7\].id.delayen1
timestamp 1665323087
transform 1 0 9108 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__einvn_8  ringosc.dstage\[7\].id.delayenb0
timestamp 1665323087
transform 1 0 7452 0 -1 13056
box -38 -48 1694 592
use sky130_fd_sc_hd__einvn_4  ringosc.dstage\[7\].id.delayenb1
timestamp 1665323087
transform 1 0 9292 0 -1 13056
box -38 -48 1050 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[7\].id.delayint0
timestamp 1665323087
transform -1 0 8740 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[8\].id.delaybuf0
timestamp 1665323087
transform 1 0 15548 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[8\].id.delaybuf1
timestamp 1665323087
transform 1 0 18216 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[8\].id.delayen0
timestamp 1665323087
transform 1 0 16744 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[8\].id.delayen1
timestamp 1665323087
transform 1 0 17480 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__einvn_8  ringosc.dstage\[8\].id.delayenb0
timestamp 1665323087
transform 1 0 14812 0 -1 13056
box -38 -48 1694 592
use sky130_fd_sc_hd__einvn_4  ringosc.dstage\[8\].id.delayenb1
timestamp 1665323087
transform 1 0 17020 0 -1 13056
box -38 -48 1050 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[8\].id.delayint0
timestamp 1665323087
transform -1 0 17848 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[9\].id.delaybuf0
timestamp 1665323087
transform 1 0 16100 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[9\].id.delaybuf1
timestamp 1665323087
transform -1 0 16468 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[9\].id.delayen0
timestamp 1665323087
transform 1 0 17756 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[9\].id.delayen1
timestamp 1665323087
transform -1 0 17756 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__einvn_8  ringosc.dstage\[9\].id.delayenb0
timestamp 1665323087
transform 1 0 16836 0 -1 11968
box -38 -48 1694 592
use sky130_fd_sc_hd__einvn_4  ringosc.dstage\[9\].id.delayenb1
timestamp 1665323087
transform 1 0 15916 0 1 10880
box -38 -48 1050 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[9\].id.delayint0
timestamp 1665323087
transform -1 0 16468 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[10\].id.delaybuf0
timestamp 1665323087
transform -1 0 18308 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[10\].id.delaybuf1
timestamp 1665323087
transform 1 0 17940 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[10\].id.delayen0
timestamp 1665323087
transform 1 0 17572 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[10\].id.delayen1
timestamp 1665323087
transform 1 0 16928 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__einvn_8  ringosc.dstage\[10\].id.delayenb0
timestamp 1665323087
transform 1 0 16652 0 1 8704
box -38 -48 1694 592
use sky130_fd_sc_hd__einvn_4  ringosc.dstage\[10\].id.delayenb1
timestamp 1665323087
transform 1 0 16744 0 1 9792
box -38 -48 1050 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[10\].id.delayint0
timestamp 1665323087
transform -1 0 16468 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[11\].id.delaybuf0
timestamp 1665323087
transform -1 0 18124 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[11\].id.delaybuf1
timestamp 1665323087
transform 1 0 17940 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[11\].id.delayen0
timestamp 1665323087
transform 1 0 16008 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[11\].id.delayen1
timestamp 1665323087
transform 1 0 16744 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__einvn_8  ringosc.dstage\[11\].id.delayenb0
timestamp 1665323087
transform 1 0 16836 0 1 7616
box -38 -48 1694 592
use sky130_fd_sc_hd__einvn_4  ringosc.dstage\[11\].id.delayenb1
timestamp 1665323087
transform 1 0 16744 0 -1 7616
box -38 -48 1050 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[11\].id.delayint0
timestamp 1665323087
transform -1 0 16468 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  ringosc.ibufp00 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform -1 0 3220 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_8  ringosc.ibufp01 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform -1 0 2668 0 -1 5440
box -38 -48 1234 592
use sky130_fd_sc_hd__clkinv_2  ringosc.ibufp10
timestamp 1665323087
transform -1 0 2300 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_8  ringosc.ibufp11
timestamp 1665323087
transform 1 0 1472 0 1 8704
box -38 -48 1234 592
use sky130_fd_sc_hd__conb_1  ringosc.iss.const1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform 1 0 17940 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__or2_2  ringosc.iss.ctrlen0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform 1 0 16008 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.iss.delaybuf0
timestamp 1665323087
transform -1 0 18124 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_2  ringosc.iss.delayen0
timestamp 1665323087
transform 1 0 17020 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__einvp_2  ringosc.iss.delayen1
timestamp 1665323087
transform 1 0 17572 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__einvn_8  ringosc.iss.delayenb0
timestamp 1665323087
transform 1 0 16836 0 -1 6528
box -38 -48 1694 592
use sky130_fd_sc_hd__einvn_4  ringosc.iss.delayenb1
timestamp 1665323087
transform 1 0 16376 0 1 6528
box -38 -48 1050 592
use sky130_fd_sc_hd__clkinv_1  ringosc.iss.delayint0
timestamp 1665323087
transform 1 0 17296 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_1  ringosc.iss.reseten0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform 1 0 17296 0 -1 4352
box -38 -48 498 592
<< labels >>
flabel metal4 s 8208 1040 8528 13648 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 16208 1040 16528 13648 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal5 s 1056 8210 18908 8530 0 FreeSans 2560 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 4208 1040 4528 13648 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 12208 1040 12528 13648 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal5 s 1056 4210 18908 4530 0 FreeSans 2560 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal5 s 1056 12210 18908 12530 0 FreeSans 2560 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal3 s 0 1232 800 1352 0 FreeSans 480 0 0 0 clockp[0]
port 2 nsew signal tristate
flabel metal3 s 0 2048 800 2168 0 FreeSans 480 0 0 0 clockp[1]
port 3 nsew signal tristate
flabel metal3 s 0 7760 800 7880 0 FreeSans 480 0 0 0 dco
port 4 nsew signal input
flabel metal3 s 0 2864 800 2984 0 FreeSans 480 0 0 0 div[0]
port 5 nsew signal input
flabel metal3 s 0 3680 800 3800 0 FreeSans 480 0 0 0 div[1]
port 6 nsew signal input
flabel metal3 s 0 4496 800 4616 0 FreeSans 480 0 0 0 div[2]
port 7 nsew signal input
flabel metal3 s 0 5312 800 5432 0 FreeSans 480 0 0 0 div[3]
port 8 nsew signal input
flabel metal3 s 0 6128 800 6248 0 FreeSans 480 0 0 0 div[4]
port 9 nsew signal input
flabel metal3 s 0 6944 800 7064 0 FreeSans 480 0 0 0 enable
port 10 nsew signal input
flabel metal3 s 0 8576 800 8696 0 FreeSans 480 0 0 0 ext_trim[0]
port 11 nsew signal input
flabel metal2 s 5538 14200 5594 15000 0 FreeSans 224 90 0 0 ext_trim[10]
port 12 nsew signal input
flabel metal2 s 7010 14200 7066 15000 0 FreeSans 224 90 0 0 ext_trim[11]
port 13 nsew signal input
flabel metal2 s 8482 14200 8538 15000 0 FreeSans 224 90 0 0 ext_trim[12]
port 14 nsew signal input
flabel metal2 s 9954 14200 10010 15000 0 FreeSans 224 90 0 0 ext_trim[13]
port 15 nsew signal input
flabel metal2 s 11426 14200 11482 15000 0 FreeSans 224 90 0 0 ext_trim[14]
port 16 nsew signal input
flabel metal2 s 12898 14200 12954 15000 0 FreeSans 224 90 0 0 ext_trim[15]
port 17 nsew signal input
flabel metal2 s 14370 14200 14426 15000 0 FreeSans 224 90 0 0 ext_trim[16]
port 18 nsew signal input
flabel metal2 s 15842 14200 15898 15000 0 FreeSans 224 90 0 0 ext_trim[17]
port 19 nsew signal input
flabel metal2 s 17314 14200 17370 15000 0 FreeSans 224 90 0 0 ext_trim[18]
port 20 nsew signal input
flabel metal2 s 18786 14200 18842 15000 0 FreeSans 224 90 0 0 ext_trim[19]
port 21 nsew signal input
flabel metal3 s 0 9392 800 9512 0 FreeSans 480 0 0 0 ext_trim[1]
port 22 nsew signal input
flabel metal3 s 19200 13472 20000 13592 0 FreeSans 480 0 0 0 ext_trim[20]
port 23 nsew signal input
flabel metal3 s 19200 11024 20000 11144 0 FreeSans 480 0 0 0 ext_trim[21]
port 24 nsew signal input
flabel metal3 s 19200 8576 20000 8696 0 FreeSans 480 0 0 0 ext_trim[22]
port 25 nsew signal input
flabel metal3 s 19200 6128 20000 6248 0 FreeSans 480 0 0 0 ext_trim[23]
port 26 nsew signal input
flabel metal3 s 19200 3680 20000 3800 0 FreeSans 480 0 0 0 ext_trim[24]
port 27 nsew signal input
flabel metal3 s 19200 1232 20000 1352 0 FreeSans 480 0 0 0 ext_trim[25]
port 28 nsew signal input
flabel metal3 s 0 10208 800 10328 0 FreeSans 480 0 0 0 ext_trim[2]
port 29 nsew signal input
flabel metal3 s 0 11024 800 11144 0 FreeSans 480 0 0 0 ext_trim[3]
port 30 nsew signal input
flabel metal3 s 0 11840 800 11960 0 FreeSans 480 0 0 0 ext_trim[4]
port 31 nsew signal input
flabel metal3 s 0 12656 800 12776 0 FreeSans 480 0 0 0 ext_trim[5]
port 32 nsew signal input
flabel metal3 s 0 13472 800 13592 0 FreeSans 480 0 0 0 ext_trim[6]
port 33 nsew signal input
flabel metal2 s 1122 14200 1178 15000 0 FreeSans 224 90 0 0 ext_trim[7]
port 34 nsew signal input
flabel metal2 s 2594 14200 2650 15000 0 FreeSans 224 90 0 0 ext_trim[8]
port 35 nsew signal input
flabel metal2 s 4066 14200 4122 15000 0 FreeSans 224 90 0 0 ext_trim[9]
port 36 nsew signal input
flabel metal2 s 14922 0 14978 800 0 FreeSans 224 90 0 0 osc
port 37 nsew signal input
flabel metal2 s 4986 0 5042 800 0 FreeSans 224 90 0 0 resetb
port 38 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 20000 15000
<< end >>
