magic
tech sky130A
magscale 1 2
timestamp 1666034820
<< viali >>
rect 3617 13481 3651 13515
rect 4261 13481 4295 13515
rect 8677 13481 8711 13515
rect 10885 13481 10919 13515
rect 13461 13481 13495 13515
rect 5549 13413 5583 13447
rect 7573 13413 7607 13447
rect 7941 13413 7975 13447
rect 9137 13413 9171 13447
rect 12633 13413 12667 13447
rect 2697 13345 2731 13379
rect 4813 13345 4847 13379
rect 6193 13345 6227 13379
rect 6469 13345 6503 13379
rect 7021 13345 7055 13379
rect 9965 13345 9999 13379
rect 12173 13345 12207 13379
rect 1685 13277 1719 13311
rect 2237 13277 2271 13311
rect 2881 13277 2915 13311
rect 3433 13277 3467 13311
rect 4353 13277 4387 13311
rect 5641 13277 5675 13311
rect 6929 13277 6963 13311
rect 7757 13277 7791 13311
rect 8073 13277 8107 13311
rect 8309 13277 8343 13311
rect 8493 13277 8527 13311
rect 9321 13277 9355 13311
rect 10701 13277 10735 13311
rect 10977 13277 11011 13311
rect 11253 13277 11287 13311
rect 11621 13277 11655 13311
rect 12357 13277 12391 13311
rect 12817 13277 12851 13311
rect 12909 13277 12943 13311
rect 13185 13277 13219 13311
rect 1501 13209 1535 13243
rect 1961 13209 1995 13243
rect 2789 13209 2823 13243
rect 3341 13209 3375 13243
rect 3893 13209 3927 13243
rect 4077 13209 4111 13243
rect 4905 13209 4939 13243
rect 5365 13209 5399 13243
rect 6101 13209 6135 13243
rect 7389 13209 7423 13243
rect 8217 13209 8251 13243
rect 8585 13209 8619 13243
rect 9781 13209 9815 13243
rect 9873 13209 9907 13243
rect 10425 13209 10459 13243
rect 10517 13209 10551 13243
rect 12081 13209 12115 13243
rect 1869 13141 1903 13175
rect 2145 13141 2179 13175
rect 4997 13141 5031 13175
rect 5089 13141 5123 13175
rect 7297 13141 7331 13175
rect 9229 13141 9263 13175
rect 11069 13141 11103 13175
rect 12449 13141 12483 13175
rect 13093 13141 13127 13175
rect 13369 13141 13403 13175
rect 3433 12869 3467 12903
rect 5273 12869 5307 12903
rect 5641 12869 5675 12903
rect 7113 12869 7147 12903
rect 7297 12869 7331 12903
rect 7573 12869 7607 12903
rect 8493 12869 8527 12903
rect 11069 12869 11103 12903
rect 11345 12869 11379 12903
rect 13093 12869 13127 12903
rect 13369 12869 13403 12903
rect 1593 12801 1627 12835
rect 1869 12801 1903 12835
rect 3341 12801 3375 12835
rect 3709 12801 3743 12835
rect 4629 12801 4663 12835
rect 5825 12801 5859 12835
rect 6009 12801 6043 12835
rect 6101 12801 6135 12835
rect 6377 12801 6411 12835
rect 7757 12801 7791 12835
rect 8304 12801 8338 12835
rect 8401 12801 8435 12835
rect 8677 12801 8711 12835
rect 8769 12801 8803 12835
rect 9689 12801 9723 12835
rect 10425 12801 10459 12835
rect 11529 12801 11563 12835
rect 12449 12801 12483 12835
rect 1777 12733 1811 12767
rect 7941 12733 7975 12767
rect 5457 12665 5491 12699
rect 10057 12665 10091 12699
rect 3617 12597 3651 12631
rect 8125 12597 8159 12631
rect 13277 12597 13311 12631
rect 4905 12393 4939 12427
rect 7205 12393 7239 12427
rect 9873 12393 9907 12427
rect 10149 12393 10183 12427
rect 10425 12393 10459 12427
rect 2973 12325 3007 12359
rect 5181 12325 5215 12359
rect 6653 12325 6687 12359
rect 1777 12189 1811 12223
rect 2053 12189 2087 12223
rect 2697 12189 2731 12223
rect 2789 12189 2823 12223
rect 3617 12189 3651 12223
rect 4721 12189 4755 12223
rect 5089 12189 5123 12223
rect 5365 12189 5399 12223
rect 6837 12189 6871 12223
rect 7337 12189 7371 12223
rect 7481 12189 7515 12223
rect 7757 12189 7791 12223
rect 7849 12189 7883 12223
rect 8033 12189 8067 12223
rect 8125 12189 8159 12223
rect 8218 12199 8252 12233
rect 8769 12189 8803 12223
rect 9229 12189 9263 12223
rect 9321 12189 9355 12223
rect 9741 12189 9775 12223
rect 10241 12189 10275 12223
rect 10609 12189 10643 12223
rect 10885 12189 10919 12223
rect 10977 12189 11011 12223
rect 11621 12189 11655 12223
rect 11897 12189 11931 12223
rect 11989 12189 12023 12223
rect 13277 12189 13311 12223
rect 1501 12121 1535 12155
rect 1685 12121 1719 12155
rect 3065 12121 3099 12155
rect 3157 12121 3191 12155
rect 3801 12121 3835 12155
rect 4077 12121 4111 12155
rect 7573 12121 7607 12155
rect 8493 12121 8527 12155
rect 9505 12121 9539 12155
rect 9597 12121 9631 12155
rect 13553 12121 13587 12155
rect 8677 12053 8711 12087
rect 9137 12053 9171 12087
rect 10793 12053 10827 12087
rect 2697 11849 2731 11883
rect 3341 11849 3375 11883
rect 7021 11849 7055 11883
rect 7113 11849 7147 11883
rect 7849 11849 7883 11883
rect 8309 11849 8343 11883
rect 2329 11781 2363 11815
rect 3709 11781 3743 11815
rect 4353 11781 4387 11815
rect 4445 11781 4479 11815
rect 7665 11781 7699 11815
rect 9689 11781 9723 11815
rect 10149 11781 10183 11815
rect 10241 11781 10275 11815
rect 10425 11781 10459 11815
rect 10793 11781 10827 11815
rect 10885 11781 10919 11815
rect 12081 11781 12115 11815
rect 13093 11781 13127 11815
rect 13277 11781 13311 11815
rect 13461 11781 13495 11815
rect 1593 11713 1627 11747
rect 2513 11713 2547 11747
rect 2789 11713 2823 11747
rect 3065 11713 3099 11747
rect 3249 11713 3283 11747
rect 3525 11713 3559 11747
rect 5365 11713 5399 11747
rect 6193 11713 6227 11747
rect 6653 11713 6687 11747
rect 6837 11713 6871 11747
rect 7225 11713 7259 11747
rect 7481 11713 7515 11747
rect 8585 11713 8619 11747
rect 8861 11713 8895 11747
rect 9045 11713 9079 11747
rect 9137 11713 9171 11747
rect 9281 11713 9315 11747
rect 9873 11713 9907 11747
rect 10057 11713 10091 11747
rect 11529 11713 11563 11747
rect 12173 11713 12207 11747
rect 2145 11645 2179 11679
rect 3893 11645 3927 11679
rect 4537 11645 4571 11679
rect 5089 11645 5123 11679
rect 5733 11645 5767 11679
rect 5917 11645 5951 11679
rect 6929 11645 6963 11679
rect 8217 11645 8251 11679
rect 8493 11645 8527 11679
rect 11345 11645 11379 11679
rect 11989 11645 12023 11679
rect 12541 11645 12575 11679
rect 2053 11577 2087 11611
rect 4629 11577 4663 11611
rect 6101 11577 6135 11611
rect 6745 11577 6779 11611
rect 8033 11577 8067 11611
rect 13001 11577 13035 11611
rect 1501 11509 1535 11543
rect 2973 11509 3007 11543
rect 5273 11509 5307 11543
rect 8777 11509 8811 11543
rect 9413 11509 9447 11543
rect 10425 11509 10459 11543
rect 10609 11509 10643 11543
rect 12265 11509 12299 11543
rect 6285 11305 6319 11339
rect 7757 11305 7791 11339
rect 10517 11305 10551 11339
rect 10885 11305 10919 11339
rect 11437 11305 11471 11339
rect 2697 11237 2731 11271
rect 5273 11237 5307 11271
rect 6101 11237 6135 11271
rect 7941 11237 7975 11271
rect 9689 11237 9723 11271
rect 12173 11237 12207 11271
rect 3065 11169 3099 11203
rect 3617 11169 3651 11203
rect 3893 11169 3927 11203
rect 6929 11169 6963 11203
rect 7205 11169 7239 11203
rect 7297 11169 7331 11203
rect 8953 11169 8987 11203
rect 10057 11169 10091 11203
rect 1409 11101 1443 11135
rect 2329 11101 2363 11135
rect 3985 11101 4019 11135
rect 5365 11101 5399 11135
rect 5917 11101 5951 11135
rect 6193 11101 6227 11135
rect 6469 11101 6503 11135
rect 6725 11101 6759 11135
rect 7019 11101 7053 11135
rect 7481 11101 7515 11135
rect 7573 11101 7607 11135
rect 8216 11101 8250 11135
rect 8309 11101 8343 11135
rect 8401 11101 8435 11135
rect 8585 11101 8619 11135
rect 9137 11101 9171 11135
rect 9275 11101 9309 11135
rect 9505 11101 9539 11135
rect 9597 11101 9631 11135
rect 9965 11101 9999 11135
rect 10241 11101 10275 11135
rect 10333 11101 10367 11135
rect 10793 11101 10827 11135
rect 11069 11101 11103 11135
rect 11621 11101 11655 11135
rect 11989 11101 12023 11135
rect 12357 11101 12391 11135
rect 13277 11101 13311 11135
rect 3157 11033 3191 11067
rect 8769 11033 8803 11067
rect 11897 11033 11931 11067
rect 13001 11033 13035 11067
rect 13553 11033 13587 11067
rect 5733 10965 5767 10999
rect 6837 10965 6871 10999
rect 11805 10965 11839 10999
rect 13369 10965 13403 10999
rect 1501 10761 1535 10795
rect 9321 10761 9355 10795
rect 11253 10761 11287 10795
rect 12541 10761 12575 10795
rect 2697 10693 2731 10727
rect 3893 10693 3927 10727
rect 4261 10693 4295 10727
rect 5089 10693 5123 10727
rect 5641 10693 5675 10727
rect 10057 10693 10091 10727
rect 10241 10693 10275 10727
rect 12173 10693 12207 10727
rect 13093 10693 13127 10727
rect 1409 10625 1443 10659
rect 1685 10625 1719 10659
rect 2513 10625 2547 10659
rect 2973 10625 3007 10659
rect 3617 10625 3651 10659
rect 4077 10625 4111 10659
rect 4353 10625 4387 10659
rect 4445 10625 4479 10659
rect 5365 10625 5399 10659
rect 5733 10625 5767 10659
rect 5917 10625 5951 10659
rect 6469 10625 6503 10659
rect 6929 10625 6963 10659
rect 7113 10625 7147 10659
rect 7297 10625 7331 10659
rect 7481 10625 7515 10659
rect 7757 10625 7791 10659
rect 7939 10625 7973 10659
rect 8126 10625 8160 10659
rect 8217 10625 8251 10659
rect 8310 10625 8344 10659
rect 8585 10625 8619 10659
rect 8677 10625 8711 10659
rect 8861 10625 8895 10659
rect 9045 10625 9079 10659
rect 9505 10625 9539 10659
rect 9597 10625 9631 10659
rect 10517 10625 10551 10659
rect 10609 10625 10643 10659
rect 10792 10625 10826 10659
rect 10885 10625 10919 10659
rect 11161 10625 11195 10659
rect 11529 10625 11563 10659
rect 11713 10625 11747 10659
rect 11943 10625 11977 10659
rect 12057 10625 12091 10659
rect 12265 10625 12299 10659
rect 12909 10625 12943 10659
rect 13185 10625 13219 10659
rect 13461 10625 13495 10659
rect 1869 10557 1903 10591
rect 2053 10557 2087 10591
rect 2605 10557 2639 10591
rect 6653 10557 6687 10591
rect 6837 10557 6871 10591
rect 9873 10557 9907 10591
rect 10977 10557 11011 10591
rect 12357 10557 12391 10591
rect 12449 10557 12483 10591
rect 12653 10557 12687 10591
rect 5457 10489 5491 10523
rect 7113 10489 7147 10523
rect 13461 10489 13495 10523
rect 6101 10421 6135 10455
rect 7573 10421 7607 10455
rect 9781 10421 9815 10455
rect 10241 10421 10275 10455
rect 1501 10217 1535 10251
rect 3985 10217 4019 10251
rect 7665 10217 7699 10251
rect 8493 10217 8527 10251
rect 9137 10217 9171 10251
rect 11897 10217 11931 10251
rect 12173 10217 12207 10251
rect 3341 10149 3375 10183
rect 5273 10149 5307 10183
rect 6469 10149 6503 10183
rect 7113 10149 7147 10183
rect 7297 10149 7331 10183
rect 8677 10149 8711 10183
rect 11069 10149 11103 10183
rect 13277 10149 13311 10183
rect 6377 10081 6411 10115
rect 10149 10081 10183 10115
rect 13369 10081 13403 10115
rect 1685 10013 1719 10047
rect 2053 10013 2087 10047
rect 3065 10013 3099 10047
rect 3801 10013 3835 10047
rect 4169 10013 4203 10047
rect 4537 10013 4571 10047
rect 4813 10013 4847 10047
rect 6009 10013 6043 10047
rect 6607 10013 6641 10047
rect 6751 10013 6785 10047
rect 7941 10013 7975 10047
rect 8217 10013 8251 10047
rect 9321 10013 9355 10047
rect 9413 10013 9447 10047
rect 9597 10013 9631 10047
rect 9689 10013 9723 10047
rect 9873 10013 9907 10047
rect 10057 10013 10091 10047
rect 10241 10023 10275 10057
rect 10885 10013 10919 10047
rect 10977 10013 11011 10047
rect 11161 10013 11195 10047
rect 11529 10013 11563 10047
rect 11621 10013 11655 10047
rect 11989 10013 12023 10047
rect 12081 10013 12115 10047
rect 12449 10013 12483 10047
rect 12541 10013 12575 10047
rect 12817 10013 12851 10047
rect 1593 9945 1627 9979
rect 4353 9945 4387 9979
rect 5365 9945 5399 9979
rect 5457 9945 5491 9979
rect 5825 9945 5859 9979
rect 6285 9945 6319 9979
rect 7573 9945 7607 9979
rect 8309 9945 8343 9979
rect 10333 9945 10367 9979
rect 13461 9945 13495 9979
rect 1869 9877 1903 9911
rect 5641 9877 5675 9911
rect 6193 9877 6227 9911
rect 8125 9877 8159 9911
rect 8493 9877 8527 9911
rect 6193 9673 6227 9707
rect 7021 9673 7055 9707
rect 7205 9673 7239 9707
rect 9689 9673 9723 9707
rect 11253 9673 11287 9707
rect 2881 9605 2915 9639
rect 7398 9605 7432 9639
rect 7803 9605 7837 9639
rect 8861 9605 8895 9639
rect 9413 9605 9447 9639
rect 10517 9605 10551 9639
rect 13185 9605 13219 9639
rect 13369 9605 13403 9639
rect 1869 9537 1903 9571
rect 2605 9537 2639 9571
rect 3157 9537 3191 9571
rect 3801 9537 3835 9571
rect 4077 9537 4111 9571
rect 4445 9537 4479 9571
rect 5917 9537 5951 9571
rect 6653 9537 6687 9571
rect 6837 9537 6871 9571
rect 7021 9537 7055 9571
rect 8217 9537 8251 9571
rect 8309 9537 8343 9571
rect 8585 9537 8619 9571
rect 8953 9537 8987 9571
rect 9045 9537 9079 9571
rect 9229 9537 9263 9571
rect 9873 9537 9907 9571
rect 10149 9537 10183 9571
rect 10333 9537 10367 9571
rect 10609 9537 10643 9571
rect 10793 9537 10827 9571
rect 11069 9537 11103 9571
rect 11713 9537 11747 9571
rect 11805 9537 11839 9571
rect 11989 9537 12023 9571
rect 12173 9537 12207 9571
rect 12449 9537 12483 9571
rect 8769 9469 8803 9503
rect 10057 9469 10091 9503
rect 5733 9401 5767 9435
rect 7941 9401 7975 9435
rect 11529 9401 11563 9435
rect 1501 9333 1535 9367
rect 2789 9333 2823 9367
rect 3893 9333 3927 9367
rect 4261 9333 4295 9367
rect 6469 9333 6503 9367
rect 7757 9333 7791 9367
rect 10701 9333 10735 9367
rect 13461 9333 13495 9367
rect 6101 9129 6135 9163
rect 6561 9129 6595 9163
rect 7481 9129 7515 9163
rect 7757 9129 7791 9163
rect 10701 9129 10735 9163
rect 11437 9129 11471 9163
rect 4629 9061 4663 9095
rect 6929 9061 6963 9095
rect 9229 9061 9263 9095
rect 11069 9061 11103 9095
rect 11157 9061 11191 9095
rect 3157 8993 3191 9027
rect 4721 8993 4755 9027
rect 7113 8993 7147 9027
rect 9777 8993 9811 9027
rect 10057 8993 10091 9027
rect 1409 8925 1443 8959
rect 3617 8925 3651 8959
rect 3893 8925 3927 8959
rect 4169 8925 4203 8959
rect 4629 8925 4663 8959
rect 5089 8925 5123 8959
rect 5733 8925 5767 8959
rect 6009 8925 6043 8959
rect 6377 8925 6411 8959
rect 6653 8925 6687 8959
rect 6929 8925 6963 8959
rect 7573 8925 7607 8959
rect 7941 8925 7975 8959
rect 8092 8925 8126 8959
rect 8217 8925 8251 8959
rect 8309 8925 8343 8959
rect 8493 8925 8527 8959
rect 8677 8925 8711 8959
rect 8953 8925 8987 8959
rect 9137 8925 9171 8959
rect 9597 8925 9631 8959
rect 9689 8925 9723 8959
rect 9873 8925 9907 8959
rect 10333 8925 10367 8959
rect 10517 8925 10551 8959
rect 10977 8925 11011 8959
rect 11253 8925 11287 8959
rect 11621 8925 11655 8959
rect 11989 8925 12023 8959
rect 13277 8925 13311 8959
rect 3801 8857 3835 8891
rect 4261 8857 4295 8891
rect 7297 8857 7331 8891
rect 8769 8857 8803 8891
rect 13553 8857 13587 8891
rect 3433 8789 3467 8823
rect 4905 8789 4939 8823
rect 10517 8789 10551 8823
rect 11805 8789 11839 8823
rect 1593 8585 1627 8619
rect 1869 8585 1903 8619
rect 2973 8585 3007 8619
rect 8953 8585 8987 8619
rect 3525 8517 3559 8551
rect 3617 8517 3651 8551
rect 5641 8517 5675 8551
rect 6193 8517 6227 8551
rect 6929 8517 6963 8551
rect 9965 8517 9999 8551
rect 10149 8517 10183 8551
rect 11713 8517 11747 8551
rect 11805 8517 11839 8551
rect 12449 8517 12483 8551
rect 13553 8517 13587 8551
rect 1409 8449 1443 8483
rect 1685 8449 1719 8483
rect 2053 8449 2087 8483
rect 2237 8449 2271 8483
rect 2329 8449 2363 8483
rect 2455 8449 2489 8483
rect 3249 8449 3283 8483
rect 4445 8449 4479 8483
rect 4813 8449 4847 8483
rect 5089 8449 5123 8483
rect 5181 8449 5215 8483
rect 5825 8449 5859 8483
rect 6101 8449 6135 8483
rect 6561 8449 6595 8483
rect 6745 8449 6779 8483
rect 7389 8449 7423 8483
rect 7665 8449 7699 8483
rect 7849 8449 7883 8483
rect 8401 8449 8435 8483
rect 8493 8449 8527 8483
rect 8861 8449 8895 8483
rect 9137 8449 9171 8483
rect 9321 8449 9355 8483
rect 9413 8449 9447 8483
rect 9597 8449 9631 8483
rect 10609 8449 10643 8483
rect 10793 8449 10827 8483
rect 11069 8449 11103 8483
rect 11253 8449 11287 8483
rect 11529 8449 11563 8483
rect 11949 8449 11983 8483
rect 12265 8449 12299 8483
rect 12541 8449 12575 8483
rect 12685 8449 12719 8483
rect 2881 8381 2915 8415
rect 3433 8381 3467 8415
rect 4077 8381 4111 8415
rect 4629 8381 4663 8415
rect 4721 8381 4755 8415
rect 5733 8381 5767 8415
rect 6377 8381 6411 8415
rect 7021 8381 7055 8415
rect 7573 8381 7607 8415
rect 13001 8381 13035 8415
rect 2697 8313 2731 8347
rect 4261 8313 4295 8347
rect 7113 8313 7147 8347
rect 7941 8313 7975 8347
rect 8217 8313 8251 8347
rect 10609 8313 10643 8347
rect 11253 8313 11287 8347
rect 12081 8313 12115 8347
rect 13461 8313 13495 8347
rect 8677 8245 8711 8279
rect 9781 8245 9815 8279
rect 10149 8245 10183 8279
rect 10333 8245 10367 8279
rect 12817 8245 12851 8279
rect 3525 8041 3559 8075
rect 5825 8041 5859 8075
rect 6193 8041 6227 8075
rect 9873 8041 9907 8075
rect 10701 8041 10735 8075
rect 13461 8041 13495 8075
rect 3065 7973 3099 8007
rect 10885 7973 10919 8007
rect 3801 7905 3835 7939
rect 5457 7905 5491 7939
rect 1685 7837 1719 7871
rect 1961 7837 1995 7871
rect 2053 7837 2087 7871
rect 2237 7837 2271 7871
rect 2421 7837 2455 7871
rect 2605 7837 2639 7871
rect 2973 7837 3007 7871
rect 3341 7837 3375 7871
rect 4076 7837 4110 7871
rect 4169 7837 4203 7871
rect 4261 7837 4295 7871
rect 4445 7837 4479 7871
rect 6009 7837 6043 7871
rect 6377 7837 6411 7871
rect 6469 7837 6503 7871
rect 7093 7837 7127 7871
rect 7389 7837 7423 7871
rect 7665 7837 7699 7871
rect 9321 7837 9355 7871
rect 9413 7837 9447 7871
rect 9689 7837 9723 7871
rect 9965 7837 9999 7871
rect 10233 7837 10267 7871
rect 11069 7837 11103 7871
rect 11253 7837 11287 7871
rect 11345 7837 11379 7871
rect 11454 7837 11488 7871
rect 11897 7837 11931 7871
rect 12081 7837 12115 7871
rect 12449 7837 12483 7871
rect 13369 7837 13403 7871
rect 1777 7769 1811 7803
rect 4905 7769 4939 7803
rect 6653 7769 6687 7803
rect 6837 7769 6871 7803
rect 8677 7769 8711 7803
rect 10333 7769 10367 7803
rect 10710 7769 10744 7803
rect 11713 7769 11747 7803
rect 13185 7769 13219 7803
rect 1501 7701 1535 7735
rect 3617 7701 3651 7735
rect 7205 7701 7239 7735
rect 7297 7701 7331 7735
rect 9137 7701 9171 7735
rect 11989 7701 12023 7735
rect 4353 7497 4387 7531
rect 6469 7497 6503 7531
rect 8033 7497 8067 7531
rect 9597 7497 9631 7531
rect 9781 7497 9815 7531
rect 9873 7497 9907 7531
rect 11529 7497 11563 7531
rect 13461 7497 13495 7531
rect 2973 7429 3007 7463
rect 3157 7429 3191 7463
rect 8401 7429 8435 7463
rect 10793 7429 10827 7463
rect 13185 7429 13219 7463
rect 1685 7361 1719 7395
rect 1869 7361 1903 7395
rect 2237 7361 2271 7395
rect 2329 7361 2363 7395
rect 2421 7361 2455 7395
rect 2513 7361 2547 7395
rect 3709 7361 3743 7395
rect 4721 7361 4755 7395
rect 4997 7361 5031 7395
rect 5181 7361 5215 7395
rect 5457 7361 5491 7395
rect 5641 7361 5675 7395
rect 5917 7361 5951 7395
rect 6561 7361 6595 7395
rect 7021 7361 7055 7395
rect 7941 7361 7975 7395
rect 8585 7361 8619 7395
rect 8953 7361 8987 7395
rect 9691 7361 9725 7395
rect 9985 7361 10019 7395
rect 10241 7361 10275 7395
rect 11897 7361 11931 7395
rect 12265 7361 12299 7395
rect 12725 7361 12759 7395
rect 13369 7361 13403 7395
rect 2053 7293 2087 7327
rect 3801 7293 3835 7327
rect 4905 7293 4939 7327
rect 7113 7293 7147 7327
rect 7757 7293 7791 7327
rect 10701 7293 10735 7327
rect 10885 7293 10919 7327
rect 13277 7293 13311 7327
rect 1777 7225 1811 7259
rect 5089 7225 5123 7259
rect 6101 7225 6135 7259
rect 8309 7225 8343 7259
rect 11253 7225 11287 7259
rect 2789 7157 2823 7191
rect 2973 7157 3007 7191
rect 4537 7157 4571 7191
rect 5549 7157 5583 7191
rect 10241 7157 10275 7191
rect 1777 6953 1811 6987
rect 4629 6953 4663 6987
rect 8493 6953 8527 6987
rect 3801 6885 3835 6919
rect 8309 6885 8343 6919
rect 10333 6885 10367 6919
rect 10421 6885 10455 6919
rect 10977 6885 11011 6919
rect 2053 6817 2087 6851
rect 2145 6817 2179 6851
rect 2973 6817 3007 6851
rect 3525 6817 3559 6851
rect 4813 6817 4847 6851
rect 6745 6817 6779 6851
rect 8677 6817 8711 6851
rect 12357 6817 12391 6851
rect 13369 6817 13403 6851
rect 1409 6749 1443 6783
rect 1961 6749 1995 6783
rect 2237 6749 2271 6783
rect 2421 6749 2455 6783
rect 2697 6749 2731 6783
rect 2789 6749 2823 6783
rect 3341 6749 3375 6783
rect 3985 6749 4019 6783
rect 4537 6749 4571 6783
rect 5089 6749 5123 6783
rect 5273 6749 5307 6783
rect 6101 6749 6135 6783
rect 6377 6749 6411 6783
rect 7205 6749 7239 6783
rect 7481 6749 7515 6783
rect 8217 6749 8251 6783
rect 9413 6749 9447 6783
rect 9689 6749 9723 6783
rect 10241 6749 10275 6783
rect 10517 6749 10551 6783
rect 10793 6749 10827 6783
rect 10885 6749 10919 6783
rect 11161 6749 11195 6783
rect 12817 6749 12851 6783
rect 13461 6749 13495 6783
rect 1593 6681 1627 6715
rect 2513 6681 2547 6715
rect 3065 6681 3099 6715
rect 4353 6681 4387 6715
rect 11529 6681 11563 6715
rect 13277 6681 13311 6715
rect 4077 6613 4111 6647
rect 4169 6613 4203 6647
rect 5457 6613 5491 6647
rect 6837 6613 6871 6647
rect 8033 6613 8067 6647
rect 10057 6613 10091 6647
rect 11345 6613 11379 6647
rect 1409 6409 1443 6443
rect 3157 6409 3191 6443
rect 6101 6409 6135 6443
rect 7389 6409 7423 6443
rect 8769 6409 8803 6443
rect 9137 6409 9171 6443
rect 9505 6409 9539 6443
rect 9965 6409 9999 6443
rect 11161 6409 11195 6443
rect 4077 6341 4111 6375
rect 4997 6341 5031 6375
rect 8033 6341 8067 6375
rect 8585 6341 8619 6375
rect 11897 6341 11931 6375
rect 2053 6273 2087 6307
rect 2605 6273 2639 6307
rect 2789 6273 2823 6307
rect 3341 6273 3375 6307
rect 3433 6273 3467 6307
rect 3617 6273 3651 6307
rect 3709 6273 3743 6307
rect 3893 6273 3927 6307
rect 4261 6273 4295 6307
rect 4813 6273 4847 6307
rect 5549 6273 5583 6307
rect 5825 6273 5859 6307
rect 6009 6273 6043 6307
rect 6745 6273 6779 6307
rect 7113 6273 7147 6307
rect 7297 6273 7331 6307
rect 9597 6273 9631 6307
rect 9963 6273 9997 6307
rect 11529 6273 11563 6307
rect 11713 6273 11747 6307
rect 11989 6273 12023 6307
rect 13461 6273 13495 6307
rect 2329 6205 2363 6239
rect 2881 6205 2915 6239
rect 5089 6205 5123 6239
rect 6653 6205 6687 6239
rect 7389 6205 7423 6239
rect 8861 6205 8895 6239
rect 10425 6205 10459 6239
rect 11161 6205 11195 6239
rect 11253 6205 11287 6239
rect 7021 6137 7055 6171
rect 10333 6137 10367 6171
rect 13277 6137 13311 6171
rect 4537 6069 4571 6103
rect 5733 6069 5767 6103
rect 6377 6069 6411 6103
rect 7849 6069 7883 6103
rect 8309 6069 8343 6103
rect 9781 6069 9815 6103
rect 10701 6069 10735 6103
rect 1501 5865 1535 5899
rect 2881 5865 2915 5899
rect 3801 5865 3835 5899
rect 7481 5865 7515 5899
rect 7757 5865 7791 5899
rect 11621 5865 11655 5899
rect 12173 5865 12207 5899
rect 13369 5865 13403 5899
rect 1777 5797 1811 5831
rect 2145 5797 2179 5831
rect 3525 5797 3559 5831
rect 4537 5797 4571 5831
rect 8585 5797 8619 5831
rect 7665 5729 7699 5763
rect 9873 5729 9907 5763
rect 11805 5729 11839 5763
rect 1409 5661 1443 5695
rect 1961 5661 1995 5695
rect 2237 5661 2271 5695
rect 2421 5661 2455 5695
rect 2605 5661 2639 5695
rect 2697 5661 2731 5695
rect 3065 5661 3099 5695
rect 3249 5661 3283 5695
rect 3617 5661 3651 5695
rect 4077 5661 4111 5695
rect 4261 5661 4295 5695
rect 4629 5661 4663 5695
rect 4721 5661 4755 5695
rect 4997 5639 5031 5673
rect 5181 5661 5215 5695
rect 5273 5661 5307 5695
rect 5366 5661 5400 5695
rect 5733 5661 5767 5695
rect 7941 5661 7975 5695
rect 8033 5661 8067 5695
rect 8401 5661 8435 5695
rect 8953 5661 8987 5695
rect 9793 5661 9827 5695
rect 11989 5661 12023 5695
rect 12357 5661 12391 5695
rect 13553 5661 13587 5695
rect 5641 5593 5675 5627
rect 6009 5593 6043 5627
rect 10149 5593 10183 5627
rect 13001 5593 13035 5627
rect 13277 5593 13311 5627
rect 4261 5525 4295 5559
rect 8217 5525 8251 5559
rect 9137 5525 9171 5559
rect 9597 5525 9631 5559
rect 1961 5321 1995 5355
rect 5273 5321 5307 5355
rect 7481 5321 7515 5355
rect 9505 5321 9539 5355
rect 10517 5321 10551 5355
rect 11253 5321 11287 5355
rect 13277 5321 13311 5355
rect 13553 5321 13587 5355
rect 2605 5253 2639 5287
rect 2789 5253 2823 5287
rect 3801 5253 3835 5287
rect 8033 5253 8067 5287
rect 11805 5253 11839 5287
rect 1777 5185 1811 5219
rect 2145 5185 2179 5219
rect 3433 5185 3467 5219
rect 6101 5185 6135 5219
rect 6193 5185 6227 5219
rect 6377 5185 6411 5219
rect 6653 5185 6687 5219
rect 7297 5185 7331 5219
rect 9965 5185 9999 5219
rect 10333 5185 10367 5219
rect 10701 5185 10735 5219
rect 10977 5185 11011 5219
rect 11253 5185 11287 5219
rect 11529 5185 11563 5219
rect 2881 5117 2915 5151
rect 3525 5117 3559 5151
rect 5917 5117 5951 5151
rect 7113 5117 7147 5151
rect 7757 5117 7791 5151
rect 2329 5049 2363 5083
rect 6837 5049 6871 5083
rect 9781 5049 9815 5083
rect 10241 5049 10275 5083
rect 1593 4981 1627 5015
rect 3249 4981 3283 5015
rect 5457 4981 5491 5015
rect 5733 4981 5767 5015
rect 6469 4981 6503 5015
rect 3249 4777 3283 4811
rect 4077 4777 4111 4811
rect 11345 4777 11379 4811
rect 3525 4709 3559 4743
rect 6745 4709 6779 4743
rect 7021 4709 7055 4743
rect 11805 4709 11839 4743
rect 1777 4641 1811 4675
rect 4445 4641 4479 4675
rect 8769 4641 8803 4675
rect 9597 4641 9631 4675
rect 1501 4573 1535 4607
rect 3433 4573 3467 4607
rect 4997 4573 5031 4607
rect 9137 4573 9171 4607
rect 11621 4573 11655 4607
rect 11713 4573 11747 4607
rect 11989 4573 12023 4607
rect 13277 4573 13311 4607
rect 3801 4505 3835 4539
rect 4629 4505 4663 4539
rect 4905 4505 4939 4539
rect 5273 4505 5307 4539
rect 8493 4505 8527 4539
rect 9873 4505 9907 4539
rect 13553 4505 13587 4539
rect 4537 4437 4571 4471
rect 9137 4437 9171 4471
rect 3249 4233 3283 4267
rect 6561 4233 6595 4267
rect 7021 4233 7055 4267
rect 10609 4233 10643 4267
rect 11253 4233 11287 4267
rect 4445 4165 4479 4199
rect 6377 4165 6411 4199
rect 13369 4165 13403 4199
rect 1685 4097 1719 4131
rect 2237 4097 2271 4131
rect 2881 4097 2915 4131
rect 3341 4097 3375 4131
rect 3525 4097 3559 4131
rect 3709 4097 3743 4131
rect 3893 4097 3927 4131
rect 4176 4097 4210 4131
rect 7021 4097 7055 4131
rect 7205 4097 7239 4131
rect 7665 4097 7699 4131
rect 9965 4097 9999 4131
rect 10057 4097 10091 4131
rect 10609 4097 10643 4131
rect 10793 4097 10827 4131
rect 11069 4097 11103 4131
rect 11161 4097 11195 4131
rect 11529 4097 11563 4131
rect 11989 4097 12023 4131
rect 12541 4097 12575 4131
rect 13001 4097 13035 4131
rect 1777 4029 1811 4063
rect 2053 4029 2087 4063
rect 2145 4029 2179 4063
rect 2697 4029 2731 4063
rect 3065 4029 3099 4063
rect 4077 4029 4111 4063
rect 7757 4029 7791 4063
rect 8033 4029 8067 4063
rect 9505 4029 9539 4063
rect 11897 4029 11931 4063
rect 12449 4029 12483 4063
rect 13093 4029 13127 4063
rect 2421 3961 2455 3995
rect 9781 3961 9815 3995
rect 1501 3893 1535 3927
rect 5917 3893 5951 3927
rect 6101 3893 6135 3927
rect 6561 3893 6595 3927
rect 6745 3893 6779 3927
rect 7481 3893 7515 3927
rect 10241 3893 10275 3927
rect 11713 3893 11747 3927
rect 13277 3893 13311 3927
rect 1409 3689 1443 3723
rect 1685 3689 1719 3723
rect 3525 3689 3559 3723
rect 6377 3689 6411 3723
rect 7867 3689 7901 3723
rect 12357 3689 12391 3723
rect 13369 3689 13403 3723
rect 5365 3621 5399 3655
rect 8677 3621 8711 3655
rect 9045 3621 9079 3655
rect 11437 3621 11471 3655
rect 2421 3553 2455 3587
rect 4721 3553 4755 3587
rect 5917 3553 5951 3587
rect 8125 3553 8159 3587
rect 8309 3553 8343 3587
rect 1869 3485 1903 3519
rect 2053 3485 2087 3519
rect 3157 3485 3191 3519
rect 3341 3485 3375 3519
rect 3893 3485 3927 3519
rect 5089 3485 5123 3519
rect 5365 3485 5399 3519
rect 5733 3485 5767 3519
rect 6101 3485 6135 3519
rect 8401 3485 8435 3519
rect 8585 3485 8619 3519
rect 9045 3485 9079 3519
rect 9321 3485 9355 3519
rect 9689 3485 9723 3519
rect 11621 3485 11655 3519
rect 11805 3485 11839 3519
rect 12265 3485 12299 3519
rect 12633 3485 12667 3519
rect 12725 3485 12759 3519
rect 13001 3485 13035 3519
rect 13369 3485 13403 3519
rect 2145 3417 2179 3451
rect 6009 3417 6043 3451
rect 9965 3417 9999 3451
rect 12081 3417 12115 3451
rect 9413 3349 9447 3383
rect 11713 3349 11747 3383
rect 12633 3349 12667 3383
rect 2237 3145 2271 3179
rect 4427 3145 4461 3179
rect 5825 3145 5859 3179
rect 6745 3145 6779 3179
rect 7941 3145 7975 3179
rect 13185 3145 13219 3179
rect 1777 3077 1811 3111
rect 4905 3077 4939 3111
rect 6929 3077 6963 3111
rect 12081 3077 12115 3111
rect 12173 3077 12207 3111
rect 1961 3009 1995 3043
rect 2329 3009 2363 3043
rect 4721 3009 4755 3043
rect 5549 3009 5583 3043
rect 5917 3009 5951 3043
rect 6009 3009 6043 3043
rect 6561 3009 6595 3043
rect 7021 3009 7055 3043
rect 7297 3009 7331 3043
rect 7573 3009 7607 3043
rect 7665 3009 7699 3043
rect 7941 3009 7975 3043
rect 8217 3009 8251 3043
rect 9229 3009 9263 3043
rect 11621 3009 11655 3043
rect 11897 3009 11931 3043
rect 12817 3009 12851 3043
rect 13369 3009 13403 3043
rect 1685 2941 1719 2975
rect 2421 2941 2455 2975
rect 2697 2941 2731 2975
rect 4169 2941 4203 2975
rect 4997 2941 5031 2975
rect 5365 2941 5399 2975
rect 6377 2941 6411 2975
rect 7389 2941 7423 2975
rect 9505 2941 9539 2975
rect 9781 2941 9815 2975
rect 11529 2941 11563 2975
rect 12173 2941 12207 2975
rect 6101 2873 6135 2907
rect 9321 2873 9355 2907
rect 11253 2873 11287 2907
rect 12633 2873 12667 2907
rect 5181 2805 5215 2839
rect 13001 2805 13035 2839
rect 2145 2601 2179 2635
rect 2697 2601 2731 2635
rect 3893 2601 3927 2635
rect 7481 2601 7515 2635
rect 12633 2601 12667 2635
rect 3525 2533 3559 2567
rect 4445 2465 4479 2499
rect 5733 2465 5767 2499
rect 7665 2465 7699 2499
rect 10885 2465 10919 2499
rect 12817 2465 12851 2499
rect 13369 2465 13403 2499
rect 1685 2397 1719 2431
rect 1961 2397 1995 2431
rect 2237 2397 2271 2431
rect 2421 2397 2455 2431
rect 2973 2397 3007 2431
rect 3157 2397 3191 2431
rect 3341 2397 3375 2431
rect 3433 2397 3467 2431
rect 4629 2397 4663 2431
rect 4997 2397 5031 2431
rect 5273 2397 5307 2431
rect 5641 2397 5675 2431
rect 7849 2397 7883 2431
rect 7941 2397 7975 2431
rect 8401 2397 8435 2431
rect 8677 2397 8711 2431
rect 9137 2397 9171 2431
rect 11437 2397 11471 2431
rect 11621 2397 11655 2431
rect 12449 2397 12483 2431
rect 13277 2397 13311 2431
rect 2605 2329 2639 2363
rect 4169 2329 4203 2363
rect 5089 2329 5123 2363
rect 6009 2329 6043 2363
rect 8493 2329 8527 2363
rect 9413 2329 9447 2363
rect 13001 2329 13035 2363
rect 1501 2261 1535 2295
rect 4353 2261 4387 2295
rect 4813 2261 4847 2295
rect 9045 2261 9079 2295
rect 12909 2261 12943 2295
rect 2237 2057 2271 2091
rect 4445 2057 4479 2091
rect 7297 2057 7331 2091
rect 7757 2057 7791 2091
rect 9597 2057 9631 2091
rect 1501 1989 1535 2023
rect 10333 1989 10367 2023
rect 10885 1989 10919 2023
rect 1685 1921 1719 1955
rect 1869 1921 1903 1955
rect 2145 1921 2179 1955
rect 2237 1921 2271 1955
rect 2421 1921 2455 1955
rect 6193 1921 6227 1955
rect 6561 1921 6595 1955
rect 7389 1921 7423 1955
rect 7573 1921 7607 1955
rect 7849 1921 7883 1955
rect 9873 1921 9907 1955
rect 9965 1921 9999 1955
rect 10241 1921 10275 1955
rect 10517 1921 10551 1955
rect 10793 1921 10827 1955
rect 11253 1921 11287 1955
rect 11529 1921 11563 1955
rect 2697 1853 2731 1887
rect 5917 1853 5951 1887
rect 6469 1853 6503 1887
rect 7113 1853 7147 1887
rect 8125 1853 8159 1887
rect 11805 1853 11839 1887
rect 6837 1785 6871 1819
rect 10057 1785 10091 1819
rect 11069 1785 11103 1819
rect 4169 1717 4203 1751
rect 13277 1717 13311 1751
rect 3893 1513 3927 1547
rect 6929 1513 6963 1547
rect 11161 1513 11195 1547
rect 13001 1513 13035 1547
rect 3525 1445 3559 1479
rect 1409 1377 1443 1411
rect 4997 1377 5031 1411
rect 5549 1377 5583 1411
rect 8401 1377 8435 1411
rect 8677 1377 8711 1411
rect 9413 1377 9447 1411
rect 9689 1377 9723 1411
rect 12081 1377 12115 1411
rect 12173 1377 12207 1411
rect 3157 1309 3191 1343
rect 3433 1309 3467 1343
rect 3617 1309 3651 1343
rect 4077 1309 4111 1343
rect 4169 1309 4203 1343
rect 4721 1309 4755 1343
rect 5733 1309 5767 1343
rect 5917 1309 5951 1343
rect 6561 1309 6595 1343
rect 6745 1309 6779 1343
rect 9045 1309 9079 1343
rect 9321 1309 9355 1343
rect 12651 1309 12685 1343
rect 12817 1309 12851 1343
rect 13185 1309 13219 1343
rect 6377 1241 6411 1275
rect 5917 1173 5951 1207
rect 6101 1173 6135 1207
rect 9229 1173 9263 1207
rect 11529 1173 11563 1207
rect 12173 1173 12207 1207
rect 13369 1173 13403 1207
<< metal1 >>
rect 3602 14288 3608 14340
rect 3660 14328 3666 14340
rect 10778 14328 10784 14340
rect 3660 14300 10784 14328
rect 3660 14288 3666 14300
rect 10778 14288 10784 14300
rect 10836 14288 10842 14340
rect 7834 14084 7840 14136
rect 7892 14124 7898 14136
rect 9766 14124 9772 14136
rect 7892 14096 9772 14124
rect 7892 14084 7898 14096
rect 9766 14084 9772 14096
rect 9824 14084 9830 14136
rect 2866 14016 2872 14068
rect 2924 14056 2930 14068
rect 6638 14056 6644 14068
rect 2924 14028 6644 14056
rect 2924 14016 2930 14028
rect 6638 14016 6644 14028
rect 6696 14016 6702 14068
rect 6454 13948 6460 14000
rect 6512 13988 6518 14000
rect 10410 13988 10416 14000
rect 6512 13960 10416 13988
rect 6512 13948 6518 13960
rect 10410 13948 10416 13960
rect 10468 13948 10474 14000
rect 3418 13880 3424 13932
rect 3476 13920 3482 13932
rect 7926 13920 7932 13932
rect 3476 13892 7932 13920
rect 3476 13880 3482 13892
rect 7926 13880 7932 13892
rect 7984 13880 7990 13932
rect 5350 13812 5356 13864
rect 5408 13852 5414 13864
rect 11698 13852 11704 13864
rect 5408 13824 11704 13852
rect 5408 13812 5414 13824
rect 11698 13812 11704 13824
rect 11756 13812 11762 13864
rect 5534 13744 5540 13796
rect 5592 13784 5598 13796
rect 9674 13784 9680 13796
rect 5592 13756 9680 13784
rect 5592 13744 5598 13756
rect 9674 13744 9680 13756
rect 9732 13784 9738 13796
rect 11238 13784 11244 13796
rect 9732 13756 11244 13784
rect 9732 13744 9738 13756
rect 11238 13744 11244 13756
rect 11296 13744 11302 13796
rect 6086 13676 6092 13728
rect 6144 13716 6150 13728
rect 8018 13716 8024 13728
rect 6144 13688 8024 13716
rect 6144 13676 6150 13688
rect 8018 13676 8024 13688
rect 8076 13716 8082 13728
rect 8570 13716 8576 13728
rect 8076 13688 8576 13716
rect 8076 13676 8082 13688
rect 8570 13676 8576 13688
rect 8628 13676 8634 13728
rect 9950 13676 9956 13728
rect 10008 13716 10014 13728
rect 10962 13716 10968 13728
rect 10008 13688 10968 13716
rect 10008 13676 10014 13688
rect 10962 13676 10968 13688
rect 11020 13676 11026 13728
rect 1104 13626 13892 13648
rect 1104 13574 4214 13626
rect 4266 13574 4278 13626
rect 4330 13574 4342 13626
rect 4394 13574 4406 13626
rect 4458 13574 4470 13626
rect 4522 13574 12214 13626
rect 12266 13574 12278 13626
rect 12330 13574 12342 13626
rect 12394 13574 12406 13626
rect 12458 13574 12470 13626
rect 12522 13574 13892 13626
rect 1104 13552 13892 13574
rect 3602 13512 3608 13524
rect 3563 13484 3608 13512
rect 3602 13472 3608 13484
rect 3660 13472 3666 13524
rect 4249 13515 4307 13521
rect 4249 13481 4261 13515
rect 4295 13512 4307 13515
rect 6086 13512 6092 13524
rect 4295 13484 6092 13512
rect 4295 13481 4307 13484
rect 4249 13475 4307 13481
rect 6086 13472 6092 13484
rect 6144 13472 6150 13524
rect 8665 13515 8723 13521
rect 8665 13512 8677 13515
rect 6196 13484 8677 13512
rect 5534 13444 5540 13456
rect 5495 13416 5540 13444
rect 5534 13404 5540 13416
rect 5592 13404 5598 13456
rect 2685 13379 2743 13385
rect 2685 13345 2697 13379
rect 2731 13376 2743 13379
rect 4801 13379 4859 13385
rect 2731 13348 3648 13376
rect 2731 13345 2743 13348
rect 2685 13339 2743 13345
rect 1670 13308 1676 13320
rect 1631 13280 1676 13308
rect 1670 13268 1676 13280
rect 1728 13268 1734 13320
rect 1854 13268 1860 13320
rect 1912 13308 1918 13320
rect 2225 13311 2283 13317
rect 2225 13308 2237 13311
rect 1912 13280 2237 13308
rect 1912 13268 1918 13280
rect 2225 13277 2237 13280
rect 2271 13277 2283 13311
rect 2866 13308 2872 13320
rect 2827 13280 2872 13308
rect 2225 13271 2283 13277
rect 2866 13268 2872 13280
rect 2924 13268 2930 13320
rect 3418 13308 3424 13320
rect 3379 13280 3424 13308
rect 3418 13268 3424 13280
rect 3476 13268 3482 13320
rect 1486 13240 1492 13252
rect 1447 13212 1492 13240
rect 1486 13200 1492 13212
rect 1544 13200 1550 13252
rect 1946 13240 1952 13252
rect 1907 13212 1952 13240
rect 1946 13200 1952 13212
rect 2004 13200 2010 13252
rect 2777 13243 2835 13249
rect 2777 13209 2789 13243
rect 2823 13240 2835 13243
rect 3142 13240 3148 13252
rect 2823 13212 3148 13240
rect 2823 13209 2835 13212
rect 2777 13203 2835 13209
rect 3142 13200 3148 13212
rect 3200 13200 3206 13252
rect 3326 13240 3332 13252
rect 3287 13212 3332 13240
rect 3326 13200 3332 13212
rect 3384 13200 3390 13252
rect 3620 13240 3648 13348
rect 4801 13345 4813 13379
rect 4847 13376 4859 13379
rect 5350 13376 5356 13388
rect 4847 13348 5356 13376
rect 4847 13345 4859 13348
rect 4801 13339 4859 13345
rect 5350 13336 5356 13348
rect 5408 13336 5414 13388
rect 6196 13385 6224 13484
rect 8665 13481 8677 13484
rect 8711 13481 8723 13515
rect 8665 13475 8723 13481
rect 10042 13472 10048 13524
rect 10100 13512 10106 13524
rect 10873 13515 10931 13521
rect 10873 13512 10885 13515
rect 10100 13484 10885 13512
rect 10100 13472 10106 13484
rect 10873 13481 10885 13484
rect 10919 13481 10931 13515
rect 10873 13475 10931 13481
rect 10962 13472 10968 13524
rect 11020 13512 11026 13524
rect 13449 13515 13507 13521
rect 13449 13512 13461 13515
rect 11020 13484 13461 13512
rect 11020 13472 11026 13484
rect 13449 13481 13461 13484
rect 13495 13481 13507 13515
rect 13449 13475 13507 13481
rect 7561 13447 7619 13453
rect 7561 13444 7573 13447
rect 7024 13416 7573 13444
rect 6181 13379 6239 13385
rect 6181 13345 6193 13379
rect 6227 13345 6239 13379
rect 6454 13376 6460 13388
rect 6415 13348 6460 13376
rect 6181 13339 6239 13345
rect 6454 13336 6460 13348
rect 6512 13336 6518 13388
rect 7024 13385 7052 13416
rect 7561 13413 7573 13416
rect 7607 13413 7619 13447
rect 7561 13407 7619 13413
rect 7650 13404 7656 13456
rect 7708 13444 7714 13456
rect 7929 13447 7987 13453
rect 7929 13444 7941 13447
rect 7708 13416 7941 13444
rect 7708 13404 7714 13416
rect 7929 13413 7941 13416
rect 7975 13413 7987 13447
rect 7929 13407 7987 13413
rect 9125 13447 9183 13453
rect 9125 13413 9137 13447
rect 9171 13444 9183 13447
rect 9171 13416 10732 13444
rect 9171 13413 9183 13416
rect 9125 13407 9183 13413
rect 7009 13379 7067 13385
rect 7009 13345 7021 13379
rect 7055 13345 7067 13379
rect 7009 13339 7067 13345
rect 7484 13348 8432 13376
rect 3694 13268 3700 13320
rect 3752 13308 3758 13320
rect 4341 13311 4399 13317
rect 4341 13308 4353 13311
rect 3752 13280 4353 13308
rect 3752 13268 3758 13280
rect 4341 13277 4353 13280
rect 4387 13277 4399 13311
rect 5626 13308 5632 13320
rect 5587 13280 5632 13308
rect 4341 13271 4399 13277
rect 5626 13268 5632 13280
rect 5684 13268 5690 13320
rect 6917 13311 6975 13317
rect 6917 13277 6929 13311
rect 6963 13308 6975 13311
rect 7098 13308 7104 13320
rect 6963 13280 7104 13308
rect 6963 13277 6975 13280
rect 6917 13271 6975 13277
rect 7098 13268 7104 13280
rect 7156 13308 7162 13320
rect 7484 13308 7512 13348
rect 7156 13280 7512 13308
rect 7156 13268 7162 13280
rect 7650 13268 7656 13320
rect 7708 13308 7714 13320
rect 7745 13311 7803 13317
rect 7745 13308 7757 13311
rect 7708 13280 7757 13308
rect 7708 13268 7714 13280
rect 7745 13277 7757 13280
rect 7791 13277 7803 13311
rect 7745 13271 7803 13277
rect 8018 13268 8024 13320
rect 8076 13317 8082 13320
rect 8076 13311 8119 13317
rect 8107 13277 8119 13311
rect 8294 13308 8300 13320
rect 8255 13280 8300 13308
rect 8076 13271 8119 13277
rect 8076 13268 8082 13271
rect 8294 13268 8300 13280
rect 8352 13268 8358 13320
rect 3881 13243 3939 13249
rect 3881 13240 3893 13243
rect 3620 13212 3893 13240
rect 1857 13175 1915 13181
rect 1857 13141 1869 13175
rect 1903 13172 1915 13175
rect 2038 13172 2044 13184
rect 1903 13144 2044 13172
rect 1903 13141 1915 13144
rect 1857 13135 1915 13141
rect 2038 13132 2044 13144
rect 2096 13132 2102 13184
rect 2133 13175 2191 13181
rect 2133 13141 2145 13175
rect 2179 13172 2191 13175
rect 3050 13172 3056 13184
rect 2179 13144 3056 13172
rect 2179 13141 2191 13144
rect 2133 13135 2191 13141
rect 3050 13132 3056 13144
rect 3108 13132 3114 13184
rect 3510 13132 3516 13184
rect 3568 13172 3574 13184
rect 3620 13172 3648 13212
rect 3881 13209 3893 13212
rect 3927 13209 3939 13243
rect 4062 13240 4068 13252
rect 4023 13212 4068 13240
rect 3881 13203 3939 13209
rect 4062 13200 4068 13212
rect 4120 13200 4126 13252
rect 4890 13200 4896 13252
rect 4948 13240 4954 13252
rect 4948 13212 4993 13240
rect 4948 13200 4954 13212
rect 5258 13200 5264 13252
rect 5316 13240 5322 13252
rect 5353 13243 5411 13249
rect 5353 13240 5365 13243
rect 5316 13212 5365 13240
rect 5316 13200 5322 13212
rect 5353 13209 5365 13212
rect 5399 13209 5411 13243
rect 5353 13203 5411 13209
rect 5810 13200 5816 13252
rect 5868 13240 5874 13252
rect 6089 13243 6147 13249
rect 6089 13240 6101 13243
rect 5868 13212 6101 13240
rect 5868 13200 5874 13212
rect 6089 13209 6101 13212
rect 6135 13209 6147 13243
rect 6089 13203 6147 13209
rect 7377 13243 7435 13249
rect 7377 13209 7389 13243
rect 7423 13240 7435 13243
rect 8202 13240 8208 13252
rect 7423 13212 8064 13240
rect 8163 13212 8208 13240
rect 7423 13209 7435 13212
rect 7377 13203 7435 13209
rect 3568 13144 3648 13172
rect 3568 13132 3574 13144
rect 4614 13132 4620 13184
rect 4672 13172 4678 13184
rect 4985 13175 5043 13181
rect 4985 13172 4997 13175
rect 4672 13144 4997 13172
rect 4672 13132 4678 13144
rect 4985 13141 4997 13144
rect 5031 13141 5043 13175
rect 4985 13135 5043 13141
rect 5074 13132 5080 13184
rect 5132 13172 5138 13184
rect 7282 13172 7288 13184
rect 5132 13144 5177 13172
rect 7243 13144 7288 13172
rect 5132 13132 5138 13144
rect 7282 13132 7288 13144
rect 7340 13172 7346 13184
rect 7650 13172 7656 13184
rect 7340 13144 7656 13172
rect 7340 13132 7346 13144
rect 7650 13132 7656 13144
rect 7708 13132 7714 13184
rect 8036 13172 8064 13212
rect 8202 13200 8208 13212
rect 8260 13200 8266 13252
rect 8404 13240 8432 13348
rect 9858 13336 9864 13388
rect 9916 13376 9922 13388
rect 9953 13379 10011 13385
rect 9953 13376 9965 13379
rect 9916 13348 9965 13376
rect 9916 13336 9922 13348
rect 9953 13345 9965 13348
rect 9999 13345 10011 13379
rect 10704 13376 10732 13416
rect 11974 13404 11980 13456
rect 12032 13444 12038 13456
rect 12621 13447 12679 13453
rect 12621 13444 12633 13447
rect 12032 13416 12633 13444
rect 12032 13404 12038 13416
rect 12621 13413 12633 13416
rect 12667 13413 12679 13447
rect 12621 13407 12679 13413
rect 12161 13379 12219 13385
rect 12161 13376 12173 13379
rect 10704 13348 12173 13376
rect 9953 13339 10011 13345
rect 12161 13345 12173 13348
rect 12207 13345 12219 13379
rect 12161 13339 12219 13345
rect 8478 13268 8484 13320
rect 8536 13308 8542 13320
rect 8536 13280 8581 13308
rect 8536 13268 8542 13280
rect 8754 13268 8760 13320
rect 8812 13308 8818 13320
rect 9309 13311 9367 13317
rect 9309 13308 9321 13311
rect 8812 13280 9321 13308
rect 8812 13268 8818 13280
rect 9309 13277 9321 13280
rect 9355 13277 9367 13311
rect 10686 13308 10692 13320
rect 10647 13280 10692 13308
rect 9309 13271 9367 13277
rect 10686 13268 10692 13280
rect 10744 13268 10750 13320
rect 10962 13308 10968 13320
rect 10923 13280 10968 13308
rect 10962 13268 10968 13280
rect 11020 13268 11026 13320
rect 11238 13308 11244 13320
rect 11199 13280 11244 13308
rect 11238 13268 11244 13280
rect 11296 13268 11302 13320
rect 11514 13268 11520 13320
rect 11572 13308 11578 13320
rect 11609 13311 11667 13317
rect 11609 13308 11621 13311
rect 11572 13280 11621 13308
rect 11572 13268 11578 13280
rect 11609 13277 11621 13280
rect 11655 13277 11667 13311
rect 11609 13271 11667 13277
rect 11698 13268 11704 13320
rect 11756 13308 11762 13320
rect 12345 13311 12403 13317
rect 12345 13308 12357 13311
rect 11756 13280 12357 13308
rect 11756 13268 11762 13280
rect 12345 13277 12357 13280
rect 12391 13277 12403 13311
rect 12345 13271 12403 13277
rect 12805 13311 12863 13317
rect 12805 13277 12817 13311
rect 12851 13277 12863 13311
rect 12805 13271 12863 13277
rect 12897 13311 12955 13317
rect 12897 13277 12909 13311
rect 12943 13277 12955 13311
rect 12897 13271 12955 13277
rect 13173 13311 13231 13317
rect 13173 13277 13185 13311
rect 13219 13308 13231 13311
rect 13446 13308 13452 13320
rect 13219 13280 13452 13308
rect 13219 13277 13231 13280
rect 13173 13271 13231 13277
rect 8573 13243 8631 13249
rect 8573 13240 8585 13243
rect 8404 13212 8585 13240
rect 8573 13209 8585 13212
rect 8619 13209 8631 13243
rect 9766 13240 9772 13252
rect 8573 13203 8631 13209
rect 9048 13212 9772 13240
rect 9048 13172 9076 13212
rect 9766 13200 9772 13212
rect 9824 13200 9830 13252
rect 9861 13243 9919 13249
rect 9861 13209 9873 13243
rect 9907 13240 9919 13243
rect 10134 13240 10140 13252
rect 9907 13212 10140 13240
rect 9907 13209 9919 13212
rect 9861 13203 9919 13209
rect 10134 13200 10140 13212
rect 10192 13200 10198 13252
rect 10226 13200 10232 13252
rect 10284 13240 10290 13252
rect 10413 13243 10471 13249
rect 10413 13240 10425 13243
rect 10284 13212 10425 13240
rect 10284 13200 10290 13212
rect 10413 13209 10425 13212
rect 10459 13209 10471 13243
rect 10413 13203 10471 13209
rect 10505 13243 10563 13249
rect 10505 13209 10517 13243
rect 10551 13209 10563 13243
rect 12066 13240 12072 13252
rect 12027 13212 12072 13240
rect 10505 13203 10563 13209
rect 9214 13172 9220 13184
rect 8036 13144 9076 13172
rect 9175 13144 9220 13172
rect 9214 13132 9220 13144
rect 9272 13132 9278 13184
rect 10520 13172 10548 13203
rect 12066 13200 12072 13212
rect 12124 13200 12130 13252
rect 11057 13175 11115 13181
rect 11057 13172 11069 13175
rect 10520 13144 11069 13172
rect 11057 13141 11069 13144
rect 11103 13141 11115 13175
rect 11057 13135 11115 13141
rect 11882 13132 11888 13184
rect 11940 13172 11946 13184
rect 12437 13175 12495 13181
rect 12437 13172 12449 13175
rect 11940 13144 12449 13172
rect 11940 13132 11946 13144
rect 12437 13141 12449 13144
rect 12483 13172 12495 13175
rect 12820 13172 12848 13271
rect 12912 13240 12940 13271
rect 13446 13268 13452 13280
rect 13504 13268 13510 13320
rect 13262 13240 13268 13252
rect 12912 13212 13268 13240
rect 13262 13200 13268 13212
rect 13320 13200 13326 13252
rect 13078 13172 13084 13184
rect 12483 13144 12848 13172
rect 13039 13144 13084 13172
rect 12483 13141 12495 13144
rect 12437 13135 12495 13141
rect 13078 13132 13084 13144
rect 13136 13132 13142 13184
rect 13354 13172 13360 13184
rect 13315 13144 13360 13172
rect 13354 13132 13360 13144
rect 13412 13132 13418 13184
rect 1104 13082 13892 13104
rect 1104 13030 8214 13082
rect 8266 13030 8278 13082
rect 8330 13030 8342 13082
rect 8394 13030 8406 13082
rect 8458 13030 8470 13082
rect 8522 13030 13892 13082
rect 1104 13008 13892 13030
rect 1762 12928 1768 12980
rect 1820 12968 1826 12980
rect 2958 12968 2964 12980
rect 1820 12940 2964 12968
rect 1820 12928 1826 12940
rect 2958 12928 2964 12940
rect 3016 12928 3022 12980
rect 3050 12928 3056 12980
rect 3108 12968 3114 12980
rect 3878 12968 3884 12980
rect 3108 12940 3884 12968
rect 3108 12928 3114 12940
rect 3878 12928 3884 12940
rect 3936 12928 3942 12980
rect 4982 12928 4988 12980
rect 5040 12968 5046 12980
rect 7466 12968 7472 12980
rect 5040 12940 7472 12968
rect 5040 12928 5046 12940
rect 7466 12928 7472 12940
rect 7524 12928 7530 12980
rect 9214 12928 9220 12980
rect 9272 12968 9278 12980
rect 11606 12968 11612 12980
rect 9272 12940 11612 12968
rect 9272 12928 9278 12940
rect 11606 12928 11612 12940
rect 11664 12928 11670 12980
rect 3421 12903 3479 12909
rect 3421 12869 3433 12903
rect 3467 12900 3479 12903
rect 3510 12900 3516 12912
rect 3467 12872 3516 12900
rect 3467 12869 3479 12872
rect 3421 12863 3479 12869
rect 3510 12860 3516 12872
rect 3568 12860 3574 12912
rect 5261 12903 5319 12909
rect 5261 12869 5273 12903
rect 5307 12900 5319 12903
rect 5350 12900 5356 12912
rect 5307 12872 5356 12900
rect 5307 12869 5319 12872
rect 5261 12863 5319 12869
rect 5350 12860 5356 12872
rect 5408 12860 5414 12912
rect 5626 12900 5632 12912
rect 5587 12872 5632 12900
rect 5626 12860 5632 12872
rect 5684 12860 5690 12912
rect 7098 12900 7104 12912
rect 7059 12872 7104 12900
rect 7098 12860 7104 12872
rect 7156 12860 7162 12912
rect 7282 12900 7288 12912
rect 7243 12872 7288 12900
rect 7282 12860 7288 12872
rect 7340 12860 7346 12912
rect 7561 12903 7619 12909
rect 7561 12869 7573 12903
rect 7607 12900 7619 12903
rect 8481 12903 8539 12909
rect 8481 12900 8493 12903
rect 7607 12872 8493 12900
rect 7607 12869 7619 12872
rect 7561 12863 7619 12869
rect 8481 12869 8493 12872
rect 8527 12900 8539 12903
rect 8938 12900 8944 12912
rect 8527 12872 8944 12900
rect 8527 12869 8539 12872
rect 8481 12863 8539 12869
rect 1581 12835 1639 12841
rect 1581 12801 1593 12835
rect 1627 12832 1639 12835
rect 1670 12832 1676 12844
rect 1627 12804 1676 12832
rect 1627 12801 1639 12804
rect 1581 12795 1639 12801
rect 1670 12792 1676 12804
rect 1728 12792 1734 12844
rect 1854 12832 1860 12844
rect 1815 12804 1860 12832
rect 1854 12792 1860 12804
rect 1912 12792 1918 12844
rect 3329 12835 3387 12841
rect 3329 12801 3341 12835
rect 3375 12801 3387 12835
rect 3694 12832 3700 12844
rect 3655 12804 3700 12832
rect 3329 12795 3387 12801
rect 1762 12764 1768 12776
rect 1675 12736 1768 12764
rect 1762 12724 1768 12736
rect 1820 12764 1826 12776
rect 3344 12764 3372 12795
rect 3694 12792 3700 12804
rect 3752 12792 3758 12844
rect 4062 12832 4068 12844
rect 3804 12804 4068 12832
rect 3804 12776 3832 12804
rect 4062 12792 4068 12804
rect 4120 12832 4126 12844
rect 4617 12835 4675 12841
rect 4617 12832 4629 12835
rect 4120 12804 4629 12832
rect 4120 12792 4126 12804
rect 4617 12801 4629 12804
rect 4663 12801 4675 12835
rect 4617 12795 4675 12801
rect 5813 12835 5871 12841
rect 5813 12801 5825 12835
rect 5859 12801 5871 12835
rect 5813 12795 5871 12801
rect 1820 12736 3372 12764
rect 1820 12724 1826 12736
rect 3344 12696 3372 12736
rect 3786 12724 3792 12776
rect 3844 12724 3850 12776
rect 5828 12764 5856 12795
rect 5902 12792 5908 12844
rect 5960 12832 5966 12844
rect 5997 12835 6055 12841
rect 5997 12832 6009 12835
rect 5960 12804 6009 12832
rect 5960 12792 5966 12804
rect 5997 12801 6009 12804
rect 6043 12801 6055 12835
rect 5997 12795 6055 12801
rect 6086 12792 6092 12844
rect 6144 12832 6150 12844
rect 6365 12835 6423 12841
rect 6144 12804 6189 12832
rect 6144 12792 6150 12804
rect 6365 12801 6377 12835
rect 6411 12832 6423 12835
rect 6454 12832 6460 12844
rect 6411 12804 6460 12832
rect 6411 12801 6423 12804
rect 6365 12795 6423 12801
rect 6454 12792 6460 12804
rect 6512 12792 6518 12844
rect 6546 12764 6552 12776
rect 5828 12736 6552 12764
rect 6546 12724 6552 12736
rect 6604 12724 6610 12776
rect 7006 12724 7012 12776
rect 7064 12764 7070 12776
rect 7576 12764 7604 12863
rect 8938 12860 8944 12872
rect 8996 12860 9002 12912
rect 10226 12860 10232 12912
rect 10284 12900 10290 12912
rect 11057 12903 11115 12909
rect 11057 12900 11069 12903
rect 10284 12872 11069 12900
rect 10284 12860 10290 12872
rect 11057 12869 11069 12872
rect 11103 12869 11115 12903
rect 11057 12863 11115 12869
rect 11238 12860 11244 12912
rect 11296 12900 11302 12912
rect 11333 12903 11391 12909
rect 11333 12900 11345 12903
rect 11296 12872 11345 12900
rect 11296 12860 11302 12872
rect 11333 12869 11345 12872
rect 11379 12869 11391 12903
rect 11333 12863 11391 12869
rect 12066 12860 12072 12912
rect 12124 12900 12130 12912
rect 13081 12903 13139 12909
rect 13081 12900 13093 12903
rect 12124 12872 13093 12900
rect 12124 12860 12130 12872
rect 13081 12869 13093 12872
rect 13127 12900 13139 12903
rect 13357 12903 13415 12909
rect 13357 12900 13369 12903
rect 13127 12872 13369 12900
rect 13127 12869 13139 12872
rect 13081 12863 13139 12869
rect 13357 12869 13369 12872
rect 13403 12869 13415 12903
rect 13357 12863 13415 12869
rect 7650 12792 7656 12844
rect 7708 12832 7714 12844
rect 7745 12835 7803 12841
rect 7745 12832 7757 12835
rect 7708 12804 7757 12832
rect 7708 12792 7714 12804
rect 7745 12801 7757 12804
rect 7791 12801 7803 12835
rect 8292 12835 8350 12841
rect 8292 12832 8304 12835
rect 7745 12795 7803 12801
rect 7852 12804 8304 12832
rect 7064 12736 7604 12764
rect 7064 12724 7070 12736
rect 3970 12696 3976 12708
rect 3344 12668 3976 12696
rect 3970 12656 3976 12668
rect 4028 12656 4034 12708
rect 5445 12699 5503 12705
rect 5445 12665 5457 12699
rect 5491 12696 5503 12699
rect 7852 12696 7880 12804
rect 8292 12801 8304 12804
rect 8338 12801 8350 12835
rect 8292 12795 8350 12801
rect 7929 12767 7987 12773
rect 7929 12733 7941 12767
rect 7975 12733 7987 12767
rect 8312 12764 8340 12795
rect 8386 12792 8392 12844
rect 8444 12832 8450 12844
rect 8444 12804 8489 12832
rect 8444 12792 8450 12804
rect 8570 12792 8576 12844
rect 8628 12832 8634 12844
rect 8665 12835 8723 12841
rect 8665 12832 8677 12835
rect 8628 12804 8677 12832
rect 8628 12792 8634 12804
rect 8665 12801 8677 12804
rect 8711 12801 8723 12835
rect 8665 12795 8723 12801
rect 8754 12792 8760 12844
rect 8812 12832 8818 12844
rect 8812 12804 8857 12832
rect 8812 12792 8818 12804
rect 9674 12792 9680 12844
rect 9732 12832 9738 12844
rect 9732 12804 9777 12832
rect 9732 12792 9738 12804
rect 9858 12792 9864 12844
rect 9916 12832 9922 12844
rect 10413 12835 10471 12841
rect 10413 12832 10425 12835
rect 9916 12804 10425 12832
rect 9916 12792 9922 12804
rect 10413 12801 10425 12804
rect 10459 12801 10471 12835
rect 11514 12832 11520 12844
rect 11475 12804 11520 12832
rect 10413 12795 10471 12801
rect 11514 12792 11520 12804
rect 11572 12792 11578 12844
rect 11882 12792 11888 12844
rect 11940 12832 11946 12844
rect 12437 12835 12495 12841
rect 12437 12832 12449 12835
rect 11940 12804 12449 12832
rect 11940 12792 11946 12804
rect 12437 12801 12449 12804
rect 12483 12801 12495 12835
rect 12437 12795 12495 12801
rect 8312 12736 12434 12764
rect 7929 12727 7987 12733
rect 5491 12668 7880 12696
rect 7944 12696 7972 12727
rect 8570 12696 8576 12708
rect 7944 12668 8576 12696
rect 5491 12665 5503 12668
rect 5445 12659 5503 12665
rect 8570 12656 8576 12668
rect 8628 12656 8634 12708
rect 9766 12656 9772 12708
rect 9824 12696 9830 12708
rect 10045 12699 10103 12705
rect 10045 12696 10057 12699
rect 9824 12668 10057 12696
rect 9824 12656 9830 12668
rect 10045 12665 10057 12668
rect 10091 12665 10103 12699
rect 12406 12696 12434 12736
rect 14366 12696 14372 12708
rect 12406 12668 14372 12696
rect 10045 12659 10103 12665
rect 14366 12656 14372 12668
rect 14424 12656 14430 12708
rect 2958 12588 2964 12640
rect 3016 12628 3022 12640
rect 3605 12631 3663 12637
rect 3605 12628 3617 12631
rect 3016 12600 3617 12628
rect 3016 12588 3022 12600
rect 3605 12597 3617 12600
rect 3651 12628 3663 12631
rect 7098 12628 7104 12640
rect 3651 12600 7104 12628
rect 3651 12597 3663 12600
rect 3605 12591 3663 12597
rect 7098 12588 7104 12600
rect 7156 12588 7162 12640
rect 7190 12588 7196 12640
rect 7248 12628 7254 12640
rect 8113 12631 8171 12637
rect 8113 12628 8125 12631
rect 7248 12600 8125 12628
rect 7248 12588 7254 12600
rect 8113 12597 8125 12600
rect 8159 12597 8171 12631
rect 8113 12591 8171 12597
rect 8294 12588 8300 12640
rect 8352 12628 8358 12640
rect 9582 12628 9588 12640
rect 8352 12600 9588 12628
rect 8352 12588 8358 12600
rect 9582 12588 9588 12600
rect 9640 12588 9646 12640
rect 13262 12628 13268 12640
rect 13223 12600 13268 12628
rect 13262 12588 13268 12600
rect 13320 12588 13326 12640
rect 1104 12538 13892 12560
rect 1104 12486 4214 12538
rect 4266 12486 4278 12538
rect 4330 12486 4342 12538
rect 4394 12486 4406 12538
rect 4458 12486 4470 12538
rect 4522 12486 12214 12538
rect 12266 12486 12278 12538
rect 12330 12486 12342 12538
rect 12394 12486 12406 12538
rect 12458 12486 12470 12538
rect 12522 12486 13892 12538
rect 1104 12464 13892 12486
rect 3326 12424 3332 12436
rect 2056 12396 3332 12424
rect 1762 12220 1768 12232
rect 1723 12192 1768 12220
rect 1762 12180 1768 12192
rect 1820 12180 1826 12232
rect 2056 12229 2084 12396
rect 3326 12384 3332 12396
rect 3384 12384 3390 12436
rect 4154 12384 4160 12436
rect 4212 12424 4218 12436
rect 4893 12427 4951 12433
rect 4893 12424 4905 12427
rect 4212 12396 4905 12424
rect 4212 12384 4218 12396
rect 4893 12393 4905 12396
rect 4939 12424 4951 12427
rect 5350 12424 5356 12436
rect 4939 12396 5356 12424
rect 4939 12393 4951 12396
rect 4893 12387 4951 12393
rect 5350 12384 5356 12396
rect 5408 12424 5414 12436
rect 5902 12424 5908 12436
rect 5408 12396 5908 12424
rect 5408 12384 5414 12396
rect 5902 12384 5908 12396
rect 5960 12384 5966 12436
rect 5994 12384 6000 12436
rect 6052 12424 6058 12436
rect 7006 12424 7012 12436
rect 6052 12396 7012 12424
rect 6052 12384 6058 12396
rect 7006 12384 7012 12396
rect 7064 12384 7070 12436
rect 7193 12427 7251 12433
rect 7193 12393 7205 12427
rect 7239 12424 7251 12427
rect 9858 12424 9864 12436
rect 7239 12396 9720 12424
rect 9819 12396 9864 12424
rect 7239 12393 7251 12396
rect 7193 12387 7251 12393
rect 2961 12359 3019 12365
rect 2961 12325 2973 12359
rect 3007 12356 3019 12359
rect 3602 12356 3608 12368
rect 3007 12328 3608 12356
rect 3007 12325 3019 12328
rect 2961 12319 3019 12325
rect 3602 12316 3608 12328
rect 3660 12316 3666 12368
rect 5166 12356 5172 12368
rect 5127 12328 5172 12356
rect 5166 12316 5172 12328
rect 5224 12316 5230 12368
rect 5810 12316 5816 12368
rect 5868 12356 5874 12368
rect 6641 12359 6699 12365
rect 6641 12356 6653 12359
rect 5868 12328 6653 12356
rect 5868 12316 5874 12328
rect 6641 12325 6653 12328
rect 6687 12325 6699 12359
rect 6641 12319 6699 12325
rect 7282 12316 7288 12368
rect 7340 12316 7346 12368
rect 7374 12316 7380 12368
rect 7432 12316 7438 12368
rect 7466 12316 7472 12368
rect 7524 12356 7530 12368
rect 8202 12356 8208 12368
rect 7524 12328 8208 12356
rect 7524 12316 7530 12328
rect 8202 12316 8208 12328
rect 8260 12316 8266 12368
rect 8846 12316 8852 12368
rect 8904 12356 8910 12368
rect 9030 12356 9036 12368
rect 8904 12328 9036 12356
rect 8904 12316 8910 12328
rect 9030 12316 9036 12328
rect 9088 12316 9094 12368
rect 9692 12356 9720 12396
rect 9858 12384 9864 12396
rect 9916 12384 9922 12436
rect 10134 12424 10140 12436
rect 10095 12396 10140 12424
rect 10134 12384 10140 12396
rect 10192 12384 10198 12436
rect 10410 12424 10416 12436
rect 10371 12396 10416 12424
rect 10410 12384 10416 12396
rect 10468 12384 10474 12436
rect 11514 12356 11520 12368
rect 9692 12328 11520 12356
rect 11514 12316 11520 12328
rect 11572 12316 11578 12368
rect 2332 12260 2820 12288
rect 2041 12223 2099 12229
rect 2041 12189 2053 12223
rect 2087 12189 2099 12223
rect 2041 12183 2099 12189
rect 2332 12164 2360 12260
rect 2682 12220 2688 12232
rect 2643 12192 2688 12220
rect 2682 12180 2688 12192
rect 2740 12180 2746 12232
rect 2792 12229 2820 12260
rect 3050 12248 3056 12300
rect 3108 12288 3114 12300
rect 6178 12288 6184 12300
rect 3108 12260 6184 12288
rect 3108 12248 3114 12260
rect 6178 12248 6184 12260
rect 6236 12248 6242 12300
rect 7300 12288 7328 12316
rect 6840 12260 7328 12288
rect 7392 12288 7420 12316
rect 7392 12260 8156 12288
rect 2777 12223 2835 12229
rect 2777 12189 2789 12223
rect 2823 12189 2835 12223
rect 2777 12183 2835 12189
rect 3605 12223 3663 12229
rect 3605 12189 3617 12223
rect 3651 12220 3663 12223
rect 4709 12223 4767 12229
rect 4709 12220 4721 12223
rect 3651 12192 4721 12220
rect 3651 12189 3663 12192
rect 3605 12183 3663 12189
rect 4709 12189 4721 12192
rect 4755 12220 4767 12223
rect 4798 12220 4804 12232
rect 4755 12192 4804 12220
rect 4755 12189 4767 12192
rect 4709 12183 4767 12189
rect 4798 12180 4804 12192
rect 4856 12180 4862 12232
rect 5077 12223 5135 12229
rect 5077 12189 5089 12223
rect 5123 12189 5135 12223
rect 5077 12183 5135 12189
rect 5353 12223 5411 12229
rect 5353 12189 5365 12223
rect 5399 12220 5411 12223
rect 5626 12220 5632 12232
rect 5399 12192 5632 12220
rect 5399 12189 5411 12192
rect 5353 12183 5411 12189
rect 1489 12155 1547 12161
rect 1489 12121 1501 12155
rect 1535 12121 1547 12155
rect 1489 12115 1547 12121
rect 1673 12155 1731 12161
rect 1673 12121 1685 12155
rect 1719 12152 1731 12155
rect 2314 12152 2320 12164
rect 1719 12124 2320 12152
rect 1719 12121 1731 12124
rect 1673 12115 1731 12121
rect 1504 12084 1532 12115
rect 2314 12112 2320 12124
rect 2372 12112 2378 12164
rect 3053 12155 3111 12161
rect 3053 12152 3065 12155
rect 2792 12124 3065 12152
rect 2792 12096 2820 12124
rect 3053 12121 3065 12124
rect 3099 12121 3111 12155
rect 3053 12115 3111 12121
rect 3145 12155 3203 12161
rect 3145 12121 3157 12155
rect 3191 12121 3203 12155
rect 3145 12115 3203 12121
rect 2498 12084 2504 12096
rect 1504 12056 2504 12084
rect 2498 12044 2504 12056
rect 2556 12044 2562 12096
rect 2774 12044 2780 12096
rect 2832 12044 2838 12096
rect 3160 12084 3188 12115
rect 3326 12112 3332 12164
rect 3384 12152 3390 12164
rect 3786 12152 3792 12164
rect 3384 12124 3792 12152
rect 3384 12112 3390 12124
rect 3786 12112 3792 12124
rect 3844 12112 3850 12164
rect 4062 12152 4068 12164
rect 4023 12124 4068 12152
rect 4062 12112 4068 12124
rect 4120 12112 4126 12164
rect 4522 12112 4528 12164
rect 4580 12152 4586 12164
rect 5092 12152 5120 12183
rect 5626 12180 5632 12192
rect 5684 12180 5690 12232
rect 6840 12229 6868 12260
rect 6825 12223 6883 12229
rect 6825 12189 6837 12223
rect 6871 12189 6883 12223
rect 6825 12183 6883 12189
rect 7098 12180 7104 12232
rect 7156 12220 7162 12232
rect 7325 12223 7383 12229
rect 7325 12220 7337 12223
rect 7156 12192 7337 12220
rect 7156 12180 7162 12192
rect 7325 12189 7337 12192
rect 7371 12189 7383 12223
rect 7466 12220 7472 12232
rect 7427 12192 7472 12220
rect 7325 12183 7383 12189
rect 7466 12180 7472 12192
rect 7524 12180 7530 12232
rect 7745 12223 7803 12229
rect 7745 12189 7757 12223
rect 7791 12220 7803 12223
rect 7837 12223 7895 12229
rect 7837 12220 7849 12223
rect 7791 12192 7849 12220
rect 7791 12189 7803 12192
rect 7745 12183 7803 12189
rect 7837 12189 7849 12192
rect 7883 12220 7895 12223
rect 7926 12220 7932 12232
rect 7883 12192 7932 12220
rect 7883 12189 7895 12192
rect 7837 12183 7895 12189
rect 7926 12180 7932 12192
rect 7984 12180 7990 12232
rect 8128 12229 8156 12260
rect 8478 12248 8484 12300
rect 8536 12288 8542 12300
rect 8536 12260 8984 12288
rect 8536 12248 8542 12260
rect 8206 12233 8264 12239
rect 8206 12232 8218 12233
rect 8252 12232 8264 12233
rect 8021 12223 8079 12229
rect 8021 12189 8033 12223
rect 8067 12189 8079 12223
rect 8021 12183 8079 12189
rect 8113 12223 8171 12229
rect 8113 12189 8125 12223
rect 8159 12189 8171 12223
rect 8113 12183 8171 12189
rect 4580 12124 5120 12152
rect 4580 12112 4586 12124
rect 5166 12112 5172 12164
rect 5224 12152 5230 12164
rect 7006 12152 7012 12164
rect 5224 12124 7012 12152
rect 5224 12112 5230 12124
rect 7006 12112 7012 12124
rect 7064 12112 7070 12164
rect 7561 12155 7619 12161
rect 7561 12121 7573 12155
rect 7607 12152 7619 12155
rect 7650 12152 7656 12164
rect 7607 12124 7656 12152
rect 7607 12121 7619 12124
rect 7561 12115 7619 12121
rect 4080 12084 4108 12112
rect 3160 12056 4108 12084
rect 6546 12044 6552 12096
rect 6604 12084 6610 12096
rect 7576 12084 7604 12115
rect 7650 12112 7656 12124
rect 7708 12152 7714 12164
rect 8036 12152 8064 12183
rect 8202 12180 8208 12232
rect 8260 12230 8266 12232
rect 8260 12202 8295 12230
rect 8260 12180 8266 12202
rect 8662 12180 8668 12232
rect 8720 12220 8726 12232
rect 8757 12223 8815 12229
rect 8757 12220 8769 12223
rect 8720 12192 8769 12220
rect 8720 12180 8726 12192
rect 8757 12189 8769 12192
rect 8803 12189 8815 12223
rect 8757 12183 8815 12189
rect 8846 12180 8852 12232
rect 8904 12180 8910 12232
rect 7708 12124 8064 12152
rect 8481 12155 8539 12161
rect 7708 12112 7714 12124
rect 8481 12121 8493 12155
rect 8527 12152 8539 12155
rect 8864 12152 8892 12180
rect 8527 12124 8892 12152
rect 8956 12152 8984 12260
rect 9122 12248 9128 12300
rect 9180 12254 9186 12300
rect 10042 12288 10048 12300
rect 9508 12260 10048 12288
rect 9180 12248 9260 12254
rect 9140 12229 9260 12248
rect 9140 12226 9275 12229
rect 9217 12223 9275 12226
rect 9217 12189 9229 12223
rect 9263 12189 9275 12223
rect 9217 12183 9275 12189
rect 9309 12223 9367 12229
rect 9309 12189 9321 12223
rect 9355 12220 9367 12223
rect 9398 12220 9404 12232
rect 9355 12192 9404 12220
rect 9355 12189 9367 12192
rect 9309 12183 9367 12189
rect 9398 12180 9404 12192
rect 9456 12180 9462 12232
rect 9508 12161 9536 12260
rect 10042 12248 10048 12260
rect 10100 12248 10106 12300
rect 10134 12248 10140 12300
rect 10192 12288 10198 12300
rect 13170 12288 13176 12300
rect 10192 12260 13176 12288
rect 10192 12248 10198 12260
rect 13170 12248 13176 12260
rect 13228 12248 13234 12300
rect 9729 12223 9787 12229
rect 9729 12189 9741 12223
rect 9775 12220 9787 12223
rect 9950 12220 9956 12232
rect 9775 12192 9956 12220
rect 9775 12189 9787 12192
rect 9729 12183 9787 12189
rect 9950 12180 9956 12192
rect 10008 12180 10014 12232
rect 10226 12220 10232 12232
rect 10187 12192 10232 12220
rect 10226 12180 10232 12192
rect 10284 12180 10290 12232
rect 10594 12220 10600 12232
rect 10555 12192 10600 12220
rect 10594 12180 10600 12192
rect 10652 12180 10658 12232
rect 10778 12180 10784 12232
rect 10836 12220 10842 12232
rect 10873 12223 10931 12229
rect 10873 12220 10885 12223
rect 10836 12192 10885 12220
rect 10836 12180 10842 12192
rect 10873 12189 10885 12192
rect 10919 12189 10931 12223
rect 10873 12183 10931 12189
rect 10965 12223 11023 12229
rect 10965 12189 10977 12223
rect 11011 12220 11023 12223
rect 11514 12220 11520 12232
rect 11011 12192 11520 12220
rect 11011 12189 11023 12192
rect 10965 12183 11023 12189
rect 11514 12180 11520 12192
rect 11572 12180 11578 12232
rect 11606 12180 11612 12232
rect 11664 12220 11670 12232
rect 11882 12220 11888 12232
rect 11664 12192 11709 12220
rect 11843 12192 11888 12220
rect 11664 12180 11670 12192
rect 11882 12180 11888 12192
rect 11940 12180 11946 12232
rect 11977 12223 12035 12229
rect 11977 12189 11989 12223
rect 12023 12189 12035 12223
rect 13262 12220 13268 12232
rect 13223 12192 13268 12220
rect 11977 12183 12035 12189
rect 9493 12155 9551 12161
rect 8956 12124 9444 12152
rect 8527 12121 8539 12124
rect 8481 12115 8539 12121
rect 6604 12056 7604 12084
rect 6604 12044 6610 12056
rect 7742 12044 7748 12096
rect 7800 12084 7806 12096
rect 8665 12087 8723 12093
rect 8665 12084 8677 12087
rect 7800 12056 8677 12084
rect 7800 12044 7806 12056
rect 8665 12053 8677 12056
rect 8711 12053 8723 12087
rect 8665 12047 8723 12053
rect 8846 12044 8852 12096
rect 8904 12084 8910 12096
rect 8956 12084 8984 12124
rect 9122 12084 9128 12096
rect 8904 12056 8984 12084
rect 9083 12056 9128 12084
rect 8904 12044 8910 12056
rect 9122 12044 9128 12056
rect 9180 12044 9186 12096
rect 9416 12084 9444 12124
rect 9493 12121 9505 12155
rect 9539 12121 9551 12155
rect 9493 12115 9551 12121
rect 9582 12112 9588 12164
rect 9640 12152 9646 12164
rect 9640 12124 9685 12152
rect 9640 12112 9646 12124
rect 10042 12112 10048 12164
rect 10100 12152 10106 12164
rect 10100 12124 10824 12152
rect 10100 12112 10106 12124
rect 10502 12084 10508 12096
rect 9416 12056 10508 12084
rect 10502 12044 10508 12056
rect 10560 12044 10566 12096
rect 10796 12093 10824 12124
rect 11330 12112 11336 12164
rect 11388 12152 11394 12164
rect 11992 12152 12020 12183
rect 13262 12180 13268 12192
rect 13320 12180 13326 12232
rect 11388 12124 12020 12152
rect 13541 12155 13599 12161
rect 11388 12112 11394 12124
rect 13541 12121 13553 12155
rect 13587 12152 13599 12155
rect 13587 12124 13952 12152
rect 13587 12121 13599 12124
rect 13541 12115 13599 12121
rect 10781 12087 10839 12093
rect 10781 12053 10793 12087
rect 10827 12084 10839 12087
rect 11882 12084 11888 12096
rect 10827 12056 11888 12084
rect 10827 12053 10839 12056
rect 10781 12047 10839 12053
rect 11882 12044 11888 12056
rect 11940 12044 11946 12096
rect 1104 11994 13892 12016
rect 1104 11942 8214 11994
rect 8266 11942 8278 11994
rect 8330 11942 8342 11994
rect 8394 11942 8406 11994
rect 8458 11942 8470 11994
rect 8522 11942 13892 11994
rect 1104 11920 13892 11942
rect 842 11840 848 11892
rect 900 11880 906 11892
rect 900 11852 2452 11880
rect 900 11840 906 11852
rect 1854 11772 1860 11824
rect 1912 11812 1918 11824
rect 2317 11815 2375 11821
rect 2317 11812 2329 11815
rect 1912 11784 2329 11812
rect 1912 11772 1918 11784
rect 2317 11781 2329 11784
rect 2363 11781 2375 11815
rect 2424 11812 2452 11852
rect 2590 11840 2596 11892
rect 2648 11880 2654 11892
rect 2685 11883 2743 11889
rect 2685 11880 2697 11883
rect 2648 11852 2697 11880
rect 2648 11840 2654 11852
rect 2685 11849 2697 11852
rect 2731 11880 2743 11883
rect 3329 11883 3387 11889
rect 3329 11880 3341 11883
rect 2731 11852 3341 11880
rect 2731 11849 2743 11852
rect 2685 11843 2743 11849
rect 3329 11849 3341 11852
rect 3375 11880 3387 11883
rect 4154 11880 4160 11892
rect 3375 11852 4160 11880
rect 3375 11849 3387 11852
rect 3329 11843 3387 11849
rect 4154 11840 4160 11852
rect 4212 11840 4218 11892
rect 5258 11880 5264 11892
rect 4356 11852 5264 11880
rect 3694 11812 3700 11824
rect 2424 11784 3280 11812
rect 3655 11784 3700 11812
rect 2317 11775 2375 11781
rect 1486 11704 1492 11756
rect 1544 11744 1550 11756
rect 1581 11747 1639 11753
rect 1581 11744 1593 11747
rect 1544 11716 1593 11744
rect 1544 11704 1550 11716
rect 1581 11713 1593 11716
rect 1627 11713 1639 11747
rect 1581 11707 1639 11713
rect 2406 11704 2412 11756
rect 2464 11744 2470 11756
rect 3252 11753 3280 11784
rect 3694 11772 3700 11784
rect 3752 11772 3758 11824
rect 4356 11821 4384 11852
rect 5258 11840 5264 11852
rect 5316 11840 5322 11892
rect 6546 11840 6552 11892
rect 6604 11880 6610 11892
rect 7009 11883 7067 11889
rect 7009 11880 7021 11883
rect 6604 11852 7021 11880
rect 6604 11840 6610 11852
rect 7009 11849 7021 11852
rect 7055 11849 7067 11883
rect 7009 11843 7067 11849
rect 7101 11883 7159 11889
rect 7101 11849 7113 11883
rect 7147 11880 7159 11883
rect 7374 11880 7380 11892
rect 7147 11852 7380 11880
rect 7147 11849 7159 11852
rect 7101 11843 7159 11849
rect 7374 11840 7380 11852
rect 7432 11840 7438 11892
rect 7466 11840 7472 11892
rect 7524 11880 7530 11892
rect 7834 11880 7840 11892
rect 7524 11852 7840 11880
rect 7524 11840 7530 11852
rect 7834 11840 7840 11852
rect 7892 11840 7898 11892
rect 8297 11883 8355 11889
rect 8297 11849 8309 11883
rect 8343 11880 8355 11883
rect 8846 11880 8852 11892
rect 8343 11852 8852 11880
rect 8343 11849 8355 11852
rect 8297 11843 8355 11849
rect 8846 11840 8852 11852
rect 8904 11840 8910 11892
rect 9122 11840 9128 11892
rect 9180 11880 9186 11892
rect 13924 11880 13952 12124
rect 9180 11852 10824 11880
rect 9180 11840 9186 11852
rect 4341 11815 4399 11821
rect 4341 11781 4353 11815
rect 4387 11781 4399 11815
rect 4341 11775 4399 11781
rect 4433 11815 4491 11821
rect 4433 11781 4445 11815
rect 4479 11812 4491 11815
rect 5074 11812 5080 11824
rect 4479 11784 5080 11812
rect 4479 11781 4491 11784
rect 4433 11775 4491 11781
rect 5074 11772 5080 11784
rect 5132 11772 5138 11824
rect 5166 11772 5172 11824
rect 5224 11812 5230 11824
rect 7653 11815 7711 11821
rect 5224 11784 7604 11812
rect 5224 11772 5230 11784
rect 2501 11747 2559 11753
rect 2501 11744 2513 11747
rect 2464 11716 2513 11744
rect 2464 11704 2470 11716
rect 2501 11713 2513 11716
rect 2547 11713 2559 11747
rect 2501 11707 2559 11713
rect 2777 11747 2835 11753
rect 2777 11713 2789 11747
rect 2823 11744 2835 11747
rect 3053 11747 3111 11753
rect 2823 11716 3004 11744
rect 2823 11713 2835 11716
rect 2777 11707 2835 11713
rect 2133 11679 2191 11685
rect 2133 11676 2145 11679
rect 1596 11648 2145 11676
rect 1596 11620 1624 11648
rect 2133 11645 2145 11648
rect 2179 11645 2191 11679
rect 2976 11676 3004 11716
rect 3053 11713 3065 11747
rect 3099 11744 3111 11747
rect 3237 11747 3295 11753
rect 3099 11716 3188 11744
rect 3099 11713 3111 11716
rect 3053 11707 3111 11713
rect 2976 11648 3096 11676
rect 2133 11639 2191 11645
rect 1578 11568 1584 11620
rect 1636 11568 1642 11620
rect 1762 11568 1768 11620
rect 1820 11608 1826 11620
rect 2041 11611 2099 11617
rect 2041 11608 2053 11611
rect 1820 11580 2053 11608
rect 1820 11568 1826 11580
rect 2041 11577 2053 11580
rect 2087 11577 2099 11611
rect 2041 11571 2099 11577
rect 1489 11543 1547 11549
rect 1489 11509 1501 11543
rect 1535 11540 1547 11543
rect 1670 11540 1676 11552
rect 1535 11512 1676 11540
rect 1535 11509 1547 11512
rect 1489 11503 1547 11509
rect 1670 11500 1676 11512
rect 1728 11500 1734 11552
rect 2958 11540 2964 11552
rect 2919 11512 2964 11540
rect 2958 11500 2964 11512
rect 3016 11500 3022 11552
rect 3068 11540 3096 11648
rect 3160 11608 3188 11716
rect 3237 11713 3249 11747
rect 3283 11744 3295 11747
rect 3418 11744 3424 11756
rect 3283 11716 3424 11744
rect 3283 11713 3295 11716
rect 3237 11707 3295 11713
rect 3418 11704 3424 11716
rect 3476 11704 3482 11756
rect 3513 11747 3571 11753
rect 3513 11713 3525 11747
rect 3559 11744 3571 11747
rect 5353 11747 5411 11753
rect 3559 11716 5212 11744
rect 3559 11713 3571 11716
rect 3513 11707 3571 11713
rect 3881 11679 3939 11685
rect 3881 11645 3893 11679
rect 3927 11676 3939 11679
rect 3970 11676 3976 11688
rect 3927 11648 3976 11676
rect 3927 11645 3939 11648
rect 3881 11639 3939 11645
rect 3970 11636 3976 11648
rect 4028 11636 4034 11688
rect 4525 11679 4583 11685
rect 4525 11645 4537 11679
rect 4571 11676 4583 11679
rect 4706 11676 4712 11688
rect 4571 11648 4712 11676
rect 4571 11645 4583 11648
rect 4525 11639 4583 11645
rect 4706 11636 4712 11648
rect 4764 11636 4770 11688
rect 4982 11636 4988 11688
rect 5040 11676 5046 11688
rect 5077 11679 5135 11685
rect 5077 11676 5089 11679
rect 5040 11648 5089 11676
rect 5040 11636 5046 11648
rect 5077 11645 5089 11648
rect 5123 11645 5135 11679
rect 5184 11676 5212 11716
rect 5353 11713 5365 11747
rect 5399 11744 5411 11747
rect 5534 11744 5540 11756
rect 5399 11716 5540 11744
rect 5399 11713 5411 11716
rect 5353 11707 5411 11713
rect 5534 11704 5540 11716
rect 5592 11704 5598 11756
rect 6181 11747 6239 11753
rect 6181 11713 6193 11747
rect 6227 11744 6239 11747
rect 6454 11744 6460 11756
rect 6227 11716 6460 11744
rect 6227 11713 6239 11716
rect 6181 11707 6239 11713
rect 6454 11704 6460 11716
rect 6512 11704 6518 11756
rect 6641 11747 6699 11753
rect 6641 11713 6653 11747
rect 6687 11713 6699 11747
rect 6822 11744 6828 11756
rect 6783 11716 6828 11744
rect 6641 11707 6699 11713
rect 5721 11679 5779 11685
rect 5721 11676 5733 11679
rect 5184 11648 5733 11676
rect 5077 11639 5135 11645
rect 5721 11645 5733 11648
rect 5767 11645 5779 11679
rect 5721 11639 5779 11645
rect 5905 11679 5963 11685
rect 5905 11645 5917 11679
rect 5951 11676 5963 11679
rect 5994 11676 6000 11688
rect 5951 11648 6000 11676
rect 5951 11645 5963 11648
rect 5905 11639 5963 11645
rect 5994 11636 6000 11648
rect 6052 11636 6058 11688
rect 4614 11608 4620 11620
rect 3160 11580 4476 11608
rect 4575 11580 4620 11608
rect 3234 11540 3240 11552
rect 3068 11512 3240 11540
rect 3234 11500 3240 11512
rect 3292 11540 3298 11552
rect 3786 11540 3792 11552
rect 3292 11512 3792 11540
rect 3292 11500 3298 11512
rect 3786 11500 3792 11512
rect 3844 11500 3850 11552
rect 4448 11540 4476 11580
rect 4614 11568 4620 11580
rect 4672 11568 4678 11620
rect 5810 11608 5816 11620
rect 5184 11580 5816 11608
rect 5184 11540 5212 11580
rect 5810 11568 5816 11580
rect 5868 11568 5874 11620
rect 6086 11608 6092 11620
rect 6047 11580 6092 11608
rect 6086 11568 6092 11580
rect 6144 11568 6150 11620
rect 4448 11512 5212 11540
rect 5261 11543 5319 11549
rect 5261 11509 5273 11543
rect 5307 11540 5319 11543
rect 5350 11540 5356 11552
rect 5307 11512 5356 11540
rect 5307 11509 5319 11512
rect 5261 11503 5319 11509
rect 5350 11500 5356 11512
rect 5408 11500 5414 11552
rect 6656 11540 6684 11707
rect 6822 11704 6828 11716
rect 6880 11704 6886 11756
rect 7098 11704 7104 11756
rect 7156 11744 7162 11756
rect 7213 11747 7271 11753
rect 7213 11744 7225 11747
rect 7156 11716 7225 11744
rect 7156 11704 7162 11716
rect 7213 11713 7225 11716
rect 7259 11713 7271 11747
rect 7213 11707 7271 11713
rect 7469 11747 7527 11753
rect 7469 11713 7481 11747
rect 7515 11713 7527 11747
rect 7576 11744 7604 11784
rect 7653 11781 7665 11815
rect 7699 11812 7711 11815
rect 7926 11812 7932 11824
rect 7699 11784 7932 11812
rect 7699 11781 7711 11784
rect 7653 11775 7711 11781
rect 7926 11772 7932 11784
rect 7984 11772 7990 11824
rect 9677 11815 9735 11821
rect 9677 11812 9689 11815
rect 8036 11784 9689 11812
rect 8036 11744 8064 11784
rect 9677 11781 9689 11784
rect 9723 11781 9735 11815
rect 10134 11812 10140 11824
rect 10095 11784 10140 11812
rect 9677 11775 9735 11781
rect 10134 11772 10140 11784
rect 10192 11772 10198 11824
rect 10226 11772 10232 11824
rect 10284 11812 10290 11824
rect 10284 11784 10329 11812
rect 10284 11772 10290 11784
rect 10410 11772 10416 11824
rect 10468 11812 10474 11824
rect 10796 11821 10824 11852
rect 10888 11852 13952 11880
rect 10888 11821 10916 11852
rect 10781 11815 10839 11821
rect 10468 11784 10513 11812
rect 10468 11772 10474 11784
rect 10781 11781 10793 11815
rect 10827 11781 10839 11815
rect 10781 11775 10839 11781
rect 10873 11815 10931 11821
rect 10873 11781 10885 11815
rect 10919 11781 10931 11815
rect 10873 11775 10931 11781
rect 11422 11772 11428 11824
rect 11480 11812 11486 11824
rect 11480 11784 11744 11812
rect 11480 11772 11486 11784
rect 8570 11744 8576 11756
rect 7576 11716 8064 11744
rect 8531 11716 8576 11744
rect 7469 11707 7527 11713
rect 6914 11676 6920 11688
rect 6748 11648 6920 11676
rect 6748 11617 6776 11648
rect 6914 11636 6920 11648
rect 6972 11636 6978 11688
rect 7484 11676 7512 11707
rect 8570 11704 8576 11716
rect 8628 11704 8634 11756
rect 8846 11704 8852 11756
rect 8904 11744 8910 11756
rect 9030 11744 9036 11756
rect 8904 11716 8949 11744
rect 8991 11716 9036 11744
rect 8904 11704 8910 11716
rect 9030 11704 9036 11716
rect 9088 11704 9094 11756
rect 9122 11704 9128 11756
rect 9180 11744 9186 11756
rect 9306 11753 9312 11756
rect 9269 11747 9312 11753
rect 9180 11716 9225 11744
rect 9180 11704 9186 11716
rect 9269 11713 9281 11747
rect 9269 11707 9312 11713
rect 9306 11704 9312 11707
rect 9364 11704 9370 11756
rect 9398 11704 9404 11756
rect 9456 11744 9462 11756
rect 9861 11747 9919 11753
rect 9861 11744 9873 11747
rect 9456 11716 9873 11744
rect 9456 11704 9462 11716
rect 9861 11713 9873 11716
rect 9907 11713 9919 11747
rect 10042 11744 10048 11756
rect 10003 11716 10048 11744
rect 9861 11707 9919 11713
rect 10042 11704 10048 11716
rect 10100 11704 10106 11756
rect 11054 11744 11060 11756
rect 10244 11716 11060 11744
rect 7926 11676 7932 11688
rect 7484 11648 7932 11676
rect 7926 11636 7932 11648
rect 7984 11636 7990 11688
rect 8205 11679 8263 11685
rect 8205 11645 8217 11679
rect 8251 11645 8263 11679
rect 8478 11676 8484 11688
rect 8439 11648 8484 11676
rect 8205 11639 8263 11645
rect 6733 11611 6791 11617
rect 6733 11577 6745 11611
rect 6779 11577 6791 11611
rect 6733 11571 6791 11577
rect 7098 11568 7104 11620
rect 7156 11608 7162 11620
rect 8021 11611 8079 11617
rect 8021 11608 8033 11611
rect 7156 11580 8033 11608
rect 7156 11568 7162 11580
rect 8021 11577 8033 11580
rect 8067 11577 8079 11611
rect 8220 11608 8248 11639
rect 8478 11636 8484 11648
rect 8536 11636 8542 11688
rect 10244 11676 10272 11716
rect 11054 11704 11060 11716
rect 11112 11704 11118 11756
rect 11514 11744 11520 11756
rect 11475 11716 11520 11744
rect 11514 11704 11520 11716
rect 11572 11704 11578 11756
rect 11716 11744 11744 11784
rect 11974 11772 11980 11824
rect 12032 11812 12038 11824
rect 12069 11815 12127 11821
rect 12069 11812 12081 11815
rect 12032 11784 12081 11812
rect 12032 11772 12038 11784
rect 12069 11781 12081 11784
rect 12115 11781 12127 11815
rect 13078 11812 13084 11824
rect 13039 11784 13084 11812
rect 12069 11775 12127 11781
rect 13078 11772 13084 11784
rect 13136 11772 13142 11824
rect 13280 11821 13308 11852
rect 13265 11815 13323 11821
rect 13265 11781 13277 11815
rect 13311 11781 13323 11815
rect 13446 11812 13452 11824
rect 13407 11784 13452 11812
rect 13265 11775 13323 11781
rect 13446 11772 13452 11784
rect 13504 11772 13510 11824
rect 12161 11747 12219 11753
rect 12161 11744 12173 11747
rect 11716 11716 12173 11744
rect 12161 11713 12173 11716
rect 12207 11713 12219 11747
rect 12161 11707 12219 11713
rect 11330 11676 11336 11688
rect 9048 11648 10272 11676
rect 10336 11648 11336 11676
rect 8294 11608 8300 11620
rect 8220 11580 8300 11608
rect 8021 11571 8079 11577
rect 8294 11568 8300 11580
rect 8352 11568 8358 11620
rect 7006 11540 7012 11552
rect 6656 11512 7012 11540
rect 7006 11500 7012 11512
rect 7064 11500 7070 11552
rect 7282 11500 7288 11552
rect 7340 11540 7346 11552
rect 7742 11540 7748 11552
rect 7340 11512 7748 11540
rect 7340 11500 7346 11512
rect 7742 11500 7748 11512
rect 7800 11500 7806 11552
rect 7834 11500 7840 11552
rect 7892 11540 7898 11552
rect 8765 11543 8823 11549
rect 8765 11540 8777 11543
rect 7892 11512 8777 11540
rect 7892 11500 7898 11512
rect 8765 11509 8777 11512
rect 8811 11540 8823 11543
rect 9048 11540 9076 11648
rect 9122 11568 9128 11620
rect 9180 11608 9186 11620
rect 9582 11608 9588 11620
rect 9180 11580 9588 11608
rect 9180 11568 9186 11580
rect 9582 11568 9588 11580
rect 9640 11568 9646 11620
rect 8811 11512 9076 11540
rect 9401 11543 9459 11549
rect 8811 11509 8823 11512
rect 8765 11503 8823 11509
rect 9401 11509 9413 11543
rect 9447 11540 9459 11543
rect 10336 11540 10364 11648
rect 11330 11636 11336 11648
rect 11388 11636 11394 11688
rect 11606 11636 11612 11688
rect 11664 11676 11670 11688
rect 11977 11679 12035 11685
rect 11977 11676 11989 11679
rect 11664 11648 11989 11676
rect 11664 11636 11670 11648
rect 11977 11645 11989 11648
rect 12023 11645 12035 11679
rect 11977 11639 12035 11645
rect 12529 11679 12587 11685
rect 12529 11645 12541 11679
rect 12575 11676 12587 11679
rect 12618 11676 12624 11688
rect 12575 11648 12624 11676
rect 12575 11645 12587 11648
rect 12529 11639 12587 11645
rect 12618 11636 12624 11648
rect 12676 11636 12682 11688
rect 10686 11568 10692 11620
rect 10744 11608 10750 11620
rect 12986 11608 12992 11620
rect 10744 11580 12992 11608
rect 10744 11568 10750 11580
rect 12986 11568 12992 11580
rect 13044 11568 13050 11620
rect 9447 11512 10364 11540
rect 10413 11543 10471 11549
rect 9447 11509 9459 11512
rect 9401 11503 9459 11509
rect 10413 11509 10425 11543
rect 10459 11540 10471 11543
rect 10502 11540 10508 11552
rect 10459 11512 10508 11540
rect 10459 11509 10471 11512
rect 10413 11503 10471 11509
rect 10502 11500 10508 11512
rect 10560 11500 10566 11552
rect 10594 11500 10600 11552
rect 10652 11540 10658 11552
rect 10870 11540 10876 11552
rect 10652 11512 10876 11540
rect 10652 11500 10658 11512
rect 10870 11500 10876 11512
rect 10928 11500 10934 11552
rect 12253 11543 12311 11549
rect 12253 11509 12265 11543
rect 12299 11540 12311 11543
rect 12710 11540 12716 11552
rect 12299 11512 12716 11540
rect 12299 11509 12311 11512
rect 12253 11503 12311 11509
rect 12710 11500 12716 11512
rect 12768 11500 12774 11552
rect 1104 11450 13892 11472
rect 1104 11398 4214 11450
rect 4266 11398 4278 11450
rect 4330 11398 4342 11450
rect 4394 11398 4406 11450
rect 4458 11398 4470 11450
rect 4522 11398 12214 11450
rect 12266 11398 12278 11450
rect 12330 11398 12342 11450
rect 12394 11398 12406 11450
rect 12458 11398 12470 11450
rect 12522 11398 13892 11450
rect 1104 11376 13892 11398
rect 3602 11336 3608 11348
rect 3160 11308 3608 11336
rect 1762 11228 1768 11280
rect 1820 11268 1826 11280
rect 2685 11271 2743 11277
rect 2685 11268 2697 11271
rect 1820 11240 2697 11268
rect 1820 11228 1826 11240
rect 2685 11237 2697 11240
rect 2731 11237 2743 11271
rect 2685 11231 2743 11237
rect 3053 11203 3111 11209
rect 3053 11169 3065 11203
rect 3099 11200 3111 11203
rect 3160 11200 3188 11308
rect 3602 11296 3608 11308
rect 3660 11296 3666 11348
rect 4798 11296 4804 11348
rect 4856 11336 4862 11348
rect 6273 11339 6331 11345
rect 6273 11336 6285 11339
rect 4856 11308 6285 11336
rect 4856 11296 4862 11308
rect 6273 11305 6285 11308
rect 6319 11305 6331 11339
rect 6273 11299 6331 11305
rect 6454 11296 6460 11348
rect 6512 11336 6518 11348
rect 7745 11339 7803 11345
rect 6512 11308 7168 11336
rect 6512 11296 6518 11308
rect 5074 11268 5080 11280
rect 3620 11240 5080 11268
rect 3620 11212 3648 11240
rect 5074 11228 5080 11240
rect 5132 11228 5138 11280
rect 5258 11268 5264 11280
rect 5219 11240 5264 11268
rect 5258 11228 5264 11240
rect 5316 11228 5322 11280
rect 6086 11268 6092 11280
rect 6047 11240 6092 11268
rect 6086 11228 6092 11240
rect 6144 11228 6150 11280
rect 6638 11268 6644 11280
rect 6380 11240 6644 11268
rect 3602 11200 3608 11212
rect 3099 11172 3188 11200
rect 3515 11172 3608 11200
rect 3099 11169 3111 11172
rect 3053 11163 3111 11169
rect 3602 11160 3608 11172
rect 3660 11160 3666 11212
rect 3881 11203 3939 11209
rect 3881 11169 3893 11203
rect 3927 11200 3939 11203
rect 6270 11200 6276 11212
rect 3927 11172 6276 11200
rect 3927 11169 3939 11172
rect 3881 11163 3939 11169
rect 6270 11160 6276 11172
rect 6328 11160 6334 11212
rect 1397 11135 1455 11141
rect 1397 11101 1409 11135
rect 1443 11132 1455 11135
rect 1486 11132 1492 11144
rect 1443 11104 1492 11132
rect 1443 11101 1455 11104
rect 1397 11095 1455 11101
rect 1486 11092 1492 11104
rect 1544 11092 1550 11144
rect 2314 11132 2320 11144
rect 2275 11104 2320 11132
rect 2314 11092 2320 11104
rect 2372 11092 2378 11144
rect 3970 11132 3976 11144
rect 3931 11104 3976 11132
rect 3970 11092 3976 11104
rect 4028 11092 4034 11144
rect 5166 11132 5172 11144
rect 4080 11104 5172 11132
rect 3145 11067 3203 11073
rect 3145 11033 3157 11067
rect 3191 11064 3203 11067
rect 3234 11064 3240 11076
rect 3191 11036 3240 11064
rect 3191 11033 3203 11036
rect 3145 11027 3203 11033
rect 3234 11024 3240 11036
rect 3292 11024 3298 11076
rect 3510 11024 3516 11076
rect 3568 11064 3574 11076
rect 4080 11064 4108 11104
rect 5166 11092 5172 11104
rect 5224 11092 5230 11144
rect 5350 11132 5356 11144
rect 5311 11104 5356 11132
rect 5350 11092 5356 11104
rect 5408 11092 5414 11144
rect 5905 11135 5963 11141
rect 5905 11101 5917 11135
rect 5951 11132 5963 11135
rect 5994 11132 6000 11144
rect 5951 11104 6000 11132
rect 5951 11101 5963 11104
rect 5905 11095 5963 11101
rect 3568 11036 4108 11064
rect 3568 11024 3574 11036
rect 4154 11024 4160 11076
rect 4212 11064 4218 11076
rect 5920 11064 5948 11095
rect 5994 11092 6000 11104
rect 6052 11092 6058 11144
rect 6181 11135 6239 11141
rect 6181 11101 6193 11135
rect 6227 11132 6239 11135
rect 6380 11132 6408 11240
rect 6638 11228 6644 11240
rect 6696 11228 6702 11280
rect 7140 11268 7168 11308
rect 7745 11305 7757 11339
rect 7791 11336 7803 11339
rect 8846 11336 8852 11348
rect 7791 11308 8852 11336
rect 7791 11305 7803 11308
rect 7745 11299 7803 11305
rect 8846 11296 8852 11308
rect 8904 11296 8910 11348
rect 9030 11296 9036 11348
rect 9088 11336 9094 11348
rect 9088 11308 9812 11336
rect 9088 11296 9094 11308
rect 7140 11240 7236 11268
rect 6917 11203 6975 11209
rect 6917 11169 6929 11203
rect 6963 11200 6975 11203
rect 7098 11200 7104 11212
rect 6963 11172 7104 11200
rect 6963 11169 6975 11172
rect 6917 11163 6975 11169
rect 7098 11160 7104 11172
rect 7156 11160 7162 11212
rect 7208 11209 7236 11240
rect 7466 11228 7472 11280
rect 7524 11228 7530 11280
rect 7929 11271 7987 11277
rect 7929 11237 7941 11271
rect 7975 11268 7987 11271
rect 8202 11268 8208 11280
rect 7975 11240 8208 11268
rect 7975 11237 7987 11240
rect 7929 11231 7987 11237
rect 8202 11228 8208 11240
rect 8260 11228 8266 11280
rect 8570 11228 8576 11280
rect 8628 11268 8634 11280
rect 9677 11271 9735 11277
rect 9677 11268 9689 11271
rect 8628 11240 9689 11268
rect 8628 11228 8634 11240
rect 9677 11237 9689 11240
rect 9723 11237 9735 11271
rect 9784 11268 9812 11308
rect 10410 11296 10416 11348
rect 10468 11336 10474 11348
rect 10505 11339 10563 11345
rect 10505 11336 10517 11339
rect 10468 11308 10517 11336
rect 10468 11296 10474 11308
rect 10505 11305 10517 11308
rect 10551 11305 10563 11339
rect 10505 11299 10563 11305
rect 10594 11296 10600 11348
rect 10652 11336 10658 11348
rect 10873 11339 10931 11345
rect 10873 11336 10885 11339
rect 10652 11308 10885 11336
rect 10652 11296 10658 11308
rect 10873 11305 10885 11308
rect 10919 11305 10931 11339
rect 10873 11299 10931 11305
rect 11425 11339 11483 11345
rect 11425 11305 11437 11339
rect 11471 11336 11483 11339
rect 11514 11336 11520 11348
rect 11471 11308 11520 11336
rect 11471 11305 11483 11308
rect 11425 11299 11483 11305
rect 11514 11296 11520 11308
rect 11572 11296 11578 11348
rect 10962 11268 10968 11280
rect 9784 11240 10968 11268
rect 9677 11231 9735 11237
rect 10962 11228 10968 11240
rect 11020 11228 11026 11280
rect 11054 11228 11060 11280
rect 11112 11268 11118 11280
rect 12161 11271 12219 11277
rect 12161 11268 12173 11271
rect 11112 11240 12173 11268
rect 11112 11228 11118 11240
rect 12161 11237 12173 11240
rect 12207 11237 12219 11271
rect 12161 11231 12219 11237
rect 7193 11203 7251 11209
rect 7193 11169 7205 11203
rect 7239 11169 7251 11203
rect 7193 11163 7251 11169
rect 7282 11160 7288 11212
rect 7340 11200 7346 11212
rect 7484 11200 7512 11228
rect 7340 11172 7385 11200
rect 7484 11172 8432 11200
rect 7340 11160 7346 11172
rect 6227 11104 6408 11132
rect 6457 11135 6515 11141
rect 6227 11101 6239 11104
rect 6181 11095 6239 11101
rect 6457 11101 6469 11135
rect 6503 11101 6515 11135
rect 6457 11095 6515 11101
rect 6713 11135 6771 11141
rect 6713 11101 6725 11135
rect 6759 11101 6771 11135
rect 6713 11095 6771 11101
rect 4212 11036 5948 11064
rect 4212 11024 4218 11036
rect 6472 11008 6500 11095
rect 6728 11064 6756 11095
rect 6822 11092 6828 11144
rect 6880 11132 6886 11144
rect 7392 11141 7512 11142
rect 7007 11135 7065 11141
rect 7007 11132 7019 11135
rect 6880 11104 7019 11132
rect 6880 11092 6886 11104
rect 7007 11101 7019 11104
rect 7053 11101 7065 11135
rect 7007 11095 7065 11101
rect 7392 11135 7527 11141
rect 7392 11114 7481 11135
rect 7190 11064 7196 11076
rect 6728 11036 7196 11064
rect 7190 11024 7196 11036
rect 7248 11024 7254 11076
rect 7392 11064 7420 11114
rect 7469 11101 7481 11114
rect 7515 11101 7527 11135
rect 7469 11095 7527 11101
rect 7561 11135 7619 11141
rect 7561 11101 7573 11135
rect 7607 11132 7619 11135
rect 7607 11104 7970 11132
rect 7607 11101 7619 11104
rect 7561 11095 7619 11101
rect 7834 11064 7840 11076
rect 7392 11036 7840 11064
rect 1486 10956 1492 11008
rect 1544 10996 1550 11008
rect 2038 10996 2044 11008
rect 1544 10968 2044 10996
rect 1544 10956 1550 10968
rect 2038 10956 2044 10968
rect 2096 10996 2102 11008
rect 2590 10996 2596 11008
rect 2096 10968 2596 10996
rect 2096 10956 2102 10968
rect 2590 10956 2596 10968
rect 2648 10956 2654 11008
rect 4246 10956 4252 11008
rect 4304 10996 4310 11008
rect 5442 10996 5448 11008
rect 4304 10968 5448 10996
rect 4304 10956 4310 10968
rect 5442 10956 5448 10968
rect 5500 10956 5506 11008
rect 5626 10956 5632 11008
rect 5684 10996 5690 11008
rect 5721 10999 5779 11005
rect 5721 10996 5733 10999
rect 5684 10968 5733 10996
rect 5684 10956 5690 10968
rect 5721 10965 5733 10968
rect 5767 10965 5779 10999
rect 5721 10959 5779 10965
rect 6454 10956 6460 11008
rect 6512 10956 6518 11008
rect 6730 10956 6736 11008
rect 6788 10996 6794 11008
rect 6825 10999 6883 11005
rect 6825 10996 6837 10999
rect 6788 10968 6837 10996
rect 6788 10956 6794 10968
rect 6825 10965 6837 10968
rect 6871 10965 6883 10999
rect 6825 10959 6883 10965
rect 7006 10956 7012 11008
rect 7064 10996 7070 11008
rect 7392 10996 7420 11036
rect 7834 11024 7840 11036
rect 7892 11024 7898 11076
rect 7942 11064 7970 11104
rect 8110 11092 8116 11144
rect 8168 11132 8174 11144
rect 8404 11141 8432 11172
rect 8478 11160 8484 11212
rect 8536 11200 8542 11212
rect 8941 11203 8999 11209
rect 8941 11200 8953 11203
rect 8536 11172 8953 11200
rect 8536 11160 8542 11172
rect 8941 11169 8953 11172
rect 8987 11169 8999 11203
rect 8941 11163 8999 11169
rect 9030 11160 9036 11212
rect 9088 11200 9094 11212
rect 9088 11172 9168 11200
rect 9088 11160 9094 11172
rect 8204 11135 8262 11141
rect 8204 11132 8216 11135
rect 8168 11104 8216 11132
rect 8168 11092 8174 11104
rect 8204 11101 8216 11104
rect 8250 11101 8262 11135
rect 8204 11095 8262 11101
rect 8297 11135 8355 11141
rect 8297 11101 8309 11135
rect 8343 11101 8355 11135
rect 8297 11095 8355 11101
rect 8389 11135 8447 11141
rect 8389 11101 8401 11135
rect 8435 11101 8447 11135
rect 8570 11132 8576 11144
rect 8531 11104 8576 11132
rect 8389 11095 8447 11101
rect 8312 11064 8340 11095
rect 8570 11092 8576 11104
rect 8628 11092 8634 11144
rect 9140 11141 9168 11172
rect 9766 11160 9772 11212
rect 9824 11200 9830 11212
rect 10045 11203 10103 11209
rect 10045 11200 10057 11203
rect 9824 11172 10057 11200
rect 9824 11160 9830 11172
rect 10045 11169 10057 11172
rect 10091 11200 10103 11203
rect 10091 11172 10824 11200
rect 10091 11169 10103 11172
rect 10045 11163 10103 11169
rect 9125 11135 9183 11141
rect 9125 11101 9137 11135
rect 9171 11101 9183 11135
rect 9125 11095 9183 11101
rect 9214 11092 9220 11144
rect 9272 11141 9278 11144
rect 9272 11135 9321 11141
rect 9272 11101 9275 11135
rect 9309 11101 9321 11135
rect 9490 11132 9496 11144
rect 9451 11104 9496 11132
rect 9272 11095 9321 11101
rect 9272 11092 9278 11095
rect 9490 11092 9496 11104
rect 9548 11092 9554 11144
rect 9585 11135 9643 11141
rect 9585 11101 9597 11135
rect 9631 11101 9643 11135
rect 9585 11095 9643 11101
rect 8662 11064 8668 11076
rect 7942 11036 8668 11064
rect 8662 11024 8668 11036
rect 8720 11024 8726 11076
rect 8757 11067 8815 11073
rect 8757 11033 8769 11067
rect 8803 11064 8815 11067
rect 8938 11064 8944 11076
rect 8803 11036 8944 11064
rect 8803 11033 8815 11036
rect 8757 11027 8815 11033
rect 7064 10968 7420 10996
rect 7064 10956 7070 10968
rect 8386 10956 8392 11008
rect 8444 10996 8450 11008
rect 8772 10996 8800 11027
rect 8938 11024 8944 11036
rect 8996 11024 9002 11076
rect 9600 11064 9628 11095
rect 9858 11092 9864 11144
rect 9916 11132 9922 11144
rect 9953 11135 10011 11141
rect 9953 11132 9965 11135
rect 9916 11104 9965 11132
rect 9916 11092 9922 11104
rect 9953 11101 9965 11104
rect 9999 11101 10011 11135
rect 10226 11132 10232 11144
rect 10187 11104 10232 11132
rect 9953 11095 10011 11101
rect 9508 11036 9628 11064
rect 9968 11064 9996 11095
rect 10226 11092 10232 11104
rect 10284 11092 10290 11144
rect 10321 11135 10379 11141
rect 10321 11101 10333 11135
rect 10367 11132 10379 11135
rect 10686 11132 10692 11144
rect 10367 11104 10692 11132
rect 10367 11101 10379 11104
rect 10321 11095 10379 11101
rect 10686 11092 10692 11104
rect 10744 11092 10750 11144
rect 10796 11141 10824 11172
rect 10888 11172 12020 11200
rect 10781 11135 10839 11141
rect 10781 11101 10793 11135
rect 10827 11101 10839 11135
rect 10781 11095 10839 11101
rect 10888 11064 10916 11172
rect 11054 11132 11060 11144
rect 11015 11104 11060 11132
rect 11054 11092 11060 11104
rect 11112 11132 11118 11144
rect 11422 11132 11428 11144
rect 11112 11104 11428 11132
rect 11112 11092 11118 11104
rect 11422 11092 11428 11104
rect 11480 11092 11486 11144
rect 11606 11132 11612 11144
rect 11567 11104 11612 11132
rect 11606 11092 11612 11104
rect 11664 11092 11670 11144
rect 11992 11141 12020 11172
rect 11977 11135 12035 11141
rect 11977 11101 11989 11135
rect 12023 11101 12035 11135
rect 11977 11095 12035 11101
rect 12345 11135 12403 11141
rect 12345 11101 12357 11135
rect 12391 11132 12403 11135
rect 12618 11132 12624 11144
rect 12391 11104 12624 11132
rect 12391 11101 12403 11104
rect 12345 11095 12403 11101
rect 12618 11092 12624 11104
rect 12676 11132 12682 11144
rect 13078 11132 13084 11144
rect 12676 11104 13084 11132
rect 12676 11092 12682 11104
rect 13078 11092 13084 11104
rect 13136 11092 13142 11144
rect 13262 11132 13268 11144
rect 13223 11104 13268 11132
rect 13262 11092 13268 11104
rect 13320 11092 13326 11144
rect 9968 11036 10916 11064
rect 8444 10968 8800 10996
rect 8444 10956 8450 10968
rect 9030 10956 9036 11008
rect 9088 10996 9094 11008
rect 9214 10996 9220 11008
rect 9088 10968 9220 10996
rect 9088 10956 9094 10968
rect 9214 10956 9220 10968
rect 9272 10996 9278 11008
rect 9508 10996 9536 11036
rect 11698 11024 11704 11076
rect 11756 11064 11762 11076
rect 11885 11067 11943 11073
rect 11885 11064 11897 11067
rect 11756 11036 11897 11064
rect 11756 11024 11762 11036
rect 11885 11033 11897 11036
rect 11931 11033 11943 11067
rect 12986 11064 12992 11076
rect 12947 11036 12992 11064
rect 11885 11027 11943 11033
rect 12986 11024 12992 11036
rect 13044 11024 13050 11076
rect 13538 11064 13544 11076
rect 13499 11036 13544 11064
rect 13538 11024 13544 11036
rect 13596 11024 13602 11076
rect 9272 10968 9536 10996
rect 11793 10999 11851 11005
rect 9272 10956 9278 10968
rect 11793 10965 11805 10999
rect 11839 10996 11851 10999
rect 11974 10996 11980 11008
rect 11839 10968 11980 10996
rect 11839 10965 11851 10968
rect 11793 10959 11851 10965
rect 11974 10956 11980 10968
rect 12032 10956 12038 11008
rect 13170 10956 13176 11008
rect 13228 10996 13234 11008
rect 13357 10999 13415 11005
rect 13357 10996 13369 10999
rect 13228 10968 13369 10996
rect 13228 10956 13234 10968
rect 13357 10965 13369 10968
rect 13403 10965 13415 10999
rect 13357 10959 13415 10965
rect 1104 10906 13892 10928
rect 1104 10854 8214 10906
rect 8266 10854 8278 10906
rect 8330 10854 8342 10906
rect 8394 10854 8406 10906
rect 8458 10854 8470 10906
rect 8522 10854 13892 10906
rect 1104 10832 13892 10854
rect 1486 10792 1492 10804
rect 1447 10764 1492 10792
rect 1486 10752 1492 10764
rect 1544 10752 1550 10804
rect 1688 10764 6408 10792
rect 1397 10659 1455 10665
rect 1397 10625 1409 10659
rect 1443 10656 1455 10659
rect 1486 10656 1492 10668
rect 1443 10628 1492 10656
rect 1443 10625 1455 10628
rect 1397 10619 1455 10625
rect 1486 10616 1492 10628
rect 1544 10616 1550 10668
rect 1688 10665 1716 10764
rect 2314 10684 2320 10736
rect 2372 10724 2378 10736
rect 2685 10727 2743 10733
rect 2685 10724 2697 10727
rect 2372 10696 2697 10724
rect 2372 10684 2378 10696
rect 2685 10693 2697 10696
rect 2731 10693 2743 10727
rect 2685 10687 2743 10693
rect 3881 10727 3939 10733
rect 3881 10693 3893 10727
rect 3927 10724 3939 10727
rect 3970 10724 3976 10736
rect 3927 10696 3976 10724
rect 3927 10693 3939 10696
rect 3881 10687 3939 10693
rect 3970 10684 3976 10696
rect 4028 10684 4034 10736
rect 4246 10724 4252 10736
rect 4207 10696 4252 10724
rect 4246 10684 4252 10696
rect 4304 10684 4310 10736
rect 4614 10684 4620 10736
rect 4672 10724 4678 10736
rect 5077 10727 5135 10733
rect 5077 10724 5089 10727
rect 4672 10696 5089 10724
rect 4672 10684 4678 10696
rect 5077 10693 5089 10696
rect 5123 10693 5135 10727
rect 5077 10687 5135 10693
rect 5629 10727 5687 10733
rect 5629 10693 5641 10727
rect 5675 10724 5687 10727
rect 6270 10724 6276 10736
rect 5675 10696 6276 10724
rect 5675 10693 5687 10696
rect 5629 10687 5687 10693
rect 6270 10684 6276 10696
rect 6328 10684 6334 10736
rect 6380 10724 6408 10764
rect 6638 10752 6644 10804
rect 6696 10792 6702 10804
rect 7006 10792 7012 10804
rect 6696 10764 7012 10792
rect 6696 10752 6702 10764
rect 7006 10752 7012 10764
rect 7064 10752 7070 10804
rect 7650 10752 7656 10804
rect 7708 10792 7714 10804
rect 7708 10764 7788 10792
rect 7708 10752 7714 10764
rect 6380 10696 7696 10724
rect 1673 10659 1731 10665
rect 1673 10625 1685 10659
rect 1719 10625 1731 10659
rect 2498 10656 2504 10668
rect 2459 10628 2504 10656
rect 1673 10619 1731 10625
rect 2498 10616 2504 10628
rect 2556 10616 2562 10668
rect 2961 10659 3019 10665
rect 2961 10625 2973 10659
rect 3007 10656 3019 10659
rect 3234 10656 3240 10668
rect 3007 10628 3240 10656
rect 3007 10625 3019 10628
rect 2961 10619 3019 10625
rect 3234 10616 3240 10628
rect 3292 10616 3298 10668
rect 3602 10656 3608 10668
rect 3563 10628 3608 10656
rect 3602 10616 3608 10628
rect 3660 10616 3666 10668
rect 4065 10659 4123 10665
rect 4065 10625 4077 10659
rect 4111 10656 4123 10659
rect 4154 10656 4160 10668
rect 4111 10628 4160 10656
rect 4111 10625 4123 10628
rect 4065 10619 4123 10625
rect 4154 10616 4160 10628
rect 4212 10616 4218 10668
rect 4338 10656 4344 10668
rect 4299 10628 4344 10656
rect 4338 10616 4344 10628
rect 4396 10616 4402 10668
rect 4433 10659 4491 10665
rect 4433 10625 4445 10659
rect 4479 10656 4491 10659
rect 4982 10656 4988 10668
rect 4479 10628 4988 10656
rect 4479 10625 4491 10628
rect 4433 10619 4491 10625
rect 4982 10616 4988 10628
rect 5040 10616 5046 10668
rect 5350 10656 5356 10668
rect 5311 10628 5356 10656
rect 5350 10616 5356 10628
rect 5408 10616 5414 10668
rect 5442 10616 5448 10668
rect 5500 10656 5506 10668
rect 5721 10659 5779 10665
rect 5721 10656 5733 10659
rect 5500 10628 5733 10656
rect 5500 10616 5506 10628
rect 5721 10625 5733 10628
rect 5767 10625 5779 10659
rect 5721 10619 5779 10625
rect 5905 10659 5963 10665
rect 5905 10625 5917 10659
rect 5951 10656 5963 10659
rect 6457 10659 6515 10665
rect 6457 10656 6469 10659
rect 5951 10628 6469 10656
rect 5951 10625 5963 10628
rect 5905 10619 5963 10625
rect 6457 10625 6469 10628
rect 6503 10625 6515 10659
rect 6457 10619 6515 10625
rect 6730 10616 6736 10668
rect 6788 10656 6794 10668
rect 6917 10659 6975 10665
rect 6917 10656 6929 10659
rect 6788 10628 6929 10656
rect 6788 10616 6794 10628
rect 6917 10625 6929 10628
rect 6963 10625 6975 10659
rect 7098 10656 7104 10668
rect 7059 10628 7104 10656
rect 6917 10619 6975 10625
rect 7098 10616 7104 10628
rect 7156 10616 7162 10668
rect 7282 10656 7288 10668
rect 7243 10628 7288 10656
rect 7282 10616 7288 10628
rect 7340 10616 7346 10668
rect 7466 10656 7472 10668
rect 7427 10628 7472 10656
rect 7466 10616 7472 10628
rect 7524 10616 7530 10668
rect 1857 10591 1915 10597
rect 1857 10557 1869 10591
rect 1903 10588 1915 10591
rect 2038 10588 2044 10600
rect 1903 10560 2044 10588
rect 1903 10557 1915 10560
rect 1857 10551 1915 10557
rect 2038 10548 2044 10560
rect 2096 10548 2102 10600
rect 2590 10588 2596 10600
rect 2551 10560 2596 10588
rect 2590 10548 2596 10560
rect 2648 10548 2654 10600
rect 6086 10548 6092 10600
rect 6144 10588 6150 10600
rect 6144 10560 6500 10588
rect 6144 10548 6150 10560
rect 3694 10480 3700 10532
rect 3752 10520 3758 10532
rect 5445 10523 5503 10529
rect 5445 10520 5457 10523
rect 3752 10492 5457 10520
rect 3752 10480 3758 10492
rect 5445 10489 5457 10492
rect 5491 10520 5503 10523
rect 5810 10520 5816 10532
rect 5491 10492 5816 10520
rect 5491 10489 5503 10492
rect 5445 10483 5503 10489
rect 5810 10480 5816 10492
rect 5868 10480 5874 10532
rect 6362 10480 6368 10532
rect 6420 10480 6426 10532
rect 6472 10520 6500 10560
rect 6546 10548 6552 10600
rect 6604 10588 6610 10600
rect 6641 10591 6699 10597
rect 6641 10588 6653 10591
rect 6604 10560 6653 10588
rect 6604 10548 6610 10560
rect 6641 10557 6653 10560
rect 6687 10557 6699 10591
rect 6641 10551 6699 10557
rect 6825 10591 6883 10597
rect 6825 10557 6837 10591
rect 6871 10588 6883 10591
rect 7668 10588 7696 10696
rect 7760 10665 7788 10764
rect 7926 10752 7932 10804
rect 7984 10792 7990 10804
rect 7984 10764 8524 10792
rect 7984 10752 7990 10764
rect 7834 10684 7840 10736
rect 7892 10724 7898 10736
rect 8496 10724 8524 10764
rect 8570 10752 8576 10804
rect 8628 10792 8634 10804
rect 9309 10795 9367 10801
rect 9309 10792 9321 10795
rect 8628 10764 9321 10792
rect 8628 10752 8634 10764
rect 9309 10761 9321 10764
rect 9355 10761 9367 10795
rect 9309 10755 9367 10761
rect 10336 10764 11192 10792
rect 8938 10724 8944 10736
rect 7892 10696 7972 10724
rect 7892 10684 7898 10696
rect 7944 10665 7972 10696
rect 8496 10696 8944 10724
rect 7745 10659 7803 10665
rect 7745 10625 7757 10659
rect 7791 10625 7803 10659
rect 7745 10619 7803 10625
rect 7927 10659 7985 10665
rect 7927 10625 7939 10659
rect 7973 10625 7985 10659
rect 8110 10656 8116 10668
rect 8072 10628 8116 10656
rect 7927 10619 7985 10625
rect 8110 10616 8116 10628
rect 8168 10616 8174 10668
rect 8205 10659 8263 10665
rect 8205 10625 8217 10659
rect 8251 10625 8263 10659
rect 8205 10619 8263 10625
rect 7834 10588 7840 10600
rect 6871 10560 7236 10588
rect 7668 10560 7840 10588
rect 6871 10557 6883 10560
rect 6825 10551 6883 10557
rect 6472 10492 6684 10520
rect 3970 10412 3976 10464
rect 4028 10452 4034 10464
rect 4338 10452 4344 10464
rect 4028 10424 4344 10452
rect 4028 10412 4034 10424
rect 4338 10412 4344 10424
rect 4396 10452 4402 10464
rect 5258 10452 5264 10464
rect 4396 10424 5264 10452
rect 4396 10412 4402 10424
rect 5258 10412 5264 10424
rect 5316 10412 5322 10464
rect 6089 10455 6147 10461
rect 6089 10421 6101 10455
rect 6135 10452 6147 10455
rect 6178 10452 6184 10464
rect 6135 10424 6184 10452
rect 6135 10421 6147 10424
rect 6089 10415 6147 10421
rect 6178 10412 6184 10424
rect 6236 10412 6242 10464
rect 6380 10452 6408 10480
rect 6546 10452 6552 10464
rect 6380 10424 6552 10452
rect 6546 10412 6552 10424
rect 6604 10412 6610 10464
rect 6656 10452 6684 10492
rect 6730 10480 6736 10532
rect 6788 10520 6794 10532
rect 7101 10523 7159 10529
rect 7101 10520 7113 10523
rect 6788 10492 7113 10520
rect 6788 10480 6794 10492
rect 7101 10489 7113 10492
rect 7147 10489 7159 10523
rect 7208 10520 7236 10560
rect 7834 10548 7840 10560
rect 7892 10548 7898 10600
rect 8221 10588 8249 10619
rect 8294 10616 8300 10668
rect 8352 10656 8358 10668
rect 8496 10656 8524 10696
rect 8938 10684 8944 10696
rect 8996 10684 9002 10736
rect 9140 10696 9628 10724
rect 8573 10659 8631 10665
rect 8573 10656 8585 10659
rect 8352 10628 8397 10656
rect 8496 10628 8585 10656
rect 8352 10616 8358 10628
rect 8573 10625 8585 10628
rect 8619 10625 8631 10659
rect 8573 10619 8631 10625
rect 8662 10616 8668 10668
rect 8720 10656 8726 10668
rect 8846 10656 8852 10668
rect 8720 10628 8765 10656
rect 8807 10628 8852 10656
rect 8720 10616 8726 10628
rect 8846 10616 8852 10628
rect 8904 10616 8910 10668
rect 9030 10656 9036 10668
rect 8991 10628 9036 10656
rect 9030 10616 9036 10628
rect 9088 10616 9094 10668
rect 8386 10588 8392 10600
rect 8221 10560 8392 10588
rect 8386 10548 8392 10560
rect 8444 10548 8450 10600
rect 7374 10520 7380 10532
rect 7208 10492 7380 10520
rect 7101 10483 7159 10489
rect 7374 10480 7380 10492
rect 7432 10520 7438 10532
rect 8110 10520 8116 10532
rect 7432 10492 8116 10520
rect 7432 10480 7438 10492
rect 8110 10480 8116 10492
rect 8168 10520 8174 10532
rect 8680 10520 8708 10616
rect 9140 10588 9168 10696
rect 9600 10665 9628 10696
rect 9674 10684 9680 10736
rect 9732 10724 9738 10736
rect 10045 10727 10103 10733
rect 10045 10724 10057 10727
rect 9732 10696 10057 10724
rect 9732 10684 9738 10696
rect 10045 10693 10057 10696
rect 10091 10693 10103 10727
rect 10226 10724 10232 10736
rect 10187 10696 10232 10724
rect 10045 10687 10103 10693
rect 10226 10684 10232 10696
rect 10284 10684 10290 10736
rect 9493 10659 9551 10665
rect 9493 10625 9505 10659
rect 9539 10625 9551 10659
rect 9493 10619 9551 10625
rect 9585 10659 9643 10665
rect 9585 10625 9597 10659
rect 9631 10656 9643 10659
rect 9766 10656 9772 10668
rect 9631 10628 9772 10656
rect 9631 10625 9643 10628
rect 9585 10619 9643 10625
rect 8168 10492 8708 10520
rect 9048 10560 9168 10588
rect 9508 10588 9536 10619
rect 9766 10616 9772 10628
rect 9824 10616 9830 10668
rect 10336 10656 10364 10764
rect 11054 10724 11060 10736
rect 10888 10696 11060 10724
rect 10502 10656 10508 10668
rect 9876 10628 10364 10656
rect 10463 10628 10508 10656
rect 9674 10588 9680 10600
rect 9508 10560 9680 10588
rect 8168 10480 8174 10492
rect 7561 10455 7619 10461
rect 7561 10452 7573 10455
rect 6656 10424 7573 10452
rect 7561 10421 7573 10424
rect 7607 10452 7619 10455
rect 9048 10452 9076 10560
rect 9674 10548 9680 10560
rect 9732 10548 9738 10600
rect 9876 10597 9904 10628
rect 10502 10616 10508 10628
rect 10560 10616 10566 10668
rect 10594 10616 10600 10668
rect 10652 10656 10658 10668
rect 10888 10665 10916 10696
rect 11054 10684 11060 10696
rect 11112 10684 11118 10736
rect 11164 10724 11192 10764
rect 11238 10752 11244 10804
rect 11296 10792 11302 10804
rect 12434 10792 12440 10804
rect 11296 10764 11341 10792
rect 11440 10764 12440 10792
rect 11296 10752 11302 10764
rect 11440 10724 11468 10764
rect 12434 10752 12440 10764
rect 12492 10752 12498 10804
rect 12529 10795 12587 10801
rect 12529 10761 12541 10795
rect 12575 10761 12587 10795
rect 12529 10755 12587 10761
rect 12158 10724 12164 10736
rect 11164 10696 11468 10724
rect 12119 10696 12164 10724
rect 11164 10665 11192 10696
rect 12158 10684 12164 10696
rect 12216 10724 12222 10736
rect 12544 10724 12572 10755
rect 13078 10724 13084 10736
rect 12216 10696 12572 10724
rect 13039 10696 13084 10724
rect 12216 10684 12222 10696
rect 13078 10684 13084 10696
rect 13136 10684 13142 10736
rect 10780 10659 10838 10665
rect 10652 10628 10697 10656
rect 10652 10616 10658 10628
rect 10780 10625 10792 10659
rect 10826 10625 10838 10659
rect 10780 10619 10838 10625
rect 10873 10659 10931 10665
rect 10873 10625 10885 10659
rect 10919 10625 10931 10659
rect 10873 10619 10931 10625
rect 11149 10659 11207 10665
rect 11149 10625 11161 10659
rect 11195 10625 11207 10659
rect 11149 10619 11207 10625
rect 9861 10591 9919 10597
rect 9861 10557 9873 10591
rect 9907 10557 9919 10591
rect 9861 10551 9919 10557
rect 10686 10548 10692 10600
rect 10744 10588 10750 10600
rect 10795 10588 10823 10619
rect 11238 10616 11244 10668
rect 11296 10656 11302 10668
rect 11517 10659 11575 10665
rect 11517 10656 11529 10659
rect 11296 10628 11529 10656
rect 11296 10616 11302 10628
rect 11517 10625 11529 10628
rect 11563 10625 11575 10659
rect 11517 10619 11575 10625
rect 11701 10659 11759 10665
rect 11701 10625 11713 10659
rect 11747 10625 11759 10659
rect 11701 10619 11759 10625
rect 10744 10560 10823 10588
rect 10965 10591 11023 10597
rect 10744 10548 10750 10560
rect 10965 10557 10977 10591
rect 11011 10557 11023 10591
rect 10965 10551 11023 10557
rect 9122 10480 9128 10532
rect 9180 10520 9186 10532
rect 10980 10520 11008 10551
rect 11054 10548 11060 10600
rect 11112 10588 11118 10600
rect 11716 10588 11744 10619
rect 11790 10616 11796 10668
rect 11848 10656 11854 10668
rect 11931 10659 11989 10665
rect 11931 10656 11943 10659
rect 11848 10628 11943 10656
rect 11848 10616 11854 10628
rect 11931 10625 11943 10628
rect 11977 10625 11989 10659
rect 11931 10619 11989 10625
rect 12045 10659 12103 10665
rect 12045 10625 12057 10659
rect 12091 10656 12103 10659
rect 12250 10656 12256 10668
rect 12091 10625 12112 10656
rect 12211 10628 12256 10656
rect 12045 10619 12112 10625
rect 12084 10588 12112 10619
rect 12250 10616 12256 10628
rect 12308 10656 12314 10668
rect 12894 10656 12900 10668
rect 12308 10628 12480 10656
rect 12855 10628 12900 10656
rect 12308 10616 12314 10628
rect 12452 10597 12480 10628
rect 12894 10616 12900 10628
rect 12952 10616 12958 10668
rect 12986 10616 12992 10668
rect 13044 10656 13050 10668
rect 13173 10659 13231 10665
rect 13173 10656 13185 10659
rect 13044 10628 13185 10656
rect 13044 10616 13050 10628
rect 13173 10625 13185 10628
rect 13219 10625 13231 10659
rect 13173 10619 13231 10625
rect 13449 10659 13507 10665
rect 13449 10625 13461 10659
rect 13495 10656 13507 10659
rect 13722 10656 13728 10668
rect 13495 10628 13728 10656
rect 13495 10625 13507 10628
rect 13449 10619 13507 10625
rect 13722 10616 13728 10628
rect 13780 10616 13786 10668
rect 11112 10560 11744 10588
rect 11900 10560 12112 10588
rect 12345 10591 12403 10597
rect 11112 10548 11118 10560
rect 11900 10532 11928 10560
rect 12345 10557 12357 10591
rect 12391 10557 12403 10591
rect 12345 10551 12403 10557
rect 12437 10591 12495 10597
rect 12437 10557 12449 10591
rect 12483 10557 12495 10591
rect 12437 10551 12495 10557
rect 12641 10591 12699 10597
rect 12641 10557 12653 10591
rect 12687 10588 12699 10591
rect 13630 10588 13636 10600
rect 12687 10560 13636 10588
rect 12687 10557 12699 10560
rect 12641 10551 12699 10557
rect 9180 10492 11008 10520
rect 9180 10480 9186 10492
rect 11882 10480 11888 10532
rect 11940 10480 11946 10532
rect 12066 10480 12072 10532
rect 12124 10520 12130 10532
rect 12360 10520 12388 10551
rect 13630 10548 13636 10560
rect 13688 10548 13694 10600
rect 12124 10492 12388 10520
rect 13449 10523 13507 10529
rect 12124 10480 12130 10492
rect 13449 10489 13461 10523
rect 13495 10489 13507 10523
rect 13449 10483 13507 10489
rect 7607 10424 9076 10452
rect 7607 10421 7619 10424
rect 7561 10415 7619 10421
rect 9766 10412 9772 10464
rect 9824 10452 9830 10464
rect 10226 10452 10232 10464
rect 9824 10424 9869 10452
rect 10187 10424 10232 10452
rect 9824 10412 9830 10424
rect 10226 10412 10232 10424
rect 10284 10412 10290 10464
rect 10962 10412 10968 10464
rect 11020 10452 11026 10464
rect 13464 10452 13492 10483
rect 11020 10424 13492 10452
rect 11020 10412 11026 10424
rect 1104 10362 13892 10384
rect 1104 10310 4214 10362
rect 4266 10310 4278 10362
rect 4330 10310 4342 10362
rect 4394 10310 4406 10362
rect 4458 10310 4470 10362
rect 4522 10310 12214 10362
rect 12266 10310 12278 10362
rect 12330 10310 12342 10362
rect 12394 10310 12406 10362
rect 12458 10310 12470 10362
rect 12522 10310 13892 10362
rect 1104 10288 13892 10310
rect 1489 10251 1547 10257
rect 1489 10217 1501 10251
rect 1535 10248 1547 10251
rect 2590 10248 2596 10260
rect 1535 10220 2596 10248
rect 1535 10217 1547 10220
rect 1489 10211 1547 10217
rect 2590 10208 2596 10220
rect 2648 10208 2654 10260
rect 3973 10251 4031 10257
rect 3973 10217 3985 10251
rect 4019 10248 4031 10251
rect 4706 10248 4712 10260
rect 4019 10220 4712 10248
rect 4019 10217 4031 10220
rect 3973 10211 4031 10217
rect 4706 10208 4712 10220
rect 4764 10208 4770 10260
rect 4798 10208 4804 10260
rect 4856 10248 4862 10260
rect 4982 10248 4988 10260
rect 4856 10220 4988 10248
rect 4856 10208 4862 10220
rect 4982 10208 4988 10220
rect 5040 10208 5046 10260
rect 6546 10208 6552 10260
rect 6604 10248 6610 10260
rect 7653 10251 7711 10257
rect 7653 10248 7665 10251
rect 6604 10220 7665 10248
rect 6604 10208 6610 10220
rect 7653 10217 7665 10220
rect 7699 10248 7711 10251
rect 8294 10248 8300 10260
rect 7699 10220 8300 10248
rect 7699 10217 7711 10220
rect 7653 10211 7711 10217
rect 8294 10208 8300 10220
rect 8352 10208 8358 10260
rect 8481 10251 8539 10257
rect 8481 10217 8493 10251
rect 8527 10248 8539 10251
rect 8570 10248 8576 10260
rect 8527 10220 8576 10248
rect 8527 10217 8539 10220
rect 8481 10211 8539 10217
rect 8570 10208 8576 10220
rect 8628 10208 8634 10260
rect 8754 10208 8760 10260
rect 8812 10248 8818 10260
rect 9125 10251 9183 10257
rect 9125 10248 9137 10251
rect 8812 10220 9137 10248
rect 8812 10208 8818 10220
rect 9125 10217 9137 10220
rect 9171 10217 9183 10251
rect 9125 10211 9183 10217
rect 9324 10220 9720 10248
rect 2498 10140 2504 10192
rect 2556 10180 2562 10192
rect 3329 10183 3387 10189
rect 3329 10180 3341 10183
rect 2556 10152 3341 10180
rect 2556 10140 2562 10152
rect 3329 10149 3341 10152
rect 3375 10149 3387 10183
rect 3329 10143 3387 10149
rect 5261 10183 5319 10189
rect 5261 10149 5273 10183
rect 5307 10180 5319 10183
rect 5534 10180 5540 10192
rect 5307 10152 5540 10180
rect 5307 10149 5319 10152
rect 5261 10143 5319 10149
rect 5534 10140 5540 10152
rect 5592 10180 5598 10192
rect 5718 10180 5724 10192
rect 5592 10152 5724 10180
rect 5592 10140 5598 10152
rect 5718 10140 5724 10152
rect 5776 10140 5782 10192
rect 6086 10140 6092 10192
rect 6144 10180 6150 10192
rect 6457 10183 6515 10189
rect 6457 10180 6469 10183
rect 6144 10152 6469 10180
rect 6144 10140 6150 10152
rect 6457 10149 6469 10152
rect 6503 10149 6515 10183
rect 6457 10143 6515 10149
rect 6730 10140 6736 10192
rect 6788 10140 6794 10192
rect 6914 10140 6920 10192
rect 6972 10180 6978 10192
rect 7101 10183 7159 10189
rect 7101 10180 7113 10183
rect 6972 10152 7113 10180
rect 6972 10140 6978 10152
rect 7101 10149 7113 10152
rect 7147 10149 7159 10183
rect 7101 10143 7159 10149
rect 7285 10183 7343 10189
rect 7285 10149 7297 10183
rect 7331 10180 7343 10183
rect 7466 10180 7472 10192
rect 7331 10152 7472 10180
rect 7331 10149 7343 10152
rect 7285 10143 7343 10149
rect 7466 10140 7472 10152
rect 7524 10140 7530 10192
rect 8386 10180 8392 10192
rect 8036 10152 8392 10180
rect 2958 10112 2964 10124
rect 1688 10084 2964 10112
rect 1688 10056 1716 10084
rect 2958 10072 2964 10084
rect 3016 10112 3022 10124
rect 3694 10112 3700 10124
rect 3016 10084 3700 10112
rect 3016 10072 3022 10084
rect 3694 10072 3700 10084
rect 3752 10072 3758 10124
rect 5350 10112 5356 10124
rect 3804 10084 5356 10112
rect 1670 10044 1676 10056
rect 1631 10016 1676 10044
rect 1670 10004 1676 10016
rect 1728 10004 1734 10056
rect 2038 10044 2044 10056
rect 1999 10016 2044 10044
rect 2038 10004 2044 10016
rect 2096 10004 2102 10056
rect 3050 10044 3056 10056
rect 3011 10016 3056 10044
rect 3050 10004 3056 10016
rect 3108 10004 3114 10056
rect 3804 10053 3832 10084
rect 5350 10072 5356 10084
rect 5408 10072 5414 10124
rect 5810 10072 5816 10124
rect 5868 10112 5874 10124
rect 6365 10115 6423 10121
rect 6365 10112 6377 10115
rect 5868 10084 6377 10112
rect 5868 10072 5874 10084
rect 6365 10081 6377 10084
rect 6411 10081 6423 10115
rect 6748 10112 6776 10140
rect 7006 10112 7012 10124
rect 6365 10075 6423 10081
rect 6610 10084 6776 10112
rect 6840 10084 7012 10112
rect 3789 10047 3847 10053
rect 3789 10013 3801 10047
rect 3835 10013 3847 10047
rect 3789 10007 3847 10013
rect 3878 10004 3884 10056
rect 3936 10044 3942 10056
rect 4157 10047 4215 10053
rect 4157 10044 4169 10047
rect 3936 10016 4169 10044
rect 3936 10004 3942 10016
rect 4157 10013 4169 10016
rect 4203 10013 4215 10047
rect 4522 10044 4528 10056
rect 4483 10016 4528 10044
rect 4157 10007 4215 10013
rect 4522 10004 4528 10016
rect 4580 10004 4586 10056
rect 4798 10044 4804 10056
rect 4759 10016 4804 10044
rect 4798 10004 4804 10016
rect 4856 10004 4862 10056
rect 5626 10004 5632 10056
rect 5684 10044 5690 10056
rect 5997 10047 6055 10053
rect 5997 10044 6009 10047
rect 5684 10016 6009 10044
rect 5684 10004 5690 10016
rect 5997 10013 6009 10016
rect 6043 10013 6055 10047
rect 5997 10007 6055 10013
rect 6086 10004 6092 10056
rect 6144 10044 6150 10056
rect 6610 10053 6638 10084
rect 6595 10047 6653 10053
rect 6595 10044 6607 10047
rect 6144 10016 6607 10044
rect 6144 10004 6150 10016
rect 6595 10013 6607 10016
rect 6641 10013 6653 10047
rect 6739 10047 6797 10053
rect 6739 10034 6751 10047
rect 6785 10034 6797 10047
rect 6595 10007 6653 10013
rect 1581 9979 1639 9985
rect 1581 9945 1593 9979
rect 1627 9976 1639 9979
rect 3142 9976 3148 9988
rect 1627 9948 3148 9976
rect 1627 9945 1639 9948
rect 1581 9939 1639 9945
rect 3142 9936 3148 9948
rect 3200 9936 3206 9988
rect 4341 9979 4399 9985
rect 4341 9945 4353 9979
rect 4387 9976 4399 9979
rect 5074 9976 5080 9988
rect 4387 9948 5080 9976
rect 4387 9945 4399 9948
rect 4341 9939 4399 9945
rect 5074 9936 5080 9948
rect 5132 9936 5138 9988
rect 5353 9979 5411 9985
rect 5353 9945 5365 9979
rect 5399 9976 5411 9979
rect 5445 9979 5503 9985
rect 5445 9976 5457 9979
rect 5399 9948 5457 9976
rect 5399 9945 5411 9948
rect 5353 9939 5411 9945
rect 5445 9945 5457 9948
rect 5491 9945 5503 9979
rect 5445 9939 5503 9945
rect 5534 9936 5540 9988
rect 5592 9976 5598 9988
rect 5813 9979 5871 9985
rect 5813 9976 5825 9979
rect 5592 9948 5825 9976
rect 5592 9936 5598 9948
rect 5813 9945 5825 9948
rect 5859 9945 5871 9979
rect 5813 9939 5871 9945
rect 6270 9936 6276 9988
rect 6328 9976 6334 9988
rect 6730 9982 6736 10034
rect 6788 10007 6797 10034
rect 6788 9982 6794 10007
rect 6328 9948 6373 9976
rect 6328 9936 6334 9948
rect 1857 9911 1915 9917
rect 1857 9877 1869 9911
rect 1903 9908 1915 9911
rect 4706 9908 4712 9920
rect 1903 9880 4712 9908
rect 1903 9877 1915 9880
rect 1857 9871 1915 9877
rect 4706 9868 4712 9880
rect 4764 9868 4770 9920
rect 5626 9908 5632 9920
rect 5587 9880 5632 9908
rect 5626 9868 5632 9880
rect 5684 9868 5690 9920
rect 6181 9911 6239 9917
rect 6181 9877 6193 9911
rect 6227 9908 6239 9911
rect 6546 9908 6552 9920
rect 6227 9880 6552 9908
rect 6227 9877 6239 9880
rect 6181 9871 6239 9877
rect 6546 9868 6552 9880
rect 6604 9868 6610 9920
rect 6730 9868 6736 9920
rect 6788 9908 6794 9920
rect 6840 9908 6868 10084
rect 7006 10072 7012 10084
rect 7064 10072 7070 10124
rect 7190 10072 7196 10124
rect 7248 10112 7254 10124
rect 7248 10084 7972 10112
rect 7248 10072 7254 10084
rect 7944 10053 7972 10084
rect 7929 10047 7987 10053
rect 7929 10013 7941 10047
rect 7975 10013 7987 10047
rect 7929 10007 7987 10013
rect 7006 9936 7012 9988
rect 7064 9976 7070 9988
rect 7561 9979 7619 9985
rect 7561 9976 7573 9979
rect 7064 9948 7573 9976
rect 7064 9936 7070 9948
rect 7561 9945 7573 9948
rect 7607 9976 7619 9979
rect 8036 9976 8064 10152
rect 8386 10140 8392 10152
rect 8444 10140 8450 10192
rect 8665 10183 8723 10189
rect 8665 10149 8677 10183
rect 8711 10180 8723 10183
rect 9214 10180 9220 10192
rect 8711 10152 9220 10180
rect 8711 10149 8723 10152
rect 8665 10143 8723 10149
rect 9214 10140 9220 10152
rect 9272 10140 9278 10192
rect 8294 10072 8300 10124
rect 8352 10112 8358 10124
rect 8352 10084 8892 10112
rect 8352 10072 8358 10084
rect 8205 10047 8263 10053
rect 8205 10013 8217 10047
rect 8251 10044 8263 10047
rect 8762 10044 8768 10056
rect 8251 10016 8768 10044
rect 8251 10013 8263 10016
rect 8205 10007 8263 10013
rect 8312 9985 8340 10016
rect 8762 10004 8768 10016
rect 8820 10004 8826 10056
rect 8864 10044 8892 10084
rect 8938 10072 8944 10124
rect 8996 10112 9002 10124
rect 9324 10112 9352 10220
rect 9582 10140 9588 10192
rect 9640 10140 9646 10192
rect 9600 10112 9628 10140
rect 8996 10084 9352 10112
rect 9416 10084 9628 10112
rect 9692 10112 9720 10220
rect 10318 10208 10324 10260
rect 10376 10248 10382 10260
rect 11882 10248 11888 10260
rect 10376 10220 11652 10248
rect 11843 10220 11888 10248
rect 10376 10208 10382 10220
rect 9858 10180 9864 10192
rect 9771 10152 9864 10180
rect 9858 10140 9864 10152
rect 9916 10180 9922 10192
rect 9916 10152 10548 10180
rect 9916 10140 9922 10152
rect 9692 10084 9808 10112
rect 8996 10072 9002 10084
rect 9416 10053 9444 10084
rect 9309 10047 9367 10053
rect 9309 10044 9321 10047
rect 8864 10016 9321 10044
rect 9309 10013 9321 10016
rect 9355 10013 9367 10047
rect 9309 10007 9367 10013
rect 9401 10047 9459 10053
rect 9401 10013 9413 10047
rect 9447 10013 9459 10047
rect 9582 10044 9588 10056
rect 9543 10016 9588 10044
rect 9401 10007 9459 10013
rect 9582 10004 9588 10016
rect 9640 10004 9646 10056
rect 9677 10047 9735 10053
rect 9677 10013 9689 10047
rect 9723 10013 9735 10047
rect 9677 10007 9735 10013
rect 7607 9948 8064 9976
rect 8297 9979 8355 9985
rect 7607 9945 7619 9948
rect 7561 9939 7619 9945
rect 8297 9945 8309 9979
rect 8343 9945 8355 9979
rect 9600 9976 9628 10004
rect 8297 9939 8355 9945
rect 8404 9948 9628 9976
rect 6788 9880 6868 9908
rect 6788 9868 6794 9880
rect 6914 9868 6920 9920
rect 6972 9908 6978 9920
rect 7282 9908 7288 9920
rect 6972 9880 7288 9908
rect 6972 9868 6978 9880
rect 7282 9868 7288 9880
rect 7340 9908 7346 9920
rect 7926 9908 7932 9920
rect 7340 9880 7932 9908
rect 7340 9868 7346 9880
rect 7926 9868 7932 9880
rect 7984 9868 7990 9920
rect 8113 9911 8171 9917
rect 8113 9877 8125 9911
rect 8159 9908 8171 9911
rect 8404 9908 8432 9948
rect 8159 9880 8432 9908
rect 8159 9877 8171 9880
rect 8113 9871 8171 9877
rect 8478 9868 8484 9920
rect 8536 9908 8542 9920
rect 9214 9908 9220 9920
rect 8536 9880 9220 9908
rect 8536 9868 8542 9880
rect 9214 9868 9220 9880
rect 9272 9868 9278 9920
rect 9692 9908 9720 10007
rect 9780 9976 9808 10084
rect 9876 10053 9904 10140
rect 9950 10072 9956 10124
rect 10008 10112 10014 10124
rect 10137 10115 10195 10121
rect 10137 10112 10149 10115
rect 10008 10084 10149 10112
rect 10008 10072 10014 10084
rect 10137 10081 10149 10084
rect 10183 10081 10195 10115
rect 10137 10075 10195 10081
rect 10244 10063 10456 10078
rect 10229 10057 10456 10063
rect 9861 10047 9919 10053
rect 9861 10013 9873 10047
rect 9907 10013 9919 10047
rect 10042 10044 10048 10056
rect 10003 10016 10048 10044
rect 9861 10007 9919 10013
rect 10042 10004 10048 10016
rect 10100 10004 10106 10056
rect 10229 10023 10241 10057
rect 10275 10056 10456 10057
rect 10275 10050 10416 10056
rect 10275 10023 10287 10050
rect 10229 10017 10287 10023
rect 10410 10004 10416 10050
rect 10468 10004 10474 10056
rect 10321 9979 10379 9985
rect 10321 9976 10333 9979
rect 9780 9948 10333 9976
rect 10321 9945 10333 9948
rect 10367 9945 10379 9979
rect 10520 9976 10548 10152
rect 10594 10140 10600 10192
rect 10652 10180 10658 10192
rect 11057 10183 11115 10189
rect 11057 10180 11069 10183
rect 10652 10152 11069 10180
rect 10652 10140 10658 10152
rect 11057 10149 11069 10152
rect 11103 10180 11115 10183
rect 11514 10180 11520 10192
rect 11103 10152 11520 10180
rect 11103 10149 11115 10152
rect 11057 10143 11115 10149
rect 11514 10140 11520 10152
rect 11572 10140 11578 10192
rect 10686 10072 10692 10124
rect 10744 10112 10750 10124
rect 11624 10112 11652 10220
rect 11882 10208 11888 10220
rect 11940 10208 11946 10260
rect 12066 10208 12072 10260
rect 12124 10248 12130 10260
rect 12161 10251 12219 10257
rect 12161 10248 12173 10251
rect 12124 10220 12173 10248
rect 12124 10208 12130 10220
rect 12161 10217 12173 10220
rect 12207 10217 12219 10251
rect 12161 10211 12219 10217
rect 13170 10140 13176 10192
rect 13228 10180 13234 10192
rect 13265 10183 13323 10189
rect 13265 10180 13277 10183
rect 13228 10152 13277 10180
rect 13228 10140 13234 10152
rect 13265 10149 13277 10152
rect 13311 10149 13323 10183
rect 13265 10143 13323 10149
rect 13354 10112 13360 10124
rect 10744 10084 11192 10112
rect 10744 10072 10750 10084
rect 10873 10047 10931 10053
rect 10873 10013 10885 10047
rect 10919 10013 10931 10047
rect 10873 10007 10931 10013
rect 10888 9976 10916 10007
rect 10962 10004 10968 10056
rect 11020 10044 11026 10056
rect 11164 10053 11192 10084
rect 11532 10084 12572 10112
rect 13315 10084 13360 10112
rect 11532 10053 11560 10084
rect 11149 10047 11207 10053
rect 11020 10016 11065 10044
rect 11020 10004 11026 10016
rect 11149 10013 11161 10047
rect 11195 10013 11207 10047
rect 11149 10007 11207 10013
rect 11517 10047 11575 10053
rect 11517 10013 11529 10047
rect 11563 10013 11575 10047
rect 11517 10007 11575 10013
rect 11609 10047 11667 10053
rect 11609 10013 11621 10047
rect 11655 10013 11667 10047
rect 11609 10007 11667 10013
rect 11977 10047 12035 10053
rect 11977 10013 11989 10047
rect 12023 10044 12035 10047
rect 12066 10044 12072 10056
rect 12023 10016 12072 10044
rect 12023 10013 12035 10016
rect 11977 10007 12035 10013
rect 11422 9976 11428 9988
rect 10520 9948 10640 9976
rect 10888 9948 11428 9976
rect 10321 9939 10379 9945
rect 10502 9908 10508 9920
rect 9692 9880 10508 9908
rect 10502 9868 10508 9880
rect 10560 9868 10566 9920
rect 10612 9908 10640 9948
rect 11422 9936 11428 9948
rect 11480 9976 11486 9988
rect 11624 9976 11652 10007
rect 12066 10004 12072 10016
rect 12124 10004 12130 10056
rect 12434 10044 12440 10056
rect 12395 10016 12440 10044
rect 12434 10004 12440 10016
rect 12492 10004 12498 10056
rect 12544 10053 12572 10084
rect 13354 10072 13360 10084
rect 13412 10072 13418 10124
rect 12529 10047 12587 10053
rect 12529 10013 12541 10047
rect 12575 10013 12587 10047
rect 12802 10044 12808 10056
rect 12763 10016 12808 10044
rect 12529 10007 12587 10013
rect 12802 10004 12808 10016
rect 12860 10004 12866 10056
rect 11480 9948 11652 9976
rect 11480 9936 11486 9948
rect 11790 9936 11796 9988
rect 11848 9976 11854 9988
rect 13449 9979 13507 9985
rect 13449 9976 13461 9979
rect 11848 9948 13461 9976
rect 11848 9936 11854 9948
rect 13449 9945 13461 9948
rect 13495 9945 13507 9979
rect 13449 9939 13507 9945
rect 11238 9908 11244 9920
rect 10612 9880 11244 9908
rect 11238 9868 11244 9880
rect 11296 9868 11302 9920
rect 1104 9818 13892 9840
rect 1104 9766 8214 9818
rect 8266 9766 8278 9818
rect 8330 9766 8342 9818
rect 8394 9766 8406 9818
rect 8458 9766 8470 9818
rect 8522 9766 13892 9818
rect 1104 9744 13892 9766
rect 6181 9707 6239 9713
rect 6181 9673 6193 9707
rect 6227 9704 6239 9707
rect 6270 9704 6276 9716
rect 6227 9676 6276 9704
rect 6227 9673 6239 9676
rect 6181 9667 6239 9673
rect 6270 9664 6276 9676
rect 6328 9664 6334 9716
rect 7009 9707 7067 9713
rect 7009 9673 7021 9707
rect 7055 9673 7067 9707
rect 7009 9667 7067 9673
rect 2869 9639 2927 9645
rect 2869 9636 2881 9639
rect 2746 9608 2881 9636
rect 1854 9568 1860 9580
rect 1815 9540 1860 9568
rect 1854 9528 1860 9540
rect 1912 9528 1918 9580
rect 2593 9571 2651 9577
rect 2593 9537 2605 9571
rect 2639 9568 2651 9571
rect 2746 9568 2774 9608
rect 2869 9605 2881 9608
rect 2915 9636 2927 9639
rect 3050 9636 3056 9648
rect 2915 9608 3056 9636
rect 2915 9605 2927 9608
rect 2869 9599 2927 9605
rect 3050 9596 3056 9608
rect 3108 9596 3114 9648
rect 3694 9596 3700 9648
rect 3752 9636 3758 9648
rect 7022 9636 7050 9667
rect 7190 9664 7196 9716
rect 7248 9704 7254 9716
rect 7248 9676 7293 9704
rect 7248 9664 7254 9676
rect 7466 9664 7472 9716
rect 7524 9704 7530 9716
rect 7524 9676 7604 9704
rect 7524 9664 7530 9676
rect 7386 9639 7444 9645
rect 7386 9636 7398 9639
rect 3752 9608 4108 9636
rect 3752 9596 3758 9608
rect 3142 9568 3148 9580
rect 2639 9540 2774 9568
rect 3055 9540 3148 9568
rect 2639 9537 2651 9540
rect 2593 9531 2651 9537
rect 3142 9528 3148 9540
rect 3200 9568 3206 9580
rect 3602 9568 3608 9580
rect 3200 9540 3608 9568
rect 3200 9528 3206 9540
rect 3602 9528 3608 9540
rect 3660 9528 3666 9580
rect 4080 9577 4108 9608
rect 4356 9608 6960 9636
rect 7022 9608 7398 9636
rect 3789 9571 3847 9577
rect 3789 9537 3801 9571
rect 3835 9537 3847 9571
rect 3789 9531 3847 9537
rect 4065 9571 4123 9577
rect 4065 9537 4077 9571
rect 4111 9537 4123 9571
rect 4065 9531 4123 9537
rect 3694 9460 3700 9512
rect 3752 9500 3758 9512
rect 3804 9500 3832 9531
rect 4356 9500 4384 9608
rect 4433 9571 4491 9577
rect 4433 9537 4445 9571
rect 4479 9568 4491 9571
rect 4798 9568 4804 9580
rect 4479 9540 4804 9568
rect 4479 9537 4491 9540
rect 4433 9531 4491 9537
rect 4798 9528 4804 9540
rect 4856 9528 4862 9580
rect 5902 9568 5908 9580
rect 5863 9540 5908 9568
rect 5902 9528 5908 9540
rect 5960 9528 5966 9580
rect 6454 9528 6460 9580
rect 6512 9568 6518 9580
rect 6641 9571 6699 9577
rect 6641 9568 6653 9571
rect 6512 9540 6653 9568
rect 6512 9528 6518 9540
rect 6641 9537 6653 9540
rect 6687 9537 6699 9571
rect 6641 9531 6699 9537
rect 6825 9571 6883 9577
rect 6825 9537 6837 9571
rect 6871 9537 6883 9571
rect 6825 9531 6883 9537
rect 3752 9472 4384 9500
rect 3752 9460 3758 9472
rect 5718 9432 5724 9444
rect 5679 9404 5724 9432
rect 5718 9392 5724 9404
rect 5776 9392 5782 9444
rect 6840 9432 6868 9531
rect 6932 9500 6960 9608
rect 7386 9605 7398 9608
rect 7432 9636 7444 9639
rect 7576 9636 7604 9676
rect 8202 9664 8208 9716
rect 8260 9704 8266 9716
rect 9677 9707 9735 9713
rect 9677 9704 9689 9707
rect 8260 9676 8984 9704
rect 8260 9664 8266 9676
rect 7432 9608 7604 9636
rect 7791 9639 7849 9645
rect 7432 9605 7444 9608
rect 7386 9599 7444 9605
rect 7791 9605 7803 9639
rect 7837 9636 7849 9639
rect 8849 9639 8907 9645
rect 8849 9636 8861 9639
rect 7837 9608 8861 9636
rect 7837 9605 7849 9608
rect 7791 9599 7849 9605
rect 8849 9605 8861 9608
rect 8895 9605 8907 9639
rect 8956 9636 8984 9676
rect 9284 9676 9689 9704
rect 8956 9608 9076 9636
rect 8849 9599 8907 9605
rect 7006 9528 7012 9580
rect 7064 9568 7070 9580
rect 8202 9568 8208 9580
rect 7064 9540 7109 9568
rect 7576 9558 8208 9568
rect 7484 9552 8208 9558
rect 7340 9540 8208 9552
rect 7064 9528 7070 9540
rect 7340 9530 7604 9540
rect 7340 9524 7512 9530
rect 8202 9528 8208 9540
rect 8260 9528 8266 9580
rect 8297 9571 8355 9577
rect 8297 9537 8309 9571
rect 8343 9568 8355 9571
rect 8386 9568 8392 9580
rect 8343 9540 8392 9568
rect 8343 9537 8355 9540
rect 8297 9531 8355 9537
rect 8386 9528 8392 9540
rect 8444 9528 8450 9580
rect 8570 9528 8576 9580
rect 8628 9568 8634 9580
rect 9048 9577 9076 9608
rect 9122 9596 9128 9648
rect 9180 9636 9186 9648
rect 9284 9636 9312 9676
rect 9677 9673 9689 9676
rect 9723 9704 9735 9707
rect 10318 9704 10324 9716
rect 9723 9676 10324 9704
rect 9723 9673 9735 9676
rect 9677 9667 9735 9673
rect 10318 9664 10324 9676
rect 10376 9664 10382 9716
rect 10428 9676 10824 9704
rect 9398 9636 9404 9648
rect 9180 9608 9312 9636
rect 9359 9608 9404 9636
rect 9180 9596 9186 9608
rect 9398 9596 9404 9608
rect 9456 9596 9462 9648
rect 10428 9636 10456 9676
rect 9692 9608 10456 9636
rect 10505 9639 10563 9645
rect 8941 9571 8999 9577
rect 8628 9540 8673 9568
rect 8628 9528 8634 9540
rect 8941 9537 8953 9571
rect 8987 9537 8999 9571
rect 8941 9531 8999 9537
rect 9033 9571 9091 9577
rect 9033 9537 9045 9571
rect 9079 9537 9091 9571
rect 9033 9531 9091 9537
rect 6932 9472 7236 9500
rect 7006 9432 7012 9444
rect 6840 9404 7012 9432
rect 7006 9392 7012 9404
rect 7064 9392 7070 9444
rect 1394 9324 1400 9376
rect 1452 9364 1458 9376
rect 1489 9367 1547 9373
rect 1489 9364 1501 9367
rect 1452 9336 1501 9364
rect 1452 9324 1458 9336
rect 1489 9333 1501 9336
rect 1535 9333 1547 9367
rect 1489 9327 1547 9333
rect 2777 9367 2835 9373
rect 2777 9333 2789 9367
rect 2823 9364 2835 9367
rect 3510 9364 3516 9376
rect 2823 9336 3516 9364
rect 2823 9333 2835 9336
rect 2777 9327 2835 9333
rect 3510 9324 3516 9336
rect 3568 9324 3574 9376
rect 3878 9364 3884 9376
rect 3839 9336 3884 9364
rect 3878 9324 3884 9336
rect 3936 9324 3942 9376
rect 4249 9367 4307 9373
rect 4249 9333 4261 9367
rect 4295 9364 4307 9367
rect 4522 9364 4528 9376
rect 4295 9336 4528 9364
rect 4295 9333 4307 9336
rect 4249 9327 4307 9333
rect 4522 9324 4528 9336
rect 4580 9364 4586 9376
rect 4982 9364 4988 9376
rect 4580 9336 4988 9364
rect 4580 9324 4586 9336
rect 4982 9324 4988 9336
rect 5040 9324 5046 9376
rect 6457 9367 6515 9373
rect 6457 9333 6469 9367
rect 6503 9364 6515 9367
rect 7098 9364 7104 9376
rect 6503 9336 7104 9364
rect 6503 9333 6515 9336
rect 6457 9327 6515 9333
rect 7098 9324 7104 9336
rect 7156 9324 7162 9376
rect 7208 9364 7236 9472
rect 7282 9460 7288 9512
rect 7340 9472 7368 9524
rect 8754 9500 8760 9512
rect 8715 9472 8760 9500
rect 7340 9460 7346 9472
rect 8754 9460 8760 9472
rect 8812 9460 8818 9512
rect 8956 9500 8984 9531
rect 9140 9500 9168 9596
rect 9217 9571 9275 9577
rect 9217 9537 9229 9571
rect 9263 9568 9275 9571
rect 9582 9568 9588 9580
rect 9263 9540 9588 9568
rect 9263 9537 9275 9540
rect 9217 9531 9275 9537
rect 9582 9528 9588 9540
rect 9640 9568 9646 9580
rect 9692 9568 9720 9608
rect 10505 9605 10517 9639
rect 10551 9636 10563 9639
rect 10686 9636 10692 9648
rect 10551 9608 10692 9636
rect 10551 9605 10563 9608
rect 10505 9599 10563 9605
rect 10686 9596 10692 9608
rect 10744 9596 10750 9648
rect 10796 9636 10824 9676
rect 10962 9664 10968 9716
rect 11020 9704 11026 9716
rect 11241 9707 11299 9713
rect 11241 9704 11253 9707
rect 11020 9676 11253 9704
rect 11020 9664 11026 9676
rect 11241 9673 11253 9676
rect 11287 9673 11299 9707
rect 11241 9667 11299 9673
rect 13170 9636 13176 9648
rect 10796 9608 12020 9636
rect 13131 9608 13176 9636
rect 9858 9568 9864 9580
rect 9640 9540 9720 9568
rect 9819 9540 9864 9568
rect 9640 9528 9646 9540
rect 9858 9528 9864 9540
rect 9916 9528 9922 9580
rect 10137 9571 10195 9577
rect 10137 9568 10149 9571
rect 9968 9540 10149 9568
rect 8956 9472 9168 9500
rect 9398 9460 9404 9512
rect 9456 9500 9462 9512
rect 9968 9500 9996 9540
rect 10137 9537 10149 9540
rect 10183 9537 10195 9571
rect 10318 9568 10324 9580
rect 10279 9540 10324 9568
rect 10137 9531 10195 9537
rect 10318 9528 10324 9540
rect 10376 9528 10382 9580
rect 10594 9568 10600 9580
rect 10555 9540 10600 9568
rect 10594 9528 10600 9540
rect 10652 9528 10658 9580
rect 10781 9571 10839 9577
rect 10781 9537 10793 9571
rect 10827 9537 10839 9571
rect 10781 9531 10839 9537
rect 11057 9571 11115 9577
rect 11057 9537 11069 9571
rect 11103 9568 11115 9571
rect 11422 9568 11428 9580
rect 11103 9540 11428 9568
rect 11103 9537 11115 9540
rect 11057 9531 11115 9537
rect 9456 9472 9996 9500
rect 10045 9503 10103 9509
rect 9456 9460 9462 9472
rect 10045 9469 10057 9503
rect 10091 9469 10103 9503
rect 10045 9463 10103 9469
rect 7834 9432 7840 9444
rect 7484 9404 7840 9432
rect 7484 9364 7512 9404
rect 7834 9392 7840 9404
rect 7892 9392 7898 9444
rect 7929 9435 7987 9441
rect 7929 9401 7941 9435
rect 7975 9432 7987 9435
rect 9490 9432 9496 9444
rect 7975 9404 9496 9432
rect 7975 9401 7987 9404
rect 7929 9395 7987 9401
rect 9490 9392 9496 9404
rect 9548 9392 9554 9444
rect 10060 9432 10088 9463
rect 10134 9432 10140 9444
rect 10060 9404 10140 9432
rect 10134 9392 10140 9404
rect 10192 9432 10198 9444
rect 10410 9432 10416 9444
rect 10192 9404 10416 9432
rect 10192 9392 10198 9404
rect 10410 9392 10416 9404
rect 10468 9392 10474 9444
rect 10796 9432 10824 9531
rect 11422 9528 11428 9540
rect 11480 9528 11486 9580
rect 11701 9571 11759 9577
rect 11701 9568 11713 9571
rect 11532 9540 11713 9568
rect 10520 9404 10824 9432
rect 7208 9336 7512 9364
rect 7650 9324 7656 9376
rect 7708 9364 7714 9376
rect 7745 9367 7803 9373
rect 7745 9364 7757 9367
rect 7708 9336 7757 9364
rect 7708 9324 7714 9336
rect 7745 9333 7757 9336
rect 7791 9333 7803 9367
rect 7745 9327 7803 9333
rect 9030 9324 9036 9376
rect 9088 9364 9094 9376
rect 10520 9364 10548 9404
rect 10686 9364 10692 9376
rect 9088 9336 10548 9364
rect 10647 9336 10692 9364
rect 9088 9324 9094 9336
rect 10686 9324 10692 9336
rect 10744 9324 10750 9376
rect 10796 9364 10824 9404
rect 10962 9392 10968 9444
rect 11020 9432 11026 9444
rect 11532 9441 11560 9540
rect 11701 9537 11713 9540
rect 11747 9537 11759 9571
rect 11701 9531 11759 9537
rect 11793 9571 11851 9577
rect 11793 9537 11805 9571
rect 11839 9568 11851 9571
rect 11882 9568 11888 9580
rect 11839 9540 11888 9568
rect 11839 9537 11851 9540
rect 11793 9531 11851 9537
rect 11882 9528 11888 9540
rect 11940 9528 11946 9580
rect 11992 9577 12020 9608
rect 13170 9596 13176 9608
rect 13228 9596 13234 9648
rect 13262 9596 13268 9648
rect 13320 9636 13326 9648
rect 13357 9639 13415 9645
rect 13357 9636 13369 9639
rect 13320 9608 13369 9636
rect 13320 9596 13326 9608
rect 13357 9605 13369 9608
rect 13403 9636 13415 9639
rect 13446 9636 13452 9648
rect 13403 9608 13452 9636
rect 13403 9605 13415 9608
rect 13357 9599 13415 9605
rect 13446 9596 13452 9608
rect 13504 9596 13510 9648
rect 11977 9571 12035 9577
rect 11977 9537 11989 9571
rect 12023 9537 12035 9571
rect 11977 9531 12035 9537
rect 12161 9571 12219 9577
rect 12161 9537 12173 9571
rect 12207 9568 12219 9571
rect 12437 9571 12495 9577
rect 12437 9568 12449 9571
rect 12207 9540 12449 9568
rect 12207 9537 12219 9540
rect 12161 9531 12219 9537
rect 12437 9537 12449 9540
rect 12483 9568 12495 9571
rect 12802 9568 12808 9580
rect 12483 9540 12808 9568
rect 12483 9537 12495 9540
rect 12437 9531 12495 9537
rect 12802 9528 12808 9540
rect 12860 9528 12866 9580
rect 11517 9435 11575 9441
rect 11517 9432 11529 9435
rect 11020 9404 11529 9432
rect 11020 9392 11026 9404
rect 11517 9401 11529 9404
rect 11563 9401 11575 9435
rect 11517 9395 11575 9401
rect 11974 9364 11980 9376
rect 10796 9336 11980 9364
rect 11974 9324 11980 9336
rect 12032 9364 12038 9376
rect 12434 9364 12440 9376
rect 12032 9336 12440 9364
rect 12032 9324 12038 9336
rect 12434 9324 12440 9336
rect 12492 9324 12498 9376
rect 13446 9364 13452 9376
rect 13407 9336 13452 9364
rect 13446 9324 13452 9336
rect 13504 9324 13510 9376
rect 1104 9274 13892 9296
rect 1104 9222 4214 9274
rect 4266 9222 4278 9274
rect 4330 9222 4342 9274
rect 4394 9222 4406 9274
rect 4458 9222 4470 9274
rect 4522 9222 12214 9274
rect 12266 9222 12278 9274
rect 12330 9222 12342 9274
rect 12394 9222 12406 9274
rect 12458 9222 12470 9274
rect 12522 9222 13892 9274
rect 1104 9200 13892 9222
rect 5810 9120 5816 9172
rect 5868 9160 5874 9172
rect 6089 9163 6147 9169
rect 6089 9160 6101 9163
rect 5868 9132 6101 9160
rect 5868 9120 5874 9132
rect 6089 9129 6101 9132
rect 6135 9129 6147 9163
rect 6089 9123 6147 9129
rect 6549 9163 6607 9169
rect 6549 9129 6561 9163
rect 6595 9160 6607 9163
rect 6822 9160 6828 9172
rect 6595 9132 6828 9160
rect 6595 9129 6607 9132
rect 6549 9123 6607 9129
rect 6822 9120 6828 9132
rect 6880 9120 6886 9172
rect 7006 9120 7012 9172
rect 7064 9160 7070 9172
rect 7374 9160 7380 9172
rect 7064 9132 7380 9160
rect 7064 9120 7070 9132
rect 7374 9120 7380 9132
rect 7432 9160 7438 9172
rect 7469 9163 7527 9169
rect 7469 9160 7481 9163
rect 7432 9132 7481 9160
rect 7432 9120 7438 9132
rect 7469 9129 7481 9132
rect 7515 9129 7527 9163
rect 7469 9123 7527 9129
rect 7650 9120 7656 9172
rect 7708 9160 7714 9172
rect 7745 9163 7803 9169
rect 7745 9160 7757 9163
rect 7708 9132 7757 9160
rect 7708 9120 7714 9132
rect 7745 9129 7757 9132
rect 7791 9129 7803 9163
rect 8938 9160 8944 9172
rect 7745 9123 7803 9129
rect 8095 9132 8944 9160
rect 4617 9095 4675 9101
rect 4617 9061 4629 9095
rect 4663 9092 4675 9095
rect 4798 9092 4804 9104
rect 4663 9064 4804 9092
rect 4663 9061 4675 9064
rect 4617 9055 4675 9061
rect 4798 9052 4804 9064
rect 4856 9052 4862 9104
rect 6917 9095 6975 9101
rect 6917 9061 6929 9095
rect 6963 9061 6975 9095
rect 6917 9055 6975 9061
rect 3145 9027 3203 9033
rect 3145 8993 3157 9027
rect 3191 9024 3203 9027
rect 3786 9024 3792 9036
rect 3191 8996 3792 9024
rect 3191 8993 3203 8996
rect 3145 8987 3203 8993
rect 3786 8984 3792 8996
rect 3844 8984 3850 9036
rect 4706 9024 4712 9036
rect 4667 8996 4712 9024
rect 4706 8984 4712 8996
rect 4764 8984 4770 9036
rect 6932 9024 6960 9055
rect 7098 9024 7104 9036
rect 5009 8996 6592 9024
rect 1394 8956 1400 8968
rect 1355 8928 1400 8956
rect 1394 8916 1400 8928
rect 1452 8916 1458 8968
rect 2958 8916 2964 8968
rect 3016 8956 3022 8968
rect 3605 8959 3663 8965
rect 3605 8956 3617 8959
rect 3016 8928 3617 8956
rect 3016 8916 3022 8928
rect 3605 8925 3617 8928
rect 3651 8925 3663 8959
rect 3878 8956 3884 8968
rect 3839 8928 3884 8956
rect 3605 8919 3663 8925
rect 3878 8916 3884 8928
rect 3936 8916 3942 8968
rect 4157 8959 4215 8965
rect 4157 8925 4169 8959
rect 4203 8956 4215 8959
rect 4617 8959 4675 8965
rect 4203 8928 4568 8956
rect 4203 8925 4215 8928
rect 4157 8919 4215 8925
rect 3789 8891 3847 8897
rect 3789 8857 3801 8891
rect 3835 8888 3847 8891
rect 4249 8891 4307 8897
rect 4249 8888 4261 8891
rect 3835 8860 4261 8888
rect 3835 8857 3847 8860
rect 3789 8851 3847 8857
rect 4249 8857 4261 8860
rect 4295 8857 4307 8891
rect 4540 8888 4568 8928
rect 4617 8925 4629 8959
rect 4663 8956 4675 8959
rect 5009 8956 5037 8996
rect 4663 8928 5037 8956
rect 5077 8959 5135 8965
rect 4663 8925 4675 8928
rect 4617 8919 4675 8925
rect 5077 8925 5089 8959
rect 5123 8956 5135 8959
rect 5534 8956 5540 8968
rect 5123 8928 5540 8956
rect 5123 8925 5135 8928
rect 5077 8919 5135 8925
rect 5534 8916 5540 8928
rect 5592 8916 5598 8968
rect 5626 8916 5632 8968
rect 5684 8956 5690 8968
rect 5721 8959 5779 8965
rect 5721 8956 5733 8959
rect 5684 8928 5733 8956
rect 5684 8916 5690 8928
rect 5721 8925 5733 8928
rect 5767 8925 5779 8959
rect 5721 8919 5779 8925
rect 5902 8916 5908 8968
rect 5960 8956 5966 8968
rect 5997 8959 6055 8965
rect 5997 8956 6009 8959
rect 5960 8928 6009 8956
rect 5960 8916 5966 8928
rect 5997 8925 6009 8928
rect 6043 8925 6055 8959
rect 5997 8919 6055 8925
rect 6270 8916 6276 8968
rect 6328 8956 6334 8968
rect 6365 8959 6423 8965
rect 6365 8956 6377 8959
rect 6328 8928 6377 8956
rect 6328 8916 6334 8928
rect 6365 8925 6377 8928
rect 6411 8925 6423 8959
rect 6365 8919 6423 8925
rect 4982 8888 4988 8900
rect 4540 8860 4988 8888
rect 4249 8851 4307 8857
rect 4982 8848 4988 8860
rect 5040 8888 5046 8900
rect 5442 8888 5448 8900
rect 5040 8860 5448 8888
rect 5040 8848 5046 8860
rect 5442 8848 5448 8860
rect 5500 8848 5506 8900
rect 6564 8888 6592 8996
rect 6656 8996 6960 9024
rect 7059 8996 7104 9024
rect 6656 8965 6684 8996
rect 7098 8984 7104 8996
rect 7156 8984 7162 9036
rect 8095 9024 8123 9132
rect 8938 9120 8944 9132
rect 8996 9120 9002 9172
rect 9858 9120 9864 9172
rect 9916 9160 9922 9172
rect 10134 9160 10140 9172
rect 9916 9132 10140 9160
rect 9916 9120 9922 9132
rect 10134 9120 10140 9132
rect 10192 9120 10198 9172
rect 10226 9120 10232 9172
rect 10284 9160 10290 9172
rect 10689 9163 10747 9169
rect 10689 9160 10701 9163
rect 10284 9132 10701 9160
rect 10284 9120 10290 9132
rect 10689 9129 10701 9132
rect 10735 9129 10747 9163
rect 10689 9123 10747 9129
rect 11425 9163 11483 9169
rect 11425 9129 11437 9163
rect 11471 9160 11483 9163
rect 11606 9160 11612 9172
rect 11471 9132 11612 9160
rect 11471 9129 11483 9132
rect 11425 9123 11483 9129
rect 11606 9120 11612 9132
rect 11664 9120 11670 9172
rect 11882 9120 11888 9172
rect 11940 9160 11946 9172
rect 12158 9160 12164 9172
rect 11940 9132 12164 9160
rect 11940 9120 11946 9132
rect 12158 9120 12164 9132
rect 12216 9120 12222 9172
rect 9217 9095 9275 9101
rect 9217 9061 9229 9095
rect 9263 9092 9275 9095
rect 9398 9092 9404 9104
rect 9263 9064 9404 9092
rect 9263 9061 9275 9064
rect 9217 9055 9275 9061
rect 7576 8996 8123 9024
rect 6641 8959 6699 8965
rect 6641 8925 6653 8959
rect 6687 8925 6699 8959
rect 6641 8919 6699 8925
rect 6730 8916 6736 8968
rect 6788 8956 6794 8968
rect 7576 8965 7604 8996
rect 6917 8959 6975 8965
rect 6917 8956 6929 8959
rect 6788 8928 6929 8956
rect 6788 8916 6794 8928
rect 6917 8925 6929 8928
rect 6963 8925 6975 8959
rect 6917 8919 6975 8925
rect 7561 8959 7619 8965
rect 7561 8925 7573 8959
rect 7607 8925 7619 8959
rect 7561 8919 7619 8925
rect 7190 8888 7196 8900
rect 6564 8860 7196 8888
rect 7190 8848 7196 8860
rect 7248 8848 7254 8900
rect 7285 8891 7343 8897
rect 7285 8857 7297 8891
rect 7331 8888 7343 8891
rect 7374 8888 7380 8900
rect 7331 8860 7380 8888
rect 7331 8857 7343 8860
rect 7285 8851 7343 8857
rect 7374 8848 7380 8860
rect 7432 8888 7438 8900
rect 7576 8888 7604 8919
rect 7834 8916 7840 8968
rect 7892 8950 7898 8968
rect 8095 8965 8123 8996
rect 8386 8984 8392 9036
rect 8444 9024 8450 9036
rect 9232 9024 9260 9055
rect 9398 9052 9404 9064
rect 9456 9052 9462 9104
rect 9674 9052 9680 9104
rect 9732 9092 9738 9104
rect 9732 9064 9904 9092
rect 9732 9052 9738 9064
rect 9765 9027 9823 9033
rect 9765 9024 9777 9027
rect 8444 8996 9260 9024
rect 9416 8996 9777 9024
rect 8444 8984 8450 8996
rect 8496 8965 8524 8996
rect 7929 8959 7987 8965
rect 7929 8950 7941 8959
rect 7892 8925 7941 8950
rect 7975 8925 7987 8959
rect 7892 8922 7987 8925
rect 7892 8916 7898 8922
rect 7929 8919 7987 8922
rect 8080 8959 8138 8965
rect 8080 8925 8092 8959
rect 8126 8956 8138 8959
rect 8205 8959 8263 8965
rect 8126 8928 8160 8956
rect 8126 8925 8138 8928
rect 8080 8919 8138 8925
rect 8205 8925 8217 8959
rect 8251 8925 8263 8959
rect 8205 8919 8263 8925
rect 8297 8959 8355 8965
rect 8297 8925 8309 8959
rect 8343 8956 8355 8959
rect 8481 8959 8539 8965
rect 8343 8928 8432 8956
rect 8343 8925 8355 8928
rect 8297 8919 8355 8925
rect 8219 8888 8247 8919
rect 7432 8860 7604 8888
rect 8036 8860 8247 8888
rect 8404 8888 8432 8928
rect 8481 8925 8493 8959
rect 8527 8956 8539 8959
rect 8665 8959 8723 8965
rect 8527 8928 8561 8956
rect 8527 8925 8539 8928
rect 8481 8919 8539 8925
rect 8665 8925 8677 8959
rect 8711 8956 8723 8959
rect 8846 8956 8852 8968
rect 8711 8928 8852 8956
rect 8711 8925 8723 8928
rect 8665 8919 8723 8925
rect 8680 8888 8708 8919
rect 8846 8916 8852 8928
rect 8904 8916 8910 8968
rect 8938 8916 8944 8968
rect 8996 8956 9002 8968
rect 8996 8928 9041 8956
rect 8996 8916 9002 8928
rect 9122 8916 9128 8968
rect 9180 8956 9186 8968
rect 9180 8928 9225 8956
rect 9180 8916 9186 8928
rect 8404 8860 8708 8888
rect 8757 8891 8815 8897
rect 7432 8848 7438 8860
rect 2774 8780 2780 8832
rect 2832 8820 2838 8832
rect 3421 8823 3479 8829
rect 3421 8820 3433 8823
rect 2832 8792 3433 8820
rect 2832 8780 2838 8792
rect 3421 8789 3433 8792
rect 3467 8789 3479 8823
rect 3421 8783 3479 8789
rect 3970 8780 3976 8832
rect 4028 8820 4034 8832
rect 4893 8823 4951 8829
rect 4893 8820 4905 8823
rect 4028 8792 4905 8820
rect 4028 8780 4034 8792
rect 4893 8789 4905 8792
rect 4939 8789 4951 8823
rect 4893 8783 4951 8789
rect 7098 8780 7104 8832
rect 7156 8820 7162 8832
rect 8036 8820 8064 8860
rect 8757 8857 8769 8891
rect 8803 8888 8815 8891
rect 9416 8888 9444 8996
rect 9765 8993 9777 8996
rect 9811 8993 9823 9027
rect 9765 8987 9823 8993
rect 9490 8916 9496 8968
rect 9548 8956 9554 8968
rect 9585 8959 9643 8965
rect 9585 8956 9597 8959
rect 9548 8928 9597 8956
rect 9548 8916 9554 8928
rect 9585 8925 9597 8928
rect 9631 8925 9643 8959
rect 9585 8919 9643 8925
rect 9677 8959 9735 8965
rect 9677 8925 9689 8959
rect 9723 8925 9735 8959
rect 9677 8919 9735 8925
rect 9692 8888 9720 8919
rect 9780 8900 9808 8987
rect 9876 8965 9904 9064
rect 10778 9052 10784 9104
rect 10836 9092 10842 9104
rect 11146 9101 11152 9104
rect 11057 9095 11115 9101
rect 11057 9092 11069 9095
rect 10836 9064 11069 9092
rect 10836 9052 10842 9064
rect 11057 9061 11069 9064
rect 11103 9061 11115 9095
rect 11057 9055 11115 9061
rect 11145 9055 11152 9101
rect 11204 9092 11210 9104
rect 11204 9064 11245 9092
rect 11146 9052 11152 9055
rect 11204 9052 11210 9064
rect 10045 9027 10103 9033
rect 10045 8993 10057 9027
rect 10091 9024 10103 9027
rect 10091 8996 12020 9024
rect 10091 8993 10103 8996
rect 10045 8987 10103 8993
rect 9861 8959 9919 8965
rect 9861 8925 9873 8959
rect 9907 8925 9919 8959
rect 9861 8919 9919 8925
rect 10226 8916 10232 8968
rect 10284 8956 10290 8968
rect 10321 8959 10379 8965
rect 10321 8956 10333 8959
rect 10284 8928 10333 8956
rect 10284 8916 10290 8928
rect 10321 8925 10333 8928
rect 10367 8925 10379 8959
rect 10321 8919 10379 8925
rect 10410 8916 10416 8968
rect 10468 8956 10474 8968
rect 10505 8959 10563 8965
rect 10505 8956 10517 8959
rect 10468 8928 10517 8956
rect 10468 8916 10474 8928
rect 10505 8925 10517 8928
rect 10551 8956 10563 8959
rect 10778 8956 10784 8968
rect 10551 8928 10784 8956
rect 10551 8925 10563 8928
rect 10505 8919 10563 8925
rect 10778 8916 10784 8928
rect 10836 8916 10842 8968
rect 10870 8916 10876 8968
rect 10928 8956 10934 8968
rect 10965 8959 11023 8965
rect 10965 8956 10977 8959
rect 10928 8928 10977 8956
rect 10928 8916 10934 8928
rect 10965 8925 10977 8928
rect 11011 8925 11023 8959
rect 10965 8919 11023 8925
rect 11054 8916 11060 8968
rect 11112 8956 11118 8968
rect 11241 8959 11299 8965
rect 11241 8956 11253 8959
rect 11112 8928 11253 8956
rect 11112 8916 11118 8928
rect 11241 8925 11253 8928
rect 11287 8925 11299 8959
rect 11241 8919 11299 8925
rect 11330 8916 11336 8968
rect 11388 8956 11394 8968
rect 11992 8965 12020 8996
rect 11609 8959 11667 8965
rect 11609 8956 11621 8959
rect 11388 8928 11621 8956
rect 11388 8916 11394 8928
rect 11609 8925 11621 8928
rect 11655 8925 11667 8959
rect 11609 8919 11667 8925
rect 11977 8959 12035 8965
rect 11977 8925 11989 8959
rect 12023 8956 12035 8959
rect 12986 8956 12992 8968
rect 12023 8928 12992 8956
rect 12023 8925 12035 8928
rect 11977 8919 12035 8925
rect 12986 8916 12992 8928
rect 13044 8916 13050 8968
rect 13262 8956 13268 8968
rect 13223 8928 13268 8956
rect 13262 8916 13268 8928
rect 13320 8916 13326 8968
rect 8803 8860 9444 8888
rect 9646 8860 9720 8888
rect 8803 8857 8815 8860
rect 8757 8851 8815 8857
rect 7156 8792 8064 8820
rect 7156 8780 7162 8792
rect 8110 8780 8116 8832
rect 8168 8820 8174 8832
rect 8294 8820 8300 8832
rect 8168 8792 8300 8820
rect 8168 8780 8174 8792
rect 8294 8780 8300 8792
rect 8352 8780 8358 8832
rect 8570 8780 8576 8832
rect 8628 8820 8634 8832
rect 9398 8820 9404 8832
rect 8628 8792 9404 8820
rect 8628 8780 8634 8792
rect 9398 8780 9404 8792
rect 9456 8820 9462 8832
rect 9646 8820 9674 8860
rect 9766 8848 9772 8900
rect 9824 8848 9830 8900
rect 10594 8848 10600 8900
rect 10652 8888 10658 8900
rect 11146 8888 11152 8900
rect 10652 8860 11152 8888
rect 10652 8848 10658 8860
rect 11146 8848 11152 8860
rect 11204 8888 11210 8900
rect 11422 8888 11428 8900
rect 11204 8860 11428 8888
rect 11204 8848 11210 8860
rect 11422 8848 11428 8860
rect 11480 8848 11486 8900
rect 13354 8848 13360 8900
rect 13412 8888 13418 8900
rect 13541 8891 13599 8897
rect 13541 8888 13553 8891
rect 13412 8860 13553 8888
rect 13412 8848 13418 8860
rect 13541 8857 13553 8860
rect 13587 8857 13599 8891
rect 13541 8851 13599 8857
rect 10502 8820 10508 8832
rect 9456 8792 9674 8820
rect 10463 8792 10508 8820
rect 9456 8780 9462 8792
rect 10502 8780 10508 8792
rect 10560 8780 10566 8832
rect 11054 8780 11060 8832
rect 11112 8820 11118 8832
rect 11793 8823 11851 8829
rect 11793 8820 11805 8823
rect 11112 8792 11805 8820
rect 11112 8780 11118 8792
rect 11793 8789 11805 8792
rect 11839 8789 11851 8823
rect 11793 8783 11851 8789
rect 12066 8780 12072 8832
rect 12124 8820 12130 8832
rect 12342 8820 12348 8832
rect 12124 8792 12348 8820
rect 12124 8780 12130 8792
rect 12342 8780 12348 8792
rect 12400 8780 12406 8832
rect 1104 8730 13892 8752
rect 1104 8678 8214 8730
rect 8266 8678 8278 8730
rect 8330 8678 8342 8730
rect 8394 8678 8406 8730
rect 8458 8678 8470 8730
rect 8522 8678 13892 8730
rect 1104 8656 13892 8678
rect 1581 8619 1639 8625
rect 1581 8585 1593 8619
rect 1627 8585 1639 8619
rect 1854 8616 1860 8628
rect 1815 8588 1860 8616
rect 1581 8579 1639 8585
rect 1596 8548 1624 8579
rect 1854 8576 1860 8588
rect 1912 8576 1918 8628
rect 2682 8616 2688 8628
rect 2148 8588 2688 8616
rect 2148 8548 2176 8588
rect 2682 8576 2688 8588
rect 2740 8576 2746 8628
rect 2866 8576 2872 8628
rect 2924 8616 2930 8628
rect 2961 8619 3019 8625
rect 2961 8616 2973 8619
rect 2924 8588 2973 8616
rect 2924 8576 2930 8588
rect 2961 8585 2973 8588
rect 3007 8585 3019 8619
rect 2961 8579 3019 8585
rect 6270 8576 6276 8628
rect 6328 8616 6334 8628
rect 6546 8616 6552 8628
rect 6328 8588 6552 8616
rect 6328 8576 6334 8588
rect 6546 8576 6552 8588
rect 6604 8576 6610 8628
rect 7006 8576 7012 8628
rect 7064 8616 7070 8628
rect 7064 8588 7788 8616
rect 7064 8576 7070 8588
rect 2590 8548 2596 8560
rect 1596 8520 2176 8548
rect 2332 8520 2596 8548
rect 1397 8483 1455 8489
rect 1397 8449 1409 8483
rect 1443 8449 1455 8483
rect 1670 8480 1676 8492
rect 1631 8452 1676 8480
rect 1397 8443 1455 8449
rect 1412 8344 1440 8443
rect 1670 8440 1676 8452
rect 1728 8440 1734 8492
rect 1762 8440 1768 8492
rect 1820 8480 1826 8492
rect 2332 8489 2360 8520
rect 2590 8508 2596 8520
rect 2648 8548 2654 8560
rect 3510 8548 3516 8560
rect 2648 8520 3280 8548
rect 3471 8520 3516 8548
rect 2648 8508 2654 8520
rect 2498 8489 2504 8492
rect 2041 8483 2099 8489
rect 2041 8480 2053 8483
rect 1820 8452 2053 8480
rect 1820 8440 1826 8452
rect 2041 8449 2053 8452
rect 2087 8449 2099 8483
rect 2041 8443 2099 8449
rect 2225 8483 2283 8489
rect 2225 8449 2237 8483
rect 2271 8449 2283 8483
rect 2225 8443 2283 8449
rect 2317 8483 2375 8489
rect 2317 8449 2329 8483
rect 2363 8449 2375 8483
rect 2317 8443 2375 8449
rect 2443 8483 2504 8489
rect 2443 8449 2455 8483
rect 2489 8449 2504 8483
rect 2443 8443 2504 8449
rect 1946 8372 1952 8424
rect 2004 8412 2010 8424
rect 2240 8412 2268 8443
rect 2498 8440 2504 8443
rect 2556 8480 2562 8492
rect 3252 8489 3280 8520
rect 3510 8508 3516 8520
rect 3568 8508 3574 8560
rect 3602 8508 3608 8560
rect 3660 8548 3666 8560
rect 5626 8548 5632 8560
rect 3660 8520 3705 8548
rect 5587 8520 5632 8548
rect 3660 8508 3666 8520
rect 5626 8508 5632 8520
rect 5684 8508 5690 8560
rect 6181 8551 6239 8557
rect 6181 8517 6193 8551
rect 6227 8548 6239 8551
rect 6638 8548 6644 8560
rect 6227 8520 6644 8548
rect 6227 8517 6239 8520
rect 6181 8511 6239 8517
rect 6638 8508 6644 8520
rect 6696 8508 6702 8560
rect 6917 8551 6975 8557
rect 6917 8517 6929 8551
rect 6963 8548 6975 8551
rect 6963 8520 7696 8548
rect 6963 8517 6975 8520
rect 6917 8511 6975 8517
rect 3237 8483 3295 8489
rect 2556 8452 3096 8480
rect 2556 8440 2562 8452
rect 2869 8415 2927 8421
rect 2869 8412 2881 8415
rect 2004 8384 2881 8412
rect 2004 8372 2010 8384
rect 2869 8381 2881 8384
rect 2915 8381 2927 8415
rect 3068 8412 3096 8452
rect 3237 8449 3249 8483
rect 3283 8449 3295 8483
rect 3237 8443 3295 8449
rect 3694 8440 3700 8492
rect 3752 8440 3758 8492
rect 3970 8440 3976 8492
rect 4028 8480 4034 8492
rect 4433 8483 4491 8489
rect 4028 8452 4200 8480
rect 4028 8440 4034 8452
rect 3421 8415 3479 8421
rect 3421 8412 3433 8415
rect 3068 8384 3433 8412
rect 2869 8375 2927 8381
rect 3421 8381 3433 8384
rect 3467 8381 3479 8415
rect 3712 8412 3740 8440
rect 4065 8415 4123 8421
rect 4065 8412 4077 8415
rect 3712 8384 4077 8412
rect 3421 8375 3479 8381
rect 4065 8381 4077 8384
rect 4111 8381 4123 8415
rect 4172 8412 4200 8452
rect 4433 8449 4445 8483
rect 4479 8480 4491 8483
rect 4522 8480 4528 8492
rect 4479 8452 4528 8480
rect 4479 8449 4491 8452
rect 4433 8443 4491 8449
rect 4522 8440 4528 8452
rect 4580 8440 4586 8492
rect 4798 8480 4804 8492
rect 4759 8452 4804 8480
rect 4798 8440 4804 8452
rect 4856 8440 4862 8492
rect 5074 8480 5080 8492
rect 5035 8452 5080 8480
rect 5074 8440 5080 8452
rect 5132 8440 5138 8492
rect 5169 8483 5227 8489
rect 5169 8449 5181 8483
rect 5215 8480 5227 8483
rect 5534 8480 5540 8492
rect 5215 8452 5540 8480
rect 5215 8449 5227 8452
rect 5169 8443 5227 8449
rect 5534 8440 5540 8452
rect 5592 8440 5598 8492
rect 5810 8480 5816 8492
rect 5771 8452 5816 8480
rect 5810 8440 5816 8452
rect 5868 8440 5874 8492
rect 6086 8480 6092 8492
rect 6047 8452 6092 8480
rect 6086 8440 6092 8452
rect 6144 8440 6150 8492
rect 6549 8483 6607 8489
rect 6549 8449 6561 8483
rect 6595 8449 6607 8483
rect 6730 8480 6736 8492
rect 6691 8452 6736 8480
rect 6549 8443 6607 8449
rect 4617 8415 4675 8421
rect 4617 8412 4629 8415
rect 4172 8384 4629 8412
rect 4065 8375 4123 8381
rect 4617 8381 4629 8384
rect 4663 8381 4675 8415
rect 4617 8375 4675 8381
rect 4706 8372 4712 8424
rect 4764 8412 4770 8424
rect 5721 8415 5779 8421
rect 4764 8384 4809 8412
rect 4764 8372 4770 8384
rect 5721 8381 5733 8415
rect 5767 8381 5779 8415
rect 5828 8412 5856 8440
rect 6365 8415 6423 8421
rect 6365 8412 6377 8415
rect 5828 8384 6377 8412
rect 5721 8375 5779 8381
rect 6365 8381 6377 8384
rect 6411 8381 6423 8415
rect 6564 8412 6592 8443
rect 6730 8440 6736 8452
rect 6788 8440 6794 8492
rect 7098 8480 7104 8492
rect 6840 8452 7104 8480
rect 6840 8412 6868 8452
rect 7098 8440 7104 8452
rect 7156 8440 7162 8492
rect 7668 8489 7696 8520
rect 7377 8483 7435 8489
rect 7377 8449 7389 8483
rect 7423 8449 7435 8483
rect 7377 8443 7435 8449
rect 7653 8483 7711 8489
rect 7653 8449 7665 8483
rect 7699 8449 7711 8483
rect 7760 8480 7788 8588
rect 7834 8576 7840 8628
rect 7892 8616 7898 8628
rect 8110 8616 8116 8628
rect 7892 8588 8116 8616
rect 7892 8576 7898 8588
rect 8110 8576 8116 8588
rect 8168 8576 8174 8628
rect 8570 8576 8576 8628
rect 8628 8616 8634 8628
rect 8941 8619 8999 8625
rect 8941 8616 8953 8619
rect 8628 8588 8953 8616
rect 8628 8576 8634 8588
rect 8941 8585 8953 8588
rect 8987 8585 8999 8619
rect 10318 8616 10324 8628
rect 8941 8579 8999 8585
rect 9048 8588 10324 8616
rect 7926 8508 7932 8560
rect 7984 8548 7990 8560
rect 9048 8548 9076 8588
rect 10318 8576 10324 8588
rect 10376 8576 10382 8628
rect 10502 8576 10508 8628
rect 10560 8616 10566 8628
rect 10560 8588 12480 8616
rect 10560 8576 10566 8588
rect 9953 8551 10011 8557
rect 9953 8548 9965 8551
rect 7984 8520 9076 8548
rect 9508 8520 9965 8548
rect 7984 8508 7990 8520
rect 8496 8489 8524 8520
rect 9508 8492 9536 8520
rect 9953 8517 9965 8520
rect 9999 8517 10011 8551
rect 9953 8511 10011 8517
rect 10137 8551 10195 8557
rect 10137 8517 10149 8551
rect 10183 8548 10195 8551
rect 10410 8548 10416 8560
rect 10183 8520 10416 8548
rect 10183 8517 10195 8520
rect 10137 8511 10195 8517
rect 10410 8508 10416 8520
rect 10468 8508 10474 8560
rect 10870 8508 10876 8560
rect 10928 8548 10934 8560
rect 12452 8557 12480 8588
rect 11701 8551 11759 8557
rect 11701 8548 11713 8551
rect 10928 8520 11713 8548
rect 10928 8508 10934 8520
rect 11701 8517 11713 8520
rect 11747 8517 11759 8551
rect 11701 8511 11759 8517
rect 11793 8551 11851 8557
rect 11793 8517 11805 8551
rect 11839 8548 11851 8551
rect 12437 8551 12495 8557
rect 11839 8520 12388 8548
rect 11839 8517 11851 8520
rect 11793 8511 11851 8517
rect 7837 8483 7895 8489
rect 7837 8480 7849 8483
rect 7760 8452 7849 8480
rect 7653 8443 7711 8449
rect 7837 8449 7849 8452
rect 7883 8449 7895 8483
rect 7837 8443 7895 8449
rect 8389 8483 8447 8489
rect 8389 8449 8401 8483
rect 8435 8449 8447 8483
rect 8389 8443 8447 8449
rect 8481 8483 8539 8489
rect 8481 8449 8493 8483
rect 8527 8449 8539 8483
rect 8481 8443 8539 8449
rect 8849 8483 8907 8489
rect 8849 8449 8861 8483
rect 8895 8480 8907 8483
rect 9030 8480 9036 8492
rect 8895 8452 9036 8480
rect 8895 8449 8907 8452
rect 8849 8443 8907 8449
rect 7006 8412 7012 8424
rect 6564 8384 6868 8412
rect 6967 8384 7012 8412
rect 6365 8375 6423 8381
rect 1412 8316 2360 8344
rect 2332 8276 2360 8316
rect 2406 8304 2412 8356
rect 2464 8344 2470 8356
rect 2685 8347 2743 8353
rect 2685 8344 2697 8347
rect 2464 8316 2697 8344
rect 2464 8304 2470 8316
rect 2685 8313 2697 8316
rect 2731 8313 2743 8347
rect 3326 8344 3332 8356
rect 2685 8307 2743 8313
rect 2792 8316 3332 8344
rect 2792 8276 2820 8316
rect 3326 8304 3332 8316
rect 3384 8304 3390 8356
rect 3694 8304 3700 8356
rect 3752 8344 3758 8356
rect 4249 8347 4307 8353
rect 4249 8344 4261 8347
rect 3752 8316 4261 8344
rect 3752 8304 3758 8316
rect 4249 8313 4261 8316
rect 4295 8313 4307 8347
rect 5736 8344 5764 8375
rect 5810 8344 5816 8356
rect 5736 8316 5816 8344
rect 4249 8307 4307 8313
rect 5810 8304 5816 8316
rect 5868 8304 5874 8356
rect 2332 8248 2820 8276
rect 6380 8276 6408 8375
rect 7006 8372 7012 8384
rect 7064 8372 7070 8424
rect 7098 8344 7104 8356
rect 7059 8316 7104 8344
rect 7098 8304 7104 8316
rect 7156 8304 7162 8356
rect 7392 8344 7420 8443
rect 7558 8412 7564 8424
rect 7519 8384 7564 8412
rect 7558 8372 7564 8384
rect 7616 8372 7622 8424
rect 7926 8344 7932 8356
rect 7392 8316 7932 8344
rect 7926 8304 7932 8316
rect 7984 8304 7990 8356
rect 8202 8344 8208 8356
rect 8163 8316 8208 8344
rect 8202 8304 8208 8316
rect 8260 8304 8266 8356
rect 8110 8276 8116 8288
rect 6380 8248 8116 8276
rect 8110 8236 8116 8248
rect 8168 8276 8174 8288
rect 8404 8276 8432 8443
rect 9030 8440 9036 8452
rect 9088 8440 9094 8492
rect 9125 8483 9183 8489
rect 9125 8449 9137 8483
rect 9171 8449 9183 8483
rect 9306 8480 9312 8492
rect 9267 8452 9312 8480
rect 9125 8443 9183 8449
rect 8662 8372 8668 8424
rect 8720 8372 8726 8424
rect 8938 8372 8944 8424
rect 8996 8412 9002 8424
rect 9140 8412 9168 8443
rect 9306 8440 9312 8452
rect 9364 8440 9370 8492
rect 9401 8483 9459 8489
rect 9401 8449 9413 8483
rect 9447 8480 9459 8483
rect 9490 8480 9496 8492
rect 9447 8452 9496 8480
rect 9447 8449 9459 8452
rect 9401 8443 9459 8449
rect 9490 8440 9496 8452
rect 9548 8440 9554 8492
rect 9585 8483 9643 8489
rect 9585 8449 9597 8483
rect 9631 8449 9643 8483
rect 9585 8443 9643 8449
rect 8996 8384 9168 8412
rect 9600 8412 9628 8443
rect 9766 8440 9772 8492
rect 9824 8480 9830 8492
rect 10597 8483 10655 8489
rect 10597 8480 10609 8483
rect 9824 8452 10609 8480
rect 9824 8440 9830 8452
rect 10597 8449 10609 8452
rect 10643 8449 10655 8483
rect 10597 8443 10655 8449
rect 10686 8440 10692 8492
rect 10744 8480 10750 8492
rect 10781 8483 10839 8489
rect 10781 8480 10793 8483
rect 10744 8452 10793 8480
rect 10744 8440 10750 8452
rect 10781 8449 10793 8452
rect 10827 8449 10839 8483
rect 11054 8480 11060 8492
rect 11015 8452 11060 8480
rect 10781 8443 10839 8449
rect 11054 8440 11060 8452
rect 11112 8440 11118 8492
rect 11146 8440 11152 8492
rect 11204 8480 11210 8492
rect 11241 8483 11299 8489
rect 11241 8480 11253 8483
rect 11204 8452 11253 8480
rect 11204 8440 11210 8452
rect 11241 8449 11253 8452
rect 11287 8449 11299 8483
rect 11514 8480 11520 8492
rect 11475 8452 11520 8480
rect 11241 8443 11299 8449
rect 11514 8440 11520 8452
rect 11572 8440 11578 8492
rect 11606 8440 11612 8492
rect 11664 8480 11670 8492
rect 11808 8480 11836 8511
rect 11664 8452 11836 8480
rect 11937 8483 11995 8489
rect 11664 8440 11670 8452
rect 11937 8449 11949 8483
rect 11983 8480 11995 8483
rect 12253 8483 12311 8489
rect 11983 8452 12204 8480
rect 11983 8449 11995 8452
rect 11937 8443 11995 8449
rect 9858 8412 9864 8424
rect 9600 8384 9864 8412
rect 8996 8372 9002 8384
rect 8680 8285 8708 8372
rect 9140 8344 9168 8384
rect 9858 8372 9864 8384
rect 9916 8372 9922 8424
rect 11422 8412 11428 8424
rect 9968 8384 11428 8412
rect 9968 8344 9996 8384
rect 11422 8372 11428 8384
rect 11480 8372 11486 8424
rect 10597 8347 10655 8353
rect 10597 8344 10609 8347
rect 9140 8316 9996 8344
rect 10152 8316 10609 8344
rect 8168 8248 8432 8276
rect 8665 8279 8723 8285
rect 8168 8236 8174 8248
rect 8665 8245 8677 8279
rect 8711 8245 8723 8279
rect 8665 8239 8723 8245
rect 9122 8236 9128 8288
rect 9180 8276 9186 8288
rect 9582 8276 9588 8288
rect 9180 8248 9588 8276
rect 9180 8236 9186 8248
rect 9582 8236 9588 8248
rect 9640 8236 9646 8288
rect 9766 8276 9772 8288
rect 9727 8248 9772 8276
rect 9766 8236 9772 8248
rect 9824 8236 9830 8288
rect 10042 8236 10048 8288
rect 10100 8276 10106 8288
rect 10152 8285 10180 8316
rect 10597 8313 10609 8316
rect 10643 8313 10655 8347
rect 11238 8344 11244 8356
rect 11199 8316 11244 8344
rect 10597 8307 10655 8313
rect 11238 8304 11244 8316
rect 11296 8304 11302 8356
rect 12066 8344 12072 8356
rect 12027 8316 12072 8344
rect 12066 8304 12072 8316
rect 12124 8304 12130 8356
rect 12176 8344 12204 8452
rect 12253 8449 12265 8483
rect 12299 8449 12311 8483
rect 12360 8480 12388 8520
rect 12437 8517 12449 8551
rect 12483 8517 12495 8551
rect 13538 8548 13544 8560
rect 13499 8520 13544 8548
rect 12437 8511 12495 8517
rect 13538 8508 13544 8520
rect 13596 8508 13602 8560
rect 12710 8489 12716 8492
rect 12529 8483 12587 8489
rect 12529 8480 12541 8483
rect 12360 8452 12541 8480
rect 12253 8443 12311 8449
rect 12529 8449 12541 8452
rect 12575 8449 12587 8483
rect 12529 8443 12587 8449
rect 12673 8483 12716 8489
rect 12673 8449 12685 8483
rect 12768 8480 12774 8492
rect 13446 8480 13452 8492
rect 12768 8452 13452 8480
rect 12673 8443 12716 8449
rect 12268 8412 12296 8443
rect 12710 8440 12716 8443
rect 12768 8440 12774 8452
rect 13446 8440 13452 8452
rect 13504 8440 13510 8492
rect 12342 8412 12348 8424
rect 12268 8384 12348 8412
rect 12342 8372 12348 8384
rect 12400 8372 12406 8424
rect 12986 8412 12992 8424
rect 12947 8384 12992 8412
rect 12986 8372 12992 8384
rect 13044 8372 13050 8424
rect 13262 8344 13268 8356
rect 12176 8316 13268 8344
rect 13262 8304 13268 8316
rect 13320 8304 13326 8356
rect 13354 8304 13360 8356
rect 13412 8344 13418 8356
rect 13449 8347 13507 8353
rect 13449 8344 13461 8347
rect 13412 8316 13461 8344
rect 13412 8304 13418 8316
rect 13449 8313 13461 8316
rect 13495 8313 13507 8347
rect 13449 8307 13507 8313
rect 10137 8279 10195 8285
rect 10137 8276 10149 8279
rect 10100 8248 10149 8276
rect 10100 8236 10106 8248
rect 10137 8245 10149 8248
rect 10183 8245 10195 8279
rect 10318 8276 10324 8288
rect 10279 8248 10324 8276
rect 10137 8239 10195 8245
rect 10318 8236 10324 8248
rect 10376 8236 10382 8288
rect 12158 8236 12164 8288
rect 12216 8276 12222 8288
rect 12618 8276 12624 8288
rect 12216 8248 12624 8276
rect 12216 8236 12222 8248
rect 12618 8236 12624 8248
rect 12676 8236 12682 8288
rect 12802 8276 12808 8288
rect 12763 8248 12808 8276
rect 12802 8236 12808 8248
rect 12860 8236 12866 8288
rect 1104 8186 13892 8208
rect 1104 8134 4214 8186
rect 4266 8134 4278 8186
rect 4330 8134 4342 8186
rect 4394 8134 4406 8186
rect 4458 8134 4470 8186
rect 4522 8134 12214 8186
rect 12266 8134 12278 8186
rect 12330 8134 12342 8186
rect 12394 8134 12406 8186
rect 12458 8134 12470 8186
rect 12522 8134 13892 8186
rect 1104 8112 13892 8134
rect 2038 8032 2044 8084
rect 2096 8072 2102 8084
rect 2590 8072 2596 8084
rect 2096 8044 2596 8072
rect 2096 8032 2102 8044
rect 2590 8032 2596 8044
rect 2648 8032 2654 8084
rect 3513 8075 3571 8081
rect 3513 8041 3525 8075
rect 3559 8072 3571 8075
rect 4890 8072 4896 8084
rect 3559 8044 4896 8072
rect 3559 8041 3571 8044
rect 3513 8035 3571 8041
rect 4890 8032 4896 8044
rect 4948 8032 4954 8084
rect 5810 8032 5816 8084
rect 5868 8072 5874 8084
rect 6181 8075 6239 8081
rect 5868 8044 5913 8072
rect 5868 8032 5874 8044
rect 6181 8041 6193 8075
rect 6227 8072 6239 8075
rect 7006 8072 7012 8084
rect 6227 8044 7012 8072
rect 6227 8041 6239 8044
rect 6181 8035 6239 8041
rect 7006 8032 7012 8044
rect 7064 8032 7070 8084
rect 7834 8032 7840 8084
rect 7892 8072 7898 8084
rect 8570 8072 8576 8084
rect 7892 8044 8576 8072
rect 7892 8032 7898 8044
rect 8570 8032 8576 8044
rect 8628 8032 8634 8084
rect 9861 8075 9919 8081
rect 9861 8041 9873 8075
rect 9907 8072 9919 8075
rect 10042 8072 10048 8084
rect 9907 8044 10048 8072
rect 9907 8041 9919 8044
rect 9861 8035 9919 8041
rect 10042 8032 10048 8044
rect 10100 8032 10106 8084
rect 10134 8032 10140 8084
rect 10192 8032 10198 8084
rect 10226 8032 10232 8084
rect 10284 8072 10290 8084
rect 10689 8075 10747 8081
rect 10284 8044 10548 8072
rect 10284 8032 10290 8044
rect 3053 8007 3111 8013
rect 3053 7973 3065 8007
rect 3099 8004 3111 8007
rect 8846 8004 8852 8016
rect 3099 7976 8852 8004
rect 3099 7973 3111 7976
rect 3053 7967 3111 7973
rect 8846 7964 8852 7976
rect 8904 7964 8910 8016
rect 10152 8004 10180 8032
rect 10410 8004 10416 8016
rect 8956 7976 10180 8004
rect 10244 7976 10416 8004
rect 1394 7896 1400 7948
rect 1452 7936 1458 7948
rect 2498 7936 2504 7948
rect 1452 7908 2504 7936
rect 1452 7896 1458 7908
rect 1670 7868 1676 7880
rect 1631 7840 1676 7868
rect 1670 7828 1676 7840
rect 1728 7828 1734 7880
rect 1946 7868 1952 7880
rect 1907 7840 1952 7868
rect 1946 7828 1952 7840
rect 2004 7828 2010 7880
rect 2038 7828 2044 7880
rect 2096 7868 2102 7880
rect 2240 7877 2268 7908
rect 2498 7896 2504 7908
rect 2556 7896 2562 7948
rect 3789 7939 3847 7945
rect 3789 7936 3801 7939
rect 2746 7908 3801 7936
rect 2225 7871 2283 7877
rect 2096 7840 2141 7868
rect 2096 7828 2102 7840
rect 2225 7837 2237 7871
rect 2271 7837 2283 7871
rect 2406 7868 2412 7880
rect 2367 7840 2412 7868
rect 2225 7831 2283 7837
rect 2406 7828 2412 7840
rect 2464 7828 2470 7880
rect 2590 7868 2596 7880
rect 2551 7840 2596 7868
rect 2590 7828 2596 7840
rect 2648 7868 2654 7880
rect 2746 7868 2774 7908
rect 3789 7905 3801 7908
rect 3835 7905 3847 7939
rect 4614 7936 4620 7948
rect 3789 7899 3847 7905
rect 4172 7908 4620 7936
rect 2648 7840 2774 7868
rect 2961 7871 3019 7877
rect 2648 7828 2654 7840
rect 2961 7837 2973 7871
rect 3007 7868 3019 7871
rect 3050 7868 3056 7880
rect 3007 7840 3056 7868
rect 3007 7837 3019 7840
rect 2961 7831 3019 7837
rect 3050 7828 3056 7840
rect 3108 7828 3114 7880
rect 3329 7871 3387 7877
rect 3329 7837 3341 7871
rect 3375 7868 3387 7871
rect 3694 7868 3700 7880
rect 3375 7840 3700 7868
rect 3375 7837 3387 7840
rect 3329 7831 3387 7837
rect 3694 7828 3700 7840
rect 3752 7828 3758 7880
rect 3970 7828 3976 7880
rect 4028 7868 4034 7880
rect 4172 7877 4200 7908
rect 4614 7896 4620 7908
rect 4672 7896 4678 7948
rect 4798 7896 4804 7948
rect 4856 7936 4862 7948
rect 5166 7936 5172 7948
rect 4856 7908 5172 7936
rect 4856 7896 4862 7908
rect 5166 7896 5172 7908
rect 5224 7936 5230 7948
rect 5445 7939 5503 7945
rect 5445 7936 5457 7939
rect 5224 7908 5457 7936
rect 5224 7896 5230 7908
rect 5445 7905 5457 7908
rect 5491 7905 5503 7939
rect 6730 7936 6736 7948
rect 5445 7899 5503 7905
rect 6380 7908 6736 7936
rect 4064 7871 4122 7877
rect 4064 7868 4076 7871
rect 4028 7840 4076 7868
rect 4028 7828 4034 7840
rect 4064 7837 4076 7840
rect 4110 7837 4122 7871
rect 4064 7831 4122 7837
rect 4157 7871 4215 7877
rect 4157 7837 4169 7871
rect 4203 7837 4215 7871
rect 4157 7831 4215 7837
rect 4246 7828 4252 7880
rect 4304 7868 4310 7880
rect 4433 7871 4491 7877
rect 4304 7840 4349 7868
rect 4304 7828 4310 7840
rect 4433 7837 4445 7871
rect 4479 7868 4491 7871
rect 4706 7868 4712 7880
rect 4479 7840 4712 7868
rect 4479 7837 4491 7840
rect 4433 7831 4491 7837
rect 4706 7828 4712 7840
rect 4764 7828 4770 7880
rect 5074 7828 5080 7880
rect 5132 7828 5138 7880
rect 5902 7828 5908 7880
rect 5960 7868 5966 7880
rect 6380 7877 6408 7908
rect 6730 7896 6736 7908
rect 6788 7896 6794 7948
rect 8202 7936 8208 7948
rect 6840 7908 8208 7936
rect 5997 7871 6055 7877
rect 5997 7868 6009 7871
rect 5960 7840 6009 7868
rect 5960 7828 5966 7840
rect 5997 7837 6009 7840
rect 6043 7837 6055 7871
rect 6365 7871 6423 7877
rect 6365 7868 6377 7871
rect 5997 7831 6055 7837
rect 6288 7840 6377 7868
rect 1762 7800 1768 7812
rect 1723 7772 1768 7800
rect 1762 7760 1768 7772
rect 1820 7760 1826 7812
rect 4890 7800 4896 7812
rect 4851 7772 4896 7800
rect 4890 7760 4896 7772
rect 4948 7760 4954 7812
rect 1486 7732 1492 7744
rect 1447 7704 1492 7732
rect 1486 7692 1492 7704
rect 1544 7692 1550 7744
rect 3605 7735 3663 7741
rect 3605 7701 3617 7735
rect 3651 7732 3663 7735
rect 4062 7732 4068 7744
rect 3651 7704 4068 7732
rect 3651 7701 3663 7704
rect 3605 7695 3663 7701
rect 4062 7692 4068 7704
rect 4120 7692 4126 7744
rect 4154 7692 4160 7744
rect 4212 7732 4218 7744
rect 6288 7732 6316 7840
rect 6365 7837 6377 7840
rect 6411 7837 6423 7871
rect 6365 7831 6423 7837
rect 6454 7828 6460 7880
rect 6512 7868 6518 7880
rect 6512 7840 6557 7868
rect 6512 7828 6518 7840
rect 6840 7812 6868 7908
rect 8202 7896 8208 7908
rect 8260 7896 8266 7948
rect 8570 7896 8576 7948
rect 8628 7936 8634 7948
rect 8956 7936 8984 7976
rect 9490 7936 9496 7948
rect 8628 7908 8984 7936
rect 9324 7908 9496 7936
rect 8628 7896 8634 7908
rect 7081 7871 7139 7877
rect 7081 7837 7093 7871
rect 7127 7868 7139 7871
rect 7282 7868 7288 7880
rect 7127 7840 7288 7868
rect 7127 7837 7139 7840
rect 7081 7831 7139 7837
rect 7282 7828 7288 7840
rect 7340 7828 7346 7880
rect 7377 7871 7435 7877
rect 7377 7837 7389 7871
rect 7423 7868 7435 7871
rect 7558 7868 7564 7880
rect 7423 7840 7564 7868
rect 7423 7837 7435 7840
rect 7377 7831 7435 7837
rect 7558 7828 7564 7840
rect 7616 7828 7622 7880
rect 7653 7871 7711 7877
rect 7653 7837 7665 7871
rect 7699 7837 7711 7871
rect 8326 7854 8892 7868
rect 7653 7831 7711 7837
rect 8312 7840 8892 7854
rect 6638 7800 6644 7812
rect 6599 7772 6644 7800
rect 6638 7760 6644 7772
rect 6696 7760 6702 7812
rect 6822 7800 6828 7812
rect 6783 7772 6828 7800
rect 6822 7760 6828 7772
rect 6880 7760 6886 7812
rect 7668 7800 7696 7831
rect 7926 7800 7932 7812
rect 7300 7772 7932 7800
rect 4212 7704 6316 7732
rect 4212 7692 4218 7704
rect 7006 7692 7012 7744
rect 7064 7732 7070 7744
rect 7300 7741 7328 7772
rect 7926 7760 7932 7772
rect 7984 7760 7990 7812
rect 8312 7800 8340 7840
rect 8036 7772 8340 7800
rect 8665 7803 8723 7809
rect 7193 7735 7251 7741
rect 7193 7732 7205 7735
rect 7064 7704 7205 7732
rect 7064 7692 7070 7704
rect 7193 7701 7205 7704
rect 7239 7701 7251 7735
rect 7193 7695 7251 7701
rect 7285 7735 7343 7741
rect 7285 7701 7297 7735
rect 7331 7701 7343 7735
rect 7285 7695 7343 7701
rect 7558 7692 7564 7744
rect 7616 7732 7622 7744
rect 8036 7732 8064 7772
rect 8665 7769 8677 7803
rect 8711 7800 8723 7803
rect 8754 7800 8760 7812
rect 8711 7772 8760 7800
rect 8711 7769 8723 7772
rect 8665 7763 8723 7769
rect 8754 7760 8760 7772
rect 8812 7760 8818 7812
rect 8864 7800 8892 7840
rect 9122 7828 9128 7880
rect 9180 7868 9186 7880
rect 9324 7877 9352 7908
rect 9490 7896 9496 7908
rect 9548 7896 9554 7948
rect 9309 7871 9367 7877
rect 9309 7868 9321 7871
rect 9180 7840 9321 7868
rect 9180 7828 9186 7840
rect 9309 7837 9321 7840
rect 9355 7837 9367 7871
rect 9309 7831 9367 7837
rect 9398 7828 9404 7880
rect 9456 7868 9462 7880
rect 9968 7877 9996 7976
rect 10244 7877 10272 7976
rect 10410 7964 10416 7976
rect 10468 7964 10474 8016
rect 9677 7871 9735 7877
rect 9456 7840 9501 7868
rect 9456 7828 9462 7840
rect 9677 7837 9689 7871
rect 9723 7837 9735 7871
rect 9677 7831 9735 7837
rect 9953 7871 10011 7877
rect 9953 7837 9965 7871
rect 9999 7837 10011 7871
rect 9953 7831 10011 7837
rect 10221 7871 10279 7877
rect 10221 7837 10233 7871
rect 10267 7837 10279 7871
rect 10520 7868 10548 8044
rect 10689 8041 10701 8075
rect 10735 8072 10747 8075
rect 12618 8072 12624 8084
rect 10735 8044 12624 8072
rect 10735 8041 10747 8044
rect 10689 8035 10747 8041
rect 12618 8032 12624 8044
rect 12676 8032 12682 8084
rect 13262 8032 13268 8084
rect 13320 8072 13326 8084
rect 13449 8075 13507 8081
rect 13449 8072 13461 8075
rect 13320 8044 13461 8072
rect 13320 8032 13326 8044
rect 13449 8041 13461 8044
rect 13495 8072 13507 8075
rect 13538 8072 13544 8084
rect 13495 8044 13544 8072
rect 13495 8041 13507 8044
rect 13449 8035 13507 8041
rect 13538 8032 13544 8044
rect 13596 8032 13602 8084
rect 10870 8004 10876 8016
rect 10831 7976 10876 8004
rect 10870 7964 10876 7976
rect 10928 7964 10934 8016
rect 11974 7964 11980 8016
rect 12032 8004 12038 8016
rect 12032 7976 12296 8004
rect 12032 7964 12038 7976
rect 12268 7948 12296 7976
rect 10686 7896 10692 7948
rect 10744 7936 10750 7948
rect 12158 7936 12164 7948
rect 10744 7908 11376 7936
rect 10744 7896 10750 7908
rect 11054 7868 11060 7880
rect 10221 7831 10279 7837
rect 10428 7840 10548 7868
rect 11015 7840 11060 7868
rect 10428 7834 10456 7840
rect 9490 7800 9496 7812
rect 8864 7772 9496 7800
rect 9490 7760 9496 7772
rect 9548 7760 9554 7812
rect 7616 7704 8064 7732
rect 7616 7692 7622 7704
rect 8202 7692 8208 7744
rect 8260 7732 8266 7744
rect 9030 7732 9036 7744
rect 8260 7704 9036 7732
rect 8260 7692 8266 7704
rect 9030 7692 9036 7704
rect 9088 7732 9094 7744
rect 9125 7735 9183 7741
rect 9125 7732 9137 7735
rect 9088 7704 9137 7732
rect 9088 7692 9094 7704
rect 9125 7701 9137 7704
rect 9171 7701 9183 7735
rect 9692 7732 9720 7831
rect 10336 7809 10456 7834
rect 11054 7828 11060 7840
rect 11112 7828 11118 7880
rect 11238 7868 11244 7880
rect 11199 7840 11244 7868
rect 11238 7828 11244 7840
rect 11296 7828 11302 7880
rect 11348 7877 11376 7908
rect 11532 7908 12164 7936
rect 11333 7871 11391 7877
rect 11333 7837 11345 7871
rect 11379 7837 11391 7871
rect 11333 7831 11391 7837
rect 11422 7828 11428 7880
rect 11480 7877 11486 7880
rect 11480 7871 11500 7877
rect 11488 7868 11500 7871
rect 11532 7868 11560 7908
rect 12158 7896 12164 7908
rect 12216 7896 12222 7948
rect 12250 7896 12256 7948
rect 12308 7896 12314 7948
rect 11488 7840 11573 7868
rect 11488 7837 11500 7840
rect 11480 7831 11500 7837
rect 11480 7828 11486 7831
rect 11606 7828 11612 7880
rect 11664 7868 11670 7880
rect 11885 7871 11943 7877
rect 11885 7868 11897 7871
rect 11664 7840 11897 7868
rect 11664 7828 11670 7840
rect 11885 7837 11897 7840
rect 11931 7837 11943 7871
rect 11885 7831 11943 7837
rect 11974 7828 11980 7880
rect 12032 7868 12038 7880
rect 12069 7871 12127 7877
rect 12069 7868 12081 7871
rect 12032 7840 12081 7868
rect 12032 7828 12038 7840
rect 12069 7837 12081 7840
rect 12115 7837 12127 7871
rect 12069 7831 12127 7837
rect 12437 7871 12495 7877
rect 12437 7837 12449 7871
rect 12483 7868 12495 7871
rect 12802 7868 12808 7880
rect 12483 7840 12808 7868
rect 12483 7837 12495 7840
rect 12437 7831 12495 7837
rect 12802 7828 12808 7840
rect 12860 7828 12866 7880
rect 13357 7871 13415 7877
rect 13357 7837 13369 7871
rect 13403 7868 13415 7871
rect 13446 7868 13452 7880
rect 13403 7840 13452 7868
rect 13403 7837 13415 7840
rect 13357 7831 13415 7837
rect 13446 7828 13452 7840
rect 13504 7828 13510 7880
rect 10321 7806 10456 7809
rect 10321 7803 10379 7806
rect 10321 7769 10333 7803
rect 10367 7769 10379 7803
rect 10686 7800 10692 7812
rect 10744 7809 10750 7812
rect 10656 7772 10692 7800
rect 10321 7763 10379 7769
rect 10686 7760 10692 7772
rect 10744 7763 10756 7809
rect 11698 7800 11704 7812
rect 11659 7772 11704 7800
rect 10744 7760 10750 7763
rect 11698 7760 11704 7772
rect 11756 7760 11762 7812
rect 11992 7800 12020 7828
rect 13170 7800 13176 7812
rect 11808 7772 12020 7800
rect 13131 7772 13176 7800
rect 9858 7732 9864 7744
rect 9692 7704 9864 7732
rect 9125 7695 9183 7701
rect 9858 7692 9864 7704
rect 9916 7732 9922 7744
rect 11808 7732 11836 7772
rect 13170 7760 13176 7772
rect 13228 7760 13234 7812
rect 11974 7732 11980 7744
rect 9916 7704 11836 7732
rect 11935 7704 11980 7732
rect 9916 7692 9922 7704
rect 11974 7692 11980 7704
rect 12032 7692 12038 7744
rect 1104 7642 13892 7664
rect 1104 7590 8214 7642
rect 8266 7590 8278 7642
rect 8330 7590 8342 7642
rect 8394 7590 8406 7642
rect 8458 7590 8470 7642
rect 8522 7590 13892 7642
rect 1104 7568 13892 7590
rect 3694 7528 3700 7540
rect 2332 7500 3700 7528
rect 1486 7420 1492 7472
rect 1544 7460 1550 7472
rect 1544 7432 2268 7460
rect 1544 7420 1550 7432
rect 1673 7395 1731 7401
rect 1673 7361 1685 7395
rect 1719 7361 1731 7395
rect 1673 7355 1731 7361
rect 1857 7395 1915 7401
rect 1857 7361 1869 7395
rect 1903 7392 1915 7395
rect 2130 7392 2136 7404
rect 1903 7364 2136 7392
rect 1903 7361 1915 7364
rect 1857 7355 1915 7361
rect 1688 7324 1716 7355
rect 2130 7352 2136 7364
rect 2188 7352 2194 7404
rect 2240 7401 2268 7432
rect 2332 7401 2360 7500
rect 3694 7488 3700 7500
rect 3752 7488 3758 7540
rect 4341 7531 4399 7537
rect 4341 7497 4353 7531
rect 4387 7528 4399 7531
rect 4614 7528 4620 7540
rect 4387 7500 4620 7528
rect 4387 7497 4399 7500
rect 4341 7491 4399 7497
rect 4614 7488 4620 7500
rect 4672 7488 4678 7540
rect 4706 7488 4712 7540
rect 4764 7528 4770 7540
rect 4764 7500 5488 7528
rect 4764 7488 4770 7500
rect 2866 7460 2872 7472
rect 2424 7432 2872 7460
rect 2424 7401 2452 7432
rect 2866 7420 2872 7432
rect 2924 7420 2930 7472
rect 2958 7420 2964 7472
rect 3016 7460 3022 7472
rect 3142 7460 3148 7472
rect 3016 7432 3061 7460
rect 3103 7432 3148 7460
rect 3016 7420 3022 7432
rect 3142 7420 3148 7432
rect 3200 7420 3206 7472
rect 4890 7460 4896 7472
rect 3712 7432 4896 7460
rect 2225 7395 2283 7401
rect 2225 7361 2237 7395
rect 2271 7361 2283 7395
rect 2225 7355 2283 7361
rect 2317 7395 2375 7401
rect 2317 7361 2329 7395
rect 2363 7361 2375 7395
rect 2317 7355 2375 7361
rect 2409 7395 2467 7401
rect 2409 7361 2421 7395
rect 2455 7361 2467 7395
rect 2409 7355 2467 7361
rect 2501 7395 2559 7401
rect 2501 7361 2513 7395
rect 2547 7392 2559 7395
rect 2590 7392 2596 7404
rect 2547 7364 2596 7392
rect 2547 7361 2559 7364
rect 2501 7355 2559 7361
rect 2590 7352 2596 7364
rect 2648 7352 2654 7404
rect 3712 7401 3740 7432
rect 4890 7420 4896 7432
rect 4948 7460 4954 7472
rect 4948 7432 5212 7460
rect 4948 7420 4954 7432
rect 3697 7395 3755 7401
rect 3697 7361 3709 7395
rect 3743 7361 3755 7395
rect 4706 7392 4712 7404
rect 4667 7364 4712 7392
rect 3697 7355 3755 7361
rect 4706 7352 4712 7364
rect 4764 7352 4770 7404
rect 5184 7401 5212 7432
rect 5460 7401 5488 7500
rect 5902 7488 5908 7540
rect 5960 7528 5966 7540
rect 6457 7531 6515 7537
rect 6457 7528 6469 7531
rect 5960 7500 6469 7528
rect 5960 7488 5966 7500
rect 6457 7497 6469 7500
rect 6503 7497 6515 7531
rect 6457 7491 6515 7497
rect 7650 7488 7656 7540
rect 7708 7528 7714 7540
rect 8021 7531 8079 7537
rect 8021 7528 8033 7531
rect 7708 7500 8033 7528
rect 7708 7488 7714 7500
rect 8021 7497 8033 7500
rect 8067 7497 8079 7531
rect 8021 7491 8079 7497
rect 9398 7488 9404 7540
rect 9456 7528 9462 7540
rect 9585 7531 9643 7537
rect 9585 7528 9597 7531
rect 9456 7500 9597 7528
rect 9456 7488 9462 7500
rect 9585 7497 9597 7500
rect 9631 7528 9643 7531
rect 9769 7531 9827 7537
rect 9769 7528 9781 7531
rect 9631 7500 9781 7528
rect 9631 7497 9643 7500
rect 9585 7491 9643 7497
rect 9769 7497 9781 7500
rect 9815 7497 9827 7531
rect 9769 7491 9827 7497
rect 9861 7531 9919 7537
rect 9861 7497 9873 7531
rect 9907 7528 9919 7531
rect 9950 7528 9956 7540
rect 9907 7500 9956 7528
rect 9907 7497 9919 7500
rect 9861 7491 9919 7497
rect 9950 7488 9956 7500
rect 10008 7488 10014 7540
rect 11422 7488 11428 7540
rect 11480 7528 11486 7540
rect 11517 7531 11575 7537
rect 11517 7528 11529 7531
rect 11480 7500 11529 7528
rect 11480 7488 11486 7500
rect 11517 7497 11529 7500
rect 11563 7497 11575 7531
rect 11517 7491 11575 7497
rect 12158 7488 12164 7540
rect 12216 7528 12222 7540
rect 13449 7531 13507 7537
rect 13449 7528 13461 7531
rect 12216 7500 13461 7528
rect 12216 7488 12222 7500
rect 13449 7497 13461 7500
rect 13495 7497 13507 7531
rect 13449 7491 13507 7497
rect 5534 7420 5540 7472
rect 5592 7460 5598 7472
rect 5592 7432 5948 7460
rect 5592 7420 5598 7432
rect 5920 7401 5948 7432
rect 6730 7420 6736 7472
rect 6788 7460 6794 7472
rect 8386 7460 8392 7472
rect 6788 7432 8064 7460
rect 8347 7432 8392 7460
rect 6788 7420 6794 7432
rect 4985 7395 5043 7401
rect 4985 7392 4997 7395
rect 4816 7364 4997 7392
rect 2041 7327 2099 7333
rect 1688 7296 1900 7324
rect 1762 7256 1768 7268
rect 1723 7228 1768 7256
rect 1762 7216 1768 7228
rect 1820 7216 1826 7268
rect 1872 7256 1900 7296
rect 2041 7293 2053 7327
rect 2087 7324 2099 7327
rect 3786 7324 3792 7336
rect 2087 7296 2544 7324
rect 3747 7296 3792 7324
rect 2087 7293 2099 7296
rect 2041 7287 2099 7293
rect 2314 7256 2320 7268
rect 1872 7228 2320 7256
rect 2314 7216 2320 7228
rect 2372 7216 2378 7268
rect 2516 7256 2544 7296
rect 3786 7284 3792 7296
rect 3844 7324 3850 7336
rect 4816 7324 4844 7364
rect 4985 7361 4997 7364
rect 5031 7361 5043 7395
rect 4985 7355 5043 7361
rect 5169 7395 5227 7401
rect 5169 7361 5181 7395
rect 5215 7361 5227 7395
rect 5169 7355 5227 7361
rect 5445 7395 5503 7401
rect 5445 7361 5457 7395
rect 5491 7361 5503 7395
rect 5445 7355 5503 7361
rect 5629 7395 5687 7401
rect 5629 7361 5641 7395
rect 5675 7361 5687 7395
rect 5629 7355 5687 7361
rect 5905 7395 5963 7401
rect 5905 7361 5917 7395
rect 5951 7361 5963 7395
rect 5905 7355 5963 7361
rect 6549 7395 6607 7401
rect 6549 7361 6561 7395
rect 6595 7361 6607 7395
rect 7006 7392 7012 7404
rect 6967 7364 7012 7392
rect 6549 7355 6607 7361
rect 3844 7296 4844 7324
rect 3844 7284 3850 7296
rect 4890 7284 4896 7336
rect 4948 7324 4954 7336
rect 5644 7324 5672 7355
rect 4948 7296 5672 7324
rect 4948 7284 4954 7296
rect 4154 7256 4160 7268
rect 2516 7228 4160 7256
rect 4154 7216 4160 7228
rect 4212 7216 4218 7268
rect 4246 7216 4252 7268
rect 4304 7256 4310 7268
rect 5077 7259 5135 7265
rect 5077 7256 5089 7259
rect 4304 7228 5089 7256
rect 4304 7216 4310 7228
rect 5077 7225 5089 7228
rect 5123 7225 5135 7259
rect 5077 7219 5135 7225
rect 2774 7148 2780 7200
rect 2832 7188 2838 7200
rect 2961 7191 3019 7197
rect 2832 7160 2877 7188
rect 2832 7148 2838 7160
rect 2961 7157 2973 7191
rect 3007 7188 3019 7191
rect 3510 7188 3516 7200
rect 3007 7160 3516 7188
rect 3007 7157 3019 7160
rect 2961 7151 3019 7157
rect 3510 7148 3516 7160
rect 3568 7148 3574 7200
rect 4525 7191 4583 7197
rect 4525 7157 4537 7191
rect 4571 7188 4583 7191
rect 4614 7188 4620 7200
rect 4571 7160 4620 7188
rect 4571 7157 4583 7160
rect 4525 7151 4583 7157
rect 4614 7148 4620 7160
rect 4672 7148 4678 7200
rect 5534 7188 5540 7200
rect 5495 7160 5540 7188
rect 5534 7148 5540 7160
rect 5592 7148 5598 7200
rect 5920 7188 5948 7355
rect 6089 7259 6147 7265
rect 6089 7225 6101 7259
rect 6135 7256 6147 7259
rect 6270 7256 6276 7268
rect 6135 7228 6276 7256
rect 6135 7225 6147 7228
rect 6089 7219 6147 7225
rect 6270 7216 6276 7228
rect 6328 7216 6334 7268
rect 6564 7256 6592 7355
rect 7006 7352 7012 7364
rect 7064 7352 7070 7404
rect 7190 7352 7196 7404
rect 7248 7392 7254 7404
rect 7929 7395 7987 7401
rect 7929 7392 7941 7395
rect 7248 7364 7941 7392
rect 7248 7352 7254 7364
rect 7929 7361 7941 7364
rect 7975 7361 7987 7395
rect 8036 7392 8064 7432
rect 8386 7420 8392 7432
rect 8444 7420 8450 7472
rect 10781 7463 10839 7469
rect 10781 7429 10793 7463
rect 10827 7429 10839 7463
rect 13170 7460 13176 7472
rect 13131 7432 13176 7460
rect 10781 7423 10839 7429
rect 8573 7395 8631 7401
rect 8573 7392 8585 7395
rect 8036 7364 8585 7392
rect 7929 7355 7987 7361
rect 8573 7361 8585 7364
rect 8619 7361 8631 7395
rect 8938 7392 8944 7404
rect 8899 7364 8944 7392
rect 8573 7355 8631 7361
rect 7098 7324 7104 7336
rect 7059 7296 7104 7324
rect 7098 7284 7104 7296
rect 7156 7284 7162 7336
rect 7742 7324 7748 7336
rect 7703 7296 7748 7324
rect 7742 7284 7748 7296
rect 7800 7284 7806 7336
rect 8588 7324 8616 7355
rect 8938 7352 8944 7364
rect 8996 7352 9002 7404
rect 9030 7352 9036 7404
rect 9088 7392 9094 7404
rect 9088 7364 9260 7392
rect 9088 7352 9094 7364
rect 9122 7324 9128 7336
rect 8588 7296 9128 7324
rect 9122 7284 9128 7296
rect 9180 7284 9186 7336
rect 9232 7324 9260 7364
rect 9674 7352 9680 7404
rect 9732 7392 9738 7404
rect 9732 7364 9777 7392
rect 9732 7352 9738 7364
rect 9858 7352 9864 7404
rect 9916 7392 9922 7404
rect 9973 7395 10031 7401
rect 9973 7392 9985 7395
rect 9916 7364 9985 7392
rect 9916 7352 9922 7364
rect 9973 7361 9985 7364
rect 10019 7361 10031 7395
rect 9973 7355 10031 7361
rect 10229 7395 10287 7401
rect 10229 7361 10241 7395
rect 10275 7361 10287 7395
rect 10229 7355 10287 7361
rect 10244 7324 10272 7355
rect 10502 7352 10508 7404
rect 10560 7392 10566 7404
rect 10796 7392 10824 7423
rect 13170 7420 13176 7432
rect 13228 7420 13234 7472
rect 11054 7392 11060 7404
rect 10560 7364 11060 7392
rect 10560 7352 10566 7364
rect 11054 7352 11060 7364
rect 11112 7392 11118 7404
rect 11606 7392 11612 7404
rect 11112 7364 11612 7392
rect 11112 7352 11118 7364
rect 11606 7352 11612 7364
rect 11664 7352 11670 7404
rect 11698 7352 11704 7404
rect 11756 7392 11762 7404
rect 11885 7395 11943 7401
rect 11885 7392 11897 7395
rect 11756 7364 11897 7392
rect 11756 7352 11762 7364
rect 11885 7361 11897 7364
rect 11931 7361 11943 7395
rect 12250 7392 12256 7404
rect 12211 7364 12256 7392
rect 11885 7355 11943 7361
rect 12250 7352 12256 7364
rect 12308 7352 12314 7404
rect 12713 7395 12771 7401
rect 12713 7361 12725 7395
rect 12759 7392 12771 7395
rect 12802 7392 12808 7404
rect 12759 7364 12808 7392
rect 12759 7361 12771 7364
rect 12713 7355 12771 7361
rect 12802 7352 12808 7364
rect 12860 7352 12866 7404
rect 13357 7395 13415 7401
rect 13357 7392 13369 7395
rect 12912 7364 13369 7392
rect 10410 7324 10416 7336
rect 9232 7296 10416 7324
rect 10410 7284 10416 7296
rect 10468 7324 10474 7336
rect 10689 7327 10747 7333
rect 10689 7324 10701 7327
rect 10468 7296 10701 7324
rect 10468 7284 10474 7296
rect 10689 7293 10701 7296
rect 10735 7293 10747 7327
rect 10689 7287 10747 7293
rect 10873 7327 10931 7333
rect 10873 7293 10885 7327
rect 10919 7324 10931 7327
rect 11146 7324 11152 7336
rect 10919 7296 11152 7324
rect 10919 7293 10931 7296
rect 10873 7287 10931 7293
rect 11146 7284 11152 7296
rect 11204 7324 11210 7336
rect 12912 7324 12940 7364
rect 13357 7361 13369 7364
rect 13403 7392 13415 7395
rect 13722 7392 13728 7404
rect 13403 7364 13728 7392
rect 13403 7361 13415 7364
rect 13357 7355 13415 7361
rect 13722 7352 13728 7364
rect 13780 7352 13786 7404
rect 13262 7324 13268 7336
rect 11204 7296 12940 7324
rect 13223 7296 13268 7324
rect 11204 7284 11210 7296
rect 13262 7284 13268 7296
rect 13320 7284 13326 7336
rect 8297 7259 8355 7265
rect 6564 7228 8248 7256
rect 6546 7188 6552 7200
rect 5920 7160 6552 7188
rect 6546 7148 6552 7160
rect 6604 7188 6610 7200
rect 6730 7188 6736 7200
rect 6604 7160 6736 7188
rect 6604 7148 6610 7160
rect 6730 7148 6736 7160
rect 6788 7148 6794 7200
rect 8220 7188 8248 7228
rect 8297 7225 8309 7259
rect 8343 7256 8355 7259
rect 11238 7256 11244 7268
rect 8343 7228 10824 7256
rect 11199 7228 11244 7256
rect 8343 7225 8355 7228
rect 8297 7219 8355 7225
rect 8846 7188 8852 7200
rect 8220 7160 8852 7188
rect 8846 7148 8852 7160
rect 8904 7148 8910 7200
rect 9490 7148 9496 7200
rect 9548 7188 9554 7200
rect 10229 7191 10287 7197
rect 10229 7188 10241 7191
rect 9548 7160 10241 7188
rect 9548 7148 9554 7160
rect 10229 7157 10241 7160
rect 10275 7157 10287 7191
rect 10796 7188 10824 7228
rect 11238 7216 11244 7228
rect 11296 7216 11302 7268
rect 13170 7256 13176 7268
rect 11900 7228 13176 7256
rect 11900 7188 11928 7228
rect 13170 7216 13176 7228
rect 13228 7216 13234 7268
rect 10796 7160 11928 7188
rect 10229 7151 10287 7157
rect 1104 7098 13892 7120
rect 1104 7046 4214 7098
rect 4266 7046 4278 7098
rect 4330 7046 4342 7098
rect 4394 7046 4406 7098
rect 4458 7046 4470 7098
rect 4522 7046 12214 7098
rect 12266 7046 12278 7098
rect 12330 7046 12342 7098
rect 12394 7046 12406 7098
rect 12458 7046 12470 7098
rect 12522 7046 13892 7098
rect 1104 7024 13892 7046
rect 1765 6987 1823 6993
rect 1765 6953 1777 6987
rect 1811 6984 1823 6987
rect 1946 6984 1952 6996
rect 1811 6956 1952 6984
rect 1811 6953 1823 6956
rect 1765 6947 1823 6953
rect 1946 6944 1952 6956
rect 2004 6944 2010 6996
rect 4617 6987 4675 6993
rect 4617 6984 4629 6987
rect 3344 6956 4629 6984
rect 2056 6888 2728 6916
rect 1578 6848 1584 6860
rect 1412 6820 1584 6848
rect 1412 6789 1440 6820
rect 1578 6808 1584 6820
rect 1636 6808 1642 6860
rect 2056 6857 2084 6888
rect 2041 6851 2099 6857
rect 2041 6817 2053 6851
rect 2087 6817 2099 6851
rect 2041 6811 2099 6817
rect 2133 6851 2191 6857
rect 2133 6817 2145 6851
rect 2179 6848 2191 6851
rect 2700 6848 2728 6888
rect 2958 6848 2964 6860
rect 2179 6820 2636 6848
rect 2700 6820 2820 6848
rect 2871 6820 2964 6848
rect 2179 6817 2191 6820
rect 2133 6811 2191 6817
rect 1397 6783 1455 6789
rect 1397 6749 1409 6783
rect 1443 6749 1455 6783
rect 1397 6743 1455 6749
rect 1486 6740 1492 6792
rect 1544 6780 1550 6792
rect 1949 6783 2007 6789
rect 1949 6780 1961 6783
rect 1544 6752 1961 6780
rect 1544 6740 1550 6752
rect 1949 6749 1961 6752
rect 1995 6749 2007 6783
rect 2222 6780 2228 6792
rect 2183 6752 2228 6780
rect 1949 6743 2007 6749
rect 2222 6740 2228 6752
rect 2280 6740 2286 6792
rect 2314 6740 2320 6792
rect 2372 6780 2378 6792
rect 2409 6783 2467 6789
rect 2409 6780 2421 6783
rect 2372 6752 2421 6780
rect 2372 6740 2378 6752
rect 2409 6749 2421 6752
rect 2455 6749 2467 6783
rect 2409 6743 2467 6749
rect 2608 6780 2636 6820
rect 2792 6792 2820 6820
rect 2958 6808 2964 6820
rect 3016 6848 3022 6860
rect 3344 6848 3372 6956
rect 4617 6953 4629 6956
rect 4663 6953 4675 6987
rect 4617 6947 4675 6953
rect 8110 6944 8116 6996
rect 8168 6984 8174 6996
rect 8481 6987 8539 6993
rect 8481 6984 8493 6987
rect 8168 6956 8493 6984
rect 8168 6944 8174 6956
rect 8481 6953 8493 6956
rect 8527 6953 8539 6987
rect 12250 6984 12256 6996
rect 8481 6947 8539 6953
rect 10428 6956 12256 6984
rect 10428 6928 10456 6956
rect 12250 6944 12256 6956
rect 12308 6944 12314 6996
rect 3786 6916 3792 6928
rect 3747 6888 3792 6916
rect 3786 6876 3792 6888
rect 3844 6876 3850 6928
rect 6362 6876 6368 6928
rect 6420 6916 6426 6928
rect 8297 6919 8355 6925
rect 8297 6916 8309 6919
rect 6420 6888 8309 6916
rect 6420 6876 6426 6888
rect 8297 6885 8309 6888
rect 8343 6885 8355 6919
rect 8297 6879 8355 6885
rect 10134 6876 10140 6928
rect 10192 6916 10198 6928
rect 10410 6925 10416 6928
rect 10321 6919 10379 6925
rect 10321 6916 10333 6919
rect 10192 6888 10333 6916
rect 10192 6876 10198 6888
rect 10321 6885 10333 6888
rect 10367 6885 10379 6919
rect 10321 6879 10379 6885
rect 10409 6879 10416 6925
rect 10468 6916 10474 6928
rect 10468 6888 10509 6916
rect 10410 6876 10416 6879
rect 10468 6876 10474 6888
rect 10870 6876 10876 6928
rect 10928 6916 10934 6928
rect 10965 6919 11023 6925
rect 10965 6916 10977 6919
rect 10928 6888 10977 6916
rect 10928 6876 10934 6888
rect 10965 6885 10977 6888
rect 11011 6885 11023 6919
rect 10965 6879 11023 6885
rect 12176 6888 12480 6916
rect 3510 6848 3516 6860
rect 3016 6820 3372 6848
rect 3471 6820 3516 6848
rect 3016 6808 3022 6820
rect 3510 6808 3516 6820
rect 3568 6848 3574 6860
rect 4801 6851 4859 6857
rect 3568 6820 4016 6848
rect 3568 6808 3574 6820
rect 2685 6783 2743 6789
rect 2685 6780 2697 6783
rect 2608 6752 2697 6780
rect 1581 6715 1639 6721
rect 1581 6681 1593 6715
rect 1627 6681 1639 6715
rect 1581 6675 1639 6681
rect 1596 6644 1624 6675
rect 2038 6672 2044 6724
rect 2096 6712 2102 6724
rect 2501 6715 2559 6721
rect 2501 6712 2513 6715
rect 2096 6684 2513 6712
rect 2096 6672 2102 6684
rect 2501 6681 2513 6684
rect 2547 6681 2559 6715
rect 2608 6712 2636 6752
rect 2685 6749 2697 6752
rect 2731 6749 2743 6783
rect 2685 6743 2743 6749
rect 2774 6740 2780 6792
rect 2832 6780 2838 6792
rect 2832 6752 2877 6780
rect 2832 6740 2838 6752
rect 3142 6740 3148 6792
rect 3200 6780 3206 6792
rect 3988 6789 4016 6820
rect 4801 6817 4813 6851
rect 4847 6848 4859 6851
rect 5534 6848 5540 6860
rect 4847 6820 5540 6848
rect 4847 6817 4859 6820
rect 4801 6811 4859 6817
rect 5534 6808 5540 6820
rect 5592 6808 5598 6860
rect 6733 6851 6791 6857
rect 6733 6817 6745 6851
rect 6779 6848 6791 6851
rect 7006 6848 7012 6860
rect 6779 6820 7012 6848
rect 6779 6817 6791 6820
rect 6733 6811 6791 6817
rect 7006 6808 7012 6820
rect 7064 6808 7070 6860
rect 7392 6820 8616 6848
rect 3329 6783 3387 6789
rect 3329 6780 3341 6783
rect 3200 6752 3341 6780
rect 3200 6740 3206 6752
rect 3329 6749 3341 6752
rect 3375 6749 3387 6783
rect 3329 6743 3387 6749
rect 3973 6783 4031 6789
rect 3973 6749 3985 6783
rect 4019 6749 4031 6783
rect 3973 6743 4031 6749
rect 4525 6783 4583 6789
rect 4525 6749 4537 6783
rect 4571 6780 4583 6783
rect 4706 6780 4712 6792
rect 4571 6752 4712 6780
rect 4571 6749 4583 6752
rect 4525 6743 4583 6749
rect 3053 6715 3111 6721
rect 3053 6712 3065 6715
rect 2608 6684 3065 6712
rect 2501 6675 2559 6681
rect 3053 6681 3065 6684
rect 3099 6681 3111 6715
rect 3053 6675 3111 6681
rect 3234 6644 3240 6656
rect 1596 6616 3240 6644
rect 3234 6604 3240 6616
rect 3292 6604 3298 6656
rect 3344 6644 3372 6743
rect 4706 6740 4712 6752
rect 4764 6740 4770 6792
rect 4890 6740 4896 6792
rect 4948 6780 4954 6792
rect 5077 6783 5135 6789
rect 5077 6780 5089 6783
rect 4948 6752 5089 6780
rect 4948 6740 4954 6752
rect 5077 6749 5089 6752
rect 5123 6749 5135 6783
rect 5077 6743 5135 6749
rect 5261 6783 5319 6789
rect 5261 6749 5273 6783
rect 5307 6780 5319 6783
rect 5626 6780 5632 6792
rect 5307 6752 5632 6780
rect 5307 6749 5319 6752
rect 5261 6743 5319 6749
rect 5626 6740 5632 6752
rect 5684 6740 5690 6792
rect 6089 6783 6147 6789
rect 6089 6749 6101 6783
rect 6135 6749 6147 6783
rect 6089 6743 6147 6749
rect 6365 6783 6423 6789
rect 6365 6749 6377 6783
rect 6411 6780 6423 6783
rect 6822 6780 6828 6792
rect 6411 6752 6828 6780
rect 6411 6749 6423 6752
rect 6365 6743 6423 6749
rect 4341 6715 4399 6721
rect 4341 6681 4353 6715
rect 4387 6712 4399 6715
rect 4614 6712 4620 6724
rect 4387 6684 4620 6712
rect 4387 6681 4399 6684
rect 4341 6675 4399 6681
rect 4614 6672 4620 6684
rect 4672 6672 4678 6724
rect 6104 6712 6132 6743
rect 6822 6740 6828 6752
rect 6880 6780 6886 6792
rect 7193 6783 7251 6789
rect 7193 6780 7205 6783
rect 6880 6752 7205 6780
rect 6880 6740 6886 6752
rect 7193 6749 7205 6752
rect 7239 6749 7251 6783
rect 7193 6743 7251 6749
rect 7392 6712 7420 6820
rect 7469 6783 7527 6789
rect 7469 6749 7481 6783
rect 7515 6749 7527 6783
rect 7469 6743 7527 6749
rect 6104 6684 7420 6712
rect 7484 6712 7512 6743
rect 7558 6740 7564 6792
rect 7616 6780 7622 6792
rect 8205 6783 8263 6789
rect 8205 6780 8217 6783
rect 7616 6752 8217 6780
rect 7616 6740 7622 6752
rect 8205 6749 8217 6752
rect 8251 6749 8263 6783
rect 8205 6743 8263 6749
rect 7650 6712 7656 6724
rect 7484 6684 7656 6712
rect 7650 6672 7656 6684
rect 7708 6712 7714 6724
rect 7834 6712 7840 6724
rect 7708 6684 7840 6712
rect 7708 6672 7714 6684
rect 7834 6672 7840 6684
rect 7892 6672 7898 6724
rect 8588 6712 8616 6820
rect 8662 6808 8668 6860
rect 8720 6848 8726 6860
rect 10888 6848 10916 6876
rect 11698 6848 11704 6860
rect 8720 6820 8765 6848
rect 10244 6820 10916 6848
rect 11072 6820 11704 6848
rect 8720 6808 8726 6820
rect 9398 6780 9404 6792
rect 9359 6752 9404 6780
rect 9398 6740 9404 6752
rect 9456 6740 9462 6792
rect 9674 6780 9680 6792
rect 9635 6752 9680 6780
rect 9674 6740 9680 6752
rect 9732 6740 9738 6792
rect 10244 6789 10272 6820
rect 10229 6783 10287 6789
rect 10229 6749 10241 6783
rect 10275 6780 10287 6783
rect 10318 6780 10324 6792
rect 10275 6752 10324 6780
rect 10275 6749 10287 6752
rect 10229 6743 10287 6749
rect 10318 6740 10324 6752
rect 10376 6740 10382 6792
rect 10505 6783 10563 6789
rect 10505 6749 10517 6783
rect 10551 6780 10563 6783
rect 10594 6780 10600 6792
rect 10551 6752 10600 6780
rect 10551 6749 10563 6752
rect 10505 6743 10563 6749
rect 10520 6712 10548 6743
rect 10594 6740 10600 6752
rect 10652 6740 10658 6792
rect 10778 6780 10784 6792
rect 10739 6752 10784 6780
rect 10778 6740 10784 6752
rect 10836 6740 10842 6792
rect 10873 6783 10931 6789
rect 10873 6749 10885 6783
rect 10919 6780 10931 6783
rect 11072 6780 11100 6820
rect 11698 6808 11704 6820
rect 11756 6808 11762 6860
rect 11790 6808 11796 6860
rect 11848 6848 11854 6860
rect 12176 6848 12204 6888
rect 11848 6820 12204 6848
rect 11848 6808 11854 6820
rect 12250 6808 12256 6860
rect 12308 6848 12314 6860
rect 12345 6851 12403 6857
rect 12345 6848 12357 6851
rect 12308 6820 12357 6848
rect 12308 6808 12314 6820
rect 12345 6817 12357 6820
rect 12391 6817 12403 6851
rect 12452 6848 12480 6888
rect 12452 6820 12940 6848
rect 12345 6811 12403 6817
rect 10919 6752 11100 6780
rect 11149 6783 11207 6789
rect 10919 6749 10931 6752
rect 10873 6743 10931 6749
rect 11149 6749 11161 6783
rect 11195 6780 11207 6783
rect 11238 6780 11244 6792
rect 11195 6752 11244 6780
rect 11195 6749 11207 6752
rect 11149 6743 11207 6749
rect 11238 6740 11244 6752
rect 11296 6740 11302 6792
rect 11974 6740 11980 6792
rect 12032 6740 12038 6792
rect 12805 6783 12863 6789
rect 12805 6749 12817 6783
rect 12851 6749 12863 6783
rect 12912 6780 12940 6820
rect 13170 6808 13176 6860
rect 13228 6848 13234 6860
rect 13357 6851 13415 6857
rect 13357 6848 13369 6851
rect 13228 6820 13369 6848
rect 13228 6808 13234 6820
rect 13357 6817 13369 6820
rect 13403 6817 13415 6851
rect 13357 6811 13415 6817
rect 13449 6783 13507 6789
rect 13449 6780 13461 6783
rect 12912 6752 13461 6780
rect 12805 6743 12863 6749
rect 13449 6749 13461 6752
rect 13495 6749 13507 6783
rect 13449 6743 13507 6749
rect 11514 6712 11520 6724
rect 8588 6684 10548 6712
rect 11475 6684 11520 6712
rect 11514 6672 11520 6684
rect 11572 6672 11578 6724
rect 12820 6712 12848 6743
rect 12406 6684 12848 6712
rect 4062 6644 4068 6656
rect 3344 6616 4068 6644
rect 4062 6604 4068 6616
rect 4120 6604 4126 6656
rect 4154 6604 4160 6656
rect 4212 6644 4218 6656
rect 5445 6647 5503 6653
rect 4212 6616 4257 6644
rect 4212 6604 4218 6616
rect 5445 6613 5457 6647
rect 5491 6644 5503 6647
rect 5534 6644 5540 6656
rect 5491 6616 5540 6644
rect 5491 6613 5503 6616
rect 5445 6607 5503 6613
rect 5534 6604 5540 6616
rect 5592 6604 5598 6656
rect 6825 6647 6883 6653
rect 6825 6613 6837 6647
rect 6871 6644 6883 6647
rect 6914 6644 6920 6656
rect 6871 6616 6920 6644
rect 6871 6613 6883 6616
rect 6825 6607 6883 6613
rect 6914 6604 6920 6616
rect 6972 6604 6978 6656
rect 8018 6644 8024 6656
rect 7979 6616 8024 6644
rect 8018 6604 8024 6616
rect 8076 6604 8082 6656
rect 9950 6604 9956 6656
rect 10008 6644 10014 6656
rect 10045 6647 10103 6653
rect 10045 6644 10057 6647
rect 10008 6616 10057 6644
rect 10008 6604 10014 6616
rect 10045 6613 10057 6616
rect 10091 6613 10103 6647
rect 10045 6607 10103 6613
rect 10410 6604 10416 6656
rect 10468 6644 10474 6656
rect 11146 6644 11152 6656
rect 10468 6616 11152 6644
rect 10468 6604 10474 6616
rect 11146 6604 11152 6616
rect 11204 6604 11210 6656
rect 11333 6647 11391 6653
rect 11333 6613 11345 6647
rect 11379 6644 11391 6647
rect 11790 6644 11796 6656
rect 11379 6616 11796 6644
rect 11379 6613 11391 6616
rect 11333 6607 11391 6613
rect 11790 6604 11796 6616
rect 11848 6604 11854 6656
rect 11974 6604 11980 6656
rect 12032 6644 12038 6656
rect 12406 6644 12434 6684
rect 13170 6672 13176 6724
rect 13228 6712 13234 6724
rect 13265 6715 13323 6721
rect 13265 6712 13277 6715
rect 13228 6684 13277 6712
rect 13228 6672 13234 6684
rect 13265 6681 13277 6684
rect 13311 6681 13323 6715
rect 13265 6675 13323 6681
rect 12032 6616 12434 6644
rect 12032 6604 12038 6616
rect 1104 6554 13892 6576
rect 1104 6502 8214 6554
rect 8266 6502 8278 6554
rect 8330 6502 8342 6554
rect 8394 6502 8406 6554
rect 8458 6502 8470 6554
rect 8522 6502 13892 6554
rect 1104 6480 13892 6502
rect 1397 6443 1455 6449
rect 1397 6409 1409 6443
rect 1443 6440 1455 6443
rect 2222 6440 2228 6452
rect 1443 6412 2228 6440
rect 1443 6409 1455 6412
rect 1397 6403 1455 6409
rect 2222 6400 2228 6412
rect 2280 6400 2286 6452
rect 3145 6443 3203 6449
rect 3145 6409 3157 6443
rect 3191 6440 3203 6443
rect 3510 6440 3516 6452
rect 3191 6412 3516 6440
rect 3191 6409 3203 6412
rect 3145 6403 3203 6409
rect 3510 6400 3516 6412
rect 3568 6400 3574 6452
rect 4154 6400 4160 6452
rect 4212 6440 4218 6452
rect 6089 6443 6147 6449
rect 6089 6440 6101 6443
rect 4212 6412 6101 6440
rect 4212 6400 4218 6412
rect 6089 6409 6101 6412
rect 6135 6409 6147 6443
rect 6089 6403 6147 6409
rect 7377 6443 7435 6449
rect 7377 6409 7389 6443
rect 7423 6440 7435 6443
rect 7742 6440 7748 6452
rect 7423 6412 7748 6440
rect 7423 6409 7435 6412
rect 7377 6403 7435 6409
rect 7742 6400 7748 6412
rect 7800 6400 7806 6452
rect 8754 6440 8760 6452
rect 8715 6412 8760 6440
rect 8754 6400 8760 6412
rect 8812 6400 8818 6452
rect 9125 6443 9183 6449
rect 9125 6409 9137 6443
rect 9171 6440 9183 6443
rect 9214 6440 9220 6452
rect 9171 6412 9220 6440
rect 9171 6409 9183 6412
rect 9125 6403 9183 6409
rect 9214 6400 9220 6412
rect 9272 6400 9278 6452
rect 9306 6400 9312 6452
rect 9364 6440 9370 6452
rect 9493 6443 9551 6449
rect 9493 6440 9505 6443
rect 9364 6412 9505 6440
rect 9364 6400 9370 6412
rect 9493 6409 9505 6412
rect 9539 6409 9551 6443
rect 9950 6440 9956 6452
rect 9911 6412 9956 6440
rect 9493 6403 9551 6409
rect 9950 6400 9956 6412
rect 10008 6400 10014 6452
rect 11149 6443 11207 6449
rect 11149 6409 11161 6443
rect 11195 6440 11207 6443
rect 11514 6440 11520 6452
rect 11195 6412 11520 6440
rect 11195 6409 11207 6412
rect 11149 6403 11207 6409
rect 11514 6400 11520 6412
rect 11572 6400 11578 6452
rect 4062 6372 4068 6384
rect 2792 6344 3648 6372
rect 4023 6344 4068 6372
rect 2792 6316 2820 6344
rect 2038 6304 2044 6316
rect 1999 6276 2044 6304
rect 2038 6264 2044 6276
rect 2096 6264 2102 6316
rect 2130 6264 2136 6316
rect 2188 6304 2194 6316
rect 2593 6307 2651 6313
rect 2593 6304 2605 6307
rect 2188 6276 2605 6304
rect 2188 6264 2194 6276
rect 2593 6273 2605 6276
rect 2639 6273 2651 6307
rect 2593 6267 2651 6273
rect 2774 6264 2780 6316
rect 2832 6304 2838 6316
rect 3326 6304 3332 6316
rect 2832 6276 2925 6304
rect 3287 6276 3332 6304
rect 2832 6264 2838 6276
rect 3326 6264 3332 6276
rect 3384 6264 3390 6316
rect 3620 6313 3648 6344
rect 4062 6332 4068 6344
rect 4120 6332 4126 6384
rect 4985 6375 5043 6381
rect 4985 6341 4997 6375
rect 5031 6372 5043 6375
rect 5074 6372 5080 6384
rect 5031 6344 5080 6372
rect 5031 6341 5043 6344
rect 4985 6335 5043 6341
rect 5074 6332 5080 6344
rect 5132 6332 5138 6384
rect 6178 6372 6184 6384
rect 5828 6344 6184 6372
rect 3421 6307 3479 6313
rect 3421 6273 3433 6307
rect 3467 6273 3479 6307
rect 3421 6267 3479 6273
rect 3605 6307 3663 6313
rect 3605 6273 3617 6307
rect 3651 6273 3663 6307
rect 3605 6267 3663 6273
rect 2317 6239 2375 6245
rect 2317 6205 2329 6239
rect 2363 6236 2375 6239
rect 2869 6239 2927 6245
rect 2869 6236 2881 6239
rect 2363 6208 2881 6236
rect 2363 6205 2375 6208
rect 2317 6199 2375 6205
rect 2869 6205 2881 6208
rect 2915 6205 2927 6239
rect 2869 6199 2927 6205
rect 3142 6196 3148 6248
rect 3200 6236 3206 6248
rect 3436 6236 3464 6267
rect 3694 6264 3700 6316
rect 3752 6304 3758 6316
rect 3752 6276 3797 6304
rect 3752 6264 3758 6276
rect 3878 6264 3884 6316
rect 3936 6304 3942 6316
rect 4246 6304 4252 6316
rect 3936 6276 3981 6304
rect 4207 6276 4252 6304
rect 3936 6264 3942 6276
rect 4246 6264 4252 6276
rect 4304 6264 4310 6316
rect 4801 6307 4859 6313
rect 4801 6273 4813 6307
rect 4847 6304 4859 6307
rect 5166 6304 5172 6316
rect 4847 6276 5172 6304
rect 4847 6273 4859 6276
rect 4801 6267 4859 6273
rect 5166 6264 5172 6276
rect 5224 6264 5230 6316
rect 5534 6304 5540 6316
rect 5495 6276 5540 6304
rect 5534 6264 5540 6276
rect 5592 6264 5598 6316
rect 5828 6313 5856 6344
rect 6178 6332 6184 6344
rect 6236 6332 6242 6384
rect 7006 6332 7012 6384
rect 7064 6372 7070 6384
rect 8021 6375 8079 6381
rect 8021 6372 8033 6375
rect 7064 6344 8033 6372
rect 7064 6332 7070 6344
rect 8021 6341 8033 6344
rect 8067 6341 8079 6375
rect 8570 6372 8576 6384
rect 8531 6344 8576 6372
rect 8021 6335 8079 6341
rect 8570 6332 8576 6344
rect 8628 6332 8634 6384
rect 11054 6372 11060 6384
rect 9600 6344 11060 6372
rect 5813 6307 5871 6313
rect 5813 6273 5825 6307
rect 5859 6273 5871 6307
rect 5813 6267 5871 6273
rect 5997 6307 6055 6313
rect 5997 6273 6009 6307
rect 6043 6273 6055 6307
rect 5997 6267 6055 6273
rect 6733 6307 6791 6313
rect 6733 6273 6745 6307
rect 6779 6304 6791 6307
rect 6914 6304 6920 6316
rect 6779 6276 6920 6304
rect 6779 6273 6791 6276
rect 6733 6267 6791 6273
rect 3200 6208 3464 6236
rect 3200 6196 3206 6208
rect 3510 6196 3516 6248
rect 3568 6236 3574 6248
rect 4154 6236 4160 6248
rect 3568 6208 4160 6236
rect 3568 6196 3574 6208
rect 4154 6196 4160 6208
rect 4212 6196 4218 6248
rect 4982 6196 4988 6248
rect 5040 6236 5046 6248
rect 5077 6239 5135 6245
rect 5077 6236 5089 6239
rect 5040 6208 5089 6236
rect 5040 6196 5046 6208
rect 5077 6205 5089 6208
rect 5123 6205 5135 6239
rect 5184 6236 5212 6264
rect 5828 6236 5856 6267
rect 5184 6208 5856 6236
rect 5077 6199 5135 6205
rect 4706 6128 4712 6180
rect 4764 6168 4770 6180
rect 6012 6168 6040 6267
rect 6914 6264 6920 6276
rect 6972 6264 6978 6316
rect 7101 6307 7159 6313
rect 7101 6273 7113 6307
rect 7147 6304 7159 6307
rect 7285 6307 7343 6313
rect 7285 6304 7297 6307
rect 7147 6276 7297 6304
rect 7147 6273 7159 6276
rect 7101 6267 7159 6273
rect 7285 6273 7297 6276
rect 7331 6304 7343 6307
rect 7742 6304 7748 6316
rect 7331 6276 7748 6304
rect 7331 6273 7343 6276
rect 7285 6267 7343 6273
rect 7742 6264 7748 6276
rect 7800 6304 7806 6316
rect 9600 6313 9628 6344
rect 11054 6332 11060 6344
rect 11112 6332 11118 6384
rect 11238 6332 11244 6384
rect 11296 6372 11302 6384
rect 11885 6375 11943 6381
rect 11885 6372 11897 6375
rect 11296 6344 11897 6372
rect 11296 6332 11302 6344
rect 11885 6341 11897 6344
rect 11931 6341 11943 6375
rect 11885 6335 11943 6341
rect 9585 6307 9643 6313
rect 7800 6276 8892 6304
rect 7800 6264 7806 6276
rect 6638 6236 6644 6248
rect 6599 6208 6644 6236
rect 6638 6196 6644 6208
rect 6696 6196 6702 6248
rect 7374 6236 7380 6248
rect 7335 6208 7380 6236
rect 7374 6196 7380 6208
rect 7432 6196 7438 6248
rect 8864 6245 8892 6276
rect 9585 6273 9597 6307
rect 9631 6273 9643 6307
rect 9951 6307 10009 6313
rect 9951 6304 9963 6307
rect 9585 6267 9643 6273
rect 9692 6276 9963 6304
rect 8849 6239 8907 6245
rect 8849 6205 8861 6239
rect 8895 6236 8907 6239
rect 9692 6236 9720 6276
rect 9951 6273 9963 6276
rect 9997 6304 10009 6307
rect 10502 6304 10508 6316
rect 9997 6276 10508 6304
rect 9997 6273 10009 6276
rect 9951 6267 10009 6273
rect 10502 6264 10508 6276
rect 10560 6304 10566 6316
rect 11517 6307 11575 6313
rect 11517 6304 11529 6307
rect 10560 6276 11529 6304
rect 10560 6264 10566 6276
rect 10410 6236 10416 6248
rect 8895 6208 9720 6236
rect 10371 6208 10416 6236
rect 8895 6205 8907 6208
rect 8849 6199 8907 6205
rect 10410 6196 10416 6208
rect 10468 6196 10474 6248
rect 11146 6236 11152 6248
rect 11107 6208 11152 6236
rect 11146 6196 11152 6208
rect 11204 6196 11210 6248
rect 11256 6245 11284 6276
rect 11517 6273 11529 6276
rect 11563 6273 11575 6307
rect 11698 6304 11704 6316
rect 11659 6276 11704 6304
rect 11517 6267 11575 6273
rect 11698 6264 11704 6276
rect 11756 6264 11762 6316
rect 11974 6304 11980 6316
rect 11887 6276 11980 6304
rect 11974 6264 11980 6276
rect 12032 6264 12038 6316
rect 13446 6304 13452 6316
rect 13407 6276 13452 6304
rect 13446 6264 13452 6276
rect 13504 6264 13510 6316
rect 11241 6239 11299 6245
rect 11241 6205 11253 6239
rect 11287 6205 11299 6239
rect 11241 6199 11299 6205
rect 11422 6196 11428 6248
rect 11480 6236 11486 6248
rect 11992 6236 12020 6264
rect 11480 6208 12020 6236
rect 11480 6196 11486 6208
rect 4764 6140 6040 6168
rect 7009 6171 7067 6177
rect 4764 6128 4770 6140
rect 7009 6137 7021 6171
rect 7055 6168 7067 6171
rect 7926 6168 7932 6180
rect 7055 6140 7932 6168
rect 7055 6137 7067 6140
rect 7009 6131 7067 6137
rect 7926 6128 7932 6140
rect 7984 6128 7990 6180
rect 9674 6128 9680 6180
rect 9732 6168 9738 6180
rect 10318 6168 10324 6180
rect 9732 6140 9904 6168
rect 10279 6140 10324 6168
rect 9732 6128 9738 6140
rect 2682 6060 2688 6112
rect 2740 6100 2746 6112
rect 4062 6100 4068 6112
rect 2740 6072 4068 6100
rect 2740 6060 2746 6072
rect 4062 6060 4068 6072
rect 4120 6060 4126 6112
rect 4154 6060 4160 6112
rect 4212 6100 4218 6112
rect 4525 6103 4583 6109
rect 4525 6100 4537 6103
rect 4212 6072 4537 6100
rect 4212 6060 4218 6072
rect 4525 6069 4537 6072
rect 4571 6069 4583 6103
rect 4525 6063 4583 6069
rect 5721 6103 5779 6109
rect 5721 6069 5733 6103
rect 5767 6100 5779 6103
rect 5810 6100 5816 6112
rect 5767 6072 5816 6100
rect 5767 6069 5779 6072
rect 5721 6063 5779 6069
rect 5810 6060 5816 6072
rect 5868 6060 5874 6112
rect 6362 6100 6368 6112
rect 6323 6072 6368 6100
rect 6362 6060 6368 6072
rect 6420 6060 6426 6112
rect 7834 6100 7840 6112
rect 7795 6072 7840 6100
rect 7834 6060 7840 6072
rect 7892 6060 7898 6112
rect 8297 6103 8355 6109
rect 8297 6069 8309 6103
rect 8343 6100 8355 6103
rect 8386 6100 8392 6112
rect 8343 6072 8392 6100
rect 8343 6069 8355 6072
rect 8297 6063 8355 6069
rect 8386 6060 8392 6072
rect 8444 6060 8450 6112
rect 9766 6100 9772 6112
rect 9727 6072 9772 6100
rect 9766 6060 9772 6072
rect 9824 6060 9830 6112
rect 9876 6100 9904 6140
rect 10318 6128 10324 6140
rect 10376 6128 10382 6180
rect 13170 6128 13176 6180
rect 13228 6168 13234 6180
rect 13265 6171 13323 6177
rect 13265 6168 13277 6171
rect 13228 6140 13277 6168
rect 13228 6128 13234 6140
rect 13265 6137 13277 6140
rect 13311 6137 13323 6171
rect 13265 6131 13323 6137
rect 10689 6103 10747 6109
rect 10689 6100 10701 6103
rect 9876 6072 10701 6100
rect 10689 6069 10701 6072
rect 10735 6069 10747 6103
rect 10689 6063 10747 6069
rect 1104 6010 13892 6032
rect 1104 5958 4214 6010
rect 4266 5958 4278 6010
rect 4330 5958 4342 6010
rect 4394 5958 4406 6010
rect 4458 5958 4470 6010
rect 4522 5958 12214 6010
rect 12266 5958 12278 6010
rect 12330 5958 12342 6010
rect 12394 5958 12406 6010
rect 12458 5958 12470 6010
rect 12522 5958 13892 6010
rect 1104 5936 13892 5958
rect 1486 5896 1492 5908
rect 1447 5868 1492 5896
rect 1486 5856 1492 5868
rect 1544 5856 1550 5908
rect 2038 5856 2044 5908
rect 2096 5896 2102 5908
rect 2096 5868 2268 5896
rect 2096 5856 2102 5868
rect 1765 5831 1823 5837
rect 1765 5797 1777 5831
rect 1811 5797 1823 5831
rect 2130 5828 2136 5840
rect 2091 5800 2136 5828
rect 1765 5791 1823 5797
rect 1780 5760 1808 5791
rect 2130 5788 2136 5800
rect 2188 5788 2194 5840
rect 2240 5828 2268 5868
rect 2774 5856 2780 5908
rect 2832 5896 2838 5908
rect 2869 5899 2927 5905
rect 2869 5896 2881 5899
rect 2832 5868 2881 5896
rect 2832 5856 2838 5868
rect 2869 5865 2881 5868
rect 2915 5865 2927 5899
rect 2869 5859 2927 5865
rect 3602 5856 3608 5908
rect 3660 5896 3666 5908
rect 3789 5899 3847 5905
rect 3789 5896 3801 5899
rect 3660 5868 3801 5896
rect 3660 5856 3666 5868
rect 3789 5865 3801 5868
rect 3835 5865 3847 5899
rect 3789 5859 3847 5865
rect 5442 5856 5448 5908
rect 5500 5896 5506 5908
rect 7469 5899 7527 5905
rect 7469 5896 7481 5899
rect 5500 5868 7481 5896
rect 5500 5856 5506 5868
rect 7469 5865 7481 5868
rect 7515 5865 7527 5899
rect 7742 5896 7748 5908
rect 7703 5868 7748 5896
rect 7469 5859 7527 5865
rect 7742 5856 7748 5868
rect 7800 5856 7806 5908
rect 7834 5856 7840 5908
rect 7892 5896 7898 5908
rect 7892 5868 8708 5896
rect 7892 5856 7898 5868
rect 3513 5831 3571 5837
rect 3513 5828 3525 5831
rect 2240 5800 3525 5828
rect 3513 5797 3525 5800
rect 3559 5797 3571 5831
rect 3513 5791 3571 5797
rect 4525 5831 4583 5837
rect 4525 5797 4537 5831
rect 4571 5828 4583 5831
rect 4706 5828 4712 5840
rect 4571 5800 4712 5828
rect 4571 5797 4583 5800
rect 4525 5791 4583 5797
rect 4706 5788 4712 5800
rect 4764 5788 4770 5840
rect 4890 5788 4896 5840
rect 4948 5828 4954 5840
rect 5460 5828 5488 5856
rect 4948 5800 5488 5828
rect 4948 5788 4954 5800
rect 5718 5788 5724 5840
rect 5776 5788 5782 5840
rect 8110 5788 8116 5840
rect 8168 5828 8174 5840
rect 8573 5831 8631 5837
rect 8573 5828 8585 5831
rect 8168 5800 8585 5828
rect 8168 5788 8174 5800
rect 8573 5797 8585 5800
rect 8619 5797 8631 5831
rect 8573 5791 8631 5797
rect 4798 5760 4804 5772
rect 1780 5732 2176 5760
rect 1394 5692 1400 5704
rect 1355 5664 1400 5692
rect 1394 5652 1400 5664
rect 1452 5652 1458 5704
rect 1949 5695 2007 5701
rect 1949 5661 1961 5695
rect 1995 5661 2007 5695
rect 1949 5655 2007 5661
rect 1964 5556 1992 5655
rect 2148 5624 2176 5732
rect 2240 5732 2728 5760
rect 2240 5701 2268 5732
rect 2225 5695 2283 5701
rect 2225 5661 2237 5695
rect 2271 5661 2283 5695
rect 2225 5655 2283 5661
rect 2409 5695 2467 5701
rect 2409 5661 2421 5695
rect 2455 5692 2467 5695
rect 2590 5692 2596 5704
rect 2455 5664 2596 5692
rect 2455 5661 2467 5664
rect 2409 5655 2467 5661
rect 2590 5652 2596 5664
rect 2648 5652 2654 5704
rect 2700 5701 2728 5732
rect 4632 5732 4804 5760
rect 2685 5695 2743 5701
rect 2685 5661 2697 5695
rect 2731 5692 2743 5695
rect 2774 5692 2780 5704
rect 2731 5664 2780 5692
rect 2731 5661 2743 5664
rect 2685 5655 2743 5661
rect 2774 5652 2780 5664
rect 2832 5652 2838 5704
rect 3053 5695 3111 5701
rect 3053 5661 3065 5695
rect 3099 5661 3111 5695
rect 3053 5655 3111 5661
rect 2498 5624 2504 5636
rect 2148 5596 2504 5624
rect 2498 5584 2504 5596
rect 2556 5584 2562 5636
rect 3068 5624 3096 5655
rect 3142 5652 3148 5704
rect 3200 5692 3206 5704
rect 3237 5695 3295 5701
rect 3237 5692 3249 5695
rect 3200 5664 3249 5692
rect 3200 5652 3206 5664
rect 3237 5661 3249 5664
rect 3283 5661 3295 5695
rect 3237 5655 3295 5661
rect 3605 5695 3663 5701
rect 3605 5661 3617 5695
rect 3651 5692 3663 5695
rect 3694 5692 3700 5704
rect 3651 5664 3700 5692
rect 3651 5661 3663 5664
rect 3605 5655 3663 5661
rect 3694 5652 3700 5664
rect 3752 5652 3758 5704
rect 4062 5692 4068 5704
rect 4023 5664 4068 5692
rect 4062 5652 4068 5664
rect 4120 5652 4126 5704
rect 4632 5701 4660 5732
rect 4798 5720 4804 5732
rect 4856 5720 4862 5772
rect 4249 5695 4307 5701
rect 4249 5661 4261 5695
rect 4295 5692 4307 5695
rect 4617 5695 4675 5701
rect 4295 5664 4568 5692
rect 4295 5661 4307 5664
rect 4249 5655 4307 5661
rect 3326 5624 3332 5636
rect 3068 5596 3332 5624
rect 3326 5584 3332 5596
rect 3384 5624 3390 5636
rect 3510 5624 3516 5636
rect 3384 5596 3516 5624
rect 3384 5584 3390 5596
rect 3510 5584 3516 5596
rect 3568 5584 3574 5636
rect 3602 5556 3608 5568
rect 1964 5528 3608 5556
rect 3602 5516 3608 5528
rect 3660 5516 3666 5568
rect 4246 5556 4252 5568
rect 4207 5528 4252 5556
rect 4246 5516 4252 5528
rect 4304 5516 4310 5568
rect 4540 5556 4568 5664
rect 4617 5661 4629 5695
rect 4663 5661 4675 5695
rect 4617 5655 4675 5661
rect 4709 5695 4767 5701
rect 4709 5661 4721 5695
rect 4755 5692 4767 5695
rect 4908 5692 4936 5788
rect 5736 5760 5764 5788
rect 7650 5760 7656 5772
rect 5276 5732 5764 5760
rect 7611 5732 7656 5760
rect 5276 5701 5304 5732
rect 7650 5720 7656 5732
rect 7708 5720 7714 5772
rect 7834 5720 7840 5772
rect 7892 5760 7898 5772
rect 7892 5732 8064 5760
rect 7892 5720 7898 5732
rect 4755 5664 4936 5692
rect 5169 5695 5227 5701
rect 4755 5661 4767 5664
rect 4709 5655 4767 5661
rect 4982 5630 4988 5682
rect 5040 5670 5046 5682
rect 5040 5642 5085 5670
rect 5169 5661 5181 5695
rect 5215 5661 5227 5695
rect 5169 5655 5227 5661
rect 5261 5695 5319 5701
rect 5261 5661 5273 5695
rect 5307 5661 5319 5695
rect 5261 5655 5319 5661
rect 5354 5695 5412 5701
rect 5354 5661 5366 5695
rect 5400 5692 5412 5695
rect 5442 5692 5448 5704
rect 5400 5664 5448 5692
rect 5400 5661 5412 5664
rect 5354 5655 5412 5661
rect 5040 5630 5046 5642
rect 5184 5624 5212 5655
rect 5442 5652 5448 5664
rect 5500 5652 5506 5704
rect 5534 5652 5540 5704
rect 5592 5692 5598 5704
rect 5721 5695 5779 5701
rect 5721 5692 5733 5695
rect 5592 5664 5733 5692
rect 5592 5652 5598 5664
rect 5721 5661 5733 5664
rect 5767 5661 5779 5695
rect 7926 5692 7932 5704
rect 7887 5664 7932 5692
rect 5721 5655 5779 5661
rect 7926 5652 7932 5664
rect 7984 5652 7990 5704
rect 8036 5701 8064 5732
rect 8021 5695 8079 5701
rect 8021 5661 8033 5695
rect 8067 5661 8079 5695
rect 8386 5692 8392 5704
rect 8347 5664 8392 5692
rect 8021 5655 8079 5661
rect 8386 5652 8392 5664
rect 8444 5652 8450 5704
rect 8680 5692 8708 5868
rect 9950 5856 9956 5908
rect 10008 5856 10014 5908
rect 11146 5856 11152 5908
rect 11204 5896 11210 5908
rect 11609 5899 11667 5905
rect 11609 5896 11621 5899
rect 11204 5868 11621 5896
rect 11204 5856 11210 5868
rect 11609 5865 11621 5868
rect 11655 5865 11667 5899
rect 11609 5859 11667 5865
rect 9861 5763 9919 5769
rect 9861 5729 9873 5763
rect 9907 5760 9919 5763
rect 9968 5760 9996 5856
rect 9907 5732 9996 5760
rect 9907 5729 9919 5732
rect 9861 5723 9919 5729
rect 11330 5720 11336 5772
rect 11388 5720 11394 5772
rect 11624 5760 11652 5859
rect 11882 5856 11888 5908
rect 11940 5896 11946 5908
rect 12161 5899 12219 5905
rect 12161 5896 12173 5899
rect 11940 5868 12173 5896
rect 11940 5856 11946 5868
rect 12161 5865 12173 5868
rect 12207 5865 12219 5899
rect 12161 5859 12219 5865
rect 13262 5856 13268 5908
rect 13320 5896 13326 5908
rect 13357 5899 13415 5905
rect 13357 5896 13369 5899
rect 13320 5868 13369 5896
rect 13320 5856 13326 5868
rect 13357 5865 13369 5868
rect 13403 5865 13415 5899
rect 13357 5859 13415 5865
rect 11793 5763 11851 5769
rect 11793 5760 11805 5763
rect 11624 5732 11805 5760
rect 11793 5729 11805 5732
rect 11839 5729 11851 5763
rect 11793 5723 11851 5729
rect 8941 5695 8999 5701
rect 8941 5692 8953 5695
rect 8680 5664 8953 5692
rect 8941 5661 8953 5664
rect 8987 5661 8999 5695
rect 8941 5655 8999 5661
rect 9674 5652 9680 5704
rect 9732 5688 9738 5704
rect 9781 5695 9839 5701
rect 9781 5688 9793 5695
rect 9732 5661 9793 5688
rect 9827 5661 9839 5695
rect 11348 5692 11376 5720
rect 11698 5692 11704 5704
rect 11348 5664 11704 5692
rect 9732 5660 9839 5661
rect 9732 5652 9738 5660
rect 9781 5655 9839 5660
rect 11698 5652 11704 5664
rect 11756 5692 11762 5704
rect 11977 5695 12035 5701
rect 11977 5692 11989 5695
rect 11756 5664 11989 5692
rect 11756 5652 11762 5664
rect 11977 5661 11989 5664
rect 12023 5661 12035 5695
rect 11977 5655 12035 5661
rect 12066 5652 12072 5704
rect 12124 5692 12130 5704
rect 12345 5695 12403 5701
rect 12345 5692 12357 5695
rect 12124 5664 12357 5692
rect 12124 5652 12130 5664
rect 12345 5661 12357 5664
rect 12391 5661 12403 5695
rect 12345 5655 12403 5661
rect 13446 5652 13452 5704
rect 13504 5692 13510 5704
rect 13541 5695 13599 5701
rect 13541 5692 13553 5695
rect 13504 5664 13553 5692
rect 13504 5652 13510 5664
rect 13541 5661 13553 5664
rect 13587 5661 13599 5695
rect 13541 5655 13599 5661
rect 5629 5627 5687 5633
rect 5184 5596 5488 5624
rect 4982 5556 4988 5568
rect 4540 5528 4988 5556
rect 4982 5516 4988 5528
rect 5040 5516 5046 5568
rect 5460 5556 5488 5596
rect 5629 5593 5641 5627
rect 5675 5624 5687 5627
rect 5997 5627 6055 5633
rect 5997 5624 6009 5627
rect 5675 5596 6009 5624
rect 5675 5593 5687 5596
rect 5629 5587 5687 5593
rect 5997 5593 6009 5596
rect 6043 5593 6055 5627
rect 5997 5587 6055 5593
rect 7006 5584 7012 5636
rect 7064 5584 7070 5636
rect 10137 5627 10195 5633
rect 10137 5593 10149 5627
rect 10183 5593 10195 5627
rect 11422 5624 11428 5636
rect 11362 5596 11428 5624
rect 10137 5587 10195 5593
rect 5810 5556 5816 5568
rect 5460 5528 5816 5556
rect 5810 5516 5816 5528
rect 5868 5516 5874 5568
rect 8018 5516 8024 5568
rect 8076 5556 8082 5568
rect 8205 5559 8263 5565
rect 8205 5556 8217 5559
rect 8076 5528 8217 5556
rect 8076 5516 8082 5528
rect 8205 5525 8217 5528
rect 8251 5525 8263 5559
rect 8205 5519 8263 5525
rect 8570 5516 8576 5568
rect 8628 5556 8634 5568
rect 9125 5559 9183 5565
rect 9125 5556 9137 5559
rect 8628 5528 9137 5556
rect 8628 5516 8634 5528
rect 9125 5525 9137 5528
rect 9171 5525 9183 5559
rect 9125 5519 9183 5525
rect 9585 5559 9643 5565
rect 9585 5525 9597 5559
rect 9631 5556 9643 5559
rect 10152 5556 10180 5587
rect 11422 5584 11428 5596
rect 11480 5584 11486 5636
rect 12986 5624 12992 5636
rect 12947 5596 12992 5624
rect 12986 5584 12992 5596
rect 13044 5584 13050 5636
rect 13262 5624 13268 5636
rect 13223 5596 13268 5624
rect 13262 5584 13268 5596
rect 13320 5584 13326 5636
rect 9631 5528 10180 5556
rect 9631 5525 9643 5528
rect 9585 5519 9643 5525
rect 1104 5466 13892 5488
rect 1104 5414 8214 5466
rect 8266 5414 8278 5466
rect 8330 5414 8342 5466
rect 8394 5414 8406 5466
rect 8458 5414 8470 5466
rect 8522 5414 13892 5466
rect 1104 5392 13892 5414
rect 1949 5355 2007 5361
rect 1949 5321 1961 5355
rect 1995 5352 2007 5355
rect 1995 5324 3648 5352
rect 1995 5321 2007 5324
rect 1949 5315 2007 5321
rect 2590 5284 2596 5296
rect 2551 5256 2596 5284
rect 2590 5244 2596 5256
rect 2648 5244 2654 5296
rect 2774 5244 2780 5296
rect 2832 5284 2838 5296
rect 3620 5284 3648 5324
rect 4798 5312 4804 5364
rect 4856 5352 4862 5364
rect 5261 5355 5319 5361
rect 5261 5352 5273 5355
rect 4856 5324 5273 5352
rect 4856 5312 4862 5324
rect 5261 5321 5273 5324
rect 5307 5321 5319 5355
rect 5261 5315 5319 5321
rect 7469 5355 7527 5361
rect 7469 5321 7481 5355
rect 7515 5352 7527 5355
rect 7834 5352 7840 5364
rect 7515 5324 7840 5352
rect 7515 5321 7527 5324
rect 7469 5315 7527 5321
rect 7834 5312 7840 5324
rect 7892 5312 7898 5364
rect 9493 5355 9551 5361
rect 9493 5321 9505 5355
rect 9539 5352 9551 5355
rect 10226 5352 10232 5364
rect 9539 5324 10232 5352
rect 9539 5321 9551 5324
rect 9493 5315 9551 5321
rect 10226 5312 10232 5324
rect 10284 5312 10290 5364
rect 10502 5352 10508 5364
rect 10463 5324 10508 5352
rect 10502 5312 10508 5324
rect 10560 5312 10566 5364
rect 11241 5355 11299 5361
rect 11241 5321 11253 5355
rect 11287 5352 11299 5355
rect 11606 5352 11612 5364
rect 11287 5324 11612 5352
rect 11287 5321 11299 5324
rect 11241 5315 11299 5321
rect 11606 5312 11612 5324
rect 11664 5312 11670 5364
rect 11698 5312 11704 5364
rect 11756 5352 11762 5364
rect 13265 5355 13323 5361
rect 13265 5352 13277 5355
rect 11756 5324 13277 5352
rect 11756 5312 11762 5324
rect 13265 5321 13277 5324
rect 13311 5321 13323 5355
rect 13265 5315 13323 5321
rect 13541 5355 13599 5361
rect 13541 5321 13553 5355
rect 13587 5352 13599 5355
rect 13630 5352 13636 5364
rect 13587 5324 13636 5352
rect 13587 5321 13599 5324
rect 13541 5315 13599 5321
rect 13630 5312 13636 5324
rect 13688 5312 13694 5364
rect 3789 5287 3847 5293
rect 3789 5284 3801 5287
rect 2832 5256 2877 5284
rect 3620 5256 3801 5284
rect 2832 5244 2838 5256
rect 3789 5253 3801 5256
rect 3835 5253 3847 5287
rect 3789 5247 3847 5253
rect 4246 5244 4252 5296
rect 4304 5244 4310 5296
rect 8018 5284 8024 5296
rect 6104 5256 6408 5284
rect 7979 5256 8024 5284
rect 1765 5219 1823 5225
rect 1765 5185 1777 5219
rect 1811 5185 1823 5219
rect 1765 5179 1823 5185
rect 2133 5219 2191 5225
rect 2133 5185 2145 5219
rect 2179 5216 2191 5219
rect 3326 5216 3332 5228
rect 2179 5188 3332 5216
rect 2179 5185 2191 5188
rect 2133 5179 2191 5185
rect 1780 5148 1808 5179
rect 3326 5176 3332 5188
rect 3384 5176 3390 5228
rect 3418 5176 3424 5228
rect 3476 5216 3482 5228
rect 3476 5188 3521 5216
rect 3476 5176 3482 5188
rect 5626 5176 5632 5228
rect 5684 5216 5690 5228
rect 6104 5225 6132 5256
rect 6089 5219 6147 5225
rect 6089 5216 6101 5219
rect 5684 5188 6101 5216
rect 5684 5176 5690 5188
rect 6089 5185 6101 5188
rect 6135 5185 6147 5219
rect 6089 5179 6147 5185
rect 6178 5176 6184 5228
rect 6236 5216 6242 5228
rect 6380 5225 6408 5256
rect 8018 5244 8024 5256
rect 8076 5244 8082 5296
rect 8662 5244 8668 5296
rect 8720 5244 8726 5296
rect 11790 5284 11796 5296
rect 11751 5256 11796 5284
rect 11790 5244 11796 5256
rect 11848 5244 11854 5296
rect 11882 5244 11888 5296
rect 11940 5284 11946 5296
rect 11940 5256 12282 5284
rect 11940 5244 11946 5256
rect 6365 5219 6423 5225
rect 6236 5188 6281 5216
rect 6236 5176 6242 5188
rect 6365 5185 6377 5219
rect 6411 5185 6423 5219
rect 6641 5219 6699 5225
rect 6641 5216 6653 5219
rect 6365 5179 6423 5185
rect 6472 5188 6653 5216
rect 2866 5148 2872 5160
rect 1780 5120 2360 5148
rect 2827 5120 2872 5148
rect 2332 5089 2360 5120
rect 2866 5108 2872 5120
rect 2924 5108 2930 5160
rect 3513 5151 3571 5157
rect 3513 5148 3525 5151
rect 3160 5120 3525 5148
rect 2317 5083 2375 5089
rect 2317 5049 2329 5083
rect 2363 5049 2375 5083
rect 2317 5043 2375 5049
rect 1581 5015 1639 5021
rect 1581 4981 1593 5015
rect 1627 5012 1639 5015
rect 1762 5012 1768 5024
rect 1627 4984 1768 5012
rect 1627 4981 1639 4984
rect 1581 4975 1639 4981
rect 1762 4972 1768 4984
rect 1820 4972 1826 5024
rect 1854 4972 1860 5024
rect 1912 5012 1918 5024
rect 3160 5012 3188 5120
rect 3513 5117 3525 5120
rect 3559 5148 3571 5151
rect 4522 5148 4528 5160
rect 3559 5120 4528 5148
rect 3559 5117 3571 5120
rect 3513 5111 3571 5117
rect 4522 5108 4528 5120
rect 4580 5108 4586 5160
rect 5258 5108 5264 5160
rect 5316 5148 5322 5160
rect 5905 5151 5963 5157
rect 5905 5148 5917 5151
rect 5316 5120 5917 5148
rect 5316 5108 5322 5120
rect 5905 5117 5917 5120
rect 5951 5117 5963 5151
rect 6196 5148 6224 5176
rect 6472 5148 6500 5188
rect 6641 5185 6653 5188
rect 6687 5185 6699 5219
rect 6641 5179 6699 5185
rect 6914 5176 6920 5228
rect 6972 5216 6978 5228
rect 7285 5219 7343 5225
rect 7285 5216 7297 5219
rect 6972 5188 7297 5216
rect 6972 5176 6978 5188
rect 7285 5185 7297 5188
rect 7331 5185 7343 5219
rect 7285 5179 7343 5185
rect 9953 5219 10011 5225
rect 9953 5185 9965 5219
rect 9999 5216 10011 5219
rect 10134 5216 10140 5228
rect 9999 5188 10140 5216
rect 9999 5185 10011 5188
rect 9953 5179 10011 5185
rect 10134 5176 10140 5188
rect 10192 5176 10198 5228
rect 10321 5219 10379 5225
rect 10321 5185 10333 5219
rect 10367 5185 10379 5219
rect 10321 5179 10379 5185
rect 10689 5219 10747 5225
rect 10689 5185 10701 5219
rect 10735 5216 10747 5219
rect 10778 5216 10784 5228
rect 10735 5188 10784 5216
rect 10735 5185 10747 5188
rect 10689 5179 10747 5185
rect 6196 5120 6500 5148
rect 5905 5111 5963 5117
rect 6730 5108 6736 5160
rect 6788 5148 6794 5160
rect 7101 5151 7159 5157
rect 7101 5148 7113 5151
rect 6788 5120 7113 5148
rect 6788 5108 6794 5120
rect 7101 5117 7113 5120
rect 7147 5117 7159 5151
rect 7742 5148 7748 5160
rect 7703 5120 7748 5148
rect 7101 5111 7159 5117
rect 7742 5108 7748 5120
rect 7800 5108 7806 5160
rect 10336 5148 10364 5179
rect 10778 5176 10784 5188
rect 10836 5176 10842 5228
rect 10965 5219 11023 5225
rect 10965 5185 10977 5219
rect 11011 5216 11023 5219
rect 11054 5216 11060 5228
rect 11011 5188 11060 5216
rect 11011 5185 11023 5188
rect 10965 5179 11023 5185
rect 11054 5176 11060 5188
rect 11112 5176 11118 5228
rect 11241 5219 11299 5225
rect 11241 5185 11253 5219
rect 11287 5216 11299 5219
rect 11330 5216 11336 5228
rect 11287 5188 11336 5216
rect 11287 5185 11299 5188
rect 11241 5179 11299 5185
rect 11330 5176 11336 5188
rect 11388 5176 11394 5228
rect 11514 5216 11520 5228
rect 11475 5188 11520 5216
rect 11514 5176 11520 5188
rect 11572 5176 11578 5228
rect 10336 5120 11376 5148
rect 6362 5080 6368 5092
rect 5460 5052 6368 5080
rect 1912 4984 3188 5012
rect 3237 5015 3295 5021
rect 1912 4972 1918 4984
rect 3237 4981 3249 5015
rect 3283 5012 3295 5015
rect 3418 5012 3424 5024
rect 3283 4984 3424 5012
rect 3283 4981 3295 4984
rect 3237 4975 3295 4981
rect 3418 4972 3424 4984
rect 3476 4972 3482 5024
rect 4154 4972 4160 5024
rect 4212 5012 4218 5024
rect 5460 5021 5488 5052
rect 6362 5040 6368 5052
rect 6420 5080 6426 5092
rect 6825 5083 6883 5089
rect 6825 5080 6837 5083
rect 6420 5052 6837 5080
rect 6420 5040 6426 5052
rect 6825 5049 6837 5052
rect 6871 5049 6883 5083
rect 6825 5043 6883 5049
rect 9122 5040 9128 5092
rect 9180 5080 9186 5092
rect 9769 5083 9827 5089
rect 9769 5080 9781 5083
rect 9180 5052 9781 5080
rect 9180 5040 9186 5052
rect 9769 5049 9781 5052
rect 9815 5049 9827 5083
rect 9769 5043 9827 5049
rect 10229 5083 10287 5089
rect 10229 5049 10241 5083
rect 10275 5080 10287 5083
rect 11146 5080 11152 5092
rect 10275 5052 11152 5080
rect 10275 5049 10287 5052
rect 10229 5043 10287 5049
rect 11146 5040 11152 5052
rect 11204 5040 11210 5092
rect 5445 5015 5503 5021
rect 5445 5012 5457 5015
rect 4212 4984 5457 5012
rect 4212 4972 4218 4984
rect 5445 4981 5457 4984
rect 5491 4981 5503 5015
rect 5445 4975 5503 4981
rect 5534 4972 5540 5024
rect 5592 5012 5598 5024
rect 5721 5015 5779 5021
rect 5721 5012 5733 5015
rect 5592 4984 5733 5012
rect 5592 4972 5598 4984
rect 5721 4981 5733 4984
rect 5767 4981 5779 5015
rect 6454 5012 6460 5024
rect 6415 4984 6460 5012
rect 5721 4975 5779 4981
rect 6454 4972 6460 4984
rect 6512 4972 6518 5024
rect 11348 5012 11376 5120
rect 12986 5012 12992 5024
rect 11348 4984 12992 5012
rect 12986 4972 12992 4984
rect 13044 4972 13050 5024
rect 1104 4922 13892 4944
rect 1104 4870 4214 4922
rect 4266 4870 4278 4922
rect 4330 4870 4342 4922
rect 4394 4870 4406 4922
rect 4458 4870 4470 4922
rect 4522 4870 12214 4922
rect 12266 4870 12278 4922
rect 12330 4870 12342 4922
rect 12394 4870 12406 4922
rect 12458 4870 12470 4922
rect 12522 4870 13892 4922
rect 1104 4848 13892 4870
rect 2774 4768 2780 4820
rect 2832 4808 2838 4820
rect 3237 4811 3295 4817
rect 3237 4808 3249 4811
rect 2832 4780 3249 4808
rect 2832 4768 2838 4780
rect 3237 4777 3249 4780
rect 3283 4777 3295 4811
rect 3237 4771 3295 4777
rect 2866 4700 2872 4752
rect 2924 4700 2930 4752
rect 1762 4672 1768 4684
rect 1723 4644 1768 4672
rect 1762 4632 1768 4644
rect 1820 4632 1826 4684
rect 2884 4672 2912 4700
rect 2884 4644 3188 4672
rect 1489 4607 1547 4613
rect 1489 4573 1501 4607
rect 1535 4573 1547 4607
rect 1489 4567 1547 4573
rect 1504 4536 1532 4567
rect 1762 4536 1768 4548
rect 1504 4508 1768 4536
rect 1762 4496 1768 4508
rect 1820 4496 1826 4548
rect 3050 4536 3056 4548
rect 2990 4508 3056 4536
rect 3050 4496 3056 4508
rect 3108 4496 3114 4548
rect 3160 4536 3188 4644
rect 3252 4604 3280 4771
rect 3326 4768 3332 4820
rect 3384 4808 3390 4820
rect 4065 4811 4123 4817
rect 4065 4808 4077 4811
rect 3384 4780 4077 4808
rect 3384 4768 3390 4780
rect 4065 4777 4077 4780
rect 4111 4777 4123 4811
rect 8754 4808 8760 4820
rect 4065 4771 4123 4777
rect 4172 4780 8760 4808
rect 3513 4743 3571 4749
rect 3513 4709 3525 4743
rect 3559 4740 3571 4743
rect 3878 4740 3884 4752
rect 3559 4712 3884 4740
rect 3559 4709 3571 4712
rect 3513 4703 3571 4709
rect 3878 4700 3884 4712
rect 3936 4700 3942 4752
rect 4062 4632 4068 4684
rect 4120 4672 4126 4684
rect 4172 4672 4200 4780
rect 8754 4768 8760 4780
rect 8812 4768 8818 4820
rect 10410 4768 10416 4820
rect 10468 4808 10474 4820
rect 11333 4811 11391 4817
rect 11333 4808 11345 4811
rect 10468 4780 11345 4808
rect 10468 4768 10474 4780
rect 11333 4777 11345 4780
rect 11379 4777 11391 4811
rect 11333 4771 11391 4777
rect 4890 4740 4896 4752
rect 4448 4712 4896 4740
rect 4448 4681 4476 4712
rect 4890 4700 4896 4712
rect 4948 4700 4954 4752
rect 6270 4700 6276 4752
rect 6328 4740 6334 4752
rect 6733 4743 6791 4749
rect 6733 4740 6745 4743
rect 6328 4712 6745 4740
rect 6328 4700 6334 4712
rect 6733 4709 6745 4712
rect 6779 4709 6791 4743
rect 6733 4703 6791 4709
rect 7009 4743 7067 4749
rect 7009 4709 7021 4743
rect 7055 4740 7067 4743
rect 7374 4740 7380 4752
rect 7055 4712 7380 4740
rect 7055 4709 7067 4712
rect 7009 4703 7067 4709
rect 7374 4700 7380 4712
rect 7432 4700 7438 4752
rect 11422 4700 11428 4752
rect 11480 4740 11486 4752
rect 11793 4743 11851 4749
rect 11793 4740 11805 4743
rect 11480 4712 11805 4740
rect 11480 4700 11486 4712
rect 11793 4709 11805 4712
rect 11839 4709 11851 4743
rect 11793 4703 11851 4709
rect 4120 4644 4200 4672
rect 4433 4675 4491 4681
rect 4120 4632 4126 4644
rect 4433 4641 4445 4675
rect 4479 4641 4491 4675
rect 4433 4635 4491 4641
rect 4706 4632 4712 4684
rect 4764 4672 4770 4684
rect 5350 4672 5356 4684
rect 4764 4644 5356 4672
rect 4764 4632 4770 4644
rect 3421 4607 3479 4613
rect 3421 4604 3433 4607
rect 3252 4576 3433 4604
rect 3421 4573 3433 4576
rect 3467 4573 3479 4607
rect 3421 4567 3479 4573
rect 4154 4564 4160 4616
rect 4212 4604 4218 4616
rect 4724 4604 4752 4632
rect 5000 4613 5028 4644
rect 5350 4632 5356 4644
rect 5408 4632 5414 4684
rect 7742 4632 7748 4684
rect 7800 4672 7806 4684
rect 8757 4675 8815 4681
rect 8757 4672 8769 4675
rect 7800 4644 8769 4672
rect 7800 4632 7806 4644
rect 8757 4641 8769 4644
rect 8803 4672 8815 4675
rect 9585 4675 9643 4681
rect 9585 4672 9597 4675
rect 8803 4644 9597 4672
rect 8803 4641 8815 4644
rect 8757 4635 8815 4641
rect 9585 4641 9597 4644
rect 9631 4672 9643 4675
rect 9950 4672 9956 4684
rect 9631 4644 9956 4672
rect 9631 4641 9643 4644
rect 9585 4635 9643 4641
rect 9950 4632 9956 4644
rect 10008 4672 10014 4684
rect 11514 4672 11520 4684
rect 10008 4644 11520 4672
rect 10008 4632 10014 4644
rect 11514 4632 11520 4644
rect 11572 4632 11578 4684
rect 4212 4576 4752 4604
rect 4985 4607 5043 4613
rect 4212 4564 4218 4576
rect 4985 4573 4997 4607
rect 5031 4573 5043 4607
rect 4985 4567 5043 4573
rect 8846 4564 8852 4616
rect 8904 4604 8910 4616
rect 9125 4607 9183 4613
rect 9125 4604 9137 4607
rect 8904 4576 9137 4604
rect 8904 4564 8910 4576
rect 9125 4573 9137 4576
rect 9171 4573 9183 4607
rect 11606 4604 11612 4616
rect 11567 4576 11612 4604
rect 9125 4567 9183 4573
rect 3789 4539 3847 4545
rect 3789 4536 3801 4539
rect 3160 4508 3801 4536
rect 3789 4505 3801 4508
rect 3835 4505 3847 4539
rect 4614 4536 4620 4548
rect 4575 4508 4620 4536
rect 3789 4499 3847 4505
rect 4614 4496 4620 4508
rect 4672 4496 4678 4548
rect 4893 4539 4951 4545
rect 4893 4505 4905 4539
rect 4939 4536 4951 4539
rect 5166 4536 5172 4548
rect 4939 4508 5172 4536
rect 4939 4505 4951 4508
rect 4893 4499 4951 4505
rect 5166 4496 5172 4508
rect 5224 4496 5230 4548
rect 5261 4539 5319 4545
rect 5261 4505 5273 4539
rect 5307 4536 5319 4539
rect 5534 4536 5540 4548
rect 5307 4508 5540 4536
rect 5307 4505 5319 4508
rect 5261 4499 5319 4505
rect 5534 4496 5540 4508
rect 5592 4496 5598 4548
rect 6914 4536 6920 4548
rect 6486 4508 6920 4536
rect 6914 4496 6920 4508
rect 6972 4496 6978 4548
rect 7926 4496 7932 4548
rect 7984 4496 7990 4548
rect 8481 4539 8539 4545
rect 8481 4505 8493 4539
rect 8527 4536 8539 4539
rect 8570 4536 8576 4548
rect 8527 4508 8576 4536
rect 8527 4505 8539 4508
rect 8481 4499 8539 4505
rect 8570 4496 8576 4508
rect 8628 4496 8634 4548
rect 9140 4536 9168 4567
rect 11606 4564 11612 4576
rect 11664 4564 11670 4616
rect 11701 4607 11759 4613
rect 11701 4573 11713 4607
rect 11747 4573 11759 4607
rect 11974 4604 11980 4616
rect 11935 4576 11980 4604
rect 11701 4567 11759 4573
rect 9140 4508 9720 4536
rect 2774 4428 2780 4480
rect 2832 4468 2838 4480
rect 3234 4468 3240 4480
rect 2832 4440 3240 4468
rect 2832 4428 2838 4440
rect 3234 4428 3240 4440
rect 3292 4428 3298 4480
rect 4525 4471 4583 4477
rect 4525 4437 4537 4471
rect 4571 4468 4583 4471
rect 4706 4468 4712 4480
rect 4571 4440 4712 4468
rect 4571 4437 4583 4440
rect 4525 4431 4583 4437
rect 4706 4428 4712 4440
rect 4764 4428 4770 4480
rect 9125 4471 9183 4477
rect 9125 4437 9137 4471
rect 9171 4468 9183 4471
rect 9214 4468 9220 4480
rect 9171 4440 9220 4468
rect 9171 4437 9183 4440
rect 9125 4431 9183 4437
rect 9214 4428 9220 4440
rect 9272 4428 9278 4480
rect 9692 4468 9720 4508
rect 9766 4496 9772 4548
rect 9824 4536 9830 4548
rect 9861 4539 9919 4545
rect 9861 4536 9873 4539
rect 9824 4508 9873 4536
rect 9824 4496 9830 4508
rect 9861 4505 9873 4508
rect 9907 4505 9919 4539
rect 9861 4499 9919 4505
rect 10594 4496 10600 4548
rect 10652 4496 10658 4548
rect 11146 4496 11152 4548
rect 11204 4536 11210 4548
rect 11422 4536 11428 4548
rect 11204 4508 11428 4536
rect 11204 4496 11210 4508
rect 11422 4496 11428 4508
rect 11480 4496 11486 4548
rect 11514 4496 11520 4548
rect 11572 4536 11578 4548
rect 11716 4536 11744 4567
rect 11974 4564 11980 4576
rect 12032 4564 12038 4616
rect 13262 4604 13268 4616
rect 13223 4576 13268 4604
rect 13262 4564 13268 4576
rect 13320 4564 13326 4616
rect 11572 4508 11744 4536
rect 13541 4539 13599 4545
rect 11572 4496 11578 4508
rect 13541 4505 13553 4539
rect 13587 4505 13599 4539
rect 13541 4499 13599 4505
rect 11790 4468 11796 4480
rect 9692 4440 11796 4468
rect 11790 4428 11796 4440
rect 11848 4468 11854 4480
rect 13078 4468 13084 4480
rect 11848 4440 13084 4468
rect 11848 4428 11854 4440
rect 13078 4428 13084 4440
rect 13136 4468 13142 4480
rect 13556 4468 13584 4499
rect 13136 4440 13584 4468
rect 13136 4428 13142 4440
rect 1104 4378 13892 4400
rect 1104 4326 8214 4378
rect 8266 4326 8278 4378
rect 8330 4326 8342 4378
rect 8394 4326 8406 4378
rect 8458 4326 8470 4378
rect 8522 4326 13892 4378
rect 1104 4304 13892 4326
rect 3050 4224 3056 4276
rect 3108 4264 3114 4276
rect 3237 4267 3295 4273
rect 3237 4264 3249 4267
rect 3108 4236 3249 4264
rect 3108 4224 3114 4236
rect 3237 4233 3249 4236
rect 3283 4233 3295 4267
rect 3237 4227 3295 4233
rect 3418 4224 3424 4276
rect 3476 4264 3482 4276
rect 3476 4236 4476 4264
rect 3476 4224 3482 4236
rect 4448 4205 4476 4236
rect 5718 4224 5724 4276
rect 5776 4264 5782 4276
rect 6549 4267 6607 4273
rect 6549 4264 6561 4267
rect 5776 4236 6561 4264
rect 5776 4224 5782 4236
rect 6549 4233 6561 4236
rect 6595 4233 6607 4267
rect 7006 4264 7012 4276
rect 6967 4236 7012 4264
rect 6549 4227 6607 4233
rect 7006 4224 7012 4236
rect 7064 4224 7070 4276
rect 7098 4224 7104 4276
rect 7156 4264 7162 4276
rect 10594 4264 10600 4276
rect 7156 4236 10088 4264
rect 10555 4236 10600 4264
rect 7156 4224 7162 4236
rect 4433 4199 4491 4205
rect 4433 4165 4445 4199
rect 4479 4165 4491 4199
rect 4433 4159 4491 4165
rect 5166 4156 5172 4208
rect 5224 4156 5230 4208
rect 6362 4196 6368 4208
rect 6323 4168 6368 4196
rect 6362 4156 6368 4168
rect 6420 4156 6426 4208
rect 6822 4156 6828 4208
rect 6880 4196 6886 4208
rect 8294 4196 8300 4208
rect 6880 4168 7328 4196
rect 6880 4156 6886 4168
rect 1673 4131 1731 4137
rect 1673 4097 1685 4131
rect 1719 4128 1731 4131
rect 1946 4128 1952 4140
rect 1719 4100 1952 4128
rect 1719 4097 1731 4100
rect 1673 4091 1731 4097
rect 1946 4088 1952 4100
rect 2004 4088 2010 4140
rect 2222 4128 2228 4140
rect 2183 4100 2228 4128
rect 2222 4088 2228 4100
rect 2280 4088 2286 4140
rect 2774 4088 2780 4140
rect 2832 4128 2838 4140
rect 2869 4131 2927 4137
rect 2869 4128 2881 4131
rect 2832 4100 2881 4128
rect 2832 4088 2838 4100
rect 2869 4097 2881 4100
rect 2915 4097 2927 4131
rect 2869 4091 2927 4097
rect 3329 4131 3387 4137
rect 3329 4097 3341 4131
rect 3375 4128 3387 4131
rect 3418 4128 3424 4140
rect 3375 4100 3424 4128
rect 3375 4097 3387 4100
rect 3329 4091 3387 4097
rect 3418 4088 3424 4100
rect 3476 4088 3482 4140
rect 3513 4131 3571 4137
rect 3513 4097 3525 4131
rect 3559 4097 3571 4131
rect 3694 4128 3700 4140
rect 3655 4100 3700 4128
rect 3513 4091 3571 4097
rect 1765 4063 1823 4069
rect 1765 4029 1777 4063
rect 1811 4029 1823 4063
rect 2038 4060 2044 4072
rect 1999 4032 2044 4060
rect 1765 4023 1823 4029
rect 1780 3992 1808 4023
rect 2038 4020 2044 4032
rect 2096 4020 2102 4072
rect 2130 4020 2136 4072
rect 2188 4060 2194 4072
rect 2685 4063 2743 4069
rect 2685 4060 2697 4063
rect 2188 4032 2233 4060
rect 2332 4032 2697 4060
rect 2188 4020 2194 4032
rect 1854 3992 1860 4004
rect 1767 3964 1860 3992
rect 1854 3952 1860 3964
rect 1912 3992 1918 4004
rect 2332 3992 2360 4032
rect 2685 4029 2697 4032
rect 2731 4029 2743 4063
rect 3050 4060 3056 4072
rect 3011 4032 3056 4060
rect 2685 4023 2743 4029
rect 3050 4020 3056 4032
rect 3108 4020 3114 4072
rect 3528 4060 3556 4091
rect 3694 4088 3700 4100
rect 3752 4088 3758 4140
rect 3881 4131 3939 4137
rect 3881 4097 3893 4131
rect 3927 4128 3939 4131
rect 3970 4128 3976 4140
rect 3927 4100 3976 4128
rect 3927 4097 3939 4100
rect 3881 4091 3939 4097
rect 3970 4088 3976 4100
rect 4028 4088 4034 4140
rect 4154 4128 4160 4140
rect 4212 4137 4218 4140
rect 4122 4100 4160 4128
rect 4154 4088 4160 4100
rect 4212 4091 4222 4137
rect 7006 4128 7012 4140
rect 6967 4100 7012 4128
rect 4212 4088 4218 4091
rect 7006 4088 7012 4100
rect 7064 4088 7070 4140
rect 7190 4128 7196 4140
rect 7151 4100 7196 4128
rect 7190 4088 7196 4100
rect 7248 4088 7254 4140
rect 7300 4128 7328 4168
rect 7760 4168 8300 4196
rect 7653 4131 7711 4137
rect 7653 4128 7665 4131
rect 7300 4100 7665 4128
rect 7653 4097 7665 4100
rect 7699 4128 7711 4131
rect 7760 4128 7788 4168
rect 8294 4156 8300 4168
rect 8352 4156 8358 4208
rect 9030 4156 9036 4208
rect 9088 4156 9094 4208
rect 10060 4137 10088 4236
rect 10594 4224 10600 4236
rect 10652 4224 10658 4276
rect 11241 4267 11299 4273
rect 11241 4233 11253 4267
rect 11287 4264 11299 4267
rect 11882 4264 11888 4276
rect 11287 4236 11888 4264
rect 11287 4233 11299 4236
rect 11241 4227 11299 4233
rect 11882 4224 11888 4236
rect 11940 4224 11946 4276
rect 11606 4196 11612 4208
rect 10612 4168 11612 4196
rect 9953 4131 10011 4137
rect 9953 4128 9965 4131
rect 7699 4100 7788 4128
rect 9232 4100 9965 4128
rect 7699 4097 7711 4100
rect 7653 4091 7711 4097
rect 4065 4063 4123 4069
rect 3528 4032 3924 4060
rect 3896 4004 3924 4032
rect 4065 4029 4077 4063
rect 4111 4060 4123 4063
rect 4111 4032 4200 4060
rect 4111 4029 4123 4032
rect 4065 4023 4123 4029
rect 1912 3964 2360 3992
rect 2409 3995 2467 4001
rect 1912 3952 1918 3964
rect 2409 3961 2421 3995
rect 2455 3992 2467 3995
rect 2958 3992 2964 4004
rect 2455 3964 2964 3992
rect 2455 3961 2467 3964
rect 2409 3955 2467 3961
rect 2958 3952 2964 3964
rect 3016 3952 3022 4004
rect 3878 3952 3884 4004
rect 3936 3952 3942 4004
rect 1486 3924 1492 3936
rect 1447 3896 1492 3924
rect 1486 3884 1492 3896
rect 1544 3884 1550 3936
rect 2314 3884 2320 3936
rect 2372 3924 2378 3936
rect 2590 3924 2596 3936
rect 2372 3896 2596 3924
rect 2372 3884 2378 3896
rect 2590 3884 2596 3896
rect 2648 3884 2654 3936
rect 4172 3924 4200 4032
rect 5442 4020 5448 4072
rect 5500 4060 5506 4072
rect 7742 4060 7748 4072
rect 5500 4032 7748 4060
rect 5500 4020 5506 4032
rect 7742 4020 7748 4032
rect 7800 4020 7806 4072
rect 8021 4063 8079 4069
rect 8021 4029 8033 4063
rect 8067 4060 8079 4063
rect 8110 4060 8116 4072
rect 8067 4032 8116 4060
rect 8067 4029 8079 4032
rect 8021 4023 8079 4029
rect 8110 4020 8116 4032
rect 8168 4020 8174 4072
rect 8386 4020 8392 4072
rect 8444 4060 8450 4072
rect 9232 4060 9260 4100
rect 9953 4097 9965 4100
rect 9999 4097 10011 4131
rect 9953 4091 10011 4097
rect 10045 4131 10103 4137
rect 10045 4097 10057 4131
rect 10091 4128 10103 4131
rect 10134 4128 10140 4140
rect 10091 4100 10140 4128
rect 10091 4097 10103 4100
rect 10045 4091 10103 4097
rect 10134 4088 10140 4100
rect 10192 4088 10198 4140
rect 10612 4137 10640 4168
rect 11606 4156 11612 4168
rect 11664 4156 11670 4208
rect 13354 4196 13360 4208
rect 13315 4168 13360 4196
rect 13354 4156 13360 4168
rect 13412 4156 13418 4208
rect 10597 4131 10655 4137
rect 10597 4097 10609 4131
rect 10643 4097 10655 4131
rect 10597 4091 10655 4097
rect 10781 4131 10839 4137
rect 10781 4097 10793 4131
rect 10827 4097 10839 4131
rect 10781 4091 10839 4097
rect 11057 4131 11115 4137
rect 11057 4097 11069 4131
rect 11103 4097 11115 4131
rect 11057 4091 11115 4097
rect 11149 4131 11207 4137
rect 11149 4097 11161 4131
rect 11195 4097 11207 4131
rect 11149 4091 11207 4097
rect 8444 4032 9260 4060
rect 9493 4063 9551 4069
rect 8444 4020 8450 4032
rect 9493 4029 9505 4063
rect 9539 4060 9551 4063
rect 9582 4060 9588 4072
rect 9539 4032 9588 4060
rect 9539 4029 9551 4032
rect 9493 4023 9551 4029
rect 9582 4020 9588 4032
rect 9640 4020 9646 4072
rect 10796 4060 10824 4091
rect 11072 4060 11100 4091
rect 9692 4032 10824 4060
rect 10888 4032 11100 4060
rect 5460 3964 6592 3992
rect 5460 3936 5488 3964
rect 5442 3924 5448 3936
rect 4172 3896 5448 3924
rect 5442 3884 5448 3896
rect 5500 3884 5506 3936
rect 5902 3924 5908 3936
rect 5863 3896 5908 3924
rect 5902 3884 5908 3896
rect 5960 3884 5966 3936
rect 6086 3924 6092 3936
rect 6047 3896 6092 3924
rect 6086 3884 6092 3896
rect 6144 3884 6150 3936
rect 6564 3933 6592 3964
rect 9692 3936 9720 4032
rect 9769 3995 9827 4001
rect 9769 3961 9781 3995
rect 9815 3992 9827 3995
rect 10502 3992 10508 4004
rect 9815 3964 10508 3992
rect 9815 3961 9827 3964
rect 9769 3955 9827 3961
rect 10502 3952 10508 3964
rect 10560 3992 10566 4004
rect 10888 3992 10916 4032
rect 11164 3992 11192 4091
rect 11330 4088 11336 4140
rect 11388 4128 11394 4140
rect 11517 4131 11575 4137
rect 11517 4128 11529 4131
rect 11388 4100 11529 4128
rect 11388 4088 11394 4100
rect 11517 4097 11529 4100
rect 11563 4097 11575 4131
rect 11517 4091 11575 4097
rect 11790 4088 11796 4140
rect 11848 4128 11854 4140
rect 11977 4131 12035 4137
rect 11977 4128 11989 4131
rect 11848 4100 11989 4128
rect 11848 4088 11854 4100
rect 11977 4097 11989 4100
rect 12023 4097 12035 4131
rect 11977 4091 12035 4097
rect 12066 4088 12072 4140
rect 12124 4128 12130 4140
rect 12529 4131 12587 4137
rect 12529 4128 12541 4131
rect 12124 4100 12541 4128
rect 12124 4088 12130 4100
rect 12529 4097 12541 4100
rect 12575 4097 12587 4131
rect 12986 4128 12992 4140
rect 12947 4100 12992 4128
rect 12529 4091 12587 4097
rect 12986 4088 12992 4100
rect 13044 4088 13050 4140
rect 11422 4020 11428 4072
rect 11480 4060 11486 4072
rect 11885 4063 11943 4069
rect 11885 4060 11897 4063
rect 11480 4032 11897 4060
rect 11480 4020 11486 4032
rect 11885 4029 11897 4032
rect 11931 4029 11943 4063
rect 11885 4023 11943 4029
rect 12437 4063 12495 4069
rect 12437 4029 12449 4063
rect 12483 4060 12495 4063
rect 12802 4060 12808 4072
rect 12483 4032 12808 4060
rect 12483 4029 12495 4032
rect 12437 4023 12495 4029
rect 11514 3992 11520 4004
rect 10560 3964 10916 3992
rect 11072 3964 11520 3992
rect 10560 3952 10566 3964
rect 6549 3927 6607 3933
rect 6549 3893 6561 3927
rect 6595 3893 6607 3927
rect 6549 3887 6607 3893
rect 6638 3884 6644 3936
rect 6696 3924 6702 3936
rect 6733 3927 6791 3933
rect 6733 3924 6745 3927
rect 6696 3896 6745 3924
rect 6696 3884 6702 3896
rect 6733 3893 6745 3896
rect 6779 3893 6791 3927
rect 6733 3887 6791 3893
rect 7469 3927 7527 3933
rect 7469 3893 7481 3927
rect 7515 3924 7527 3927
rect 8110 3924 8116 3936
rect 7515 3896 8116 3924
rect 7515 3893 7527 3896
rect 7469 3887 7527 3893
rect 8110 3884 8116 3896
rect 8168 3884 8174 3936
rect 9674 3884 9680 3936
rect 9732 3924 9738 3936
rect 10229 3927 10287 3933
rect 10229 3924 10241 3927
rect 9732 3896 10241 3924
rect 9732 3884 9738 3896
rect 10229 3893 10241 3896
rect 10275 3924 10287 3927
rect 11072 3924 11100 3964
rect 11514 3952 11520 3964
rect 11572 3952 11578 4004
rect 12066 3952 12072 4004
rect 12124 3992 12130 4004
rect 12452 3992 12480 4023
rect 12802 4020 12808 4032
rect 12860 4020 12866 4072
rect 13081 4063 13139 4069
rect 13081 4029 13093 4063
rect 13127 4060 13139 4063
rect 13170 4060 13176 4072
rect 13127 4032 13176 4060
rect 13127 4029 13139 4032
rect 13081 4023 13139 4029
rect 13170 4020 13176 4032
rect 13228 4020 13234 4072
rect 12124 3964 12480 3992
rect 12124 3952 12130 3964
rect 11698 3924 11704 3936
rect 10275 3896 11100 3924
rect 11659 3896 11704 3924
rect 10275 3893 10287 3896
rect 10229 3887 10287 3893
rect 11698 3884 11704 3896
rect 11756 3884 11762 3936
rect 13265 3927 13323 3933
rect 13265 3893 13277 3927
rect 13311 3924 13323 3927
rect 13446 3924 13452 3936
rect 13311 3896 13452 3924
rect 13311 3893 13323 3896
rect 13265 3887 13323 3893
rect 13446 3884 13452 3896
rect 13504 3884 13510 3936
rect 1104 3834 13892 3856
rect 1104 3782 4214 3834
rect 4266 3782 4278 3834
rect 4330 3782 4342 3834
rect 4394 3782 4406 3834
rect 4458 3782 4470 3834
rect 4522 3782 12214 3834
rect 12266 3782 12278 3834
rect 12330 3782 12342 3834
rect 12394 3782 12406 3834
rect 12458 3782 12470 3834
rect 12522 3782 13892 3834
rect 1104 3760 13892 3782
rect 1394 3720 1400 3732
rect 1355 3692 1400 3720
rect 1394 3680 1400 3692
rect 1452 3680 1458 3732
rect 1670 3720 1676 3732
rect 1631 3692 1676 3720
rect 1670 3680 1676 3692
rect 1728 3680 1734 3732
rect 3326 3680 3332 3732
rect 3384 3720 3390 3732
rect 3513 3723 3571 3729
rect 3513 3720 3525 3723
rect 3384 3692 3525 3720
rect 3384 3680 3390 3692
rect 3513 3689 3525 3692
rect 3559 3689 3571 3723
rect 3513 3683 3571 3689
rect 5074 3680 5080 3732
rect 5132 3720 5138 3732
rect 5902 3720 5908 3732
rect 5132 3692 5908 3720
rect 5132 3680 5138 3692
rect 5902 3680 5908 3692
rect 5960 3680 5966 3732
rect 5994 3680 6000 3732
rect 6052 3720 6058 3732
rect 6362 3720 6368 3732
rect 6052 3692 6368 3720
rect 6052 3680 6058 3692
rect 6362 3680 6368 3692
rect 6420 3680 6426 3732
rect 7098 3720 7104 3732
rect 6472 3692 7104 3720
rect 1486 3612 1492 3664
rect 1544 3652 1550 3664
rect 2682 3652 2688 3664
rect 1544 3624 2688 3652
rect 1544 3612 1550 3624
rect 2682 3612 2688 3624
rect 2740 3612 2746 3664
rect 3418 3612 3424 3664
rect 3476 3652 3482 3664
rect 4890 3652 4896 3664
rect 3476 3624 4896 3652
rect 3476 3612 3482 3624
rect 4890 3612 4896 3624
rect 4948 3612 4954 3664
rect 5166 3612 5172 3664
rect 5224 3652 5230 3664
rect 5353 3655 5411 3661
rect 5353 3652 5365 3655
rect 5224 3624 5365 3652
rect 5224 3612 5230 3624
rect 5353 3621 5365 3624
rect 5399 3621 5411 3655
rect 6472 3652 6500 3692
rect 7098 3680 7104 3692
rect 7156 3680 7162 3732
rect 7855 3723 7913 3729
rect 7855 3689 7867 3723
rect 7901 3720 7913 3723
rect 11698 3720 11704 3732
rect 7901 3692 11704 3720
rect 7901 3689 7913 3692
rect 7855 3683 7913 3689
rect 11698 3680 11704 3692
rect 11756 3680 11762 3732
rect 11974 3680 11980 3732
rect 12032 3720 12038 3732
rect 12345 3723 12403 3729
rect 12345 3720 12357 3723
rect 12032 3692 12357 3720
rect 12032 3680 12038 3692
rect 12345 3689 12357 3692
rect 12391 3689 12403 3723
rect 12345 3683 12403 3689
rect 13078 3680 13084 3732
rect 13136 3720 13142 3732
rect 13357 3723 13415 3729
rect 13357 3720 13369 3723
rect 13136 3692 13369 3720
rect 13136 3680 13142 3692
rect 13357 3689 13369 3692
rect 13403 3689 13415 3723
rect 13357 3683 13415 3689
rect 8662 3652 8668 3664
rect 5353 3615 5411 3621
rect 5552 3624 6500 3652
rect 8623 3624 8668 3652
rect 2409 3587 2467 3593
rect 2409 3553 2421 3587
rect 2455 3584 2467 3587
rect 2774 3584 2780 3596
rect 2455 3556 2780 3584
rect 2455 3553 2467 3556
rect 2409 3547 2467 3553
rect 2774 3544 2780 3556
rect 2832 3544 2838 3596
rect 4709 3587 4767 3593
rect 4709 3553 4721 3587
rect 4755 3584 4767 3587
rect 5442 3584 5448 3596
rect 4755 3556 5448 3584
rect 4755 3553 4767 3556
rect 4709 3547 4767 3553
rect 5442 3544 5448 3556
rect 5500 3544 5506 3596
rect 1854 3516 1860 3528
rect 1815 3488 1860 3516
rect 1854 3476 1860 3488
rect 1912 3476 1918 3528
rect 2038 3516 2044 3528
rect 1999 3488 2044 3516
rect 2038 3476 2044 3488
rect 2096 3476 2102 3528
rect 3142 3516 3148 3528
rect 3103 3488 3148 3516
rect 3142 3476 3148 3488
rect 3200 3476 3206 3528
rect 3329 3519 3387 3525
rect 3329 3485 3341 3519
rect 3375 3516 3387 3519
rect 3510 3516 3516 3528
rect 3375 3488 3516 3516
rect 3375 3485 3387 3488
rect 3329 3479 3387 3485
rect 3510 3476 3516 3488
rect 3568 3516 3574 3528
rect 3881 3519 3939 3525
rect 3881 3516 3893 3519
rect 3568 3488 3893 3516
rect 3568 3476 3574 3488
rect 3881 3485 3893 3488
rect 3927 3485 3939 3519
rect 3881 3479 3939 3485
rect 3970 3476 3976 3528
rect 4028 3516 4034 3528
rect 5077 3519 5135 3525
rect 5077 3516 5089 3519
rect 4028 3488 4278 3516
rect 4908 3488 5089 3516
rect 4028 3476 4034 3488
rect 2130 3448 2136 3460
rect 2091 3420 2136 3448
rect 2130 3408 2136 3420
rect 2188 3408 2194 3460
rect 2314 3408 2320 3460
rect 2372 3448 2378 3460
rect 4062 3448 4068 3460
rect 2372 3420 4068 3448
rect 2372 3408 2378 3420
rect 4062 3408 4068 3420
rect 4120 3408 4126 3460
rect 1946 3340 1952 3392
rect 2004 3380 2010 3392
rect 3326 3380 3332 3392
rect 2004 3352 3332 3380
rect 2004 3340 2010 3352
rect 3326 3340 3332 3352
rect 3384 3340 3390 3392
rect 3694 3340 3700 3392
rect 3752 3380 3758 3392
rect 3878 3380 3884 3392
rect 3752 3352 3884 3380
rect 3752 3340 3758 3352
rect 3878 3340 3884 3352
rect 3936 3380 3942 3392
rect 4908 3380 4936 3488
rect 5077 3485 5089 3488
rect 5123 3485 5135 3519
rect 5077 3479 5135 3485
rect 5353 3519 5411 3525
rect 5353 3485 5365 3519
rect 5399 3516 5411 3519
rect 5552 3516 5580 3624
rect 8662 3612 8668 3624
rect 8720 3612 8726 3664
rect 9030 3652 9036 3664
rect 8991 3624 9036 3652
rect 9030 3612 9036 3624
rect 9088 3612 9094 3664
rect 9674 3652 9680 3664
rect 9232 3624 9680 3652
rect 5902 3584 5908 3596
rect 5863 3556 5908 3584
rect 5902 3544 5908 3556
rect 5960 3584 5966 3596
rect 6638 3584 6644 3596
rect 5960 3556 6644 3584
rect 5960 3544 5966 3556
rect 6638 3544 6644 3556
rect 6696 3544 6702 3596
rect 7742 3544 7748 3596
rect 7800 3584 7806 3596
rect 8113 3587 8171 3593
rect 8113 3584 8125 3587
rect 7800 3556 8125 3584
rect 7800 3544 7806 3556
rect 8113 3553 8125 3556
rect 8159 3553 8171 3587
rect 8113 3547 8171 3553
rect 8297 3587 8355 3593
rect 8297 3553 8309 3587
rect 8343 3584 8355 3587
rect 8754 3584 8760 3596
rect 8343 3556 8760 3584
rect 8343 3553 8355 3556
rect 8297 3547 8355 3553
rect 8754 3544 8760 3556
rect 8812 3544 8818 3596
rect 9122 3584 9128 3596
rect 8864 3556 9128 3584
rect 5399 3488 5580 3516
rect 5721 3519 5779 3525
rect 5399 3485 5411 3488
rect 5353 3479 5411 3485
rect 5721 3485 5733 3519
rect 5767 3516 5779 3519
rect 5810 3516 5816 3528
rect 5767 3488 5816 3516
rect 5767 3485 5779 3488
rect 5721 3479 5779 3485
rect 4982 3408 4988 3460
rect 5040 3448 5046 3460
rect 5368 3448 5396 3479
rect 5810 3476 5816 3488
rect 5868 3476 5874 3528
rect 6089 3519 6147 3525
rect 6089 3516 6101 3519
rect 5920 3488 6101 3516
rect 5040 3420 5396 3448
rect 5040 3408 5046 3420
rect 5534 3408 5540 3460
rect 5592 3448 5598 3460
rect 5920 3448 5948 3488
rect 6089 3485 6101 3488
rect 6135 3516 6147 3519
rect 6454 3516 6460 3528
rect 6135 3488 6460 3516
rect 6135 3485 6147 3488
rect 6089 3479 6147 3485
rect 6454 3476 6460 3488
rect 6512 3476 6518 3528
rect 8202 3476 8208 3528
rect 8260 3516 8266 3528
rect 8389 3519 8447 3525
rect 8389 3516 8401 3519
rect 8260 3488 8401 3516
rect 8260 3476 8266 3488
rect 8389 3485 8401 3488
rect 8435 3485 8447 3519
rect 8570 3516 8576 3528
rect 8531 3488 8576 3516
rect 8389 3479 8447 3485
rect 5592 3420 5948 3448
rect 5997 3451 6055 3457
rect 5592 3408 5598 3420
rect 5997 3417 6009 3451
rect 6043 3417 6055 3451
rect 7558 3448 7564 3460
rect 7406 3420 7564 3448
rect 5997 3411 6055 3417
rect 3936 3352 4936 3380
rect 6012 3380 6040 3411
rect 7558 3408 7564 3420
rect 7616 3408 7622 3460
rect 8404 3448 8432 3479
rect 8570 3476 8576 3488
rect 8628 3516 8634 3528
rect 8864 3516 8892 3556
rect 9122 3544 9128 3556
rect 9180 3544 9186 3596
rect 9030 3516 9036 3528
rect 8628 3488 8892 3516
rect 8991 3488 9036 3516
rect 8628 3476 8634 3488
rect 9030 3476 9036 3488
rect 9088 3516 9094 3528
rect 9232 3516 9260 3624
rect 9674 3612 9680 3624
rect 9732 3612 9738 3664
rect 11238 3612 11244 3664
rect 11296 3652 11302 3664
rect 11425 3655 11483 3661
rect 11425 3652 11437 3655
rect 11296 3624 11437 3652
rect 11296 3612 11302 3624
rect 11425 3621 11437 3624
rect 11471 3621 11483 3655
rect 11425 3615 11483 3621
rect 11514 3612 11520 3664
rect 11572 3652 11578 3664
rect 11572 3624 11836 3652
rect 11572 3612 11578 3624
rect 9324 3556 11652 3584
rect 9324 3525 9352 3556
rect 11624 3528 11652 3556
rect 9088 3488 9260 3516
rect 9309 3519 9367 3525
rect 9088 3476 9094 3488
rect 9309 3485 9321 3519
rect 9355 3485 9367 3519
rect 9309 3479 9367 3485
rect 9324 3448 9352 3479
rect 9490 3476 9496 3528
rect 9548 3516 9554 3528
rect 9677 3519 9735 3525
rect 9677 3516 9689 3519
rect 9548 3488 9689 3516
rect 9548 3476 9554 3488
rect 9677 3485 9689 3488
rect 9723 3485 9735 3519
rect 11606 3516 11612 3528
rect 11567 3488 11612 3516
rect 9677 3479 9735 3485
rect 11606 3476 11612 3488
rect 11664 3476 11670 3528
rect 11808 3525 11836 3624
rect 12894 3584 12900 3596
rect 12636 3556 12900 3584
rect 11793 3519 11851 3525
rect 11793 3485 11805 3519
rect 11839 3485 11851 3519
rect 11793 3479 11851 3485
rect 11974 3476 11980 3528
rect 12032 3516 12038 3528
rect 12636 3525 12664 3556
rect 12894 3544 12900 3556
rect 12952 3544 12958 3596
rect 12253 3519 12311 3525
rect 12253 3516 12265 3519
rect 12032 3488 12265 3516
rect 12032 3476 12038 3488
rect 12253 3485 12265 3488
rect 12299 3516 12311 3519
rect 12621 3519 12679 3525
rect 12299 3488 12434 3516
rect 12299 3485 12311 3488
rect 12253 3479 12311 3485
rect 8404 3420 9352 3448
rect 9953 3451 10011 3457
rect 9953 3417 9965 3451
rect 9999 3448 10011 3451
rect 10042 3448 10048 3460
rect 9999 3420 10048 3448
rect 9999 3417 10011 3420
rect 9953 3411 10011 3417
rect 10042 3408 10048 3420
rect 10100 3408 10106 3460
rect 12066 3448 12072 3460
rect 11178 3420 11744 3448
rect 12027 3420 12072 3448
rect 6270 3380 6276 3392
rect 6012 3352 6276 3380
rect 3936 3340 3942 3352
rect 6270 3340 6276 3352
rect 6328 3340 6334 3392
rect 6822 3340 6828 3392
rect 6880 3380 6886 3392
rect 8754 3380 8760 3392
rect 6880 3352 8760 3380
rect 6880 3340 6886 3352
rect 8754 3340 8760 3352
rect 8812 3340 8818 3392
rect 9122 3340 9128 3392
rect 9180 3380 9186 3392
rect 11716 3389 11744 3420
rect 12066 3408 12072 3420
rect 12124 3408 12130 3460
rect 12406 3448 12434 3488
rect 12621 3485 12633 3519
rect 12667 3485 12679 3519
rect 12621 3479 12679 3485
rect 12713 3519 12771 3525
rect 12713 3485 12725 3519
rect 12759 3516 12771 3519
rect 12989 3519 13047 3525
rect 12989 3516 13001 3519
rect 12759 3488 13001 3516
rect 12759 3485 12771 3488
rect 12713 3479 12771 3485
rect 12989 3485 13001 3488
rect 13035 3485 13047 3519
rect 13354 3516 13360 3528
rect 13315 3488 13360 3516
rect 12989 3479 13047 3485
rect 12728 3448 12756 3479
rect 13354 3476 13360 3488
rect 13412 3476 13418 3528
rect 12406 3420 12756 3448
rect 9401 3383 9459 3389
rect 9401 3380 9413 3383
rect 9180 3352 9413 3380
rect 9180 3340 9186 3352
rect 9401 3349 9413 3352
rect 9447 3349 9459 3383
rect 9401 3343 9459 3349
rect 11701 3383 11759 3389
rect 11701 3349 11713 3383
rect 11747 3349 11759 3383
rect 11701 3343 11759 3349
rect 11790 3340 11796 3392
rect 11848 3380 11854 3392
rect 12621 3383 12679 3389
rect 12621 3380 12633 3383
rect 11848 3352 12633 3380
rect 11848 3340 11854 3352
rect 12621 3349 12633 3352
rect 12667 3349 12679 3383
rect 12621 3343 12679 3349
rect 1104 3290 13892 3312
rect 1104 3238 8214 3290
rect 8266 3238 8278 3290
rect 8330 3238 8342 3290
rect 8394 3238 8406 3290
rect 8458 3238 8470 3290
rect 8522 3238 13892 3290
rect 1104 3216 13892 3238
rect 2038 3176 2044 3188
rect 1780 3148 2044 3176
rect 1780 3117 1808 3148
rect 2038 3136 2044 3148
rect 2096 3136 2102 3188
rect 2225 3179 2283 3185
rect 2225 3145 2237 3179
rect 2271 3176 2283 3179
rect 2590 3176 2596 3188
rect 2271 3148 2596 3176
rect 2271 3145 2283 3148
rect 2225 3139 2283 3145
rect 2590 3136 2596 3148
rect 2648 3136 2654 3188
rect 3326 3136 3332 3188
rect 3384 3176 3390 3188
rect 4415 3179 4473 3185
rect 4415 3176 4427 3179
rect 3384 3148 4427 3176
rect 3384 3136 3390 3148
rect 4415 3145 4427 3148
rect 4461 3145 4473 3179
rect 5810 3176 5816 3188
rect 5771 3148 5816 3176
rect 4415 3139 4473 3145
rect 5810 3136 5816 3148
rect 5868 3136 5874 3188
rect 6733 3179 6791 3185
rect 6733 3145 6745 3179
rect 6779 3176 6791 3179
rect 6822 3176 6828 3188
rect 6779 3148 6828 3176
rect 6779 3145 6791 3148
rect 6733 3139 6791 3145
rect 6822 3136 6828 3148
rect 6880 3136 6886 3188
rect 7926 3176 7932 3188
rect 7887 3148 7932 3176
rect 7926 3136 7932 3148
rect 7984 3136 7990 3188
rect 8570 3176 8576 3188
rect 8036 3148 8576 3176
rect 1765 3111 1823 3117
rect 1765 3077 1777 3111
rect 1811 3077 1823 3111
rect 2774 3108 2780 3120
rect 1765 3071 1823 3077
rect 1964 3080 2780 3108
rect 1964 3049 1992 3080
rect 2774 3068 2780 3080
rect 2832 3068 2838 3120
rect 3418 3068 3424 3120
rect 3476 3068 3482 3120
rect 4893 3111 4951 3117
rect 4893 3108 4905 3111
rect 4172 3080 4905 3108
rect 1949 3043 2007 3049
rect 1949 3009 1961 3043
rect 1995 3009 2007 3043
rect 2314 3040 2320 3052
rect 2275 3012 2320 3040
rect 1949 3003 2007 3009
rect 2314 3000 2320 3012
rect 2372 3000 2378 3052
rect 1673 2975 1731 2981
rect 1673 2941 1685 2975
rect 1719 2941 1731 2975
rect 1673 2935 1731 2941
rect 1688 2836 1716 2935
rect 1762 2932 1768 2984
rect 1820 2972 1826 2984
rect 2406 2972 2412 2984
rect 1820 2944 2412 2972
rect 1820 2932 1826 2944
rect 2406 2932 2412 2944
rect 2464 2932 2470 2984
rect 2682 2972 2688 2984
rect 2643 2944 2688 2972
rect 2682 2932 2688 2944
rect 2740 2932 2746 2984
rect 3970 2932 3976 2984
rect 4028 2972 4034 2984
rect 4172 2981 4200 3080
rect 4893 3077 4905 3080
rect 4939 3077 4951 3111
rect 4893 3071 4951 3077
rect 5166 3068 5172 3120
rect 5224 3108 5230 3120
rect 6086 3108 6092 3120
rect 5224 3080 6092 3108
rect 5224 3068 5230 3080
rect 4706 3040 4712 3052
rect 4619 3012 4712 3040
rect 4706 3000 4712 3012
rect 4764 3040 4770 3052
rect 5442 3040 5448 3052
rect 4764 3012 5448 3040
rect 4764 3000 4770 3012
rect 5442 3000 5448 3012
rect 5500 3040 5506 3052
rect 5537 3043 5595 3049
rect 5537 3040 5549 3043
rect 5500 3012 5549 3040
rect 5500 3000 5506 3012
rect 5537 3009 5549 3012
rect 5583 3009 5595 3043
rect 5902 3040 5908 3052
rect 5863 3012 5908 3040
rect 5537 3003 5595 3009
rect 5902 3000 5908 3012
rect 5960 3000 5966 3052
rect 6012 3049 6040 3080
rect 6086 3068 6092 3080
rect 6144 3068 6150 3120
rect 6914 3108 6920 3120
rect 6875 3080 6920 3108
rect 6914 3068 6920 3080
rect 6972 3068 6978 3120
rect 7374 3068 7380 3120
rect 7432 3108 7438 3120
rect 8036 3108 8064 3148
rect 8570 3136 8576 3148
rect 8628 3136 8634 3188
rect 8754 3136 8760 3188
rect 8812 3176 8818 3188
rect 11054 3176 11060 3188
rect 8812 3148 11060 3176
rect 8812 3136 8818 3148
rect 11054 3136 11060 3148
rect 11112 3136 11118 3188
rect 11790 3176 11796 3188
rect 11164 3148 11796 3176
rect 7432 3080 8064 3108
rect 7432 3068 7438 3080
rect 5997 3043 6055 3049
rect 5997 3009 6009 3043
rect 6043 3009 6055 3043
rect 5997 3003 6055 3009
rect 6270 3000 6276 3052
rect 6328 3040 6334 3052
rect 6549 3043 6607 3049
rect 6549 3040 6561 3043
rect 6328 3012 6561 3040
rect 6328 3000 6334 3012
rect 6549 3009 6561 3012
rect 6595 3009 6607 3043
rect 7006 3040 7012 3052
rect 6967 3012 7012 3040
rect 6549 3003 6607 3009
rect 7006 3000 7012 3012
rect 7064 3000 7070 3052
rect 7190 3000 7196 3052
rect 7248 3040 7254 3052
rect 7576 3049 7604 3080
rect 7285 3043 7343 3049
rect 7285 3040 7297 3043
rect 7248 3012 7297 3040
rect 7248 3000 7254 3012
rect 7285 3009 7297 3012
rect 7331 3040 7343 3043
rect 7561 3043 7619 3049
rect 7331 3012 7512 3040
rect 7331 3009 7343 3012
rect 7285 3003 7343 3009
rect 4157 2975 4215 2981
rect 4157 2972 4169 2975
rect 4028 2944 4169 2972
rect 4028 2932 4034 2944
rect 4157 2941 4169 2944
rect 4203 2941 4215 2975
rect 4157 2935 4215 2941
rect 4614 2932 4620 2984
rect 4672 2972 4678 2984
rect 4985 2975 5043 2981
rect 4985 2972 4997 2975
rect 4672 2944 4997 2972
rect 4672 2932 4678 2944
rect 4985 2941 4997 2944
rect 5031 2972 5043 2975
rect 5074 2972 5080 2984
rect 5031 2944 5080 2972
rect 5031 2941 5043 2944
rect 4985 2935 5043 2941
rect 5074 2932 5080 2944
rect 5132 2932 5138 2984
rect 5353 2975 5411 2981
rect 5353 2941 5365 2975
rect 5399 2972 5411 2975
rect 5718 2972 5724 2984
rect 5399 2944 5724 2972
rect 5399 2941 5411 2944
rect 5353 2935 5411 2941
rect 5718 2932 5724 2944
rect 5776 2932 5782 2984
rect 6365 2975 6423 2981
rect 6365 2941 6377 2975
rect 6411 2972 6423 2975
rect 6730 2972 6736 2984
rect 6411 2944 6736 2972
rect 6411 2941 6423 2944
rect 6365 2935 6423 2941
rect 6089 2907 6147 2913
rect 6089 2904 6101 2907
rect 3896 2876 6101 2904
rect 3896 2836 3924 2876
rect 6089 2873 6101 2876
rect 6135 2873 6147 2907
rect 6089 2867 6147 2873
rect 1688 2808 3924 2836
rect 4154 2796 4160 2848
rect 4212 2836 4218 2848
rect 5166 2836 5172 2848
rect 4212 2808 5172 2836
rect 4212 2796 4218 2808
rect 5166 2796 5172 2808
rect 5224 2796 5230 2848
rect 5258 2796 5264 2848
rect 5316 2836 5322 2848
rect 6380 2836 6408 2935
rect 6730 2932 6736 2944
rect 6788 2932 6794 2984
rect 5316 2808 6408 2836
rect 7024 2836 7052 3000
rect 7374 2972 7380 2984
rect 7335 2944 7380 2972
rect 7374 2932 7380 2944
rect 7432 2932 7438 2984
rect 7484 2904 7512 3012
rect 7561 3009 7573 3043
rect 7607 3009 7619 3043
rect 7561 3003 7619 3009
rect 7653 3043 7711 3049
rect 7653 3009 7665 3043
rect 7699 3009 7711 3043
rect 7870 3040 7898 3080
rect 8110 3068 8116 3120
rect 8168 3108 8174 3120
rect 11164 3108 11192 3148
rect 11790 3136 11796 3148
rect 11848 3136 11854 3188
rect 11882 3136 11888 3188
rect 11940 3176 11946 3188
rect 12894 3176 12900 3188
rect 11940 3148 12900 3176
rect 11940 3136 11946 3148
rect 12894 3136 12900 3148
rect 12952 3136 12958 3188
rect 13170 3176 13176 3188
rect 13131 3148 13176 3176
rect 13170 3136 13176 3148
rect 13228 3136 13234 3188
rect 8168 3080 8248 3108
rect 10994 3080 11192 3108
rect 8168 3068 8174 3080
rect 8220 3049 8248 3080
rect 11238 3068 11244 3120
rect 11296 3108 11302 3120
rect 12069 3111 12127 3117
rect 12069 3108 12081 3111
rect 11296 3080 12081 3108
rect 11296 3068 11302 3080
rect 12069 3077 12081 3080
rect 12115 3077 12127 3111
rect 12069 3071 12127 3077
rect 12161 3111 12219 3117
rect 12161 3077 12173 3111
rect 12207 3077 12219 3111
rect 12161 3071 12219 3077
rect 7929 3043 7987 3049
rect 7929 3040 7941 3043
rect 7870 3012 7941 3040
rect 7653 3003 7711 3009
rect 7929 3009 7941 3012
rect 7975 3009 7987 3043
rect 7929 3003 7987 3009
rect 8205 3043 8263 3049
rect 8205 3009 8217 3043
rect 8251 3009 8263 3043
rect 9214 3040 9220 3052
rect 9175 3012 9220 3040
rect 8205 3003 8263 3009
rect 7668 2972 7696 3003
rect 8220 2972 8248 3003
rect 9214 3000 9220 3012
rect 9272 3000 9278 3052
rect 11054 3000 11060 3052
rect 11112 3040 11118 3052
rect 11609 3043 11667 3049
rect 11609 3040 11621 3043
rect 11112 3012 11621 3040
rect 11112 3000 11118 3012
rect 11609 3009 11621 3012
rect 11655 3009 11667 3043
rect 11882 3040 11888 3052
rect 11843 3012 11888 3040
rect 11609 3003 11667 3009
rect 7668 2944 8248 2972
rect 8294 2932 8300 2984
rect 8352 2972 8358 2984
rect 9490 2972 9496 2984
rect 8352 2944 9496 2972
rect 8352 2932 8358 2944
rect 8018 2904 8024 2916
rect 7484 2876 8024 2904
rect 8018 2864 8024 2876
rect 8076 2864 8082 2916
rect 9030 2904 9036 2916
rect 8128 2876 9036 2904
rect 8128 2836 8156 2876
rect 9030 2864 9036 2876
rect 9088 2864 9094 2916
rect 9214 2864 9220 2916
rect 9272 2904 9278 2916
rect 9324 2913 9352 2944
rect 9490 2932 9496 2944
rect 9548 2932 9554 2984
rect 9769 2975 9827 2981
rect 9769 2941 9781 2975
rect 9815 2972 9827 2975
rect 11514 2972 11520 2984
rect 9815 2944 11192 2972
rect 11475 2944 11520 2972
rect 9815 2941 9827 2944
rect 9769 2935 9827 2941
rect 9309 2907 9367 2913
rect 9309 2904 9321 2907
rect 9272 2876 9321 2904
rect 9272 2864 9278 2876
rect 9309 2873 9321 2876
rect 9355 2873 9367 2907
rect 9309 2867 9367 2873
rect 7024 2808 8156 2836
rect 5316 2796 5322 2808
rect 8202 2796 8208 2848
rect 8260 2836 8266 2848
rect 10502 2836 10508 2848
rect 8260 2808 10508 2836
rect 8260 2796 8266 2808
rect 10502 2796 10508 2808
rect 10560 2796 10566 2848
rect 11164 2836 11192 2944
rect 11514 2932 11520 2944
rect 11572 2932 11578 2984
rect 11624 2972 11652 3003
rect 11882 3000 11888 3012
rect 11940 3000 11946 3052
rect 12176 3040 12204 3071
rect 12805 3043 12863 3049
rect 12805 3040 12817 3043
rect 12084 3012 12204 3040
rect 12636 3012 12817 3040
rect 11974 2972 11980 2984
rect 11624 2944 11980 2972
rect 11974 2932 11980 2944
rect 12032 2932 12038 2984
rect 11241 2907 11299 2913
rect 11241 2873 11253 2907
rect 11287 2904 11299 2907
rect 11882 2904 11888 2916
rect 11287 2876 11888 2904
rect 11287 2873 11299 2876
rect 11241 2867 11299 2873
rect 11882 2864 11888 2876
rect 11940 2904 11946 2916
rect 12084 2904 12112 3012
rect 12158 2932 12164 2984
rect 12216 2972 12222 2984
rect 12216 2944 12261 2972
rect 12216 2932 12222 2944
rect 12636 2913 12664 3012
rect 12805 3009 12817 3012
rect 12851 3009 12863 3043
rect 12805 3003 12863 3009
rect 13262 3000 13268 3052
rect 13320 3040 13326 3052
rect 13357 3043 13415 3049
rect 13357 3040 13369 3043
rect 13320 3012 13369 3040
rect 13320 3000 13326 3012
rect 13357 3009 13369 3012
rect 13403 3009 13415 3043
rect 13357 3003 13415 3009
rect 11940 2876 12112 2904
rect 12621 2907 12679 2913
rect 11940 2864 11946 2876
rect 12621 2873 12633 2907
rect 12667 2873 12679 2907
rect 12621 2867 12679 2873
rect 12989 2839 13047 2845
rect 12989 2836 13001 2839
rect 11164 2808 13001 2836
rect 12989 2805 13001 2808
rect 13035 2805 13047 2839
rect 12989 2799 13047 2805
rect 1104 2746 13892 2768
rect 1104 2694 4214 2746
rect 4266 2694 4278 2746
rect 4330 2694 4342 2746
rect 4394 2694 4406 2746
rect 4458 2694 4470 2746
rect 4522 2694 12214 2746
rect 12266 2694 12278 2746
rect 12330 2694 12342 2746
rect 12394 2694 12406 2746
rect 12458 2694 12470 2746
rect 12522 2694 13892 2746
rect 1104 2672 13892 2694
rect 2130 2632 2136 2644
rect 2091 2604 2136 2632
rect 2130 2592 2136 2604
rect 2188 2592 2194 2644
rect 2222 2592 2228 2644
rect 2280 2632 2286 2644
rect 2685 2635 2743 2641
rect 2685 2632 2697 2635
rect 2280 2604 2697 2632
rect 2280 2592 2286 2604
rect 2685 2601 2697 2604
rect 2731 2601 2743 2635
rect 2685 2595 2743 2601
rect 3418 2592 3424 2644
rect 3476 2632 3482 2644
rect 3476 2604 3556 2632
rect 3476 2592 3482 2604
rect 2038 2524 2044 2576
rect 2096 2564 2102 2576
rect 3528 2573 3556 2604
rect 3602 2592 3608 2644
rect 3660 2632 3666 2644
rect 3881 2635 3939 2641
rect 3881 2632 3893 2635
rect 3660 2604 3893 2632
rect 3660 2592 3666 2604
rect 3881 2601 3893 2604
rect 3927 2601 3939 2635
rect 3881 2595 3939 2601
rect 4062 2592 4068 2644
rect 4120 2632 4126 2644
rect 7469 2635 7527 2641
rect 7469 2632 7481 2635
rect 4120 2604 7481 2632
rect 4120 2592 4126 2604
rect 7469 2601 7481 2604
rect 7515 2601 7527 2635
rect 7469 2595 7527 2601
rect 7742 2592 7748 2644
rect 7800 2632 7806 2644
rect 9122 2632 9128 2644
rect 7800 2604 9128 2632
rect 7800 2592 7806 2604
rect 9122 2592 9128 2604
rect 9180 2592 9186 2644
rect 10134 2632 10140 2644
rect 9232 2604 10140 2632
rect 3513 2567 3571 2573
rect 2096 2536 3372 2564
rect 2096 2524 2102 2536
rect 2314 2456 2320 2508
rect 2372 2456 2378 2508
rect 3344 2496 3372 2536
rect 3513 2533 3525 2567
rect 3559 2533 3571 2567
rect 3513 2527 3571 2533
rect 4356 2536 5856 2564
rect 3694 2496 3700 2508
rect 3344 2468 3700 2496
rect 1670 2428 1676 2440
rect 1631 2400 1676 2428
rect 1670 2388 1676 2400
rect 1728 2388 1734 2440
rect 1946 2428 1952 2440
rect 1907 2400 1952 2428
rect 1946 2388 1952 2400
rect 2004 2388 2010 2440
rect 2225 2431 2283 2437
rect 2225 2397 2237 2431
rect 2271 2428 2283 2431
rect 2332 2428 2360 2456
rect 2271 2400 2360 2428
rect 2409 2431 2467 2437
rect 2271 2397 2283 2400
rect 2225 2391 2283 2397
rect 2409 2397 2421 2431
rect 2455 2397 2467 2431
rect 2409 2391 2467 2397
rect 2424 2360 2452 2391
rect 2958 2388 2964 2440
rect 3016 2428 3022 2440
rect 3142 2428 3148 2440
rect 3016 2400 3061 2428
rect 3103 2400 3148 2428
rect 3016 2388 3022 2400
rect 3142 2388 3148 2400
rect 3200 2388 3206 2440
rect 3344 2437 3372 2468
rect 3694 2456 3700 2468
rect 3752 2456 3758 2508
rect 3329 2431 3387 2437
rect 3329 2397 3341 2431
rect 3375 2397 3387 2431
rect 3329 2391 3387 2397
rect 3421 2431 3479 2437
rect 3421 2397 3433 2431
rect 3467 2428 3479 2431
rect 4356 2428 4384 2536
rect 4433 2499 4491 2505
rect 4433 2465 4445 2499
rect 4479 2496 4491 2499
rect 5074 2496 5080 2508
rect 4479 2468 5080 2496
rect 4479 2465 4491 2468
rect 4433 2459 4491 2465
rect 5074 2456 5080 2468
rect 5132 2456 5138 2508
rect 5350 2456 5356 2508
rect 5408 2496 5414 2508
rect 5534 2496 5540 2508
rect 5408 2468 5540 2496
rect 5408 2456 5414 2468
rect 5534 2456 5540 2468
rect 5592 2496 5598 2508
rect 5721 2499 5779 2505
rect 5721 2496 5733 2499
rect 5592 2468 5733 2496
rect 5592 2456 5598 2468
rect 5721 2465 5733 2468
rect 5767 2465 5779 2499
rect 5828 2496 5856 2536
rect 7098 2524 7104 2576
rect 7156 2564 7162 2576
rect 9232 2564 9260 2604
rect 10134 2592 10140 2604
rect 10192 2592 10198 2644
rect 12618 2632 12624 2644
rect 12579 2604 12624 2632
rect 12618 2592 12624 2604
rect 12676 2592 12682 2644
rect 7156 2536 9260 2564
rect 7156 2524 7162 2536
rect 7282 2496 7288 2508
rect 5828 2468 7288 2496
rect 5721 2459 5779 2465
rect 7282 2456 7288 2468
rect 7340 2456 7346 2508
rect 7558 2456 7564 2508
rect 7616 2496 7622 2508
rect 7653 2499 7711 2505
rect 7653 2496 7665 2499
rect 7616 2468 7665 2496
rect 7616 2456 7622 2468
rect 7653 2465 7665 2468
rect 7699 2465 7711 2499
rect 8478 2496 8484 2508
rect 7653 2459 7711 2465
rect 7852 2468 8484 2496
rect 3467 2400 4384 2428
rect 4617 2431 4675 2437
rect 3467 2397 3479 2400
rect 3421 2391 3479 2397
rect 4617 2397 4629 2431
rect 4663 2428 4675 2431
rect 4890 2428 4896 2440
rect 4663 2400 4896 2428
rect 4663 2397 4675 2400
rect 4617 2391 4675 2397
rect 2593 2363 2651 2369
rect 2593 2360 2605 2363
rect 2424 2332 2605 2360
rect 2593 2329 2605 2332
rect 2639 2360 2651 2363
rect 2774 2360 2780 2372
rect 2639 2332 2780 2360
rect 2639 2329 2651 2332
rect 2593 2323 2651 2329
rect 2774 2320 2780 2332
rect 2832 2320 2838 2372
rect 3436 2360 3464 2391
rect 4890 2388 4896 2400
rect 4948 2388 4954 2440
rect 4985 2431 5043 2437
rect 4985 2397 4997 2431
rect 5031 2397 5043 2431
rect 5258 2428 5264 2440
rect 5219 2400 5264 2428
rect 4985 2391 5043 2397
rect 4154 2360 4160 2372
rect 3344 2332 3464 2360
rect 4067 2332 4160 2360
rect 1489 2295 1547 2301
rect 1489 2261 1501 2295
rect 1535 2292 1547 2295
rect 1670 2292 1676 2304
rect 1535 2264 1676 2292
rect 1535 2261 1547 2264
rect 1489 2255 1547 2261
rect 1670 2252 1676 2264
rect 1728 2252 1734 2304
rect 2130 2252 2136 2304
rect 2188 2292 2194 2304
rect 3344 2292 3372 2332
rect 4154 2320 4160 2332
rect 4212 2360 4218 2372
rect 5000 2360 5028 2391
rect 5258 2388 5264 2400
rect 5316 2388 5322 2440
rect 5626 2428 5632 2440
rect 5587 2400 5632 2428
rect 5626 2388 5632 2400
rect 5684 2388 5690 2440
rect 7466 2388 7472 2440
rect 7524 2428 7530 2440
rect 7852 2437 7880 2468
rect 8478 2456 8484 2468
rect 8536 2456 8542 2508
rect 10873 2499 10931 2505
rect 10873 2496 10885 2499
rect 8680 2468 10885 2496
rect 7837 2431 7895 2437
rect 7837 2428 7849 2431
rect 7524 2400 7849 2428
rect 7524 2388 7530 2400
rect 7837 2397 7849 2400
rect 7883 2397 7895 2431
rect 7837 2391 7895 2397
rect 7929 2431 7987 2437
rect 7929 2397 7941 2431
rect 7975 2428 7987 2431
rect 8018 2428 8024 2440
rect 7975 2400 8024 2428
rect 7975 2397 7987 2400
rect 7929 2391 7987 2397
rect 4212 2332 5028 2360
rect 4212 2320 4218 2332
rect 5000 2304 5028 2332
rect 5077 2363 5135 2369
rect 5077 2329 5089 2363
rect 5123 2360 5135 2363
rect 5997 2363 6055 2369
rect 5997 2360 6009 2363
rect 5123 2332 6009 2360
rect 5123 2329 5135 2332
rect 5077 2323 5135 2329
rect 5997 2329 6009 2332
rect 6043 2329 6055 2363
rect 7282 2360 7288 2372
rect 7222 2332 7288 2360
rect 5997 2323 6055 2329
rect 7282 2320 7288 2332
rect 7340 2320 7346 2372
rect 7650 2320 7656 2372
rect 7708 2360 7714 2372
rect 7944 2360 7972 2391
rect 8018 2388 8024 2400
rect 8076 2388 8082 2440
rect 8389 2431 8447 2437
rect 8389 2397 8401 2431
rect 8435 2428 8447 2431
rect 8570 2428 8576 2440
rect 8435 2400 8576 2428
rect 8435 2397 8447 2400
rect 8389 2391 8447 2397
rect 8570 2388 8576 2400
rect 8628 2388 8634 2440
rect 8680 2437 8708 2468
rect 10873 2465 10885 2468
rect 10919 2496 10931 2499
rect 10919 2468 11744 2496
rect 10919 2465 10931 2468
rect 10873 2459 10931 2465
rect 8665 2431 8723 2437
rect 8665 2397 8677 2431
rect 8711 2397 8723 2431
rect 9122 2428 9128 2440
rect 9083 2400 9128 2428
rect 8665 2391 8723 2397
rect 9122 2388 9128 2400
rect 9180 2388 9186 2440
rect 11422 2428 11428 2440
rect 11383 2400 11428 2428
rect 11422 2388 11428 2400
rect 11480 2388 11486 2440
rect 11606 2428 11612 2440
rect 11567 2400 11612 2428
rect 11606 2388 11612 2400
rect 11664 2388 11670 2440
rect 7708 2332 7972 2360
rect 8481 2363 8539 2369
rect 7708 2320 7714 2332
rect 8481 2329 8493 2363
rect 8527 2360 8539 2363
rect 9401 2363 9459 2369
rect 9401 2360 9413 2363
rect 8527 2332 9413 2360
rect 8527 2329 8539 2332
rect 8481 2323 8539 2329
rect 9401 2329 9413 2332
rect 9447 2329 9459 2363
rect 11514 2360 11520 2372
rect 10626 2332 11520 2360
rect 9401 2323 9459 2329
rect 11514 2320 11520 2332
rect 11572 2320 11578 2372
rect 11716 2360 11744 2468
rect 11882 2456 11888 2508
rect 11940 2496 11946 2508
rect 12805 2499 12863 2505
rect 12805 2496 12817 2499
rect 11940 2468 12817 2496
rect 11940 2456 11946 2468
rect 12805 2465 12817 2468
rect 12851 2465 12863 2499
rect 13354 2496 13360 2508
rect 13315 2468 13360 2496
rect 12805 2459 12863 2465
rect 13354 2456 13360 2468
rect 13412 2456 13418 2508
rect 12437 2431 12495 2437
rect 12437 2397 12449 2431
rect 12483 2428 12495 2431
rect 13170 2428 13176 2440
rect 12483 2400 13176 2428
rect 12483 2397 12495 2400
rect 12437 2391 12495 2397
rect 13170 2388 13176 2400
rect 13228 2428 13234 2440
rect 13265 2431 13323 2437
rect 13265 2428 13277 2431
rect 13228 2400 13277 2428
rect 13228 2388 13234 2400
rect 13265 2397 13277 2400
rect 13311 2397 13323 2431
rect 13265 2391 13323 2397
rect 12066 2360 12072 2372
rect 11716 2332 12072 2360
rect 12066 2320 12072 2332
rect 12124 2360 12130 2372
rect 12989 2363 13047 2369
rect 12989 2360 13001 2363
rect 12124 2332 13001 2360
rect 12124 2320 12130 2332
rect 12989 2329 13001 2332
rect 13035 2329 13047 2363
rect 12989 2323 13047 2329
rect 2188 2264 3372 2292
rect 4341 2295 4399 2301
rect 2188 2252 2194 2264
rect 4341 2261 4353 2295
rect 4387 2292 4399 2295
rect 4430 2292 4436 2304
rect 4387 2264 4436 2292
rect 4387 2261 4399 2264
rect 4341 2255 4399 2261
rect 4430 2252 4436 2264
rect 4488 2252 4494 2304
rect 4801 2295 4859 2301
rect 4801 2261 4813 2295
rect 4847 2292 4859 2295
rect 4890 2292 4896 2304
rect 4847 2264 4896 2292
rect 4847 2261 4859 2264
rect 4801 2255 4859 2261
rect 4890 2252 4896 2264
rect 4948 2252 4954 2304
rect 4982 2252 4988 2304
rect 5040 2292 5046 2304
rect 5718 2292 5724 2304
rect 5040 2264 5724 2292
rect 5040 2252 5046 2264
rect 5718 2252 5724 2264
rect 5776 2252 5782 2304
rect 9033 2295 9091 2301
rect 9033 2261 9045 2295
rect 9079 2292 9091 2295
rect 9674 2292 9680 2304
rect 9079 2264 9680 2292
rect 9079 2261 9091 2264
rect 9033 2255 9091 2261
rect 9674 2252 9680 2264
rect 9732 2252 9738 2304
rect 11974 2252 11980 2304
rect 12032 2292 12038 2304
rect 12897 2295 12955 2301
rect 12897 2292 12909 2295
rect 12032 2264 12909 2292
rect 12032 2252 12038 2264
rect 12897 2261 12909 2264
rect 12943 2261 12955 2295
rect 12897 2255 12955 2261
rect 1104 2202 13892 2224
rect 1104 2150 8214 2202
rect 8266 2150 8278 2202
rect 8330 2150 8342 2202
rect 8394 2150 8406 2202
rect 8458 2150 8470 2202
rect 8522 2150 13892 2202
rect 1104 2128 13892 2150
rect 2225 2091 2283 2097
rect 2225 2057 2237 2091
rect 2271 2057 2283 2091
rect 2225 2051 2283 2057
rect 4433 2091 4491 2097
rect 4433 2057 4445 2091
rect 4479 2088 4491 2091
rect 4614 2088 4620 2100
rect 4479 2060 4620 2088
rect 4479 2057 4491 2060
rect 4433 2051 4491 2057
rect 1489 2023 1547 2029
rect 1489 1989 1501 2023
rect 1535 2020 1547 2023
rect 1946 2020 1952 2032
rect 1535 1992 1952 2020
rect 1535 1989 1547 1992
rect 1489 1983 1547 1989
rect 1946 1980 1952 1992
rect 2004 1980 2010 2032
rect 2240 2020 2268 2051
rect 4614 2048 4620 2060
rect 4672 2048 4678 2100
rect 4890 2048 4896 2100
rect 4948 2088 4954 2100
rect 6638 2088 6644 2100
rect 4948 2060 6644 2088
rect 4948 2048 4954 2060
rect 6638 2048 6644 2060
rect 6696 2048 6702 2100
rect 7282 2088 7288 2100
rect 7243 2060 7288 2088
rect 7282 2048 7288 2060
rect 7340 2048 7346 2100
rect 7742 2088 7748 2100
rect 7703 2060 7748 2088
rect 7742 2048 7748 2060
rect 7800 2048 7806 2100
rect 9585 2091 9643 2097
rect 9585 2057 9597 2091
rect 9631 2088 9643 2091
rect 9674 2088 9680 2100
rect 9631 2060 9680 2088
rect 9631 2057 9643 2060
rect 9585 2051 9643 2057
rect 9674 2048 9680 2060
rect 9732 2088 9738 2100
rect 11606 2088 11612 2100
rect 9732 2060 11612 2088
rect 9732 2048 9738 2060
rect 11606 2048 11612 2060
rect 11664 2048 11670 2100
rect 2240 1992 3174 2020
rect 5442 1980 5448 2032
rect 5500 1980 5506 2032
rect 5626 1980 5632 2032
rect 5684 2020 5690 2032
rect 8110 2020 8116 2032
rect 5684 1992 8116 2020
rect 5684 1980 5690 1992
rect 1670 1952 1676 1964
rect 1631 1924 1676 1952
rect 1670 1912 1676 1924
rect 1728 1912 1734 1964
rect 1857 1955 1915 1961
rect 1857 1921 1869 1955
rect 1903 1921 1915 1955
rect 2130 1952 2136 1964
rect 2091 1924 2136 1952
rect 1857 1915 1915 1921
rect 1872 1748 1900 1915
rect 2130 1912 2136 1924
rect 2188 1912 2194 1964
rect 2225 1955 2283 1961
rect 2225 1921 2237 1955
rect 2271 1921 2283 1955
rect 2406 1952 2412 1964
rect 2367 1924 2412 1952
rect 2225 1915 2283 1921
rect 2038 1844 2044 1896
rect 2096 1884 2102 1896
rect 2240 1884 2268 1915
rect 2406 1912 2412 1924
rect 2464 1912 2470 1964
rect 6196 1961 6224 1992
rect 6181 1955 6239 1961
rect 6181 1921 6193 1955
rect 6227 1921 6239 1955
rect 6546 1952 6552 1964
rect 6507 1924 6552 1952
rect 6181 1915 6239 1921
rect 6546 1912 6552 1924
rect 6604 1912 6610 1964
rect 6638 1912 6644 1964
rect 6696 1952 6702 1964
rect 6840 1952 6960 1958
rect 7377 1955 7435 1961
rect 7377 1952 7389 1955
rect 6696 1930 7389 1952
rect 6696 1924 6868 1930
rect 6932 1924 7389 1930
rect 6696 1912 6702 1924
rect 7377 1921 7389 1924
rect 7423 1952 7435 1955
rect 7466 1952 7472 1964
rect 7423 1924 7472 1952
rect 7423 1921 7435 1924
rect 7377 1915 7435 1921
rect 7466 1912 7472 1924
rect 7524 1912 7530 1964
rect 7561 1955 7619 1961
rect 7561 1921 7573 1955
rect 7607 1952 7619 1955
rect 7650 1952 7656 1964
rect 7607 1924 7656 1952
rect 7607 1921 7619 1924
rect 7561 1915 7619 1921
rect 7650 1912 7656 1924
rect 7708 1912 7714 1964
rect 7852 1961 7880 1992
rect 8110 1980 8116 1992
rect 8168 1980 8174 2032
rect 9784 1992 9996 2020
rect 7837 1955 7895 1961
rect 7837 1921 7849 1955
rect 7883 1921 7895 1955
rect 7837 1915 7895 1921
rect 9214 1912 9220 1964
rect 9272 1912 9278 1964
rect 9784 1952 9812 1992
rect 9968 1961 9996 1992
rect 10134 1980 10140 2032
rect 10192 2020 10198 2032
rect 10321 2023 10379 2029
rect 10321 2020 10333 2023
rect 10192 1992 10333 2020
rect 10192 1980 10198 1992
rect 10321 1989 10333 1992
rect 10367 1989 10379 2023
rect 10321 1983 10379 1989
rect 10873 2023 10931 2029
rect 10873 1989 10885 2023
rect 10919 2020 10931 2023
rect 10919 1992 12282 2020
rect 10919 1989 10931 1992
rect 10873 1983 10931 1989
rect 9646 1924 9812 1952
rect 9861 1955 9919 1961
rect 2682 1884 2688 1896
rect 2096 1856 2268 1884
rect 2643 1856 2688 1884
rect 2096 1844 2102 1856
rect 2682 1844 2688 1856
rect 2740 1844 2746 1896
rect 5905 1887 5963 1893
rect 5905 1853 5917 1887
rect 5951 1884 5963 1887
rect 5951 1856 6408 1884
rect 5951 1853 5963 1856
rect 5905 1847 5963 1853
rect 6380 1816 6408 1856
rect 6454 1844 6460 1896
rect 6512 1884 6518 1896
rect 6512 1856 6557 1884
rect 6512 1844 6518 1856
rect 6730 1844 6736 1896
rect 6788 1884 6794 1896
rect 7101 1887 7159 1893
rect 7101 1884 7113 1887
rect 6788 1856 7113 1884
rect 6788 1844 6794 1856
rect 7101 1853 7113 1856
rect 7147 1853 7159 1887
rect 7101 1847 7159 1853
rect 6825 1819 6883 1825
rect 6825 1816 6837 1819
rect 6380 1788 6837 1816
rect 6825 1785 6837 1788
rect 6871 1785 6883 1819
rect 6825 1779 6883 1785
rect 4157 1751 4215 1757
rect 4157 1748 4169 1751
rect 1872 1720 4169 1748
rect 4157 1717 4169 1720
rect 4203 1748 4215 1751
rect 4430 1748 4436 1760
rect 4203 1720 4436 1748
rect 4203 1717 4215 1720
rect 4157 1711 4215 1717
rect 4430 1708 4436 1720
rect 4488 1748 4494 1760
rect 4614 1748 4620 1760
rect 4488 1720 4620 1748
rect 4488 1708 4494 1720
rect 4614 1708 4620 1720
rect 4672 1708 4678 1760
rect 7116 1748 7144 1847
rect 7190 1844 7196 1896
rect 7248 1884 7254 1896
rect 8113 1887 8171 1893
rect 8113 1884 8125 1887
rect 7248 1856 8125 1884
rect 7248 1844 7254 1856
rect 8113 1853 8125 1856
rect 8159 1853 8171 1887
rect 8113 1847 8171 1853
rect 8662 1844 8668 1896
rect 8720 1884 8726 1896
rect 9646 1884 9674 1924
rect 9861 1921 9873 1955
rect 9907 1921 9919 1955
rect 9861 1915 9919 1921
rect 9953 1955 10011 1961
rect 9953 1921 9965 1955
rect 9999 1921 10011 1955
rect 10226 1952 10232 1964
rect 10187 1924 10232 1952
rect 9953 1915 10011 1921
rect 8720 1856 9674 1884
rect 8720 1844 8726 1856
rect 9306 1776 9312 1828
rect 9364 1816 9370 1828
rect 9876 1816 9904 1915
rect 10226 1912 10232 1924
rect 10284 1912 10290 1964
rect 10502 1952 10508 1964
rect 10463 1924 10508 1952
rect 10502 1912 10508 1924
rect 10560 1912 10566 1964
rect 10781 1955 10839 1961
rect 10781 1921 10793 1955
rect 10827 1952 10839 1955
rect 11054 1952 11060 1964
rect 10827 1924 11060 1952
rect 10827 1921 10839 1924
rect 10781 1915 10839 1921
rect 11054 1912 11060 1924
rect 11112 1912 11118 1964
rect 11238 1952 11244 1964
rect 11199 1924 11244 1952
rect 11238 1912 11244 1924
rect 11296 1912 11302 1964
rect 11514 1952 11520 1964
rect 11475 1924 11520 1952
rect 11514 1912 11520 1924
rect 11572 1912 11578 1964
rect 11793 1887 11851 1893
rect 11793 1853 11805 1887
rect 11839 1884 11851 1887
rect 12986 1884 12992 1896
rect 11839 1856 12992 1884
rect 11839 1853 11851 1856
rect 11793 1847 11851 1853
rect 12986 1844 12992 1856
rect 13044 1844 13050 1896
rect 9364 1788 9904 1816
rect 10045 1819 10103 1825
rect 9364 1776 9370 1788
rect 10045 1785 10057 1819
rect 10091 1816 10103 1819
rect 10134 1816 10140 1828
rect 10091 1788 10140 1816
rect 10091 1785 10103 1788
rect 10045 1779 10103 1785
rect 10134 1776 10140 1788
rect 10192 1776 10198 1828
rect 11057 1819 11115 1825
rect 11057 1785 11069 1819
rect 11103 1785 11115 1819
rect 11057 1779 11115 1785
rect 8570 1748 8576 1760
rect 7116 1720 8576 1748
rect 8570 1708 8576 1720
rect 8628 1748 8634 1760
rect 11072 1748 11100 1779
rect 8628 1720 11100 1748
rect 8628 1708 8634 1720
rect 11974 1708 11980 1760
rect 12032 1748 12038 1760
rect 13265 1751 13323 1757
rect 13265 1748 13277 1751
rect 12032 1720 13277 1748
rect 12032 1708 12038 1720
rect 13265 1717 13277 1720
rect 13311 1717 13323 1751
rect 13265 1711 13323 1717
rect 1104 1658 13892 1680
rect 1104 1606 4214 1658
rect 4266 1606 4278 1658
rect 4330 1606 4342 1658
rect 4394 1606 4406 1658
rect 4458 1606 4470 1658
rect 4522 1606 12214 1658
rect 12266 1606 12278 1658
rect 12330 1606 12342 1658
rect 12394 1606 12406 1658
rect 12458 1606 12470 1658
rect 12522 1606 13892 1658
rect 1104 1584 13892 1606
rect 3142 1504 3148 1556
rect 3200 1544 3206 1556
rect 3881 1547 3939 1553
rect 3881 1544 3893 1547
rect 3200 1516 3893 1544
rect 3200 1504 3206 1516
rect 3881 1513 3893 1516
rect 3927 1513 3939 1547
rect 3881 1507 3939 1513
rect 3970 1504 3976 1556
rect 4028 1544 4034 1556
rect 6917 1547 6975 1553
rect 4028 1516 4844 1544
rect 4028 1504 4034 1516
rect 3510 1476 3516 1488
rect 3471 1448 3516 1476
rect 3510 1436 3516 1448
rect 3568 1436 3574 1488
rect 4816 1476 4844 1516
rect 5184 1516 6592 1544
rect 5184 1476 5212 1516
rect 4816 1448 5212 1476
rect 6564 1476 6592 1516
rect 6917 1513 6929 1547
rect 6963 1544 6975 1547
rect 7190 1544 7196 1556
rect 6963 1516 7196 1544
rect 6963 1513 6975 1516
rect 6917 1507 6975 1513
rect 7190 1504 7196 1516
rect 7248 1504 7254 1556
rect 7742 1544 7748 1556
rect 7300 1516 7748 1544
rect 7300 1476 7328 1516
rect 7742 1504 7748 1516
rect 7800 1504 7806 1556
rect 9766 1544 9772 1556
rect 8588 1516 9772 1544
rect 6564 1448 7328 1476
rect 1394 1408 1400 1420
rect 1355 1380 1400 1408
rect 1394 1368 1400 1380
rect 1452 1368 1458 1420
rect 2774 1368 2780 1420
rect 2832 1408 2838 1420
rect 3970 1408 3976 1420
rect 2832 1380 3976 1408
rect 2832 1368 2838 1380
rect 3970 1368 3976 1380
rect 4028 1368 4034 1420
rect 4982 1408 4988 1420
rect 4943 1380 4988 1408
rect 4982 1368 4988 1380
rect 5040 1368 5046 1420
rect 5537 1411 5595 1417
rect 5537 1377 5549 1411
rect 5583 1408 5595 1411
rect 6454 1408 6460 1420
rect 5583 1380 6460 1408
rect 5583 1377 5595 1380
rect 5537 1371 5595 1377
rect 6454 1368 6460 1380
rect 6512 1368 6518 1420
rect 7650 1408 7656 1420
rect 7208 1380 7656 1408
rect 2406 1300 2412 1352
rect 2464 1340 2470 1352
rect 3145 1343 3203 1349
rect 3145 1340 3157 1343
rect 2464 1312 3157 1340
rect 2464 1300 2470 1312
rect 3145 1309 3157 1312
rect 3191 1309 3203 1343
rect 3418 1340 3424 1352
rect 3379 1312 3424 1340
rect 3145 1303 3203 1309
rect 3418 1300 3424 1312
rect 3476 1300 3482 1352
rect 3602 1340 3608 1352
rect 3563 1312 3608 1340
rect 3602 1300 3608 1312
rect 3660 1300 3666 1352
rect 4065 1343 4123 1349
rect 4065 1309 4077 1343
rect 4111 1309 4123 1343
rect 4065 1303 4123 1309
rect 4080 1272 4108 1303
rect 4154 1300 4160 1352
rect 4212 1340 4218 1352
rect 4706 1340 4712 1352
rect 4212 1312 4257 1340
rect 4667 1312 4712 1340
rect 4212 1300 4218 1312
rect 4706 1300 4712 1312
rect 4764 1300 4770 1352
rect 5721 1343 5779 1349
rect 5721 1340 5733 1343
rect 4816 1312 5733 1340
rect 4614 1272 4620 1284
rect 4080 1244 4620 1272
rect 4614 1232 4620 1244
rect 4672 1272 4678 1284
rect 4816 1272 4844 1312
rect 5721 1309 5733 1312
rect 5767 1309 5779 1343
rect 5721 1303 5779 1309
rect 5810 1300 5816 1352
rect 5868 1340 5874 1352
rect 5905 1343 5963 1349
rect 5905 1340 5917 1343
rect 5868 1312 5917 1340
rect 5868 1300 5874 1312
rect 5905 1309 5917 1312
rect 5951 1309 5963 1343
rect 5905 1303 5963 1309
rect 6549 1343 6607 1349
rect 6549 1309 6561 1343
rect 6595 1340 6607 1343
rect 6638 1340 6644 1352
rect 6595 1312 6644 1340
rect 6595 1309 6607 1312
rect 6549 1303 6607 1309
rect 6638 1300 6644 1312
rect 6696 1300 6702 1352
rect 6733 1343 6791 1349
rect 6733 1309 6745 1343
rect 6779 1340 6791 1343
rect 7208 1340 7236 1380
rect 7650 1368 7656 1380
rect 7708 1368 7714 1420
rect 8389 1411 8447 1417
rect 8389 1377 8401 1411
rect 8435 1408 8447 1411
rect 8588 1408 8616 1516
rect 9766 1504 9772 1516
rect 9824 1544 9830 1556
rect 10962 1544 10968 1556
rect 9824 1516 10968 1544
rect 9824 1504 9830 1516
rect 10962 1504 10968 1516
rect 11020 1504 11026 1556
rect 11149 1547 11207 1553
rect 11149 1513 11161 1547
rect 11195 1544 11207 1547
rect 11422 1544 11428 1556
rect 11195 1516 11428 1544
rect 11195 1513 11207 1516
rect 11149 1507 11207 1513
rect 11422 1504 11428 1516
rect 11480 1504 11486 1556
rect 12986 1544 12992 1556
rect 12947 1516 12992 1544
rect 12986 1504 12992 1516
rect 13044 1504 13050 1556
rect 11882 1436 11888 1488
rect 11940 1476 11946 1488
rect 11940 1448 12204 1476
rect 11940 1436 11946 1448
rect 8435 1380 8616 1408
rect 8665 1411 8723 1417
rect 8435 1377 8447 1380
rect 8389 1371 8447 1377
rect 8665 1377 8677 1411
rect 8711 1408 8723 1411
rect 9401 1411 9459 1417
rect 9401 1408 9413 1411
rect 8711 1380 9413 1408
rect 8711 1377 8723 1380
rect 8665 1371 8723 1377
rect 9401 1377 9413 1380
rect 9447 1377 9459 1411
rect 9674 1408 9680 1420
rect 9635 1380 9680 1408
rect 9401 1371 9459 1377
rect 6779 1312 7236 1340
rect 6779 1309 6791 1312
rect 6733 1303 6791 1309
rect 4672 1244 4844 1272
rect 4672 1232 4678 1244
rect 5442 1232 5448 1284
rect 5500 1272 5506 1284
rect 6365 1275 6423 1281
rect 6365 1272 6377 1275
rect 5500 1244 6377 1272
rect 5500 1232 5506 1244
rect 6365 1241 6377 1244
rect 6411 1241 6423 1275
rect 6365 1235 6423 1241
rect 7374 1232 7380 1284
rect 7432 1232 7438 1284
rect 8110 1232 8116 1284
rect 8168 1272 8174 1284
rect 8680 1272 8708 1371
rect 9674 1368 9680 1380
rect 9732 1368 9738 1420
rect 11238 1368 11244 1420
rect 11296 1408 11302 1420
rect 12176 1417 12204 1448
rect 12069 1411 12127 1417
rect 12069 1408 12081 1411
rect 11296 1380 12081 1408
rect 11296 1368 11302 1380
rect 12069 1377 12081 1380
rect 12115 1377 12127 1411
rect 12069 1371 12127 1377
rect 12161 1411 12219 1417
rect 12161 1377 12173 1411
rect 12207 1377 12219 1411
rect 12161 1371 12219 1377
rect 8754 1300 8760 1352
rect 8812 1340 8818 1352
rect 9033 1343 9091 1349
rect 9033 1340 9045 1343
rect 8812 1312 9045 1340
rect 8812 1300 8818 1312
rect 9033 1309 9045 1312
rect 9079 1309 9091 1343
rect 9306 1340 9312 1352
rect 9267 1312 9312 1340
rect 9033 1303 9091 1309
rect 9306 1300 9312 1312
rect 9364 1300 9370 1352
rect 8168 1244 8708 1272
rect 8168 1232 8174 1244
rect 10134 1232 10140 1284
rect 10192 1232 10198 1284
rect 12084 1272 12112 1371
rect 12639 1343 12697 1349
rect 12639 1309 12651 1343
rect 12685 1340 12697 1343
rect 12805 1343 12863 1349
rect 12805 1340 12817 1343
rect 12685 1312 12817 1340
rect 12685 1309 12697 1312
rect 12639 1303 12697 1309
rect 12805 1309 12817 1312
rect 12851 1309 12863 1343
rect 13170 1340 13176 1352
rect 13131 1312 13176 1340
rect 12805 1303 12863 1309
rect 13170 1300 13176 1312
rect 13228 1300 13234 1352
rect 12084 1244 13400 1272
rect 5902 1204 5908 1216
rect 5863 1176 5908 1204
rect 5902 1164 5908 1176
rect 5960 1164 5966 1216
rect 6086 1204 6092 1216
rect 6047 1176 6092 1204
rect 6086 1164 6092 1176
rect 6144 1164 6150 1216
rect 9214 1204 9220 1216
rect 9175 1176 9220 1204
rect 9214 1164 9220 1176
rect 9272 1164 9278 1216
rect 11514 1204 11520 1216
rect 11475 1176 11520 1204
rect 11514 1164 11520 1176
rect 11572 1164 11578 1216
rect 11974 1164 11980 1216
rect 12032 1204 12038 1216
rect 13372 1213 13400 1244
rect 12161 1207 12219 1213
rect 12161 1204 12173 1207
rect 12032 1176 12173 1204
rect 12032 1164 12038 1176
rect 12161 1173 12173 1176
rect 12207 1173 12219 1207
rect 12161 1167 12219 1173
rect 13357 1207 13415 1213
rect 13357 1173 13369 1207
rect 13403 1173 13415 1207
rect 13357 1167 13415 1173
rect 1104 1114 13892 1136
rect 1104 1062 8214 1114
rect 8266 1062 8278 1114
rect 8330 1062 8342 1114
rect 8394 1062 8406 1114
rect 8458 1062 8470 1114
rect 8522 1062 13892 1114
rect 1104 1040 13892 1062
rect 2958 960 2964 1012
rect 3016 1000 3022 1012
rect 5902 1000 5908 1012
rect 3016 972 5908 1000
rect 3016 960 3022 972
rect 5902 960 5908 972
rect 5960 1000 5966 1012
rect 10226 1000 10232 1012
rect 5960 972 10232 1000
rect 5960 960 5966 972
rect 10226 960 10232 972
rect 10284 960 10290 1012
rect 3418 892 3424 944
rect 3476 932 3482 944
rect 11514 932 11520 944
rect 3476 904 11520 932
rect 3476 892 3482 904
rect 11514 892 11520 904
rect 11572 892 11578 944
rect 3602 824 3608 876
rect 3660 864 3666 876
rect 6086 864 6092 876
rect 3660 836 6092 864
rect 3660 824 3666 836
rect 6086 824 6092 836
rect 6144 824 6150 876
<< via1 >>
rect 3608 14288 3660 14340
rect 10784 14288 10836 14340
rect 7840 14084 7892 14136
rect 9772 14084 9824 14136
rect 2872 14016 2924 14068
rect 6644 14016 6696 14068
rect 6460 13948 6512 14000
rect 10416 13948 10468 14000
rect 3424 13880 3476 13932
rect 7932 13880 7984 13932
rect 5356 13812 5408 13864
rect 11704 13812 11756 13864
rect 5540 13744 5592 13796
rect 9680 13744 9732 13796
rect 11244 13744 11296 13796
rect 6092 13676 6144 13728
rect 8024 13676 8076 13728
rect 8576 13676 8628 13728
rect 9956 13676 10008 13728
rect 10968 13676 11020 13728
rect 4214 13574 4266 13626
rect 4278 13574 4330 13626
rect 4342 13574 4394 13626
rect 4406 13574 4458 13626
rect 4470 13574 4522 13626
rect 12214 13574 12266 13626
rect 12278 13574 12330 13626
rect 12342 13574 12394 13626
rect 12406 13574 12458 13626
rect 12470 13574 12522 13626
rect 3608 13515 3660 13524
rect 3608 13481 3617 13515
rect 3617 13481 3651 13515
rect 3651 13481 3660 13515
rect 3608 13472 3660 13481
rect 6092 13472 6144 13524
rect 5540 13447 5592 13456
rect 5540 13413 5549 13447
rect 5549 13413 5583 13447
rect 5583 13413 5592 13447
rect 5540 13404 5592 13413
rect 1676 13311 1728 13320
rect 1676 13277 1685 13311
rect 1685 13277 1719 13311
rect 1719 13277 1728 13311
rect 1676 13268 1728 13277
rect 1860 13268 1912 13320
rect 2872 13311 2924 13320
rect 2872 13277 2881 13311
rect 2881 13277 2915 13311
rect 2915 13277 2924 13311
rect 2872 13268 2924 13277
rect 3424 13311 3476 13320
rect 3424 13277 3433 13311
rect 3433 13277 3467 13311
rect 3467 13277 3476 13311
rect 3424 13268 3476 13277
rect 1492 13243 1544 13252
rect 1492 13209 1501 13243
rect 1501 13209 1535 13243
rect 1535 13209 1544 13243
rect 1492 13200 1544 13209
rect 1952 13243 2004 13252
rect 1952 13209 1961 13243
rect 1961 13209 1995 13243
rect 1995 13209 2004 13243
rect 1952 13200 2004 13209
rect 3148 13200 3200 13252
rect 3332 13243 3384 13252
rect 3332 13209 3341 13243
rect 3341 13209 3375 13243
rect 3375 13209 3384 13243
rect 3332 13200 3384 13209
rect 5356 13336 5408 13388
rect 10048 13472 10100 13524
rect 10968 13472 11020 13524
rect 6460 13379 6512 13388
rect 6460 13345 6469 13379
rect 6469 13345 6503 13379
rect 6503 13345 6512 13379
rect 6460 13336 6512 13345
rect 7656 13404 7708 13456
rect 3700 13268 3752 13320
rect 5632 13311 5684 13320
rect 5632 13277 5641 13311
rect 5641 13277 5675 13311
rect 5675 13277 5684 13311
rect 5632 13268 5684 13277
rect 7104 13268 7156 13320
rect 7656 13268 7708 13320
rect 8024 13311 8076 13320
rect 8024 13277 8073 13311
rect 8073 13277 8076 13311
rect 8300 13311 8352 13320
rect 8024 13268 8076 13277
rect 8300 13277 8309 13311
rect 8309 13277 8343 13311
rect 8343 13277 8352 13311
rect 8300 13268 8352 13277
rect 2044 13132 2096 13184
rect 3056 13132 3108 13184
rect 3516 13132 3568 13184
rect 4068 13243 4120 13252
rect 4068 13209 4077 13243
rect 4077 13209 4111 13243
rect 4111 13209 4120 13243
rect 4068 13200 4120 13209
rect 4896 13243 4948 13252
rect 4896 13209 4905 13243
rect 4905 13209 4939 13243
rect 4939 13209 4948 13243
rect 4896 13200 4948 13209
rect 5264 13200 5316 13252
rect 5816 13200 5868 13252
rect 8208 13243 8260 13252
rect 4620 13132 4672 13184
rect 5080 13175 5132 13184
rect 5080 13141 5089 13175
rect 5089 13141 5123 13175
rect 5123 13141 5132 13175
rect 7288 13175 7340 13184
rect 5080 13132 5132 13141
rect 7288 13141 7297 13175
rect 7297 13141 7331 13175
rect 7331 13141 7340 13175
rect 7288 13132 7340 13141
rect 7656 13132 7708 13184
rect 8208 13209 8217 13243
rect 8217 13209 8251 13243
rect 8251 13209 8260 13243
rect 8208 13200 8260 13209
rect 9864 13336 9916 13388
rect 11980 13404 12032 13456
rect 8484 13311 8536 13320
rect 8484 13277 8493 13311
rect 8493 13277 8527 13311
rect 8527 13277 8536 13311
rect 8484 13268 8536 13277
rect 8760 13268 8812 13320
rect 10692 13311 10744 13320
rect 10692 13277 10701 13311
rect 10701 13277 10735 13311
rect 10735 13277 10744 13311
rect 10692 13268 10744 13277
rect 10968 13311 11020 13320
rect 10968 13277 10977 13311
rect 10977 13277 11011 13311
rect 11011 13277 11020 13311
rect 10968 13268 11020 13277
rect 11244 13311 11296 13320
rect 11244 13277 11253 13311
rect 11253 13277 11287 13311
rect 11287 13277 11296 13311
rect 11244 13268 11296 13277
rect 11520 13268 11572 13320
rect 11704 13268 11756 13320
rect 9772 13243 9824 13252
rect 9772 13209 9781 13243
rect 9781 13209 9815 13243
rect 9815 13209 9824 13243
rect 9772 13200 9824 13209
rect 10140 13200 10192 13252
rect 10232 13200 10284 13252
rect 12072 13243 12124 13252
rect 9220 13175 9272 13184
rect 9220 13141 9229 13175
rect 9229 13141 9263 13175
rect 9263 13141 9272 13175
rect 9220 13132 9272 13141
rect 12072 13209 12081 13243
rect 12081 13209 12115 13243
rect 12115 13209 12124 13243
rect 12072 13200 12124 13209
rect 11888 13132 11940 13184
rect 13452 13268 13504 13320
rect 13268 13200 13320 13252
rect 13084 13175 13136 13184
rect 13084 13141 13093 13175
rect 13093 13141 13127 13175
rect 13127 13141 13136 13175
rect 13084 13132 13136 13141
rect 13360 13175 13412 13184
rect 13360 13141 13369 13175
rect 13369 13141 13403 13175
rect 13403 13141 13412 13175
rect 13360 13132 13412 13141
rect 8214 13030 8266 13082
rect 8278 13030 8330 13082
rect 8342 13030 8394 13082
rect 8406 13030 8458 13082
rect 8470 13030 8522 13082
rect 1768 12928 1820 12980
rect 2964 12928 3016 12980
rect 3056 12928 3108 12980
rect 3884 12928 3936 12980
rect 4988 12928 5040 12980
rect 7472 12928 7524 12980
rect 9220 12928 9272 12980
rect 11612 12928 11664 12980
rect 3516 12860 3568 12912
rect 5356 12860 5408 12912
rect 5632 12903 5684 12912
rect 5632 12869 5641 12903
rect 5641 12869 5675 12903
rect 5675 12869 5684 12903
rect 5632 12860 5684 12869
rect 7104 12903 7156 12912
rect 7104 12869 7113 12903
rect 7113 12869 7147 12903
rect 7147 12869 7156 12903
rect 7104 12860 7156 12869
rect 7288 12903 7340 12912
rect 7288 12869 7297 12903
rect 7297 12869 7331 12903
rect 7331 12869 7340 12903
rect 7288 12860 7340 12869
rect 1676 12792 1728 12844
rect 1860 12835 1912 12844
rect 1860 12801 1869 12835
rect 1869 12801 1903 12835
rect 1903 12801 1912 12835
rect 1860 12792 1912 12801
rect 3700 12835 3752 12844
rect 1768 12767 1820 12776
rect 1768 12733 1777 12767
rect 1777 12733 1811 12767
rect 1811 12733 1820 12767
rect 3700 12801 3709 12835
rect 3709 12801 3743 12835
rect 3743 12801 3752 12835
rect 3700 12792 3752 12801
rect 4068 12792 4120 12844
rect 1768 12724 1820 12733
rect 3792 12724 3844 12776
rect 5908 12792 5960 12844
rect 6092 12835 6144 12844
rect 6092 12801 6101 12835
rect 6101 12801 6135 12835
rect 6135 12801 6144 12835
rect 6092 12792 6144 12801
rect 6460 12792 6512 12844
rect 6552 12724 6604 12776
rect 7012 12724 7064 12776
rect 8944 12860 8996 12912
rect 10232 12860 10284 12912
rect 11244 12860 11296 12912
rect 12072 12860 12124 12912
rect 7656 12792 7708 12844
rect 3976 12656 4028 12708
rect 8392 12835 8444 12844
rect 8392 12801 8401 12835
rect 8401 12801 8435 12835
rect 8435 12801 8444 12835
rect 8392 12792 8444 12801
rect 8576 12792 8628 12844
rect 8760 12835 8812 12844
rect 8760 12801 8769 12835
rect 8769 12801 8803 12835
rect 8803 12801 8812 12835
rect 8760 12792 8812 12801
rect 9680 12835 9732 12844
rect 9680 12801 9689 12835
rect 9689 12801 9723 12835
rect 9723 12801 9732 12835
rect 9680 12792 9732 12801
rect 9864 12792 9916 12844
rect 11520 12835 11572 12844
rect 11520 12801 11529 12835
rect 11529 12801 11563 12835
rect 11563 12801 11572 12835
rect 11520 12792 11572 12801
rect 11888 12792 11940 12844
rect 8576 12656 8628 12708
rect 9772 12656 9824 12708
rect 14372 12656 14424 12708
rect 2964 12588 3016 12640
rect 7104 12588 7156 12640
rect 7196 12588 7248 12640
rect 8300 12588 8352 12640
rect 9588 12588 9640 12640
rect 13268 12631 13320 12640
rect 13268 12597 13277 12631
rect 13277 12597 13311 12631
rect 13311 12597 13320 12631
rect 13268 12588 13320 12597
rect 4214 12486 4266 12538
rect 4278 12486 4330 12538
rect 4342 12486 4394 12538
rect 4406 12486 4458 12538
rect 4470 12486 4522 12538
rect 12214 12486 12266 12538
rect 12278 12486 12330 12538
rect 12342 12486 12394 12538
rect 12406 12486 12458 12538
rect 12470 12486 12522 12538
rect 1768 12223 1820 12232
rect 1768 12189 1777 12223
rect 1777 12189 1811 12223
rect 1811 12189 1820 12223
rect 1768 12180 1820 12189
rect 3332 12384 3384 12436
rect 4160 12384 4212 12436
rect 5356 12384 5408 12436
rect 5908 12384 5960 12436
rect 6000 12384 6052 12436
rect 7012 12384 7064 12436
rect 9864 12427 9916 12436
rect 3608 12316 3660 12368
rect 5172 12359 5224 12368
rect 5172 12325 5181 12359
rect 5181 12325 5215 12359
rect 5215 12325 5224 12359
rect 5172 12316 5224 12325
rect 5816 12316 5868 12368
rect 7288 12316 7340 12368
rect 7380 12316 7432 12368
rect 7472 12316 7524 12368
rect 8208 12316 8260 12368
rect 8852 12316 8904 12368
rect 9036 12316 9088 12368
rect 9864 12393 9873 12427
rect 9873 12393 9907 12427
rect 9907 12393 9916 12427
rect 9864 12384 9916 12393
rect 10140 12427 10192 12436
rect 10140 12393 10149 12427
rect 10149 12393 10183 12427
rect 10183 12393 10192 12427
rect 10140 12384 10192 12393
rect 10416 12427 10468 12436
rect 10416 12393 10425 12427
rect 10425 12393 10459 12427
rect 10459 12393 10468 12427
rect 10416 12384 10468 12393
rect 11520 12316 11572 12368
rect 2688 12223 2740 12232
rect 2688 12189 2697 12223
rect 2697 12189 2731 12223
rect 2731 12189 2740 12223
rect 2688 12180 2740 12189
rect 3056 12248 3108 12300
rect 6184 12248 6236 12300
rect 4804 12180 4856 12232
rect 2320 12112 2372 12164
rect 2504 12044 2556 12096
rect 2780 12044 2832 12096
rect 3332 12112 3384 12164
rect 3792 12155 3844 12164
rect 3792 12121 3801 12155
rect 3801 12121 3835 12155
rect 3835 12121 3844 12155
rect 3792 12112 3844 12121
rect 4068 12155 4120 12164
rect 4068 12121 4077 12155
rect 4077 12121 4111 12155
rect 4111 12121 4120 12155
rect 4068 12112 4120 12121
rect 4528 12112 4580 12164
rect 5632 12180 5684 12232
rect 7104 12180 7156 12232
rect 7472 12223 7524 12232
rect 7472 12189 7481 12223
rect 7481 12189 7515 12223
rect 7515 12189 7524 12223
rect 7472 12180 7524 12189
rect 7932 12180 7984 12232
rect 8484 12248 8536 12300
rect 5172 12112 5224 12164
rect 7012 12112 7064 12164
rect 6552 12044 6604 12096
rect 7656 12112 7708 12164
rect 8208 12199 8218 12232
rect 8218 12199 8252 12232
rect 8252 12199 8260 12232
rect 8208 12180 8260 12199
rect 8668 12180 8720 12232
rect 8852 12180 8904 12232
rect 9128 12248 9180 12300
rect 9404 12180 9456 12232
rect 10048 12248 10100 12300
rect 10140 12248 10192 12300
rect 13176 12248 13228 12300
rect 9956 12180 10008 12232
rect 10232 12223 10284 12232
rect 10232 12189 10241 12223
rect 10241 12189 10275 12223
rect 10275 12189 10284 12223
rect 10232 12180 10284 12189
rect 10600 12223 10652 12232
rect 10600 12189 10609 12223
rect 10609 12189 10643 12223
rect 10643 12189 10652 12223
rect 10600 12180 10652 12189
rect 10784 12180 10836 12232
rect 11520 12180 11572 12232
rect 11612 12223 11664 12232
rect 11612 12189 11621 12223
rect 11621 12189 11655 12223
rect 11655 12189 11664 12223
rect 11888 12223 11940 12232
rect 11612 12180 11664 12189
rect 11888 12189 11897 12223
rect 11897 12189 11931 12223
rect 11931 12189 11940 12223
rect 11888 12180 11940 12189
rect 13268 12223 13320 12232
rect 7748 12044 7800 12096
rect 8852 12044 8904 12096
rect 9128 12087 9180 12096
rect 9128 12053 9137 12087
rect 9137 12053 9171 12087
rect 9171 12053 9180 12087
rect 9128 12044 9180 12053
rect 9588 12155 9640 12164
rect 9588 12121 9597 12155
rect 9597 12121 9631 12155
rect 9631 12121 9640 12155
rect 9588 12112 9640 12121
rect 10048 12112 10100 12164
rect 10508 12044 10560 12096
rect 11336 12112 11388 12164
rect 13268 12189 13277 12223
rect 13277 12189 13311 12223
rect 13311 12189 13320 12223
rect 13268 12180 13320 12189
rect 11888 12044 11940 12096
rect 8214 11942 8266 11994
rect 8278 11942 8330 11994
rect 8342 11942 8394 11994
rect 8406 11942 8458 11994
rect 8470 11942 8522 11994
rect 848 11840 900 11892
rect 1860 11772 1912 11824
rect 2596 11840 2648 11892
rect 4160 11840 4212 11892
rect 3700 11815 3752 11824
rect 1492 11704 1544 11756
rect 2412 11704 2464 11756
rect 3700 11781 3709 11815
rect 3709 11781 3743 11815
rect 3743 11781 3752 11815
rect 3700 11772 3752 11781
rect 5264 11840 5316 11892
rect 6552 11840 6604 11892
rect 7380 11840 7432 11892
rect 7472 11840 7524 11892
rect 7840 11883 7892 11892
rect 7840 11849 7849 11883
rect 7849 11849 7883 11883
rect 7883 11849 7892 11883
rect 7840 11840 7892 11849
rect 8852 11840 8904 11892
rect 9128 11840 9180 11892
rect 5080 11772 5132 11824
rect 5172 11772 5224 11824
rect 1584 11568 1636 11620
rect 1768 11568 1820 11620
rect 1676 11500 1728 11552
rect 2964 11543 3016 11552
rect 2964 11509 2973 11543
rect 2973 11509 3007 11543
rect 3007 11509 3016 11543
rect 2964 11500 3016 11509
rect 3424 11704 3476 11756
rect 3976 11636 4028 11688
rect 4712 11636 4764 11688
rect 4988 11636 5040 11688
rect 5540 11704 5592 11756
rect 6460 11704 6512 11756
rect 6828 11747 6880 11756
rect 6000 11636 6052 11688
rect 4620 11611 4672 11620
rect 3240 11500 3292 11552
rect 3792 11500 3844 11552
rect 4620 11577 4629 11611
rect 4629 11577 4663 11611
rect 4663 11577 4672 11611
rect 4620 11568 4672 11577
rect 5816 11568 5868 11620
rect 6092 11611 6144 11620
rect 6092 11577 6101 11611
rect 6101 11577 6135 11611
rect 6135 11577 6144 11611
rect 6092 11568 6144 11577
rect 5356 11500 5408 11552
rect 6828 11713 6837 11747
rect 6837 11713 6871 11747
rect 6871 11713 6880 11747
rect 6828 11704 6880 11713
rect 7104 11704 7156 11756
rect 7932 11772 7984 11824
rect 10140 11815 10192 11824
rect 10140 11781 10149 11815
rect 10149 11781 10183 11815
rect 10183 11781 10192 11815
rect 10140 11772 10192 11781
rect 10232 11815 10284 11824
rect 10232 11781 10241 11815
rect 10241 11781 10275 11815
rect 10275 11781 10284 11815
rect 10232 11772 10284 11781
rect 10416 11815 10468 11824
rect 10416 11781 10425 11815
rect 10425 11781 10459 11815
rect 10459 11781 10468 11815
rect 10416 11772 10468 11781
rect 11428 11772 11480 11824
rect 8576 11747 8628 11756
rect 6920 11679 6972 11688
rect 6920 11645 6929 11679
rect 6929 11645 6963 11679
rect 6963 11645 6972 11679
rect 6920 11636 6972 11645
rect 8576 11713 8585 11747
rect 8585 11713 8619 11747
rect 8619 11713 8628 11747
rect 8576 11704 8628 11713
rect 8852 11747 8904 11756
rect 8852 11713 8861 11747
rect 8861 11713 8895 11747
rect 8895 11713 8904 11747
rect 9036 11747 9088 11756
rect 8852 11704 8904 11713
rect 9036 11713 9045 11747
rect 9045 11713 9079 11747
rect 9079 11713 9088 11747
rect 9036 11704 9088 11713
rect 9128 11747 9180 11756
rect 9128 11713 9137 11747
rect 9137 11713 9171 11747
rect 9171 11713 9180 11747
rect 9312 11747 9364 11756
rect 9128 11704 9180 11713
rect 9312 11713 9315 11747
rect 9315 11713 9364 11747
rect 9312 11704 9364 11713
rect 9404 11704 9456 11756
rect 10048 11747 10100 11756
rect 10048 11713 10057 11747
rect 10057 11713 10091 11747
rect 10091 11713 10100 11747
rect 10048 11704 10100 11713
rect 7932 11636 7984 11688
rect 8484 11679 8536 11688
rect 7104 11568 7156 11620
rect 8484 11645 8493 11679
rect 8493 11645 8527 11679
rect 8527 11645 8536 11679
rect 8484 11636 8536 11645
rect 11060 11704 11112 11756
rect 11520 11747 11572 11756
rect 11520 11713 11529 11747
rect 11529 11713 11563 11747
rect 11563 11713 11572 11747
rect 11520 11704 11572 11713
rect 11980 11772 12032 11824
rect 13084 11815 13136 11824
rect 13084 11781 13093 11815
rect 13093 11781 13127 11815
rect 13127 11781 13136 11815
rect 13084 11772 13136 11781
rect 13452 11815 13504 11824
rect 13452 11781 13461 11815
rect 13461 11781 13495 11815
rect 13495 11781 13504 11815
rect 13452 11772 13504 11781
rect 11336 11679 11388 11688
rect 8300 11568 8352 11620
rect 7012 11500 7064 11552
rect 7288 11500 7340 11552
rect 7748 11500 7800 11552
rect 7840 11500 7892 11552
rect 9128 11568 9180 11620
rect 9588 11568 9640 11620
rect 11336 11645 11345 11679
rect 11345 11645 11379 11679
rect 11379 11645 11388 11679
rect 11336 11636 11388 11645
rect 11612 11636 11664 11688
rect 12624 11636 12676 11688
rect 10692 11568 10744 11620
rect 12992 11611 13044 11620
rect 12992 11577 13001 11611
rect 13001 11577 13035 11611
rect 13035 11577 13044 11611
rect 12992 11568 13044 11577
rect 10508 11500 10560 11552
rect 10600 11543 10652 11552
rect 10600 11509 10609 11543
rect 10609 11509 10643 11543
rect 10643 11509 10652 11543
rect 10600 11500 10652 11509
rect 10876 11500 10928 11552
rect 12716 11500 12768 11552
rect 4214 11398 4266 11450
rect 4278 11398 4330 11450
rect 4342 11398 4394 11450
rect 4406 11398 4458 11450
rect 4470 11398 4522 11450
rect 12214 11398 12266 11450
rect 12278 11398 12330 11450
rect 12342 11398 12394 11450
rect 12406 11398 12458 11450
rect 12470 11398 12522 11450
rect 1768 11228 1820 11280
rect 3608 11296 3660 11348
rect 4804 11296 4856 11348
rect 6460 11296 6512 11348
rect 5080 11228 5132 11280
rect 5264 11271 5316 11280
rect 5264 11237 5273 11271
rect 5273 11237 5307 11271
rect 5307 11237 5316 11271
rect 5264 11228 5316 11237
rect 6092 11271 6144 11280
rect 6092 11237 6101 11271
rect 6101 11237 6135 11271
rect 6135 11237 6144 11271
rect 6092 11228 6144 11237
rect 3608 11203 3660 11212
rect 3608 11169 3617 11203
rect 3617 11169 3651 11203
rect 3651 11169 3660 11203
rect 3608 11160 3660 11169
rect 6276 11160 6328 11212
rect 1492 11092 1544 11144
rect 2320 11135 2372 11144
rect 2320 11101 2329 11135
rect 2329 11101 2363 11135
rect 2363 11101 2372 11135
rect 2320 11092 2372 11101
rect 3976 11135 4028 11144
rect 3976 11101 3985 11135
rect 3985 11101 4019 11135
rect 4019 11101 4028 11135
rect 3976 11092 4028 11101
rect 3240 11024 3292 11076
rect 3516 11024 3568 11076
rect 5172 11092 5224 11144
rect 5356 11135 5408 11144
rect 5356 11101 5365 11135
rect 5365 11101 5399 11135
rect 5399 11101 5408 11135
rect 5356 11092 5408 11101
rect 4160 11024 4212 11076
rect 6000 11092 6052 11144
rect 6644 11228 6696 11280
rect 8852 11296 8904 11348
rect 9036 11296 9088 11348
rect 7104 11160 7156 11212
rect 7472 11228 7524 11280
rect 8208 11228 8260 11280
rect 8576 11228 8628 11280
rect 10416 11296 10468 11348
rect 10600 11296 10652 11348
rect 11520 11296 11572 11348
rect 10968 11228 11020 11280
rect 11060 11228 11112 11280
rect 7288 11203 7340 11212
rect 7288 11169 7297 11203
rect 7297 11169 7331 11203
rect 7331 11169 7340 11203
rect 7288 11160 7340 11169
rect 6828 11092 6880 11144
rect 7196 11024 7248 11076
rect 1492 10956 1544 11008
rect 2044 10956 2096 11008
rect 2596 10956 2648 11008
rect 4252 10956 4304 11008
rect 5448 10956 5500 11008
rect 5632 10956 5684 11008
rect 6460 10956 6512 11008
rect 6736 10956 6788 11008
rect 7012 10956 7064 11008
rect 7840 11024 7892 11076
rect 8116 11092 8168 11144
rect 8484 11160 8536 11212
rect 9036 11160 9088 11212
rect 8576 11135 8628 11144
rect 8576 11101 8585 11135
rect 8585 11101 8619 11135
rect 8619 11101 8628 11135
rect 8576 11092 8628 11101
rect 9772 11160 9824 11212
rect 9220 11092 9272 11144
rect 9496 11135 9548 11144
rect 9496 11101 9505 11135
rect 9505 11101 9539 11135
rect 9539 11101 9548 11135
rect 9496 11092 9548 11101
rect 8668 11024 8720 11076
rect 8392 10956 8444 11008
rect 8944 11024 8996 11076
rect 9864 11092 9916 11144
rect 10232 11135 10284 11144
rect 10232 11101 10241 11135
rect 10241 11101 10275 11135
rect 10275 11101 10284 11135
rect 10232 11092 10284 11101
rect 10692 11092 10744 11144
rect 11060 11135 11112 11144
rect 11060 11101 11069 11135
rect 11069 11101 11103 11135
rect 11103 11101 11112 11135
rect 11060 11092 11112 11101
rect 11428 11092 11480 11144
rect 11612 11135 11664 11144
rect 11612 11101 11621 11135
rect 11621 11101 11655 11135
rect 11655 11101 11664 11135
rect 11612 11092 11664 11101
rect 12624 11092 12676 11144
rect 13084 11092 13136 11144
rect 13268 11135 13320 11144
rect 13268 11101 13277 11135
rect 13277 11101 13311 11135
rect 13311 11101 13320 11135
rect 13268 11092 13320 11101
rect 9036 10956 9088 11008
rect 9220 10956 9272 11008
rect 11704 11024 11756 11076
rect 12992 11067 13044 11076
rect 12992 11033 13001 11067
rect 13001 11033 13035 11067
rect 13035 11033 13044 11067
rect 12992 11024 13044 11033
rect 13544 11067 13596 11076
rect 13544 11033 13553 11067
rect 13553 11033 13587 11067
rect 13587 11033 13596 11067
rect 13544 11024 13596 11033
rect 11980 10956 12032 11008
rect 13176 10956 13228 11008
rect 8214 10854 8266 10906
rect 8278 10854 8330 10906
rect 8342 10854 8394 10906
rect 8406 10854 8458 10906
rect 8470 10854 8522 10906
rect 1492 10795 1544 10804
rect 1492 10761 1501 10795
rect 1501 10761 1535 10795
rect 1535 10761 1544 10795
rect 1492 10752 1544 10761
rect 1492 10616 1544 10668
rect 2320 10684 2372 10736
rect 3976 10684 4028 10736
rect 4252 10727 4304 10736
rect 4252 10693 4261 10727
rect 4261 10693 4295 10727
rect 4295 10693 4304 10727
rect 4252 10684 4304 10693
rect 4620 10684 4672 10736
rect 6276 10684 6328 10736
rect 6644 10752 6696 10804
rect 7012 10752 7064 10804
rect 7656 10752 7708 10804
rect 2504 10659 2556 10668
rect 2504 10625 2513 10659
rect 2513 10625 2547 10659
rect 2547 10625 2556 10659
rect 2504 10616 2556 10625
rect 3240 10616 3292 10668
rect 3608 10659 3660 10668
rect 3608 10625 3617 10659
rect 3617 10625 3651 10659
rect 3651 10625 3660 10659
rect 3608 10616 3660 10625
rect 4160 10616 4212 10668
rect 4344 10659 4396 10668
rect 4344 10625 4353 10659
rect 4353 10625 4387 10659
rect 4387 10625 4396 10659
rect 4344 10616 4396 10625
rect 4988 10616 5040 10668
rect 5356 10659 5408 10668
rect 5356 10625 5365 10659
rect 5365 10625 5399 10659
rect 5399 10625 5408 10659
rect 5356 10616 5408 10625
rect 5448 10616 5500 10668
rect 6736 10616 6788 10668
rect 7104 10659 7156 10668
rect 7104 10625 7113 10659
rect 7113 10625 7147 10659
rect 7147 10625 7156 10659
rect 7104 10616 7156 10625
rect 7288 10659 7340 10668
rect 7288 10625 7297 10659
rect 7297 10625 7331 10659
rect 7331 10625 7340 10659
rect 7288 10616 7340 10625
rect 7472 10659 7524 10668
rect 7472 10625 7481 10659
rect 7481 10625 7515 10659
rect 7515 10625 7524 10659
rect 7472 10616 7524 10625
rect 2044 10591 2096 10600
rect 2044 10557 2053 10591
rect 2053 10557 2087 10591
rect 2087 10557 2096 10591
rect 2044 10548 2096 10557
rect 2596 10591 2648 10600
rect 2596 10557 2605 10591
rect 2605 10557 2639 10591
rect 2639 10557 2648 10591
rect 2596 10548 2648 10557
rect 6092 10548 6144 10600
rect 3700 10480 3752 10532
rect 5816 10480 5868 10532
rect 6368 10480 6420 10532
rect 6552 10548 6604 10600
rect 7932 10752 7984 10804
rect 7840 10684 7892 10736
rect 8576 10752 8628 10804
rect 8116 10659 8168 10668
rect 8116 10625 8126 10659
rect 8126 10625 8160 10659
rect 8160 10625 8168 10659
rect 8116 10616 8168 10625
rect 3976 10412 4028 10464
rect 4344 10412 4396 10464
rect 5264 10412 5316 10464
rect 6184 10412 6236 10464
rect 6552 10412 6604 10464
rect 6736 10480 6788 10532
rect 7840 10548 7892 10600
rect 8300 10659 8352 10668
rect 8300 10625 8310 10659
rect 8310 10625 8344 10659
rect 8344 10625 8352 10659
rect 8944 10684 8996 10736
rect 8300 10616 8352 10625
rect 8668 10659 8720 10668
rect 8668 10625 8677 10659
rect 8677 10625 8711 10659
rect 8711 10625 8720 10659
rect 8852 10659 8904 10668
rect 8668 10616 8720 10625
rect 8852 10625 8861 10659
rect 8861 10625 8895 10659
rect 8895 10625 8904 10659
rect 8852 10616 8904 10625
rect 9036 10659 9088 10668
rect 9036 10625 9045 10659
rect 9045 10625 9079 10659
rect 9079 10625 9088 10659
rect 9036 10616 9088 10625
rect 8392 10548 8444 10600
rect 7380 10480 7432 10532
rect 8116 10480 8168 10532
rect 9680 10684 9732 10736
rect 10232 10727 10284 10736
rect 10232 10693 10241 10727
rect 10241 10693 10275 10727
rect 10275 10693 10284 10727
rect 10232 10684 10284 10693
rect 9772 10616 9824 10668
rect 10508 10659 10560 10668
rect 9680 10548 9732 10600
rect 10508 10625 10517 10659
rect 10517 10625 10551 10659
rect 10551 10625 10560 10659
rect 10508 10616 10560 10625
rect 10600 10659 10652 10668
rect 10600 10625 10609 10659
rect 10609 10625 10643 10659
rect 10643 10625 10652 10659
rect 11060 10684 11112 10736
rect 11244 10795 11296 10804
rect 11244 10761 11253 10795
rect 11253 10761 11287 10795
rect 11287 10761 11296 10795
rect 11244 10752 11296 10761
rect 12440 10752 12492 10804
rect 12164 10727 12216 10736
rect 12164 10693 12173 10727
rect 12173 10693 12207 10727
rect 12207 10693 12216 10727
rect 13084 10727 13136 10736
rect 12164 10684 12216 10693
rect 13084 10693 13093 10727
rect 13093 10693 13127 10727
rect 13127 10693 13136 10727
rect 13084 10684 13136 10693
rect 10600 10616 10652 10625
rect 10692 10548 10744 10600
rect 11244 10616 11296 10668
rect 9128 10480 9180 10532
rect 11060 10548 11112 10600
rect 11796 10616 11848 10668
rect 12256 10659 12308 10668
rect 12256 10625 12265 10659
rect 12265 10625 12299 10659
rect 12299 10625 12308 10659
rect 12900 10659 12952 10668
rect 12256 10616 12308 10625
rect 12900 10625 12909 10659
rect 12909 10625 12943 10659
rect 12943 10625 12952 10659
rect 12900 10616 12952 10625
rect 12992 10616 13044 10668
rect 13728 10616 13780 10668
rect 11888 10480 11940 10532
rect 12072 10480 12124 10532
rect 13636 10548 13688 10600
rect 9772 10455 9824 10464
rect 9772 10421 9781 10455
rect 9781 10421 9815 10455
rect 9815 10421 9824 10455
rect 10232 10455 10284 10464
rect 9772 10412 9824 10421
rect 10232 10421 10241 10455
rect 10241 10421 10275 10455
rect 10275 10421 10284 10455
rect 10232 10412 10284 10421
rect 10968 10412 11020 10464
rect 4214 10310 4266 10362
rect 4278 10310 4330 10362
rect 4342 10310 4394 10362
rect 4406 10310 4458 10362
rect 4470 10310 4522 10362
rect 12214 10310 12266 10362
rect 12278 10310 12330 10362
rect 12342 10310 12394 10362
rect 12406 10310 12458 10362
rect 12470 10310 12522 10362
rect 2596 10208 2648 10260
rect 4712 10208 4764 10260
rect 4804 10208 4856 10260
rect 4988 10208 5040 10260
rect 6552 10208 6604 10260
rect 8300 10208 8352 10260
rect 8576 10208 8628 10260
rect 8760 10208 8812 10260
rect 2504 10140 2556 10192
rect 5540 10140 5592 10192
rect 5724 10140 5776 10192
rect 6092 10140 6144 10192
rect 6736 10140 6788 10192
rect 6920 10140 6972 10192
rect 7472 10140 7524 10192
rect 2964 10072 3016 10124
rect 3700 10072 3752 10124
rect 1676 10047 1728 10056
rect 1676 10013 1685 10047
rect 1685 10013 1719 10047
rect 1719 10013 1728 10047
rect 1676 10004 1728 10013
rect 2044 10047 2096 10056
rect 2044 10013 2053 10047
rect 2053 10013 2087 10047
rect 2087 10013 2096 10047
rect 2044 10004 2096 10013
rect 3056 10047 3108 10056
rect 3056 10013 3065 10047
rect 3065 10013 3099 10047
rect 3099 10013 3108 10047
rect 3056 10004 3108 10013
rect 5356 10072 5408 10124
rect 5816 10072 5868 10124
rect 3884 10004 3936 10056
rect 4528 10047 4580 10056
rect 4528 10013 4537 10047
rect 4537 10013 4571 10047
rect 4571 10013 4580 10047
rect 4528 10004 4580 10013
rect 4804 10047 4856 10056
rect 4804 10013 4813 10047
rect 4813 10013 4847 10047
rect 4847 10013 4856 10047
rect 4804 10004 4856 10013
rect 5632 10004 5684 10056
rect 6092 10004 6144 10056
rect 3148 9936 3200 9988
rect 5080 9936 5132 9988
rect 5540 9936 5592 9988
rect 6276 9979 6328 9988
rect 6276 9945 6285 9979
rect 6285 9945 6319 9979
rect 6319 9945 6328 9979
rect 6736 10013 6751 10034
rect 6751 10013 6785 10034
rect 6785 10013 6788 10034
rect 6736 9982 6788 10013
rect 6276 9936 6328 9945
rect 4712 9868 4764 9920
rect 5632 9911 5684 9920
rect 5632 9877 5641 9911
rect 5641 9877 5675 9911
rect 5675 9877 5684 9911
rect 5632 9868 5684 9877
rect 6552 9868 6604 9920
rect 6736 9868 6788 9920
rect 7012 10072 7064 10124
rect 7196 10072 7248 10124
rect 7012 9936 7064 9988
rect 8392 10140 8444 10192
rect 9220 10140 9272 10192
rect 8300 10072 8352 10124
rect 8768 10004 8820 10056
rect 8944 10072 8996 10124
rect 9588 10140 9640 10192
rect 10324 10208 10376 10260
rect 11888 10251 11940 10260
rect 9864 10140 9916 10192
rect 9588 10047 9640 10056
rect 9588 10013 9597 10047
rect 9597 10013 9631 10047
rect 9631 10013 9640 10047
rect 9588 10004 9640 10013
rect 6920 9868 6972 9920
rect 7288 9868 7340 9920
rect 7932 9868 7984 9920
rect 8484 9911 8536 9920
rect 8484 9877 8493 9911
rect 8493 9877 8527 9911
rect 8527 9877 8536 9911
rect 8484 9868 8536 9877
rect 9220 9868 9272 9920
rect 9956 10072 10008 10124
rect 10048 10047 10100 10056
rect 10048 10013 10057 10047
rect 10057 10013 10091 10047
rect 10091 10013 10100 10047
rect 10048 10004 10100 10013
rect 10416 10004 10468 10056
rect 10600 10140 10652 10192
rect 11520 10140 11572 10192
rect 10692 10072 10744 10124
rect 11888 10217 11897 10251
rect 11897 10217 11931 10251
rect 11931 10217 11940 10251
rect 11888 10208 11940 10217
rect 12072 10208 12124 10260
rect 13176 10140 13228 10192
rect 13360 10115 13412 10124
rect 10968 10047 11020 10056
rect 10968 10013 10977 10047
rect 10977 10013 11011 10047
rect 11011 10013 11020 10047
rect 10968 10004 11020 10013
rect 12072 10047 12124 10056
rect 10508 9868 10560 9920
rect 11428 9936 11480 9988
rect 12072 10013 12081 10047
rect 12081 10013 12115 10047
rect 12115 10013 12124 10047
rect 12072 10004 12124 10013
rect 12440 10047 12492 10056
rect 12440 10013 12449 10047
rect 12449 10013 12483 10047
rect 12483 10013 12492 10047
rect 12440 10004 12492 10013
rect 13360 10081 13369 10115
rect 13369 10081 13403 10115
rect 13403 10081 13412 10115
rect 13360 10072 13412 10081
rect 12808 10047 12860 10056
rect 12808 10013 12817 10047
rect 12817 10013 12851 10047
rect 12851 10013 12860 10047
rect 12808 10004 12860 10013
rect 11796 9936 11848 9988
rect 11244 9868 11296 9920
rect 8214 9766 8266 9818
rect 8278 9766 8330 9818
rect 8342 9766 8394 9818
rect 8406 9766 8458 9818
rect 8470 9766 8522 9818
rect 6276 9664 6328 9716
rect 1860 9571 1912 9580
rect 1860 9537 1869 9571
rect 1869 9537 1903 9571
rect 1903 9537 1912 9571
rect 1860 9528 1912 9537
rect 3056 9596 3108 9648
rect 3700 9596 3752 9648
rect 7196 9707 7248 9716
rect 7196 9673 7205 9707
rect 7205 9673 7239 9707
rect 7239 9673 7248 9707
rect 7196 9664 7248 9673
rect 7472 9664 7524 9716
rect 3148 9571 3200 9580
rect 3148 9537 3157 9571
rect 3157 9537 3191 9571
rect 3191 9537 3200 9571
rect 3148 9528 3200 9537
rect 3608 9528 3660 9580
rect 3700 9460 3752 9512
rect 4804 9528 4856 9580
rect 5908 9571 5960 9580
rect 5908 9537 5917 9571
rect 5917 9537 5951 9571
rect 5951 9537 5960 9571
rect 5908 9528 5960 9537
rect 6460 9528 6512 9580
rect 5724 9435 5776 9444
rect 5724 9401 5733 9435
rect 5733 9401 5767 9435
rect 5767 9401 5776 9435
rect 5724 9392 5776 9401
rect 8208 9664 8260 9716
rect 7012 9571 7064 9580
rect 7012 9537 7021 9571
rect 7021 9537 7055 9571
rect 7055 9537 7064 9571
rect 8208 9571 8260 9580
rect 7012 9528 7064 9537
rect 8208 9537 8217 9571
rect 8217 9537 8251 9571
rect 8251 9537 8260 9571
rect 8208 9528 8260 9537
rect 8392 9528 8444 9580
rect 8576 9571 8628 9580
rect 8576 9537 8585 9571
rect 8585 9537 8619 9571
rect 8619 9537 8628 9571
rect 9128 9596 9180 9648
rect 10324 9664 10376 9716
rect 9404 9639 9456 9648
rect 9404 9605 9413 9639
rect 9413 9605 9447 9639
rect 9447 9605 9456 9639
rect 9404 9596 9456 9605
rect 8576 9528 8628 9537
rect 7012 9392 7064 9444
rect 1400 9324 1452 9376
rect 3516 9324 3568 9376
rect 3884 9367 3936 9376
rect 3884 9333 3893 9367
rect 3893 9333 3927 9367
rect 3927 9333 3936 9367
rect 3884 9324 3936 9333
rect 4528 9324 4580 9376
rect 4988 9324 5040 9376
rect 7104 9324 7156 9376
rect 7288 9460 7340 9512
rect 8760 9503 8812 9512
rect 8760 9469 8769 9503
rect 8769 9469 8803 9503
rect 8803 9469 8812 9503
rect 8760 9460 8812 9469
rect 9588 9528 9640 9580
rect 10692 9596 10744 9648
rect 10968 9664 11020 9716
rect 13176 9639 13228 9648
rect 9864 9571 9916 9580
rect 9864 9537 9873 9571
rect 9873 9537 9907 9571
rect 9907 9537 9916 9571
rect 9864 9528 9916 9537
rect 9404 9460 9456 9512
rect 10324 9571 10376 9580
rect 10324 9537 10333 9571
rect 10333 9537 10367 9571
rect 10367 9537 10376 9571
rect 10324 9528 10376 9537
rect 10600 9571 10652 9580
rect 10600 9537 10609 9571
rect 10609 9537 10643 9571
rect 10643 9537 10652 9571
rect 10600 9528 10652 9537
rect 7840 9392 7892 9444
rect 9496 9392 9548 9444
rect 10140 9392 10192 9444
rect 10416 9392 10468 9444
rect 11428 9528 11480 9580
rect 7656 9324 7708 9376
rect 9036 9324 9088 9376
rect 10692 9367 10744 9376
rect 10692 9333 10701 9367
rect 10701 9333 10735 9367
rect 10735 9333 10744 9367
rect 10692 9324 10744 9333
rect 10968 9392 11020 9444
rect 11888 9528 11940 9580
rect 13176 9605 13185 9639
rect 13185 9605 13219 9639
rect 13219 9605 13228 9639
rect 13176 9596 13228 9605
rect 13268 9596 13320 9648
rect 13452 9596 13504 9648
rect 12808 9528 12860 9580
rect 11980 9324 12032 9376
rect 12440 9324 12492 9376
rect 13452 9367 13504 9376
rect 13452 9333 13461 9367
rect 13461 9333 13495 9367
rect 13495 9333 13504 9367
rect 13452 9324 13504 9333
rect 4214 9222 4266 9274
rect 4278 9222 4330 9274
rect 4342 9222 4394 9274
rect 4406 9222 4458 9274
rect 4470 9222 4522 9274
rect 12214 9222 12266 9274
rect 12278 9222 12330 9274
rect 12342 9222 12394 9274
rect 12406 9222 12458 9274
rect 12470 9222 12522 9274
rect 5816 9120 5868 9172
rect 6828 9120 6880 9172
rect 7012 9120 7064 9172
rect 7380 9120 7432 9172
rect 7656 9120 7708 9172
rect 4804 9052 4856 9104
rect 3792 8984 3844 9036
rect 4712 9027 4764 9036
rect 4712 8993 4721 9027
rect 4721 8993 4755 9027
rect 4755 8993 4764 9027
rect 4712 8984 4764 8993
rect 7104 9027 7156 9036
rect 1400 8959 1452 8968
rect 1400 8925 1409 8959
rect 1409 8925 1443 8959
rect 1443 8925 1452 8959
rect 1400 8916 1452 8925
rect 2964 8916 3016 8968
rect 3884 8959 3936 8968
rect 3884 8925 3893 8959
rect 3893 8925 3927 8959
rect 3927 8925 3936 8959
rect 3884 8916 3936 8925
rect 5540 8916 5592 8968
rect 5632 8916 5684 8968
rect 5908 8916 5960 8968
rect 6276 8916 6328 8968
rect 4988 8848 5040 8900
rect 5448 8848 5500 8900
rect 7104 8993 7113 9027
rect 7113 8993 7147 9027
rect 7147 8993 7156 9027
rect 7104 8984 7156 8993
rect 8944 9120 8996 9172
rect 9864 9120 9916 9172
rect 10140 9120 10192 9172
rect 10232 9120 10284 9172
rect 11612 9120 11664 9172
rect 11888 9120 11940 9172
rect 12164 9120 12216 9172
rect 6736 8916 6788 8968
rect 7196 8848 7248 8900
rect 7380 8848 7432 8900
rect 7840 8916 7892 8968
rect 8392 8984 8444 9036
rect 9404 9052 9456 9104
rect 9680 9052 9732 9104
rect 8852 8916 8904 8968
rect 8944 8959 8996 8968
rect 8944 8925 8953 8959
rect 8953 8925 8987 8959
rect 8987 8925 8996 8959
rect 8944 8916 8996 8925
rect 9128 8959 9180 8968
rect 9128 8925 9137 8959
rect 9137 8925 9171 8959
rect 9171 8925 9180 8959
rect 9128 8916 9180 8925
rect 2780 8780 2832 8832
rect 3976 8780 4028 8832
rect 7104 8780 7156 8832
rect 9496 8916 9548 8968
rect 10784 9052 10836 9104
rect 11152 9095 11204 9104
rect 11152 9061 11157 9095
rect 11157 9061 11191 9095
rect 11191 9061 11204 9095
rect 11152 9052 11204 9061
rect 10232 8916 10284 8968
rect 10416 8916 10468 8968
rect 10784 8916 10836 8968
rect 10876 8916 10928 8968
rect 11060 8916 11112 8968
rect 11336 8916 11388 8968
rect 12992 8916 13044 8968
rect 13268 8959 13320 8968
rect 13268 8925 13277 8959
rect 13277 8925 13311 8959
rect 13311 8925 13320 8959
rect 13268 8916 13320 8925
rect 8116 8780 8168 8832
rect 8300 8780 8352 8832
rect 8576 8780 8628 8832
rect 9404 8780 9456 8832
rect 9772 8848 9824 8900
rect 10600 8848 10652 8900
rect 11152 8848 11204 8900
rect 11428 8848 11480 8900
rect 13360 8848 13412 8900
rect 10508 8823 10560 8832
rect 10508 8789 10517 8823
rect 10517 8789 10551 8823
rect 10551 8789 10560 8823
rect 10508 8780 10560 8789
rect 11060 8780 11112 8832
rect 12072 8780 12124 8832
rect 12348 8780 12400 8832
rect 8214 8678 8266 8730
rect 8278 8678 8330 8730
rect 8342 8678 8394 8730
rect 8406 8678 8458 8730
rect 8470 8678 8522 8730
rect 1860 8619 1912 8628
rect 1860 8585 1869 8619
rect 1869 8585 1903 8619
rect 1903 8585 1912 8619
rect 1860 8576 1912 8585
rect 2688 8576 2740 8628
rect 2872 8576 2924 8628
rect 6276 8576 6328 8628
rect 6552 8576 6604 8628
rect 7012 8576 7064 8628
rect 1676 8483 1728 8492
rect 1676 8449 1685 8483
rect 1685 8449 1719 8483
rect 1719 8449 1728 8483
rect 1676 8440 1728 8449
rect 1768 8440 1820 8492
rect 2596 8508 2648 8560
rect 3516 8551 3568 8560
rect 1952 8372 2004 8424
rect 2504 8440 2556 8492
rect 3516 8517 3525 8551
rect 3525 8517 3559 8551
rect 3559 8517 3568 8551
rect 3516 8508 3568 8517
rect 3608 8551 3660 8560
rect 3608 8517 3617 8551
rect 3617 8517 3651 8551
rect 3651 8517 3660 8551
rect 5632 8551 5684 8560
rect 3608 8508 3660 8517
rect 5632 8517 5641 8551
rect 5641 8517 5675 8551
rect 5675 8517 5684 8551
rect 5632 8508 5684 8517
rect 6644 8508 6696 8560
rect 3700 8440 3752 8492
rect 3976 8440 4028 8492
rect 4528 8440 4580 8492
rect 4804 8483 4856 8492
rect 4804 8449 4813 8483
rect 4813 8449 4847 8483
rect 4847 8449 4856 8483
rect 4804 8440 4856 8449
rect 5080 8483 5132 8492
rect 5080 8449 5089 8483
rect 5089 8449 5123 8483
rect 5123 8449 5132 8483
rect 5080 8440 5132 8449
rect 5540 8440 5592 8492
rect 5816 8483 5868 8492
rect 5816 8449 5825 8483
rect 5825 8449 5859 8483
rect 5859 8449 5868 8483
rect 5816 8440 5868 8449
rect 6092 8483 6144 8492
rect 6092 8449 6101 8483
rect 6101 8449 6135 8483
rect 6135 8449 6144 8483
rect 6092 8440 6144 8449
rect 6736 8483 6788 8492
rect 4712 8415 4764 8424
rect 4712 8381 4721 8415
rect 4721 8381 4755 8415
rect 4755 8381 4764 8415
rect 4712 8372 4764 8381
rect 6736 8449 6745 8483
rect 6745 8449 6779 8483
rect 6779 8449 6788 8483
rect 6736 8440 6788 8449
rect 7104 8440 7156 8492
rect 7840 8576 7892 8628
rect 8116 8576 8168 8628
rect 8576 8576 8628 8628
rect 7932 8508 7984 8560
rect 10324 8576 10376 8628
rect 10508 8576 10560 8628
rect 10416 8508 10468 8560
rect 10876 8508 10928 8560
rect 7012 8415 7064 8424
rect 2412 8304 2464 8356
rect 3332 8304 3384 8356
rect 3700 8304 3752 8356
rect 5816 8304 5868 8356
rect 7012 8381 7021 8415
rect 7021 8381 7055 8415
rect 7055 8381 7064 8415
rect 7012 8372 7064 8381
rect 7104 8347 7156 8356
rect 7104 8313 7113 8347
rect 7113 8313 7147 8347
rect 7147 8313 7156 8347
rect 7104 8304 7156 8313
rect 7564 8415 7616 8424
rect 7564 8381 7573 8415
rect 7573 8381 7607 8415
rect 7607 8381 7616 8415
rect 7564 8372 7616 8381
rect 7932 8347 7984 8356
rect 7932 8313 7941 8347
rect 7941 8313 7975 8347
rect 7975 8313 7984 8347
rect 7932 8304 7984 8313
rect 8208 8347 8260 8356
rect 8208 8313 8217 8347
rect 8217 8313 8251 8347
rect 8251 8313 8260 8347
rect 8208 8304 8260 8313
rect 8116 8236 8168 8288
rect 9036 8440 9088 8492
rect 9312 8483 9364 8492
rect 8668 8372 8720 8424
rect 8944 8372 8996 8424
rect 9312 8449 9321 8483
rect 9321 8449 9355 8483
rect 9355 8449 9364 8483
rect 9312 8440 9364 8449
rect 9496 8440 9548 8492
rect 9772 8440 9824 8492
rect 10692 8440 10744 8492
rect 11060 8483 11112 8492
rect 11060 8449 11069 8483
rect 11069 8449 11103 8483
rect 11103 8449 11112 8483
rect 11060 8440 11112 8449
rect 11152 8440 11204 8492
rect 11520 8483 11572 8492
rect 11520 8449 11529 8483
rect 11529 8449 11563 8483
rect 11563 8449 11572 8483
rect 11520 8440 11572 8449
rect 11612 8440 11664 8492
rect 9864 8372 9916 8424
rect 11428 8372 11480 8424
rect 9128 8236 9180 8288
rect 9588 8236 9640 8288
rect 9772 8279 9824 8288
rect 9772 8245 9781 8279
rect 9781 8245 9815 8279
rect 9815 8245 9824 8279
rect 9772 8236 9824 8245
rect 10048 8236 10100 8288
rect 11244 8347 11296 8356
rect 11244 8313 11253 8347
rect 11253 8313 11287 8347
rect 11287 8313 11296 8347
rect 11244 8304 11296 8313
rect 12072 8347 12124 8356
rect 12072 8313 12081 8347
rect 12081 8313 12115 8347
rect 12115 8313 12124 8347
rect 12072 8304 12124 8313
rect 13544 8551 13596 8560
rect 13544 8517 13553 8551
rect 13553 8517 13587 8551
rect 13587 8517 13596 8551
rect 13544 8508 13596 8517
rect 12716 8483 12768 8492
rect 12716 8449 12719 8483
rect 12719 8449 12768 8483
rect 12716 8440 12768 8449
rect 13452 8440 13504 8492
rect 12348 8372 12400 8424
rect 12992 8415 13044 8424
rect 12992 8381 13001 8415
rect 13001 8381 13035 8415
rect 13035 8381 13044 8415
rect 12992 8372 13044 8381
rect 13268 8304 13320 8356
rect 13360 8304 13412 8356
rect 10324 8279 10376 8288
rect 10324 8245 10333 8279
rect 10333 8245 10367 8279
rect 10367 8245 10376 8279
rect 10324 8236 10376 8245
rect 12164 8236 12216 8288
rect 12624 8236 12676 8288
rect 12808 8279 12860 8288
rect 12808 8245 12817 8279
rect 12817 8245 12851 8279
rect 12851 8245 12860 8279
rect 12808 8236 12860 8245
rect 4214 8134 4266 8186
rect 4278 8134 4330 8186
rect 4342 8134 4394 8186
rect 4406 8134 4458 8186
rect 4470 8134 4522 8186
rect 12214 8134 12266 8186
rect 12278 8134 12330 8186
rect 12342 8134 12394 8186
rect 12406 8134 12458 8186
rect 12470 8134 12522 8186
rect 2044 8032 2096 8084
rect 2596 8032 2648 8084
rect 4896 8032 4948 8084
rect 5816 8075 5868 8084
rect 5816 8041 5825 8075
rect 5825 8041 5859 8075
rect 5859 8041 5868 8075
rect 5816 8032 5868 8041
rect 7012 8032 7064 8084
rect 7840 8032 7892 8084
rect 8576 8032 8628 8084
rect 10048 8032 10100 8084
rect 10140 8032 10192 8084
rect 10232 8032 10284 8084
rect 8852 7964 8904 8016
rect 1400 7896 1452 7948
rect 1676 7871 1728 7880
rect 1676 7837 1685 7871
rect 1685 7837 1719 7871
rect 1719 7837 1728 7871
rect 1676 7828 1728 7837
rect 1952 7871 2004 7880
rect 1952 7837 1961 7871
rect 1961 7837 1995 7871
rect 1995 7837 2004 7871
rect 1952 7828 2004 7837
rect 2044 7871 2096 7880
rect 2044 7837 2053 7871
rect 2053 7837 2087 7871
rect 2087 7837 2096 7871
rect 2504 7896 2556 7948
rect 2044 7828 2096 7837
rect 2412 7871 2464 7880
rect 2412 7837 2421 7871
rect 2421 7837 2455 7871
rect 2455 7837 2464 7871
rect 2412 7828 2464 7837
rect 2596 7871 2648 7880
rect 2596 7837 2605 7871
rect 2605 7837 2639 7871
rect 2639 7837 2648 7871
rect 2596 7828 2648 7837
rect 3056 7828 3108 7880
rect 3700 7828 3752 7880
rect 3976 7828 4028 7880
rect 4620 7896 4672 7948
rect 4804 7896 4856 7948
rect 5172 7896 5224 7948
rect 4252 7871 4304 7880
rect 4252 7837 4261 7871
rect 4261 7837 4295 7871
rect 4295 7837 4304 7871
rect 4252 7828 4304 7837
rect 4712 7828 4764 7880
rect 5080 7828 5132 7880
rect 5908 7828 5960 7880
rect 6736 7896 6788 7948
rect 1768 7803 1820 7812
rect 1768 7769 1777 7803
rect 1777 7769 1811 7803
rect 1811 7769 1820 7803
rect 1768 7760 1820 7769
rect 4896 7803 4948 7812
rect 4896 7769 4905 7803
rect 4905 7769 4939 7803
rect 4939 7769 4948 7803
rect 4896 7760 4948 7769
rect 1492 7735 1544 7744
rect 1492 7701 1501 7735
rect 1501 7701 1535 7735
rect 1535 7701 1544 7735
rect 1492 7692 1544 7701
rect 4068 7692 4120 7744
rect 4160 7692 4212 7744
rect 6460 7871 6512 7880
rect 6460 7837 6469 7871
rect 6469 7837 6503 7871
rect 6503 7837 6512 7871
rect 6460 7828 6512 7837
rect 8208 7896 8260 7948
rect 8576 7896 8628 7948
rect 7288 7828 7340 7880
rect 7564 7828 7616 7880
rect 6644 7803 6696 7812
rect 6644 7769 6653 7803
rect 6653 7769 6687 7803
rect 6687 7769 6696 7803
rect 6644 7760 6696 7769
rect 6828 7803 6880 7812
rect 6828 7769 6837 7803
rect 6837 7769 6871 7803
rect 6871 7769 6880 7803
rect 6828 7760 6880 7769
rect 7012 7692 7064 7744
rect 7932 7760 7984 7812
rect 7564 7692 7616 7744
rect 8760 7760 8812 7812
rect 9128 7828 9180 7880
rect 9496 7896 9548 7948
rect 9404 7871 9456 7880
rect 9404 7837 9413 7871
rect 9413 7837 9447 7871
rect 9447 7837 9456 7871
rect 10416 7964 10468 8016
rect 9404 7828 9456 7837
rect 12624 8032 12676 8084
rect 13268 8032 13320 8084
rect 13544 8032 13596 8084
rect 10876 8007 10928 8016
rect 10876 7973 10885 8007
rect 10885 7973 10919 8007
rect 10919 7973 10928 8007
rect 10876 7964 10928 7973
rect 11980 7964 12032 8016
rect 10692 7896 10744 7948
rect 11060 7871 11112 7880
rect 9496 7760 9548 7812
rect 8208 7692 8260 7744
rect 9036 7692 9088 7744
rect 11060 7837 11069 7871
rect 11069 7837 11103 7871
rect 11103 7837 11112 7871
rect 11060 7828 11112 7837
rect 11244 7871 11296 7880
rect 11244 7837 11253 7871
rect 11253 7837 11287 7871
rect 11287 7837 11296 7871
rect 11244 7828 11296 7837
rect 11428 7871 11480 7880
rect 11428 7837 11454 7871
rect 11454 7837 11480 7871
rect 12164 7896 12216 7948
rect 12256 7896 12308 7948
rect 11428 7828 11480 7837
rect 11612 7828 11664 7880
rect 11980 7828 12032 7880
rect 12808 7828 12860 7880
rect 13452 7828 13504 7880
rect 10692 7803 10744 7812
rect 10692 7769 10710 7803
rect 10710 7769 10744 7803
rect 10692 7760 10744 7769
rect 11704 7803 11756 7812
rect 11704 7769 11713 7803
rect 11713 7769 11747 7803
rect 11747 7769 11756 7803
rect 11704 7760 11756 7769
rect 13176 7803 13228 7812
rect 9864 7692 9916 7744
rect 13176 7769 13185 7803
rect 13185 7769 13219 7803
rect 13219 7769 13228 7803
rect 13176 7760 13228 7769
rect 11980 7735 12032 7744
rect 11980 7701 11989 7735
rect 11989 7701 12023 7735
rect 12023 7701 12032 7735
rect 11980 7692 12032 7701
rect 8214 7590 8266 7642
rect 8278 7590 8330 7642
rect 8342 7590 8394 7642
rect 8406 7590 8458 7642
rect 8470 7590 8522 7642
rect 1492 7420 1544 7472
rect 2136 7352 2188 7404
rect 3700 7488 3752 7540
rect 4620 7488 4672 7540
rect 4712 7488 4764 7540
rect 2872 7420 2924 7472
rect 2964 7463 3016 7472
rect 2964 7429 2973 7463
rect 2973 7429 3007 7463
rect 3007 7429 3016 7463
rect 3148 7463 3200 7472
rect 2964 7420 3016 7429
rect 3148 7429 3157 7463
rect 3157 7429 3191 7463
rect 3191 7429 3200 7463
rect 3148 7420 3200 7429
rect 2596 7352 2648 7404
rect 4896 7420 4948 7472
rect 4712 7395 4764 7404
rect 4712 7361 4721 7395
rect 4721 7361 4755 7395
rect 4755 7361 4764 7395
rect 4712 7352 4764 7361
rect 5908 7488 5960 7540
rect 7656 7488 7708 7540
rect 9404 7488 9456 7540
rect 9956 7488 10008 7540
rect 11428 7488 11480 7540
rect 12164 7488 12216 7540
rect 5540 7420 5592 7472
rect 6736 7420 6788 7472
rect 8392 7463 8444 7472
rect 1768 7259 1820 7268
rect 1768 7225 1777 7259
rect 1777 7225 1811 7259
rect 1811 7225 1820 7259
rect 1768 7216 1820 7225
rect 3792 7327 3844 7336
rect 2320 7216 2372 7268
rect 3792 7293 3801 7327
rect 3801 7293 3835 7327
rect 3835 7293 3844 7327
rect 7012 7395 7064 7404
rect 3792 7284 3844 7293
rect 4896 7327 4948 7336
rect 4896 7293 4905 7327
rect 4905 7293 4939 7327
rect 4939 7293 4948 7327
rect 4896 7284 4948 7293
rect 4160 7216 4212 7268
rect 4252 7216 4304 7268
rect 2780 7191 2832 7200
rect 2780 7157 2789 7191
rect 2789 7157 2823 7191
rect 2823 7157 2832 7191
rect 2780 7148 2832 7157
rect 3516 7148 3568 7200
rect 4620 7148 4672 7200
rect 5540 7191 5592 7200
rect 5540 7157 5549 7191
rect 5549 7157 5583 7191
rect 5583 7157 5592 7191
rect 5540 7148 5592 7157
rect 6276 7216 6328 7268
rect 7012 7361 7021 7395
rect 7021 7361 7055 7395
rect 7055 7361 7064 7395
rect 7012 7352 7064 7361
rect 7196 7352 7248 7404
rect 8392 7429 8401 7463
rect 8401 7429 8435 7463
rect 8435 7429 8444 7463
rect 8392 7420 8444 7429
rect 13176 7463 13228 7472
rect 8944 7395 8996 7404
rect 7104 7327 7156 7336
rect 7104 7293 7113 7327
rect 7113 7293 7147 7327
rect 7147 7293 7156 7327
rect 7104 7284 7156 7293
rect 7748 7327 7800 7336
rect 7748 7293 7757 7327
rect 7757 7293 7791 7327
rect 7791 7293 7800 7327
rect 7748 7284 7800 7293
rect 8944 7361 8953 7395
rect 8953 7361 8987 7395
rect 8987 7361 8996 7395
rect 8944 7352 8996 7361
rect 9036 7352 9088 7404
rect 9128 7284 9180 7336
rect 9680 7395 9732 7404
rect 9680 7361 9691 7395
rect 9691 7361 9725 7395
rect 9725 7361 9732 7395
rect 9680 7352 9732 7361
rect 9864 7352 9916 7404
rect 10508 7352 10560 7404
rect 13176 7429 13185 7463
rect 13185 7429 13219 7463
rect 13219 7429 13228 7463
rect 13176 7420 13228 7429
rect 11060 7352 11112 7404
rect 11612 7352 11664 7404
rect 11704 7352 11756 7404
rect 12256 7395 12308 7404
rect 12256 7361 12265 7395
rect 12265 7361 12299 7395
rect 12299 7361 12308 7395
rect 12256 7352 12308 7361
rect 12808 7352 12860 7404
rect 10416 7284 10468 7336
rect 11152 7284 11204 7336
rect 13728 7352 13780 7404
rect 13268 7327 13320 7336
rect 13268 7293 13277 7327
rect 13277 7293 13311 7327
rect 13311 7293 13320 7327
rect 13268 7284 13320 7293
rect 6552 7148 6604 7200
rect 6736 7148 6788 7200
rect 11244 7259 11296 7268
rect 8852 7148 8904 7200
rect 9496 7148 9548 7200
rect 11244 7225 11253 7259
rect 11253 7225 11287 7259
rect 11287 7225 11296 7259
rect 11244 7216 11296 7225
rect 13176 7216 13228 7268
rect 4214 7046 4266 7098
rect 4278 7046 4330 7098
rect 4342 7046 4394 7098
rect 4406 7046 4458 7098
rect 4470 7046 4522 7098
rect 12214 7046 12266 7098
rect 12278 7046 12330 7098
rect 12342 7046 12394 7098
rect 12406 7046 12458 7098
rect 12470 7046 12522 7098
rect 1952 6944 2004 6996
rect 1584 6808 1636 6860
rect 2964 6851 3016 6860
rect 1492 6740 1544 6792
rect 2228 6783 2280 6792
rect 2228 6749 2237 6783
rect 2237 6749 2271 6783
rect 2271 6749 2280 6783
rect 2228 6740 2280 6749
rect 2320 6740 2372 6792
rect 2964 6817 2973 6851
rect 2973 6817 3007 6851
rect 3007 6817 3016 6851
rect 8116 6944 8168 6996
rect 12256 6944 12308 6996
rect 3792 6919 3844 6928
rect 3792 6885 3801 6919
rect 3801 6885 3835 6919
rect 3835 6885 3844 6919
rect 3792 6876 3844 6885
rect 6368 6876 6420 6928
rect 10140 6876 10192 6928
rect 10416 6919 10468 6928
rect 10416 6885 10421 6919
rect 10421 6885 10455 6919
rect 10455 6885 10468 6919
rect 10416 6876 10468 6885
rect 10876 6876 10928 6928
rect 3516 6851 3568 6860
rect 2964 6808 3016 6817
rect 3516 6817 3525 6851
rect 3525 6817 3559 6851
rect 3559 6817 3568 6851
rect 3516 6808 3568 6817
rect 2044 6672 2096 6724
rect 2780 6783 2832 6792
rect 2780 6749 2789 6783
rect 2789 6749 2823 6783
rect 2823 6749 2832 6783
rect 2780 6740 2832 6749
rect 3148 6740 3200 6792
rect 5540 6808 5592 6860
rect 7012 6808 7064 6860
rect 3240 6604 3292 6656
rect 4712 6740 4764 6792
rect 4896 6740 4948 6792
rect 5632 6740 5684 6792
rect 4620 6672 4672 6724
rect 6828 6740 6880 6792
rect 7564 6740 7616 6792
rect 7656 6672 7708 6724
rect 7840 6672 7892 6724
rect 8668 6851 8720 6860
rect 8668 6817 8677 6851
rect 8677 6817 8711 6851
rect 8711 6817 8720 6851
rect 8668 6808 8720 6817
rect 9404 6783 9456 6792
rect 9404 6749 9413 6783
rect 9413 6749 9447 6783
rect 9447 6749 9456 6783
rect 9404 6740 9456 6749
rect 9680 6783 9732 6792
rect 9680 6749 9689 6783
rect 9689 6749 9723 6783
rect 9723 6749 9732 6783
rect 9680 6740 9732 6749
rect 10324 6740 10376 6792
rect 10600 6740 10652 6792
rect 10784 6783 10836 6792
rect 10784 6749 10793 6783
rect 10793 6749 10827 6783
rect 10827 6749 10836 6783
rect 10784 6740 10836 6749
rect 11704 6808 11756 6860
rect 11796 6808 11848 6860
rect 12256 6808 12308 6860
rect 11244 6740 11296 6792
rect 11980 6740 12032 6792
rect 13176 6808 13228 6860
rect 11520 6715 11572 6724
rect 11520 6681 11529 6715
rect 11529 6681 11563 6715
rect 11563 6681 11572 6715
rect 11520 6672 11572 6681
rect 4068 6647 4120 6656
rect 4068 6613 4077 6647
rect 4077 6613 4111 6647
rect 4111 6613 4120 6647
rect 4068 6604 4120 6613
rect 4160 6647 4212 6656
rect 4160 6613 4169 6647
rect 4169 6613 4203 6647
rect 4203 6613 4212 6647
rect 4160 6604 4212 6613
rect 5540 6604 5592 6656
rect 6920 6604 6972 6656
rect 8024 6647 8076 6656
rect 8024 6613 8033 6647
rect 8033 6613 8067 6647
rect 8067 6613 8076 6647
rect 8024 6604 8076 6613
rect 9956 6604 10008 6656
rect 10416 6604 10468 6656
rect 11152 6604 11204 6656
rect 11796 6604 11848 6656
rect 11980 6604 12032 6656
rect 13176 6672 13228 6724
rect 8214 6502 8266 6554
rect 8278 6502 8330 6554
rect 8342 6502 8394 6554
rect 8406 6502 8458 6554
rect 8470 6502 8522 6554
rect 2228 6400 2280 6452
rect 3516 6400 3568 6452
rect 4160 6400 4212 6452
rect 7748 6400 7800 6452
rect 8760 6443 8812 6452
rect 8760 6409 8769 6443
rect 8769 6409 8803 6443
rect 8803 6409 8812 6443
rect 8760 6400 8812 6409
rect 9220 6400 9272 6452
rect 9312 6400 9364 6452
rect 9956 6443 10008 6452
rect 9956 6409 9965 6443
rect 9965 6409 9999 6443
rect 9999 6409 10008 6443
rect 9956 6400 10008 6409
rect 11520 6400 11572 6452
rect 4068 6375 4120 6384
rect 2044 6307 2096 6316
rect 2044 6273 2053 6307
rect 2053 6273 2087 6307
rect 2087 6273 2096 6307
rect 2044 6264 2096 6273
rect 2136 6264 2188 6316
rect 2780 6307 2832 6316
rect 2780 6273 2789 6307
rect 2789 6273 2823 6307
rect 2823 6273 2832 6307
rect 3332 6307 3384 6316
rect 2780 6264 2832 6273
rect 3332 6273 3341 6307
rect 3341 6273 3375 6307
rect 3375 6273 3384 6307
rect 3332 6264 3384 6273
rect 4068 6341 4077 6375
rect 4077 6341 4111 6375
rect 4111 6341 4120 6375
rect 4068 6332 4120 6341
rect 5080 6332 5132 6384
rect 3148 6196 3200 6248
rect 3700 6307 3752 6316
rect 3700 6273 3709 6307
rect 3709 6273 3743 6307
rect 3743 6273 3752 6307
rect 3700 6264 3752 6273
rect 3884 6307 3936 6316
rect 3884 6273 3893 6307
rect 3893 6273 3927 6307
rect 3927 6273 3936 6307
rect 4252 6307 4304 6316
rect 3884 6264 3936 6273
rect 4252 6273 4261 6307
rect 4261 6273 4295 6307
rect 4295 6273 4304 6307
rect 4252 6264 4304 6273
rect 5172 6264 5224 6316
rect 5540 6307 5592 6316
rect 5540 6273 5549 6307
rect 5549 6273 5583 6307
rect 5583 6273 5592 6307
rect 5540 6264 5592 6273
rect 6184 6332 6236 6384
rect 7012 6332 7064 6384
rect 8576 6375 8628 6384
rect 8576 6341 8585 6375
rect 8585 6341 8619 6375
rect 8619 6341 8628 6375
rect 8576 6332 8628 6341
rect 3516 6196 3568 6248
rect 4160 6196 4212 6248
rect 4988 6196 5040 6248
rect 4712 6128 4764 6180
rect 6920 6264 6972 6316
rect 7748 6264 7800 6316
rect 11060 6332 11112 6384
rect 11244 6332 11296 6384
rect 6644 6239 6696 6248
rect 6644 6205 6653 6239
rect 6653 6205 6687 6239
rect 6687 6205 6696 6239
rect 6644 6196 6696 6205
rect 7380 6239 7432 6248
rect 7380 6205 7389 6239
rect 7389 6205 7423 6239
rect 7423 6205 7432 6239
rect 7380 6196 7432 6205
rect 10508 6264 10560 6316
rect 10416 6239 10468 6248
rect 10416 6205 10425 6239
rect 10425 6205 10459 6239
rect 10459 6205 10468 6239
rect 10416 6196 10468 6205
rect 11152 6239 11204 6248
rect 11152 6205 11161 6239
rect 11161 6205 11195 6239
rect 11195 6205 11204 6239
rect 11152 6196 11204 6205
rect 11704 6307 11756 6316
rect 11704 6273 11713 6307
rect 11713 6273 11747 6307
rect 11747 6273 11756 6307
rect 11704 6264 11756 6273
rect 11980 6307 12032 6316
rect 11980 6273 11989 6307
rect 11989 6273 12023 6307
rect 12023 6273 12032 6307
rect 11980 6264 12032 6273
rect 13452 6307 13504 6316
rect 13452 6273 13461 6307
rect 13461 6273 13495 6307
rect 13495 6273 13504 6307
rect 13452 6264 13504 6273
rect 11428 6196 11480 6248
rect 7932 6128 7984 6180
rect 9680 6128 9732 6180
rect 10324 6171 10376 6180
rect 2688 6060 2740 6112
rect 4068 6060 4120 6112
rect 4160 6060 4212 6112
rect 5816 6060 5868 6112
rect 6368 6103 6420 6112
rect 6368 6069 6377 6103
rect 6377 6069 6411 6103
rect 6411 6069 6420 6103
rect 6368 6060 6420 6069
rect 7840 6103 7892 6112
rect 7840 6069 7849 6103
rect 7849 6069 7883 6103
rect 7883 6069 7892 6103
rect 7840 6060 7892 6069
rect 8392 6060 8444 6112
rect 9772 6103 9824 6112
rect 9772 6069 9781 6103
rect 9781 6069 9815 6103
rect 9815 6069 9824 6103
rect 9772 6060 9824 6069
rect 10324 6137 10333 6171
rect 10333 6137 10367 6171
rect 10367 6137 10376 6171
rect 10324 6128 10376 6137
rect 13176 6128 13228 6180
rect 4214 5958 4266 6010
rect 4278 5958 4330 6010
rect 4342 5958 4394 6010
rect 4406 5958 4458 6010
rect 4470 5958 4522 6010
rect 12214 5958 12266 6010
rect 12278 5958 12330 6010
rect 12342 5958 12394 6010
rect 12406 5958 12458 6010
rect 12470 5958 12522 6010
rect 1492 5899 1544 5908
rect 1492 5865 1501 5899
rect 1501 5865 1535 5899
rect 1535 5865 1544 5899
rect 1492 5856 1544 5865
rect 2044 5856 2096 5908
rect 2136 5831 2188 5840
rect 2136 5797 2145 5831
rect 2145 5797 2179 5831
rect 2179 5797 2188 5831
rect 2136 5788 2188 5797
rect 2780 5856 2832 5908
rect 3608 5856 3660 5908
rect 5448 5856 5500 5908
rect 7748 5899 7800 5908
rect 7748 5865 7757 5899
rect 7757 5865 7791 5899
rect 7791 5865 7800 5899
rect 7748 5856 7800 5865
rect 7840 5856 7892 5908
rect 4712 5788 4764 5840
rect 4896 5788 4948 5840
rect 5724 5788 5776 5840
rect 8116 5788 8168 5840
rect 1400 5695 1452 5704
rect 1400 5661 1409 5695
rect 1409 5661 1443 5695
rect 1443 5661 1452 5695
rect 1400 5652 1452 5661
rect 2596 5695 2648 5704
rect 2596 5661 2605 5695
rect 2605 5661 2639 5695
rect 2639 5661 2648 5695
rect 2596 5652 2648 5661
rect 2780 5652 2832 5704
rect 2504 5584 2556 5636
rect 3148 5652 3200 5704
rect 3700 5652 3752 5704
rect 4068 5695 4120 5704
rect 4068 5661 4077 5695
rect 4077 5661 4111 5695
rect 4111 5661 4120 5695
rect 4068 5652 4120 5661
rect 4804 5720 4856 5772
rect 3332 5584 3384 5636
rect 3516 5584 3568 5636
rect 3608 5516 3660 5568
rect 4252 5559 4304 5568
rect 4252 5525 4261 5559
rect 4261 5525 4295 5559
rect 4295 5525 4304 5559
rect 4252 5516 4304 5525
rect 7656 5763 7708 5772
rect 7656 5729 7665 5763
rect 7665 5729 7699 5763
rect 7699 5729 7708 5763
rect 7656 5720 7708 5729
rect 7840 5720 7892 5772
rect 4988 5673 5040 5682
rect 4988 5639 4997 5673
rect 4997 5639 5031 5673
rect 5031 5639 5040 5673
rect 4988 5630 5040 5639
rect 5448 5652 5500 5704
rect 5540 5652 5592 5704
rect 7932 5695 7984 5704
rect 7932 5661 7941 5695
rect 7941 5661 7975 5695
rect 7975 5661 7984 5695
rect 7932 5652 7984 5661
rect 8392 5695 8444 5704
rect 8392 5661 8401 5695
rect 8401 5661 8435 5695
rect 8435 5661 8444 5695
rect 8392 5652 8444 5661
rect 9956 5856 10008 5908
rect 11152 5856 11204 5908
rect 11336 5720 11388 5772
rect 11888 5856 11940 5908
rect 13268 5856 13320 5908
rect 9680 5652 9732 5704
rect 11704 5652 11756 5704
rect 12072 5652 12124 5704
rect 13452 5652 13504 5704
rect 4988 5516 5040 5568
rect 7012 5584 7064 5636
rect 5816 5516 5868 5568
rect 8024 5516 8076 5568
rect 8576 5516 8628 5568
rect 11428 5584 11480 5636
rect 12992 5627 13044 5636
rect 12992 5593 13001 5627
rect 13001 5593 13035 5627
rect 13035 5593 13044 5627
rect 12992 5584 13044 5593
rect 13268 5627 13320 5636
rect 13268 5593 13277 5627
rect 13277 5593 13311 5627
rect 13311 5593 13320 5627
rect 13268 5584 13320 5593
rect 8214 5414 8266 5466
rect 8278 5414 8330 5466
rect 8342 5414 8394 5466
rect 8406 5414 8458 5466
rect 8470 5414 8522 5466
rect 2596 5287 2648 5296
rect 2596 5253 2605 5287
rect 2605 5253 2639 5287
rect 2639 5253 2648 5287
rect 2596 5244 2648 5253
rect 2780 5287 2832 5296
rect 2780 5253 2789 5287
rect 2789 5253 2823 5287
rect 2823 5253 2832 5287
rect 4804 5312 4856 5364
rect 7840 5312 7892 5364
rect 10232 5312 10284 5364
rect 10508 5355 10560 5364
rect 10508 5321 10517 5355
rect 10517 5321 10551 5355
rect 10551 5321 10560 5355
rect 10508 5312 10560 5321
rect 11612 5312 11664 5364
rect 11704 5312 11756 5364
rect 13636 5312 13688 5364
rect 2780 5244 2832 5253
rect 4252 5244 4304 5296
rect 8024 5287 8076 5296
rect 3332 5176 3384 5228
rect 3424 5219 3476 5228
rect 3424 5185 3433 5219
rect 3433 5185 3467 5219
rect 3467 5185 3476 5219
rect 3424 5176 3476 5185
rect 5632 5176 5684 5228
rect 6184 5219 6236 5228
rect 6184 5185 6193 5219
rect 6193 5185 6227 5219
rect 6227 5185 6236 5219
rect 8024 5253 8033 5287
rect 8033 5253 8067 5287
rect 8067 5253 8076 5287
rect 8024 5244 8076 5253
rect 8668 5244 8720 5296
rect 11796 5287 11848 5296
rect 11796 5253 11805 5287
rect 11805 5253 11839 5287
rect 11839 5253 11848 5287
rect 11796 5244 11848 5253
rect 11888 5244 11940 5296
rect 6184 5176 6236 5185
rect 2872 5151 2924 5160
rect 2872 5117 2881 5151
rect 2881 5117 2915 5151
rect 2915 5117 2924 5151
rect 2872 5108 2924 5117
rect 1768 4972 1820 5024
rect 1860 4972 1912 5024
rect 4528 5108 4580 5160
rect 5264 5108 5316 5160
rect 6920 5176 6972 5228
rect 10140 5176 10192 5228
rect 6736 5108 6788 5160
rect 7748 5151 7800 5160
rect 7748 5117 7757 5151
rect 7757 5117 7791 5151
rect 7791 5117 7800 5151
rect 7748 5108 7800 5117
rect 10784 5176 10836 5228
rect 11060 5176 11112 5228
rect 11336 5176 11388 5228
rect 11520 5219 11572 5228
rect 11520 5185 11529 5219
rect 11529 5185 11563 5219
rect 11563 5185 11572 5219
rect 11520 5176 11572 5185
rect 3424 4972 3476 5024
rect 4160 4972 4212 5024
rect 6368 5040 6420 5092
rect 9128 5040 9180 5092
rect 11152 5040 11204 5092
rect 5540 4972 5592 5024
rect 6460 5015 6512 5024
rect 6460 4981 6469 5015
rect 6469 4981 6503 5015
rect 6503 4981 6512 5015
rect 6460 4972 6512 4981
rect 12992 4972 13044 5024
rect 4214 4870 4266 4922
rect 4278 4870 4330 4922
rect 4342 4870 4394 4922
rect 4406 4870 4458 4922
rect 4470 4870 4522 4922
rect 12214 4870 12266 4922
rect 12278 4870 12330 4922
rect 12342 4870 12394 4922
rect 12406 4870 12458 4922
rect 12470 4870 12522 4922
rect 2780 4768 2832 4820
rect 2872 4700 2924 4752
rect 1768 4675 1820 4684
rect 1768 4641 1777 4675
rect 1777 4641 1811 4675
rect 1811 4641 1820 4675
rect 1768 4632 1820 4641
rect 1768 4496 1820 4548
rect 3056 4496 3108 4548
rect 3332 4768 3384 4820
rect 3884 4700 3936 4752
rect 4068 4632 4120 4684
rect 8760 4768 8812 4820
rect 10416 4768 10468 4820
rect 4896 4700 4948 4752
rect 6276 4700 6328 4752
rect 7380 4700 7432 4752
rect 11428 4700 11480 4752
rect 4712 4632 4764 4684
rect 4160 4564 4212 4616
rect 5356 4632 5408 4684
rect 7748 4632 7800 4684
rect 9956 4632 10008 4684
rect 11520 4632 11572 4684
rect 8852 4564 8904 4616
rect 11612 4607 11664 4616
rect 4620 4539 4672 4548
rect 4620 4505 4629 4539
rect 4629 4505 4663 4539
rect 4663 4505 4672 4539
rect 4620 4496 4672 4505
rect 5172 4496 5224 4548
rect 5540 4496 5592 4548
rect 6920 4496 6972 4548
rect 7932 4496 7984 4548
rect 8576 4496 8628 4548
rect 11612 4573 11621 4607
rect 11621 4573 11655 4607
rect 11655 4573 11664 4607
rect 11612 4564 11664 4573
rect 11980 4607 12032 4616
rect 2780 4428 2832 4480
rect 3240 4428 3292 4480
rect 4712 4428 4764 4480
rect 9220 4428 9272 4480
rect 9772 4496 9824 4548
rect 10600 4496 10652 4548
rect 11152 4496 11204 4548
rect 11428 4496 11480 4548
rect 11520 4496 11572 4548
rect 11980 4573 11989 4607
rect 11989 4573 12023 4607
rect 12023 4573 12032 4607
rect 11980 4564 12032 4573
rect 13268 4607 13320 4616
rect 13268 4573 13277 4607
rect 13277 4573 13311 4607
rect 13311 4573 13320 4607
rect 13268 4564 13320 4573
rect 11796 4428 11848 4480
rect 13084 4428 13136 4480
rect 8214 4326 8266 4378
rect 8278 4326 8330 4378
rect 8342 4326 8394 4378
rect 8406 4326 8458 4378
rect 8470 4326 8522 4378
rect 3056 4224 3108 4276
rect 3424 4224 3476 4276
rect 5724 4224 5776 4276
rect 7012 4267 7064 4276
rect 7012 4233 7021 4267
rect 7021 4233 7055 4267
rect 7055 4233 7064 4267
rect 7012 4224 7064 4233
rect 7104 4224 7156 4276
rect 10600 4267 10652 4276
rect 5172 4156 5224 4208
rect 6368 4199 6420 4208
rect 6368 4165 6377 4199
rect 6377 4165 6411 4199
rect 6411 4165 6420 4199
rect 6368 4156 6420 4165
rect 6828 4156 6880 4208
rect 1952 4088 2004 4140
rect 2228 4131 2280 4140
rect 2228 4097 2237 4131
rect 2237 4097 2271 4131
rect 2271 4097 2280 4131
rect 2228 4088 2280 4097
rect 2780 4088 2832 4140
rect 3424 4088 3476 4140
rect 3700 4131 3752 4140
rect 2044 4063 2096 4072
rect 2044 4029 2053 4063
rect 2053 4029 2087 4063
rect 2087 4029 2096 4063
rect 2044 4020 2096 4029
rect 2136 4063 2188 4072
rect 2136 4029 2145 4063
rect 2145 4029 2179 4063
rect 2179 4029 2188 4063
rect 2136 4020 2188 4029
rect 1860 3952 1912 4004
rect 3056 4063 3108 4072
rect 3056 4029 3065 4063
rect 3065 4029 3099 4063
rect 3099 4029 3108 4063
rect 3056 4020 3108 4029
rect 3700 4097 3709 4131
rect 3709 4097 3743 4131
rect 3743 4097 3752 4131
rect 3700 4088 3752 4097
rect 3976 4088 4028 4140
rect 4160 4131 4212 4140
rect 4160 4097 4176 4131
rect 4176 4097 4210 4131
rect 4210 4097 4212 4131
rect 4160 4088 4212 4097
rect 7012 4131 7064 4140
rect 7012 4097 7021 4131
rect 7021 4097 7055 4131
rect 7055 4097 7064 4131
rect 7012 4088 7064 4097
rect 7196 4131 7248 4140
rect 7196 4097 7205 4131
rect 7205 4097 7239 4131
rect 7239 4097 7248 4131
rect 7196 4088 7248 4097
rect 8300 4156 8352 4208
rect 9036 4156 9088 4208
rect 10600 4233 10609 4267
rect 10609 4233 10643 4267
rect 10643 4233 10652 4267
rect 10600 4224 10652 4233
rect 11888 4224 11940 4276
rect 2964 3952 3016 4004
rect 3884 3952 3936 4004
rect 1492 3927 1544 3936
rect 1492 3893 1501 3927
rect 1501 3893 1535 3927
rect 1535 3893 1544 3927
rect 1492 3884 1544 3893
rect 2320 3884 2372 3936
rect 2596 3884 2648 3936
rect 5448 4020 5500 4072
rect 7748 4063 7800 4072
rect 7748 4029 7757 4063
rect 7757 4029 7791 4063
rect 7791 4029 7800 4063
rect 7748 4020 7800 4029
rect 8116 4020 8168 4072
rect 8392 4020 8444 4072
rect 10140 4088 10192 4140
rect 11612 4156 11664 4208
rect 13360 4199 13412 4208
rect 13360 4165 13369 4199
rect 13369 4165 13403 4199
rect 13403 4165 13412 4199
rect 13360 4156 13412 4165
rect 9588 4020 9640 4072
rect 5448 3884 5500 3936
rect 5908 3927 5960 3936
rect 5908 3893 5917 3927
rect 5917 3893 5951 3927
rect 5951 3893 5960 3927
rect 5908 3884 5960 3893
rect 6092 3927 6144 3936
rect 6092 3893 6101 3927
rect 6101 3893 6135 3927
rect 6135 3893 6144 3927
rect 6092 3884 6144 3893
rect 10508 3952 10560 4004
rect 11336 4088 11388 4140
rect 11796 4088 11848 4140
rect 12072 4088 12124 4140
rect 12992 4131 13044 4140
rect 12992 4097 13001 4131
rect 13001 4097 13035 4131
rect 13035 4097 13044 4131
rect 12992 4088 13044 4097
rect 11428 4020 11480 4072
rect 6644 3884 6696 3936
rect 8116 3884 8168 3936
rect 9680 3884 9732 3936
rect 11520 3952 11572 4004
rect 12072 3952 12124 4004
rect 12808 4020 12860 4072
rect 13176 4020 13228 4072
rect 11704 3927 11756 3936
rect 11704 3893 11713 3927
rect 11713 3893 11747 3927
rect 11747 3893 11756 3927
rect 11704 3884 11756 3893
rect 13452 3884 13504 3936
rect 4214 3782 4266 3834
rect 4278 3782 4330 3834
rect 4342 3782 4394 3834
rect 4406 3782 4458 3834
rect 4470 3782 4522 3834
rect 12214 3782 12266 3834
rect 12278 3782 12330 3834
rect 12342 3782 12394 3834
rect 12406 3782 12458 3834
rect 12470 3782 12522 3834
rect 1400 3723 1452 3732
rect 1400 3689 1409 3723
rect 1409 3689 1443 3723
rect 1443 3689 1452 3723
rect 1400 3680 1452 3689
rect 1676 3723 1728 3732
rect 1676 3689 1685 3723
rect 1685 3689 1719 3723
rect 1719 3689 1728 3723
rect 1676 3680 1728 3689
rect 3332 3680 3384 3732
rect 5080 3680 5132 3732
rect 5908 3680 5960 3732
rect 6000 3680 6052 3732
rect 6368 3723 6420 3732
rect 6368 3689 6377 3723
rect 6377 3689 6411 3723
rect 6411 3689 6420 3723
rect 6368 3680 6420 3689
rect 1492 3612 1544 3664
rect 2688 3612 2740 3664
rect 3424 3612 3476 3664
rect 4896 3612 4948 3664
rect 5172 3612 5224 3664
rect 7104 3680 7156 3732
rect 11704 3680 11756 3732
rect 11980 3680 12032 3732
rect 13084 3680 13136 3732
rect 8668 3655 8720 3664
rect 2780 3544 2832 3596
rect 5448 3544 5500 3596
rect 1860 3519 1912 3528
rect 1860 3485 1869 3519
rect 1869 3485 1903 3519
rect 1903 3485 1912 3519
rect 1860 3476 1912 3485
rect 2044 3519 2096 3528
rect 2044 3485 2053 3519
rect 2053 3485 2087 3519
rect 2087 3485 2096 3519
rect 2044 3476 2096 3485
rect 3148 3519 3200 3528
rect 3148 3485 3157 3519
rect 3157 3485 3191 3519
rect 3191 3485 3200 3519
rect 3148 3476 3200 3485
rect 3516 3476 3568 3528
rect 3976 3476 4028 3528
rect 2136 3451 2188 3460
rect 2136 3417 2145 3451
rect 2145 3417 2179 3451
rect 2179 3417 2188 3451
rect 2136 3408 2188 3417
rect 2320 3408 2372 3460
rect 4068 3408 4120 3460
rect 1952 3340 2004 3392
rect 3332 3340 3384 3392
rect 3700 3340 3752 3392
rect 3884 3340 3936 3392
rect 8668 3621 8677 3655
rect 8677 3621 8711 3655
rect 8711 3621 8720 3655
rect 8668 3612 8720 3621
rect 9036 3655 9088 3664
rect 9036 3621 9045 3655
rect 9045 3621 9079 3655
rect 9079 3621 9088 3655
rect 9036 3612 9088 3621
rect 5908 3587 5960 3596
rect 5908 3553 5917 3587
rect 5917 3553 5951 3587
rect 5951 3553 5960 3587
rect 5908 3544 5960 3553
rect 6644 3544 6696 3596
rect 7748 3544 7800 3596
rect 8760 3544 8812 3596
rect 4988 3408 5040 3460
rect 5816 3476 5868 3528
rect 5540 3408 5592 3460
rect 6460 3476 6512 3528
rect 8208 3476 8260 3528
rect 8576 3519 8628 3528
rect 7564 3408 7616 3460
rect 8576 3485 8585 3519
rect 8585 3485 8619 3519
rect 8619 3485 8628 3519
rect 9128 3544 9180 3596
rect 9036 3519 9088 3528
rect 8576 3476 8628 3485
rect 9036 3485 9045 3519
rect 9045 3485 9079 3519
rect 9079 3485 9088 3519
rect 9680 3612 9732 3664
rect 11244 3612 11296 3664
rect 11520 3612 11572 3664
rect 9036 3476 9088 3485
rect 9496 3476 9548 3528
rect 11612 3519 11664 3528
rect 11612 3485 11621 3519
rect 11621 3485 11655 3519
rect 11655 3485 11664 3519
rect 11612 3476 11664 3485
rect 11980 3476 12032 3528
rect 12900 3544 12952 3596
rect 10048 3408 10100 3460
rect 12072 3451 12124 3460
rect 6276 3340 6328 3392
rect 6828 3340 6880 3392
rect 8760 3340 8812 3392
rect 9128 3340 9180 3392
rect 12072 3417 12081 3451
rect 12081 3417 12115 3451
rect 12115 3417 12124 3451
rect 12072 3408 12124 3417
rect 13360 3519 13412 3528
rect 13360 3485 13369 3519
rect 13369 3485 13403 3519
rect 13403 3485 13412 3519
rect 13360 3476 13412 3485
rect 11796 3340 11848 3392
rect 8214 3238 8266 3290
rect 8278 3238 8330 3290
rect 8342 3238 8394 3290
rect 8406 3238 8458 3290
rect 8470 3238 8522 3290
rect 2044 3136 2096 3188
rect 2596 3136 2648 3188
rect 3332 3136 3384 3188
rect 5816 3179 5868 3188
rect 5816 3145 5825 3179
rect 5825 3145 5859 3179
rect 5859 3145 5868 3179
rect 5816 3136 5868 3145
rect 6828 3136 6880 3188
rect 7932 3179 7984 3188
rect 7932 3145 7941 3179
rect 7941 3145 7975 3179
rect 7975 3145 7984 3179
rect 7932 3136 7984 3145
rect 2780 3068 2832 3120
rect 3424 3068 3476 3120
rect 2320 3043 2372 3052
rect 2320 3009 2329 3043
rect 2329 3009 2363 3043
rect 2363 3009 2372 3043
rect 2320 3000 2372 3009
rect 1768 2932 1820 2984
rect 2412 2975 2464 2984
rect 2412 2941 2421 2975
rect 2421 2941 2455 2975
rect 2455 2941 2464 2975
rect 2412 2932 2464 2941
rect 2688 2975 2740 2984
rect 2688 2941 2697 2975
rect 2697 2941 2731 2975
rect 2731 2941 2740 2975
rect 2688 2932 2740 2941
rect 3976 2932 4028 2984
rect 5172 3068 5224 3120
rect 4712 3043 4764 3052
rect 4712 3009 4721 3043
rect 4721 3009 4755 3043
rect 4755 3009 4764 3043
rect 4712 3000 4764 3009
rect 5448 3000 5500 3052
rect 5908 3043 5960 3052
rect 5908 3009 5917 3043
rect 5917 3009 5951 3043
rect 5951 3009 5960 3043
rect 5908 3000 5960 3009
rect 6092 3068 6144 3120
rect 6920 3111 6972 3120
rect 6920 3077 6929 3111
rect 6929 3077 6963 3111
rect 6963 3077 6972 3111
rect 6920 3068 6972 3077
rect 7380 3068 7432 3120
rect 8576 3136 8628 3188
rect 8760 3136 8812 3188
rect 11060 3136 11112 3188
rect 6276 3000 6328 3052
rect 7012 3043 7064 3052
rect 7012 3009 7021 3043
rect 7021 3009 7055 3043
rect 7055 3009 7064 3043
rect 7012 3000 7064 3009
rect 7196 3000 7248 3052
rect 4620 2932 4672 2984
rect 5080 2932 5132 2984
rect 5724 2932 5776 2984
rect 4160 2796 4212 2848
rect 5172 2839 5224 2848
rect 5172 2805 5181 2839
rect 5181 2805 5215 2839
rect 5215 2805 5224 2839
rect 5172 2796 5224 2805
rect 5264 2796 5316 2848
rect 6736 2932 6788 2984
rect 7380 2975 7432 2984
rect 7380 2941 7389 2975
rect 7389 2941 7423 2975
rect 7423 2941 7432 2975
rect 7380 2932 7432 2941
rect 8116 3068 8168 3120
rect 11796 3136 11848 3188
rect 11888 3136 11940 3188
rect 12900 3136 12952 3188
rect 13176 3179 13228 3188
rect 13176 3145 13185 3179
rect 13185 3145 13219 3179
rect 13219 3145 13228 3179
rect 13176 3136 13228 3145
rect 11244 3068 11296 3120
rect 9220 3043 9272 3052
rect 9220 3009 9229 3043
rect 9229 3009 9263 3043
rect 9263 3009 9272 3043
rect 9220 3000 9272 3009
rect 11060 3000 11112 3052
rect 11888 3043 11940 3052
rect 8300 2932 8352 2984
rect 9496 2975 9548 2984
rect 8024 2864 8076 2916
rect 9036 2864 9088 2916
rect 9220 2864 9272 2916
rect 9496 2941 9505 2975
rect 9505 2941 9539 2975
rect 9539 2941 9548 2975
rect 9496 2932 9548 2941
rect 11520 2975 11572 2984
rect 8208 2796 8260 2848
rect 10508 2796 10560 2848
rect 11520 2941 11529 2975
rect 11529 2941 11563 2975
rect 11563 2941 11572 2975
rect 11520 2932 11572 2941
rect 11888 3009 11897 3043
rect 11897 3009 11931 3043
rect 11931 3009 11940 3043
rect 11888 3000 11940 3009
rect 11980 2932 12032 2984
rect 11888 2864 11940 2916
rect 12164 2975 12216 2984
rect 12164 2941 12173 2975
rect 12173 2941 12207 2975
rect 12207 2941 12216 2975
rect 12164 2932 12216 2941
rect 13268 3000 13320 3052
rect 4214 2694 4266 2746
rect 4278 2694 4330 2746
rect 4342 2694 4394 2746
rect 4406 2694 4458 2746
rect 4470 2694 4522 2746
rect 12214 2694 12266 2746
rect 12278 2694 12330 2746
rect 12342 2694 12394 2746
rect 12406 2694 12458 2746
rect 12470 2694 12522 2746
rect 2136 2635 2188 2644
rect 2136 2601 2145 2635
rect 2145 2601 2179 2635
rect 2179 2601 2188 2635
rect 2136 2592 2188 2601
rect 2228 2592 2280 2644
rect 3424 2592 3476 2644
rect 2044 2524 2096 2576
rect 3608 2592 3660 2644
rect 4068 2592 4120 2644
rect 7748 2592 7800 2644
rect 9128 2592 9180 2644
rect 2320 2456 2372 2508
rect 1676 2431 1728 2440
rect 1676 2397 1685 2431
rect 1685 2397 1719 2431
rect 1719 2397 1728 2431
rect 1676 2388 1728 2397
rect 1952 2431 2004 2440
rect 1952 2397 1961 2431
rect 1961 2397 1995 2431
rect 1995 2397 2004 2431
rect 1952 2388 2004 2397
rect 2964 2431 3016 2440
rect 2964 2397 2973 2431
rect 2973 2397 3007 2431
rect 3007 2397 3016 2431
rect 3148 2431 3200 2440
rect 2964 2388 3016 2397
rect 3148 2397 3157 2431
rect 3157 2397 3191 2431
rect 3191 2397 3200 2431
rect 3148 2388 3200 2397
rect 3700 2456 3752 2508
rect 5080 2456 5132 2508
rect 5356 2456 5408 2508
rect 5540 2456 5592 2508
rect 7104 2524 7156 2576
rect 10140 2592 10192 2644
rect 12624 2635 12676 2644
rect 12624 2601 12633 2635
rect 12633 2601 12667 2635
rect 12667 2601 12676 2635
rect 12624 2592 12676 2601
rect 7288 2456 7340 2508
rect 7564 2456 7616 2508
rect 2780 2320 2832 2372
rect 4896 2388 4948 2440
rect 5264 2431 5316 2440
rect 4160 2363 4212 2372
rect 1676 2252 1728 2304
rect 2136 2252 2188 2304
rect 4160 2329 4169 2363
rect 4169 2329 4203 2363
rect 4203 2329 4212 2363
rect 5264 2397 5273 2431
rect 5273 2397 5307 2431
rect 5307 2397 5316 2431
rect 5264 2388 5316 2397
rect 5632 2431 5684 2440
rect 5632 2397 5641 2431
rect 5641 2397 5675 2431
rect 5675 2397 5684 2431
rect 5632 2388 5684 2397
rect 7472 2388 7524 2440
rect 8484 2456 8536 2508
rect 4160 2320 4212 2329
rect 7288 2320 7340 2372
rect 7656 2320 7708 2372
rect 8024 2388 8076 2440
rect 8576 2388 8628 2440
rect 9128 2431 9180 2440
rect 9128 2397 9137 2431
rect 9137 2397 9171 2431
rect 9171 2397 9180 2431
rect 9128 2388 9180 2397
rect 11428 2431 11480 2440
rect 11428 2397 11437 2431
rect 11437 2397 11471 2431
rect 11471 2397 11480 2431
rect 11428 2388 11480 2397
rect 11612 2431 11664 2440
rect 11612 2397 11621 2431
rect 11621 2397 11655 2431
rect 11655 2397 11664 2431
rect 11612 2388 11664 2397
rect 11520 2320 11572 2372
rect 11888 2456 11940 2508
rect 13360 2499 13412 2508
rect 13360 2465 13369 2499
rect 13369 2465 13403 2499
rect 13403 2465 13412 2499
rect 13360 2456 13412 2465
rect 13176 2388 13228 2440
rect 12072 2320 12124 2372
rect 4436 2252 4488 2304
rect 4896 2252 4948 2304
rect 4988 2252 5040 2304
rect 5724 2252 5776 2304
rect 9680 2252 9732 2304
rect 11980 2252 12032 2304
rect 8214 2150 8266 2202
rect 8278 2150 8330 2202
rect 8342 2150 8394 2202
rect 8406 2150 8458 2202
rect 8470 2150 8522 2202
rect 1952 1980 2004 2032
rect 4620 2048 4672 2100
rect 4896 2048 4948 2100
rect 6644 2048 6696 2100
rect 7288 2091 7340 2100
rect 7288 2057 7297 2091
rect 7297 2057 7331 2091
rect 7331 2057 7340 2091
rect 7288 2048 7340 2057
rect 7748 2091 7800 2100
rect 7748 2057 7757 2091
rect 7757 2057 7791 2091
rect 7791 2057 7800 2091
rect 7748 2048 7800 2057
rect 9680 2048 9732 2100
rect 11612 2048 11664 2100
rect 5448 1980 5500 2032
rect 5632 1980 5684 2032
rect 1676 1955 1728 1964
rect 1676 1921 1685 1955
rect 1685 1921 1719 1955
rect 1719 1921 1728 1955
rect 1676 1912 1728 1921
rect 2136 1955 2188 1964
rect 2136 1921 2145 1955
rect 2145 1921 2179 1955
rect 2179 1921 2188 1955
rect 2136 1912 2188 1921
rect 2412 1955 2464 1964
rect 2044 1844 2096 1896
rect 2412 1921 2421 1955
rect 2421 1921 2455 1955
rect 2455 1921 2464 1955
rect 2412 1912 2464 1921
rect 6552 1955 6604 1964
rect 6552 1921 6561 1955
rect 6561 1921 6595 1955
rect 6595 1921 6604 1955
rect 6552 1912 6604 1921
rect 6644 1912 6696 1964
rect 7472 1912 7524 1964
rect 7656 1912 7708 1964
rect 8116 1980 8168 2032
rect 9220 1912 9272 1964
rect 10140 1980 10192 2032
rect 2688 1887 2740 1896
rect 2688 1853 2697 1887
rect 2697 1853 2731 1887
rect 2731 1853 2740 1887
rect 2688 1844 2740 1853
rect 6460 1887 6512 1896
rect 6460 1853 6469 1887
rect 6469 1853 6503 1887
rect 6503 1853 6512 1887
rect 6460 1844 6512 1853
rect 6736 1844 6788 1896
rect 4436 1708 4488 1760
rect 4620 1708 4672 1760
rect 7196 1844 7248 1896
rect 8668 1844 8720 1896
rect 10232 1955 10284 1964
rect 9312 1776 9364 1828
rect 10232 1921 10241 1955
rect 10241 1921 10275 1955
rect 10275 1921 10284 1955
rect 10232 1912 10284 1921
rect 10508 1955 10560 1964
rect 10508 1921 10517 1955
rect 10517 1921 10551 1955
rect 10551 1921 10560 1955
rect 10508 1912 10560 1921
rect 11060 1912 11112 1964
rect 11244 1955 11296 1964
rect 11244 1921 11253 1955
rect 11253 1921 11287 1955
rect 11287 1921 11296 1955
rect 11244 1912 11296 1921
rect 11520 1955 11572 1964
rect 11520 1921 11529 1955
rect 11529 1921 11563 1955
rect 11563 1921 11572 1955
rect 11520 1912 11572 1921
rect 12992 1844 13044 1896
rect 10140 1776 10192 1828
rect 8576 1708 8628 1760
rect 11980 1708 12032 1760
rect 4214 1606 4266 1658
rect 4278 1606 4330 1658
rect 4342 1606 4394 1658
rect 4406 1606 4458 1658
rect 4470 1606 4522 1658
rect 12214 1606 12266 1658
rect 12278 1606 12330 1658
rect 12342 1606 12394 1658
rect 12406 1606 12458 1658
rect 12470 1606 12522 1658
rect 3148 1504 3200 1556
rect 3976 1504 4028 1556
rect 3516 1479 3568 1488
rect 3516 1445 3525 1479
rect 3525 1445 3559 1479
rect 3559 1445 3568 1479
rect 3516 1436 3568 1445
rect 7196 1504 7248 1556
rect 7748 1504 7800 1556
rect 1400 1411 1452 1420
rect 1400 1377 1409 1411
rect 1409 1377 1443 1411
rect 1443 1377 1452 1411
rect 1400 1368 1452 1377
rect 2780 1368 2832 1420
rect 3976 1368 4028 1420
rect 4988 1411 5040 1420
rect 4988 1377 4997 1411
rect 4997 1377 5031 1411
rect 5031 1377 5040 1411
rect 4988 1368 5040 1377
rect 6460 1368 6512 1420
rect 2412 1300 2464 1352
rect 3424 1343 3476 1352
rect 3424 1309 3433 1343
rect 3433 1309 3467 1343
rect 3467 1309 3476 1343
rect 3424 1300 3476 1309
rect 3608 1343 3660 1352
rect 3608 1309 3617 1343
rect 3617 1309 3651 1343
rect 3651 1309 3660 1343
rect 3608 1300 3660 1309
rect 4160 1343 4212 1352
rect 4160 1309 4169 1343
rect 4169 1309 4203 1343
rect 4203 1309 4212 1343
rect 4712 1343 4764 1352
rect 4160 1300 4212 1309
rect 4712 1309 4721 1343
rect 4721 1309 4755 1343
rect 4755 1309 4764 1343
rect 4712 1300 4764 1309
rect 4620 1232 4672 1284
rect 5816 1300 5868 1352
rect 6644 1300 6696 1352
rect 7656 1368 7708 1420
rect 9772 1504 9824 1556
rect 10968 1504 11020 1556
rect 11428 1504 11480 1556
rect 12992 1547 13044 1556
rect 12992 1513 13001 1547
rect 13001 1513 13035 1547
rect 13035 1513 13044 1547
rect 12992 1504 13044 1513
rect 11888 1436 11940 1488
rect 9680 1411 9732 1420
rect 5448 1232 5500 1284
rect 7380 1232 7432 1284
rect 8116 1232 8168 1284
rect 9680 1377 9689 1411
rect 9689 1377 9723 1411
rect 9723 1377 9732 1411
rect 9680 1368 9732 1377
rect 11244 1368 11296 1420
rect 8760 1300 8812 1352
rect 9312 1343 9364 1352
rect 9312 1309 9321 1343
rect 9321 1309 9355 1343
rect 9355 1309 9364 1343
rect 9312 1300 9364 1309
rect 10140 1232 10192 1284
rect 13176 1343 13228 1352
rect 13176 1309 13185 1343
rect 13185 1309 13219 1343
rect 13219 1309 13228 1343
rect 13176 1300 13228 1309
rect 5908 1207 5960 1216
rect 5908 1173 5917 1207
rect 5917 1173 5951 1207
rect 5951 1173 5960 1207
rect 5908 1164 5960 1173
rect 6092 1207 6144 1216
rect 6092 1173 6101 1207
rect 6101 1173 6135 1207
rect 6135 1173 6144 1207
rect 6092 1164 6144 1173
rect 9220 1207 9272 1216
rect 9220 1173 9229 1207
rect 9229 1173 9263 1207
rect 9263 1173 9272 1207
rect 9220 1164 9272 1173
rect 11520 1207 11572 1216
rect 11520 1173 11529 1207
rect 11529 1173 11563 1207
rect 11563 1173 11572 1207
rect 11520 1164 11572 1173
rect 11980 1164 12032 1216
rect 8214 1062 8266 1114
rect 8278 1062 8330 1114
rect 8342 1062 8394 1114
rect 8406 1062 8458 1114
rect 8470 1062 8522 1114
rect 2964 960 3016 1012
rect 5908 960 5960 1012
rect 10232 960 10284 1012
rect 3424 892 3476 944
rect 11520 892 11572 944
rect 3608 824 3660 876
rect 6092 824 6144 876
<< metal2 >>
rect 570 14362 626 15000
rect 570 14334 888 14362
rect 570 14200 626 14334
rect 860 11898 888 14334
rect 1674 14200 1730 15000
rect 2870 14200 2926 15000
rect 3238 14512 3294 14521
rect 3238 14447 3294 14456
rect 1688 14090 1716 14200
rect 1688 14062 1808 14090
rect 2884 14074 2912 14200
rect 1674 13424 1730 13433
rect 1674 13359 1730 13368
rect 1688 13326 1716 13359
rect 1676 13320 1728 13326
rect 1676 13262 1728 13268
rect 1492 13252 1544 13258
rect 1492 13194 1544 13200
rect 1398 12608 1454 12617
rect 1398 12543 1454 12552
rect 848 11892 900 11898
rect 848 11834 900 11840
rect 1412 10656 1440 12543
rect 1504 11762 1532 13194
rect 1780 12986 1808 14062
rect 2872 14068 2924 14074
rect 2872 14010 2924 14016
rect 1950 13560 2006 13569
rect 1950 13495 2006 13504
rect 1860 13320 1912 13326
rect 1860 13262 1912 13268
rect 1768 12980 1820 12986
rect 1768 12922 1820 12928
rect 1872 12850 1900 13262
rect 1964 13258 1992 13495
rect 2872 13320 2924 13326
rect 2870 13288 2872 13297
rect 2924 13288 2926 13297
rect 1952 13252 2004 13258
rect 2870 13223 2926 13232
rect 3148 13252 3200 13258
rect 1952 13194 2004 13200
rect 1964 12889 1992 13194
rect 2044 13184 2096 13190
rect 2044 13126 2096 13132
rect 1950 12880 2006 12889
rect 1676 12844 1728 12850
rect 1676 12786 1728 12792
rect 1860 12844 1912 12850
rect 1950 12815 2006 12824
rect 1860 12786 1912 12792
rect 1492 11756 1544 11762
rect 1492 11698 1544 11704
rect 1504 11150 1532 11698
rect 1688 11642 1716 12786
rect 1768 12776 1820 12782
rect 1768 12718 1820 12724
rect 1780 12238 1808 12718
rect 1768 12232 1820 12238
rect 1768 12174 1820 12180
rect 1872 11830 1900 12786
rect 1860 11824 1912 11830
rect 1860 11766 1912 11772
rect 1688 11626 1808 11642
rect 1584 11620 1636 11626
rect 1688 11620 1820 11626
rect 1688 11614 1768 11620
rect 1584 11562 1636 11568
rect 1768 11562 1820 11568
rect 1492 11144 1544 11150
rect 1492 11086 1544 11092
rect 1492 11008 1544 11014
rect 1492 10950 1544 10956
rect 1504 10810 1532 10950
rect 1492 10804 1544 10810
rect 1492 10746 1544 10752
rect 1492 10668 1544 10674
rect 1412 10628 1492 10656
rect 1492 10610 1544 10616
rect 1400 9376 1452 9382
rect 1400 9318 1452 9324
rect 1412 8974 1440 9318
rect 1400 8968 1452 8974
rect 1504 8945 1532 10610
rect 1400 8910 1452 8916
rect 1490 8936 1546 8945
rect 1490 8871 1546 8880
rect 1400 7948 1452 7954
rect 1400 7890 1452 7896
rect 1412 5710 1440 7890
rect 1492 7744 1544 7750
rect 1492 7686 1544 7692
rect 1504 7478 1532 7686
rect 1492 7472 1544 7478
rect 1492 7414 1544 7420
rect 1596 6866 1624 11562
rect 1676 11552 1728 11558
rect 1676 11494 1728 11500
rect 1688 10062 1716 11494
rect 1780 11286 1808 11562
rect 1768 11280 1820 11286
rect 1768 11222 1820 11228
rect 1676 10056 1728 10062
rect 1676 9998 1728 10004
rect 1780 9874 1808 11222
rect 2056 11014 2084 13126
rect 2884 12730 2912 13223
rect 3148 13194 3200 13200
rect 3056 13184 3108 13190
rect 3056 13126 3108 13132
rect 3068 12986 3096 13126
rect 2964 12980 3016 12986
rect 2964 12922 3016 12928
rect 3056 12980 3108 12986
rect 3056 12922 3108 12928
rect 2700 12702 2912 12730
rect 2700 12238 2728 12702
rect 2976 12646 3004 12922
rect 2964 12640 3016 12646
rect 2964 12582 3016 12588
rect 3056 12300 3108 12306
rect 3056 12242 3108 12248
rect 2688 12232 2740 12238
rect 2688 12174 2740 12180
rect 2320 12164 2372 12170
rect 2320 12106 2372 12112
rect 2332 11150 2360 12106
rect 2504 12096 2556 12102
rect 2504 12038 2556 12044
rect 2780 12096 2832 12102
rect 2780 12038 2832 12044
rect 2410 11792 2466 11801
rect 2410 11727 2412 11736
rect 2464 11727 2466 11736
rect 2412 11698 2464 11704
rect 2320 11144 2372 11150
rect 2320 11086 2372 11092
rect 2044 11008 2096 11014
rect 2044 10950 2096 10956
rect 2332 10742 2360 11086
rect 2320 10736 2372 10742
rect 2320 10678 2372 10684
rect 2516 10674 2544 12038
rect 2792 11914 2820 12038
rect 2596 11892 2648 11898
rect 2596 11834 2648 11840
rect 2700 11886 2820 11914
rect 2608 11014 2636 11834
rect 2700 11642 2728 11886
rect 3068 11665 3096 12242
rect 3054 11656 3110 11665
rect 2700 11614 2820 11642
rect 2596 11008 2648 11014
rect 2596 10950 2648 10956
rect 2504 10668 2556 10674
rect 2504 10610 2556 10616
rect 2044 10600 2096 10606
rect 2044 10542 2096 10548
rect 2056 10062 2084 10542
rect 2516 10198 2544 10610
rect 2596 10600 2648 10606
rect 2596 10542 2648 10548
rect 2608 10266 2636 10542
rect 2596 10260 2648 10266
rect 2596 10202 2648 10208
rect 2504 10192 2556 10198
rect 2504 10134 2556 10140
rect 2044 10056 2096 10062
rect 2044 9998 2096 10004
rect 1688 9846 1808 9874
rect 1688 8498 1716 9846
rect 1860 9580 1912 9586
rect 1860 9522 1912 9528
rect 1872 8634 1900 9522
rect 2792 8922 2820 11614
rect 3054 11591 3110 11600
rect 2964 11552 3016 11558
rect 3016 11500 3096 11506
rect 2964 11494 3096 11500
rect 2976 11478 3096 11494
rect 2964 10124 3016 10130
rect 2964 10066 3016 10072
rect 2976 8974 3004 10066
rect 3068 10062 3096 11478
rect 3160 10849 3188 13194
rect 3252 11558 3280 14447
rect 3974 14362 4030 15000
rect 3608 14340 3660 14346
rect 3608 14282 3660 14288
rect 3896 14334 4030 14362
rect 3424 13932 3476 13938
rect 3424 13874 3476 13880
rect 3436 13326 3464 13874
rect 3620 13530 3648 14282
rect 3608 13524 3660 13530
rect 3608 13466 3660 13472
rect 3424 13320 3476 13326
rect 3424 13262 3476 13268
rect 3700 13320 3752 13326
rect 3700 13262 3752 13268
rect 3332 13252 3384 13258
rect 3332 13194 3384 13200
rect 3344 12442 3372 13194
rect 3516 13184 3568 13190
rect 3516 13126 3568 13132
rect 3528 12918 3556 13126
rect 3516 12912 3568 12918
rect 3516 12854 3568 12860
rect 3712 12850 3740 13262
rect 3896 12986 3924 14334
rect 3974 14200 4030 14334
rect 5170 14200 5226 15000
rect 6274 14200 6330 15000
rect 7470 14200 7526 15000
rect 8574 14200 8630 15000
rect 9770 14362 9826 15000
rect 10874 14362 10930 15000
rect 12070 14362 12126 15000
rect 9770 14334 9996 14362
rect 10796 14346 10930 14362
rect 9770 14200 9826 14334
rect 4214 13628 4522 13637
rect 4214 13626 4220 13628
rect 4276 13626 4300 13628
rect 4356 13626 4380 13628
rect 4436 13626 4460 13628
rect 4516 13626 4522 13628
rect 4276 13574 4278 13626
rect 4458 13574 4460 13626
rect 4214 13572 4220 13574
rect 4276 13572 4300 13574
rect 4356 13572 4380 13574
rect 4436 13572 4460 13574
rect 4516 13572 4522 13574
rect 4214 13563 4522 13572
rect 4068 13252 4120 13258
rect 4068 13194 4120 13200
rect 4896 13252 4948 13258
rect 4896 13194 4948 13200
rect 3884 12980 3936 12986
rect 3884 12922 3936 12928
rect 3700 12844 3752 12850
rect 3700 12786 3752 12792
rect 3332 12436 3384 12442
rect 3384 12406 3556 12434
rect 3332 12378 3384 12384
rect 3332 12164 3384 12170
rect 3332 12106 3384 12112
rect 3240 11552 3292 11558
rect 3240 11494 3292 11500
rect 3240 11076 3292 11082
rect 3240 11018 3292 11024
rect 3146 10840 3202 10849
rect 3146 10775 3202 10784
rect 3252 10674 3280 11018
rect 3240 10668 3292 10674
rect 3240 10610 3292 10616
rect 3056 10056 3108 10062
rect 3056 9998 3108 10004
rect 3068 9654 3096 9998
rect 3148 9988 3200 9994
rect 3148 9930 3200 9936
rect 3056 9648 3108 9654
rect 3056 9590 3108 9596
rect 3160 9586 3188 9930
rect 3148 9580 3200 9586
rect 3148 9522 3200 9528
rect 2700 8894 2820 8922
rect 2964 8968 3016 8974
rect 2964 8910 3016 8916
rect 2700 8634 2728 8894
rect 2780 8832 2832 8838
rect 2780 8774 2832 8780
rect 1860 8628 1912 8634
rect 1860 8570 1912 8576
rect 2688 8628 2740 8634
rect 2688 8570 2740 8576
rect 2596 8560 2648 8566
rect 2596 8502 2648 8508
rect 1676 8492 1728 8498
rect 1676 8434 1728 8440
rect 1768 8492 1820 8498
rect 1768 8434 1820 8440
rect 2504 8492 2556 8498
rect 2504 8434 2556 8440
rect 1676 7880 1728 7886
rect 1676 7822 1728 7828
rect 1584 6860 1636 6866
rect 1584 6802 1636 6808
rect 1492 6792 1544 6798
rect 1492 6734 1544 6740
rect 1504 5914 1532 6734
rect 1492 5908 1544 5914
rect 1492 5850 1544 5856
rect 1400 5704 1452 5710
rect 1400 5646 1452 5652
rect 1412 5137 1440 5646
rect 1398 5128 1454 5137
rect 1398 5063 1454 5072
rect 1412 3738 1440 5063
rect 1492 3936 1544 3942
rect 1492 3878 1544 3884
rect 1400 3732 1452 3738
rect 1400 3674 1452 3680
rect 1504 3670 1532 3878
rect 1688 3738 1716 7822
rect 1780 7818 1808 8434
rect 1952 8424 2004 8430
rect 1952 8366 2004 8372
rect 1964 7886 1992 8366
rect 2412 8356 2464 8362
rect 2412 8298 2464 8304
rect 2044 8084 2096 8090
rect 2044 8026 2096 8032
rect 2056 7886 2084 8026
rect 2424 7886 2452 8298
rect 2516 7954 2544 8434
rect 2608 8090 2636 8502
rect 2596 8084 2648 8090
rect 2596 8026 2648 8032
rect 2504 7948 2556 7954
rect 2504 7890 2556 7896
rect 1952 7880 2004 7886
rect 1952 7822 2004 7828
rect 2044 7880 2096 7886
rect 2044 7822 2096 7828
rect 2412 7880 2464 7886
rect 2412 7822 2464 7828
rect 2596 7880 2648 7886
rect 2596 7822 2648 7828
rect 1768 7812 1820 7818
rect 1768 7754 1820 7760
rect 1780 7274 1808 7754
rect 1768 7268 1820 7274
rect 1768 7210 1820 7216
rect 1964 7002 1992 7822
rect 1952 6996 2004 7002
rect 1952 6938 2004 6944
rect 2056 6730 2084 7822
rect 2608 7410 2636 7822
rect 2136 7404 2188 7410
rect 2136 7346 2188 7352
rect 2596 7404 2648 7410
rect 2596 7346 2648 7352
rect 2148 6780 2176 7346
rect 2792 7290 2820 8774
rect 2872 8628 2924 8634
rect 2872 8570 2924 8576
rect 2884 7478 2912 8570
rect 2976 7993 3004 8910
rect 2962 7984 3018 7993
rect 2962 7919 3018 7928
rect 3056 7880 3108 7886
rect 3056 7822 3108 7828
rect 2872 7472 2924 7478
rect 2872 7414 2924 7420
rect 2964 7472 3016 7478
rect 2964 7414 3016 7420
rect 2320 7268 2372 7274
rect 2320 7210 2372 7216
rect 2700 7262 2820 7290
rect 2332 6798 2360 7210
rect 2228 6792 2280 6798
rect 2148 6752 2228 6780
rect 2228 6734 2280 6740
rect 2320 6792 2372 6798
rect 2320 6734 2372 6740
rect 2044 6724 2096 6730
rect 2044 6666 2096 6672
rect 2240 6458 2268 6734
rect 2228 6452 2280 6458
rect 2228 6394 2280 6400
rect 2044 6316 2096 6322
rect 2044 6258 2096 6264
rect 2136 6316 2188 6322
rect 2136 6258 2188 6264
rect 2056 5914 2084 6258
rect 2044 5908 2096 5914
rect 2044 5850 2096 5856
rect 2148 5846 2176 6258
rect 2136 5840 2188 5846
rect 2136 5782 2188 5788
rect 1768 5024 1820 5030
rect 1768 4966 1820 4972
rect 1860 5024 1912 5030
rect 1860 4966 1912 4972
rect 1780 4690 1808 4966
rect 1768 4684 1820 4690
rect 1768 4626 1820 4632
rect 1768 4548 1820 4554
rect 1872 4536 1900 4966
rect 1820 4508 1900 4536
rect 1768 4490 1820 4496
rect 1676 3732 1728 3738
rect 1676 3674 1728 3680
rect 1492 3664 1544 3670
rect 1492 3606 1544 3612
rect 1780 2990 1808 4490
rect 1952 4140 2004 4146
rect 1952 4082 2004 4088
rect 2228 4140 2280 4146
rect 2228 4082 2280 4088
rect 1860 4004 1912 4010
rect 1860 3946 1912 3952
rect 1872 3534 1900 3946
rect 1860 3528 1912 3534
rect 1860 3470 1912 3476
rect 1964 3398 1992 4082
rect 2044 4072 2096 4078
rect 2044 4014 2096 4020
rect 2136 4072 2188 4078
rect 2136 4014 2188 4020
rect 2056 3534 2084 4014
rect 2044 3528 2096 3534
rect 2044 3470 2096 3476
rect 1952 3392 2004 3398
rect 1952 3334 2004 3340
rect 2056 3194 2084 3470
rect 2148 3466 2176 4014
rect 2136 3460 2188 3466
rect 2136 3402 2188 3408
rect 2044 3188 2096 3194
rect 2044 3130 2096 3136
rect 1768 2984 1820 2990
rect 1768 2926 1820 2932
rect 2148 2650 2176 3402
rect 2240 2650 2268 4082
rect 2332 3942 2360 6734
rect 2594 6216 2650 6225
rect 2594 6151 2650 6160
rect 2608 5710 2636 6151
rect 2700 6118 2728 7262
rect 2780 7200 2832 7206
rect 2780 7142 2832 7148
rect 2792 6798 2820 7142
rect 2870 7032 2926 7041
rect 2870 6967 2926 6976
rect 2780 6792 2832 6798
rect 2780 6734 2832 6740
rect 2780 6316 2832 6322
rect 2780 6258 2832 6264
rect 2688 6112 2740 6118
rect 2688 6054 2740 6060
rect 2792 5914 2820 6258
rect 2780 5908 2832 5914
rect 2780 5850 2832 5856
rect 2884 5794 2912 6967
rect 2976 6866 3004 7414
rect 2964 6860 3016 6866
rect 2964 6802 3016 6808
rect 2962 6080 3018 6089
rect 2962 6015 3018 6024
rect 2700 5766 2912 5794
rect 2596 5704 2648 5710
rect 2596 5646 2648 5652
rect 2504 5636 2556 5642
rect 2504 5578 2556 5584
rect 2320 3936 2372 3942
rect 2320 3878 2372 3884
rect 2320 3460 2372 3466
rect 2320 3402 2372 3408
rect 2332 3058 2360 3402
rect 2320 3052 2372 3058
rect 2320 2994 2372 3000
rect 2412 2984 2464 2990
rect 2412 2926 2464 2932
rect 2136 2644 2188 2650
rect 2136 2586 2188 2592
rect 2228 2644 2280 2650
rect 2228 2586 2280 2592
rect 2044 2576 2096 2582
rect 2044 2518 2096 2524
rect 2318 2544 2374 2553
rect 1676 2440 1728 2446
rect 1674 2408 1676 2417
rect 1952 2440 2004 2446
rect 1728 2408 1730 2417
rect 1952 2382 2004 2388
rect 1674 2343 1730 2352
rect 1676 2304 1728 2310
rect 1676 2246 1728 2252
rect 1688 2009 1716 2246
rect 1964 2038 1992 2382
rect 1952 2032 2004 2038
rect 1674 2000 1730 2009
rect 1952 1974 2004 1980
rect 1674 1935 1676 1944
rect 1728 1935 1730 1944
rect 1676 1906 1728 1912
rect 2056 1902 2084 2518
rect 2318 2479 2320 2488
rect 2372 2479 2374 2488
rect 2320 2450 2372 2456
rect 2136 2304 2188 2310
rect 2136 2246 2188 2252
rect 2148 1970 2176 2246
rect 2424 1970 2452 2926
rect 2516 2774 2544 5578
rect 2608 5302 2636 5646
rect 2596 5296 2648 5302
rect 2596 5238 2648 5244
rect 2700 4706 2728 5766
rect 2780 5704 2832 5710
rect 2780 5646 2832 5652
rect 2792 5302 2820 5646
rect 2780 5296 2832 5302
rect 2780 5238 2832 5244
rect 2870 5264 2926 5273
rect 2792 4826 2820 5238
rect 2870 5199 2926 5208
rect 2884 5166 2912 5199
rect 2872 5160 2924 5166
rect 2872 5102 2924 5108
rect 2976 4842 3004 6015
rect 2780 4820 2832 4826
rect 2780 4762 2832 4768
rect 2884 4814 3004 4842
rect 2884 4758 2912 4814
rect 2872 4752 2924 4758
rect 2700 4678 2820 4706
rect 3068 4706 3096 7822
rect 3148 7472 3200 7478
rect 3148 7414 3200 7420
rect 3160 6798 3188 7414
rect 3148 6792 3200 6798
rect 3148 6734 3200 6740
rect 3252 6662 3280 10610
rect 3344 8362 3372 12106
rect 3424 11756 3476 11762
rect 3424 11698 3476 11704
rect 3332 8356 3384 8362
rect 3332 8298 3384 8304
rect 3240 6656 3292 6662
rect 3240 6598 3292 6604
rect 3436 6474 3464 11698
rect 3528 11082 3556 12406
rect 3608 12368 3660 12374
rect 3608 12310 3660 12316
rect 3620 11354 3648 12310
rect 3712 11830 3740 12786
rect 3792 12776 3844 12782
rect 3792 12718 3844 12724
rect 3804 12170 3832 12718
rect 3792 12164 3844 12170
rect 3792 12106 3844 12112
rect 3700 11824 3752 11830
rect 3700 11766 3752 11772
rect 3792 11552 3844 11558
rect 3792 11494 3844 11500
rect 3608 11348 3660 11354
rect 3608 11290 3660 11296
rect 3608 11212 3660 11218
rect 3608 11154 3660 11160
rect 3516 11076 3568 11082
rect 3516 11018 3568 11024
rect 3620 10674 3648 11154
rect 3608 10668 3660 10674
rect 3608 10610 3660 10616
rect 3700 10532 3752 10538
rect 3700 10474 3752 10480
rect 3712 10130 3740 10474
rect 3700 10124 3752 10130
rect 3700 10066 3752 10072
rect 3712 9654 3740 10066
rect 3700 9648 3752 9654
rect 3700 9590 3752 9596
rect 3608 9580 3660 9586
rect 3608 9522 3660 9528
rect 3516 9376 3568 9382
rect 3516 9318 3568 9324
rect 3528 8566 3556 9318
rect 3620 8566 3648 9522
rect 3700 9512 3752 9518
rect 3700 9454 3752 9460
rect 3516 8560 3568 8566
rect 3516 8502 3568 8508
rect 3608 8560 3660 8566
rect 3608 8502 3660 8508
rect 3712 8498 3740 9454
rect 3804 9217 3832 11494
rect 3896 10062 3924 12922
rect 4080 12850 4108 13194
rect 4620 13184 4672 13190
rect 4620 13126 4672 13132
rect 4068 12844 4120 12850
rect 4068 12786 4120 12792
rect 3976 12708 4028 12714
rect 3976 12650 4028 12656
rect 3988 12073 4016 12650
rect 4214 12540 4522 12549
rect 4214 12538 4220 12540
rect 4276 12538 4300 12540
rect 4356 12538 4380 12540
rect 4436 12538 4460 12540
rect 4516 12538 4522 12540
rect 4276 12486 4278 12538
rect 4458 12486 4460 12538
rect 4214 12484 4220 12486
rect 4276 12484 4300 12486
rect 4356 12484 4380 12486
rect 4436 12484 4460 12486
rect 4516 12484 4522 12486
rect 4214 12475 4522 12484
rect 4160 12436 4212 12442
rect 4160 12378 4212 12384
rect 4068 12164 4120 12170
rect 4068 12106 4120 12112
rect 3974 12064 4030 12073
rect 3974 11999 4030 12008
rect 3976 11688 4028 11694
rect 3976 11630 4028 11636
rect 3988 11150 4016 11630
rect 3976 11144 4028 11150
rect 3976 11086 4028 11092
rect 3988 10742 4016 11086
rect 3976 10736 4028 10742
rect 3976 10678 4028 10684
rect 3976 10464 4028 10470
rect 3976 10406 4028 10412
rect 3884 10056 3936 10062
rect 3884 9998 3936 10004
rect 3988 9761 4016 10406
rect 3974 9752 4030 9761
rect 3974 9687 4030 9696
rect 3884 9376 3936 9382
rect 3884 9318 3936 9324
rect 3790 9208 3846 9217
rect 3790 9143 3846 9152
rect 3792 9036 3844 9042
rect 3792 8978 3844 8984
rect 3700 8492 3752 8498
rect 3700 8434 3752 8440
rect 3700 8356 3752 8362
rect 3700 8298 3752 8304
rect 3606 7984 3662 7993
rect 3606 7919 3662 7928
rect 3516 7200 3568 7206
rect 3516 7142 3568 7148
rect 3528 6866 3556 7142
rect 3516 6860 3568 6866
rect 3516 6802 3568 6808
rect 3252 6446 3464 6474
rect 3528 6458 3556 6802
rect 3516 6452 3568 6458
rect 3148 6248 3200 6254
rect 3148 6190 3200 6196
rect 3160 5710 3188 6190
rect 3148 5704 3200 5710
rect 3148 5646 3200 5652
rect 2872 4694 2924 4700
rect 2792 4486 2820 4678
rect 2976 4678 3096 4706
rect 2780 4480 2832 4486
rect 2780 4422 2832 4428
rect 2780 4140 2832 4146
rect 2780 4082 2832 4088
rect 2596 3936 2648 3942
rect 2596 3878 2648 3884
rect 2608 3194 2636 3878
rect 2688 3664 2740 3670
rect 2688 3606 2740 3612
rect 2596 3188 2648 3194
rect 2596 3130 2648 3136
rect 2700 2990 2728 3606
rect 2792 3602 2820 4082
rect 2976 4010 3004 4678
rect 3056 4548 3108 4554
rect 3056 4490 3108 4496
rect 3068 4282 3096 4490
rect 3056 4276 3108 4282
rect 3056 4218 3108 4224
rect 3056 4072 3108 4078
rect 3056 4014 3108 4020
rect 2964 4004 3016 4010
rect 2964 3946 3016 3952
rect 2780 3596 2832 3602
rect 2780 3538 2832 3544
rect 2792 3126 2820 3538
rect 3068 3233 3096 4014
rect 3160 3534 3188 5646
rect 3252 4706 3280 6446
rect 3516 6394 3568 6400
rect 3332 6316 3384 6322
rect 3332 6258 3384 6264
rect 3344 5642 3372 6258
rect 3516 6248 3568 6254
rect 3436 6208 3516 6236
rect 3332 5636 3384 5642
rect 3332 5578 3384 5584
rect 3436 5234 3464 6208
rect 3516 6190 3568 6196
rect 3620 5914 3648 7919
rect 3712 7886 3740 8298
rect 3700 7880 3752 7886
rect 3700 7822 3752 7828
rect 3712 7546 3740 7822
rect 3700 7540 3752 7546
rect 3700 7482 3752 7488
rect 3804 7426 3832 8978
rect 3896 8974 3924 9318
rect 3884 8968 3936 8974
rect 3884 8910 3936 8916
rect 3896 8809 3924 8910
rect 3976 8832 4028 8838
rect 3882 8800 3938 8809
rect 3976 8774 4028 8780
rect 3882 8735 3938 8744
rect 3988 8498 4016 8774
rect 3976 8492 4028 8498
rect 3976 8434 4028 8440
rect 3988 7886 4016 8434
rect 3976 7880 4028 7886
rect 3976 7822 4028 7828
rect 3712 7398 3832 7426
rect 3712 6474 3740 7398
rect 3792 7336 3844 7342
rect 3792 7278 3844 7284
rect 3804 6934 3832 7278
rect 3792 6928 3844 6934
rect 3792 6870 3844 6876
rect 3712 6446 3832 6474
rect 3700 6316 3752 6322
rect 3700 6258 3752 6264
rect 3608 5908 3660 5914
rect 3608 5850 3660 5856
rect 3712 5710 3740 6258
rect 3700 5704 3752 5710
rect 3700 5646 3752 5652
rect 3516 5636 3568 5642
rect 3516 5578 3568 5584
rect 3332 5228 3384 5234
rect 3332 5170 3384 5176
rect 3424 5228 3476 5234
rect 3424 5170 3476 5176
rect 3344 4826 3372 5170
rect 3424 5024 3476 5030
rect 3424 4966 3476 4972
rect 3332 4820 3384 4826
rect 3332 4762 3384 4768
rect 3252 4678 3372 4706
rect 3240 4480 3292 4486
rect 3240 4422 3292 4428
rect 3148 3528 3200 3534
rect 3148 3470 3200 3476
rect 3054 3224 3110 3233
rect 3054 3159 3110 3168
rect 2780 3120 2832 3126
rect 2780 3062 2832 3068
rect 2688 2984 2740 2990
rect 2688 2926 2740 2932
rect 2516 2746 2636 2774
rect 2136 1964 2188 1970
rect 2136 1906 2188 1912
rect 2412 1964 2464 1970
rect 2412 1906 2464 1912
rect 2044 1896 2096 1902
rect 2044 1838 2096 1844
rect 1400 1420 1452 1426
rect 1400 1362 1452 1368
rect 1412 513 1440 1362
rect 2424 1358 2452 1906
rect 2608 1884 2636 2746
rect 3160 2446 3188 3470
rect 2964 2440 3016 2446
rect 2964 2382 3016 2388
rect 3148 2440 3200 2446
rect 3148 2382 3200 2388
rect 2780 2372 2832 2378
rect 2780 2314 2832 2320
rect 2792 2281 2820 2314
rect 2778 2272 2834 2281
rect 2778 2207 2834 2216
rect 2688 1896 2740 1902
rect 2608 1856 2688 1884
rect 2688 1838 2740 1844
rect 2792 1426 2820 2207
rect 2780 1420 2832 1426
rect 2780 1362 2832 1368
rect 2412 1352 2464 1358
rect 2412 1294 2464 1300
rect 2976 1018 3004 2382
rect 3160 1562 3188 2382
rect 3148 1556 3200 1562
rect 3148 1498 3200 1504
rect 3252 1340 3280 4422
rect 3344 3738 3372 4678
rect 3436 4282 3464 4966
rect 3424 4276 3476 4282
rect 3424 4218 3476 4224
rect 3424 4140 3476 4146
rect 3424 4082 3476 4088
rect 3332 3732 3384 3738
rect 3332 3674 3384 3680
rect 3436 3670 3464 4082
rect 3424 3664 3476 3670
rect 3424 3606 3476 3612
rect 3332 3392 3384 3398
rect 3436 3380 3464 3606
rect 3528 3534 3556 5578
rect 3608 5568 3660 5574
rect 3608 5510 3660 5516
rect 3516 3528 3568 3534
rect 3516 3470 3568 3476
rect 3436 3352 3556 3380
rect 3332 3334 3384 3340
rect 3344 3194 3372 3334
rect 3332 3188 3384 3194
rect 3332 3130 3384 3136
rect 3424 3120 3476 3126
rect 3424 3062 3476 3068
rect 3436 2650 3464 3062
rect 3424 2644 3476 2650
rect 3424 2586 3476 2592
rect 3528 1494 3556 3352
rect 3620 2650 3648 5510
rect 3712 4146 3740 5646
rect 3700 4140 3752 4146
rect 3700 4082 3752 4088
rect 3700 3392 3752 3398
rect 3700 3334 3752 3340
rect 3608 2644 3660 2650
rect 3608 2586 3660 2592
rect 3712 2514 3740 3334
rect 3804 2774 3832 6446
rect 3884 6316 3936 6322
rect 3884 6258 3936 6264
rect 3896 4758 3924 6258
rect 3988 6089 4016 7822
rect 4080 7750 4108 12106
rect 4172 11898 4200 12378
rect 4528 12164 4580 12170
rect 4528 12106 4580 12112
rect 4160 11892 4212 11898
rect 4160 11834 4212 11840
rect 4540 11665 4568 12106
rect 4526 11656 4582 11665
rect 4632 11626 4660 13126
rect 4804 12232 4856 12238
rect 4804 12174 4856 12180
rect 4712 11688 4764 11694
rect 4712 11630 4764 11636
rect 4526 11591 4582 11600
rect 4620 11620 4672 11626
rect 4620 11562 4672 11568
rect 4214 11452 4522 11461
rect 4214 11450 4220 11452
rect 4276 11450 4300 11452
rect 4356 11450 4380 11452
rect 4436 11450 4460 11452
rect 4516 11450 4522 11452
rect 4276 11398 4278 11450
rect 4458 11398 4460 11450
rect 4214 11396 4220 11398
rect 4276 11396 4300 11398
rect 4356 11396 4380 11398
rect 4436 11396 4460 11398
rect 4516 11396 4522 11398
rect 4214 11387 4522 11396
rect 4160 11076 4212 11082
rect 4160 11018 4212 11024
rect 4172 10674 4200 11018
rect 4252 11008 4304 11014
rect 4252 10950 4304 10956
rect 4264 10742 4292 10950
rect 4632 10742 4660 11562
rect 4252 10736 4304 10742
rect 4252 10678 4304 10684
rect 4620 10736 4672 10742
rect 4620 10678 4672 10684
rect 4160 10668 4212 10674
rect 4160 10610 4212 10616
rect 4344 10668 4396 10674
rect 4344 10610 4396 10616
rect 4356 10470 4384 10610
rect 4344 10464 4396 10470
rect 4344 10406 4396 10412
rect 4214 10364 4522 10373
rect 4214 10362 4220 10364
rect 4276 10362 4300 10364
rect 4356 10362 4380 10364
rect 4436 10362 4460 10364
rect 4516 10362 4522 10364
rect 4276 10310 4278 10362
rect 4458 10310 4460 10362
rect 4214 10308 4220 10310
rect 4276 10308 4300 10310
rect 4356 10308 4380 10310
rect 4436 10308 4460 10310
rect 4516 10308 4522 10310
rect 4214 10299 4522 10308
rect 4724 10266 4752 11630
rect 4816 11354 4844 12174
rect 4804 11348 4856 11354
rect 4804 11290 4856 11296
rect 4802 11248 4858 11257
rect 4802 11183 4858 11192
rect 4816 10266 4844 11183
rect 4712 10260 4764 10266
rect 4712 10202 4764 10208
rect 4804 10260 4856 10266
rect 4804 10202 4856 10208
rect 4528 10056 4580 10062
rect 4804 10056 4856 10062
rect 4528 9998 4580 10004
rect 4710 10024 4766 10033
rect 4540 9382 4568 9998
rect 4804 9998 4856 10004
rect 4710 9959 4766 9968
rect 4724 9926 4752 9959
rect 4712 9920 4764 9926
rect 4712 9862 4764 9868
rect 4528 9376 4580 9382
rect 4528 9318 4580 9324
rect 4214 9276 4522 9285
rect 4214 9274 4220 9276
rect 4276 9274 4300 9276
rect 4356 9274 4380 9276
rect 4436 9274 4460 9276
rect 4516 9274 4522 9276
rect 4276 9222 4278 9274
rect 4458 9222 4460 9274
rect 4214 9220 4220 9222
rect 4276 9220 4300 9222
rect 4356 9220 4380 9222
rect 4436 9220 4460 9222
rect 4516 9220 4522 9222
rect 4214 9211 4522 9220
rect 4724 9042 4752 9862
rect 4816 9586 4844 9998
rect 4804 9580 4856 9586
rect 4804 9522 4856 9528
rect 4816 9110 4844 9522
rect 4804 9104 4856 9110
rect 4804 9046 4856 9052
rect 4712 9036 4764 9042
rect 4712 8978 4764 8984
rect 4528 8492 4580 8498
rect 4804 8492 4856 8498
rect 4580 8452 4660 8480
rect 4528 8434 4580 8440
rect 4214 8188 4522 8197
rect 4214 8186 4220 8188
rect 4276 8186 4300 8188
rect 4356 8186 4380 8188
rect 4436 8186 4460 8188
rect 4516 8186 4522 8188
rect 4276 8134 4278 8186
rect 4458 8134 4460 8186
rect 4214 8132 4220 8134
rect 4276 8132 4300 8134
rect 4356 8132 4380 8134
rect 4436 8132 4460 8134
rect 4516 8132 4522 8134
rect 4214 8123 4522 8132
rect 4632 7954 4660 8452
rect 4804 8434 4856 8440
rect 4712 8424 4764 8430
rect 4712 8366 4764 8372
rect 4620 7948 4672 7954
rect 4620 7890 4672 7896
rect 4252 7880 4304 7886
rect 4252 7822 4304 7828
rect 4068 7744 4120 7750
rect 4068 7686 4120 7692
rect 4160 7744 4212 7750
rect 4160 7686 4212 7692
rect 4172 7274 4200 7686
rect 4264 7274 4292 7822
rect 4632 7546 4660 7890
rect 4724 7886 4752 8366
rect 4816 7954 4844 8434
rect 4908 8090 4936 13194
rect 5080 13184 5132 13190
rect 5080 13126 5132 13132
rect 4988 12980 5040 12986
rect 4988 12922 5040 12928
rect 5000 11694 5028 12922
rect 5092 11830 5120 13126
rect 5184 12374 5212 14200
rect 5356 13864 5408 13870
rect 5356 13806 5408 13812
rect 5368 13394 5396 13806
rect 5540 13796 5592 13802
rect 5540 13738 5592 13744
rect 5552 13462 5580 13738
rect 6092 13728 6144 13734
rect 6092 13670 6144 13676
rect 6104 13530 6132 13670
rect 6092 13524 6144 13530
rect 6092 13466 6144 13472
rect 5540 13456 5592 13462
rect 5540 13398 5592 13404
rect 5356 13388 5408 13394
rect 5356 13330 5408 13336
rect 5264 13252 5316 13258
rect 5264 13194 5316 13200
rect 5172 12368 5224 12374
rect 5172 12310 5224 12316
rect 5184 12170 5212 12310
rect 5172 12164 5224 12170
rect 5172 12106 5224 12112
rect 5276 11898 5304 13194
rect 5368 12918 5396 13330
rect 5632 13320 5684 13326
rect 5632 13262 5684 13268
rect 5644 12918 5672 13262
rect 5816 13252 5868 13258
rect 5816 13194 5868 13200
rect 5356 12912 5408 12918
rect 5356 12854 5408 12860
rect 5632 12912 5684 12918
rect 5632 12854 5684 12860
rect 5356 12436 5408 12442
rect 5356 12378 5408 12384
rect 5264 11892 5316 11898
rect 5264 11834 5316 11840
rect 5080 11824 5132 11830
rect 5080 11766 5132 11772
rect 5172 11824 5224 11830
rect 5172 11766 5224 11772
rect 4988 11688 5040 11694
rect 4988 11630 5040 11636
rect 5000 10674 5028 11630
rect 5080 11280 5132 11286
rect 5184 11268 5212 11766
rect 5276 11286 5304 11834
rect 5368 11642 5396 12378
rect 5644 12238 5672 12854
rect 5828 12374 5856 13194
rect 5908 12844 5960 12850
rect 5908 12786 5960 12792
rect 6092 12844 6144 12850
rect 6092 12786 6144 12792
rect 5920 12442 5948 12786
rect 5908 12436 5960 12442
rect 5908 12378 5960 12384
rect 6000 12436 6052 12442
rect 6104 12434 6132 12786
rect 6104 12406 6224 12434
rect 6000 12378 6052 12384
rect 5816 12368 5868 12374
rect 5816 12310 5868 12316
rect 5632 12232 5684 12238
rect 5632 12174 5684 12180
rect 5540 11756 5592 11762
rect 5540 11698 5592 11704
rect 5368 11614 5488 11642
rect 5356 11552 5408 11558
rect 5356 11494 5408 11500
rect 5132 11240 5212 11268
rect 5264 11280 5316 11286
rect 5080 11222 5132 11228
rect 5264 11222 5316 11228
rect 5368 11150 5396 11494
rect 5172 11144 5224 11150
rect 5172 11086 5224 11092
rect 5356 11144 5408 11150
rect 5356 11086 5408 11092
rect 4988 10668 5040 10674
rect 4988 10610 5040 10616
rect 4988 10260 5040 10266
rect 4988 10202 5040 10208
rect 5000 9382 5028 10202
rect 5080 9988 5132 9994
rect 5080 9930 5132 9936
rect 4988 9376 5040 9382
rect 4988 9318 5040 9324
rect 5000 8906 5028 9318
rect 4988 8900 5040 8906
rect 4988 8842 5040 8848
rect 5092 8673 5120 9930
rect 5078 8664 5134 8673
rect 5078 8599 5134 8608
rect 5080 8492 5132 8498
rect 5080 8434 5132 8440
rect 4896 8084 4948 8090
rect 4896 8026 4948 8032
rect 4804 7948 4856 7954
rect 4804 7890 4856 7896
rect 5092 7886 5120 8434
rect 5184 8129 5212 11086
rect 5368 10674 5396 11086
rect 5460 11014 5488 11614
rect 5448 11008 5500 11014
rect 5448 10950 5500 10956
rect 5460 10674 5488 10950
rect 5356 10668 5408 10674
rect 5356 10610 5408 10616
rect 5448 10668 5500 10674
rect 5448 10610 5500 10616
rect 5264 10464 5316 10470
rect 5264 10406 5316 10412
rect 5170 8120 5226 8129
rect 5170 8055 5226 8064
rect 5172 7948 5224 7954
rect 5172 7890 5224 7896
rect 4712 7880 4764 7886
rect 4712 7822 4764 7828
rect 5080 7880 5132 7886
rect 5080 7822 5132 7828
rect 4896 7812 4948 7818
rect 4896 7754 4948 7760
rect 4620 7540 4672 7546
rect 4620 7482 4672 7488
rect 4712 7540 4764 7546
rect 4712 7482 4764 7488
rect 4724 7410 4752 7482
rect 4908 7478 4936 7754
rect 4896 7472 4948 7478
rect 4896 7414 4948 7420
rect 4712 7404 4764 7410
rect 4764 7364 4844 7392
rect 4712 7346 4764 7352
rect 4160 7268 4212 7274
rect 4160 7210 4212 7216
rect 4252 7268 4304 7274
rect 4252 7210 4304 7216
rect 4620 7200 4672 7206
rect 4620 7142 4672 7148
rect 4214 7100 4522 7109
rect 4214 7098 4220 7100
rect 4276 7098 4300 7100
rect 4356 7098 4380 7100
rect 4436 7098 4460 7100
rect 4516 7098 4522 7100
rect 4276 7046 4278 7098
rect 4458 7046 4460 7098
rect 4214 7044 4220 7046
rect 4276 7044 4300 7046
rect 4356 7044 4380 7046
rect 4436 7044 4460 7046
rect 4516 7044 4522 7046
rect 4214 7035 4522 7044
rect 4632 6730 4660 7142
rect 4712 6792 4764 6798
rect 4712 6734 4764 6740
rect 4620 6724 4672 6730
rect 4620 6666 4672 6672
rect 4068 6656 4120 6662
rect 4068 6598 4120 6604
rect 4160 6656 4212 6662
rect 4160 6598 4212 6604
rect 4080 6390 4108 6598
rect 4172 6458 4200 6598
rect 4160 6452 4212 6458
rect 4160 6394 4212 6400
rect 4068 6384 4120 6390
rect 4068 6326 4120 6332
rect 4252 6316 4304 6322
rect 4252 6258 4304 6264
rect 4160 6248 4212 6254
rect 4264 6225 4292 6258
rect 4160 6190 4212 6196
rect 4250 6216 4306 6225
rect 4172 6118 4200 6190
rect 4724 6186 4752 6734
rect 4250 6151 4306 6160
rect 4712 6180 4764 6186
rect 4712 6122 4764 6128
rect 4068 6112 4120 6118
rect 3974 6080 4030 6089
rect 4068 6054 4120 6060
rect 4160 6112 4212 6118
rect 4160 6054 4212 6060
rect 3974 6015 4030 6024
rect 4080 5710 4108 6054
rect 4214 6012 4522 6021
rect 4214 6010 4220 6012
rect 4276 6010 4300 6012
rect 4356 6010 4380 6012
rect 4436 6010 4460 6012
rect 4516 6010 4522 6012
rect 4276 5958 4278 6010
rect 4458 5958 4460 6010
rect 4214 5956 4220 5958
rect 4276 5956 4300 5958
rect 4356 5956 4380 5958
rect 4436 5956 4460 5958
rect 4516 5956 4522 5958
rect 4214 5947 4522 5956
rect 4724 5846 4752 6122
rect 4712 5840 4764 5846
rect 4712 5782 4764 5788
rect 4816 5778 4844 7364
rect 4896 7336 4948 7342
rect 4896 7278 4948 7284
rect 4908 6798 4936 7278
rect 4896 6792 4948 6798
rect 4896 6734 4948 6740
rect 4908 5846 4936 6734
rect 5092 6390 5120 7822
rect 5080 6384 5132 6390
rect 5080 6326 5132 6332
rect 4988 6248 5040 6254
rect 4988 6190 5040 6196
rect 4896 5840 4948 5846
rect 4896 5782 4948 5788
rect 4804 5772 4856 5778
rect 4804 5714 4856 5720
rect 4068 5704 4120 5710
rect 3988 5664 4068 5692
rect 3884 4752 3936 4758
rect 3884 4694 3936 4700
rect 3988 4264 4016 5664
rect 4068 5646 4120 5652
rect 4252 5568 4304 5574
rect 4252 5510 4304 5516
rect 4264 5302 4292 5510
rect 4816 5370 4844 5714
rect 4804 5364 4856 5370
rect 4540 5324 4752 5352
rect 4252 5296 4304 5302
rect 4252 5238 4304 5244
rect 4540 5166 4568 5324
rect 4618 5264 4674 5273
rect 4618 5199 4674 5208
rect 4528 5160 4580 5166
rect 4066 5128 4122 5137
rect 4122 5086 4200 5114
rect 4528 5102 4580 5108
rect 4066 5063 4122 5072
rect 4172 5030 4200 5086
rect 4160 5024 4212 5030
rect 4160 4966 4212 4972
rect 4214 4924 4522 4933
rect 4214 4922 4220 4924
rect 4276 4922 4300 4924
rect 4356 4922 4380 4924
rect 4436 4922 4460 4924
rect 4516 4922 4522 4924
rect 4276 4870 4278 4922
rect 4458 4870 4460 4922
rect 4214 4868 4220 4870
rect 4276 4868 4300 4870
rect 4356 4868 4380 4870
rect 4436 4868 4460 4870
rect 4516 4868 4522 4870
rect 4214 4859 4522 4868
rect 4068 4684 4120 4690
rect 4068 4626 4120 4632
rect 3896 4236 4016 4264
rect 3896 4010 3924 4236
rect 4080 4185 4108 4626
rect 4160 4616 4212 4622
rect 4160 4558 4212 4564
rect 4066 4176 4122 4185
rect 3976 4140 4028 4146
rect 4172 4146 4200 4558
rect 4632 4554 4660 5199
rect 4724 4690 4752 5324
rect 4804 5306 4856 5312
rect 4712 4684 4764 4690
rect 4712 4626 4764 4632
rect 4816 4570 4844 5306
rect 4908 4758 4936 5782
rect 5000 5688 5028 6190
rect 4988 5682 5040 5688
rect 4986 5672 4988 5681
rect 5040 5672 5042 5681
rect 4986 5607 5042 5616
rect 4988 5568 5040 5574
rect 4988 5510 5040 5516
rect 4896 4752 4948 4758
rect 4896 4694 4948 4700
rect 4620 4548 4672 4554
rect 4620 4490 4672 4496
rect 4724 4542 4844 4570
rect 4066 4111 4122 4120
rect 4160 4140 4212 4146
rect 3976 4082 4028 4088
rect 3884 4004 3936 4010
rect 3884 3946 3936 3952
rect 3896 3398 3924 3946
rect 3988 3534 4016 4082
rect 3976 3528 4028 3534
rect 3976 3470 4028 3476
rect 3884 3392 3936 3398
rect 3884 3334 3936 3340
rect 3988 2990 4016 3470
rect 4080 3466 4108 4111
rect 4160 4082 4212 4088
rect 4214 3836 4522 3845
rect 4214 3834 4220 3836
rect 4276 3834 4300 3836
rect 4356 3834 4380 3836
rect 4436 3834 4460 3836
rect 4516 3834 4522 3836
rect 4276 3782 4278 3834
rect 4458 3782 4460 3834
rect 4214 3780 4220 3782
rect 4276 3780 4300 3782
rect 4356 3780 4380 3782
rect 4436 3780 4460 3782
rect 4516 3780 4522 3782
rect 4214 3771 4522 3780
rect 4068 3460 4120 3466
rect 4068 3402 4120 3408
rect 4066 3224 4122 3233
rect 4066 3159 4122 3168
rect 3976 2984 4028 2990
rect 3976 2926 4028 2932
rect 4080 2938 4108 3159
rect 4632 2990 4660 4490
rect 4724 4486 4752 4542
rect 4712 4480 4764 4486
rect 4712 4422 4764 4428
rect 4896 3664 4948 3670
rect 4896 3606 4948 3612
rect 4908 3448 4936 3606
rect 5000 3466 5028 5510
rect 5092 3738 5120 6326
rect 5184 6322 5212 7890
rect 5172 6316 5224 6322
rect 5172 6258 5224 6264
rect 5276 5658 5304 10406
rect 5368 10130 5396 10610
rect 5552 10198 5580 11698
rect 5828 11626 5856 12310
rect 5906 11792 5962 11801
rect 5906 11727 5962 11736
rect 5816 11620 5868 11626
rect 5816 11562 5868 11568
rect 5632 11008 5684 11014
rect 5632 10950 5684 10956
rect 5540 10192 5592 10198
rect 5540 10134 5592 10140
rect 5356 10124 5408 10130
rect 5356 10066 5408 10072
rect 5644 10062 5672 10950
rect 5816 10532 5868 10538
rect 5816 10474 5868 10480
rect 5724 10192 5776 10198
rect 5724 10134 5776 10140
rect 5632 10056 5684 10062
rect 5632 9998 5684 10004
rect 5540 9988 5592 9994
rect 5540 9930 5592 9936
rect 5552 8974 5580 9930
rect 5632 9920 5684 9926
rect 5632 9862 5684 9868
rect 5644 8974 5672 9862
rect 5736 9450 5764 10134
rect 5828 10130 5856 10474
rect 5920 10418 5948 11727
rect 6012 11694 6040 12378
rect 6196 12306 6224 12406
rect 6184 12300 6236 12306
rect 6184 12242 6236 12248
rect 6000 11688 6052 11694
rect 6000 11630 6052 11636
rect 6012 11150 6040 11630
rect 6092 11620 6144 11626
rect 6092 11562 6144 11568
rect 6104 11286 6132 11562
rect 6092 11280 6144 11286
rect 6092 11222 6144 11228
rect 6000 11144 6052 11150
rect 6000 11086 6052 11092
rect 6104 10606 6132 11222
rect 6092 10600 6144 10606
rect 6196 10588 6224 12242
rect 6288 11218 6316 14200
rect 6644 14068 6696 14074
rect 6644 14010 6696 14016
rect 6460 14000 6512 14006
rect 6460 13942 6512 13948
rect 6472 13394 6500 13942
rect 6460 13388 6512 13394
rect 6460 13330 6512 13336
rect 6472 12850 6500 13330
rect 6460 12844 6512 12850
rect 6460 12786 6512 12792
rect 6552 12776 6604 12782
rect 6552 12718 6604 12724
rect 6564 12102 6592 12718
rect 6552 12096 6604 12102
rect 6552 12038 6604 12044
rect 6564 11898 6592 12038
rect 6552 11892 6604 11898
rect 6552 11834 6604 11840
rect 6460 11756 6512 11762
rect 6460 11698 6512 11704
rect 6472 11354 6500 11698
rect 6460 11348 6512 11354
rect 6460 11290 6512 11296
rect 6472 11257 6500 11290
rect 6458 11248 6514 11257
rect 6276 11212 6328 11218
rect 6458 11183 6514 11192
rect 6276 11154 6328 11160
rect 6288 10742 6316 11154
rect 6460 11008 6512 11014
rect 6458 10976 6460 10985
rect 6512 10976 6514 10985
rect 6458 10911 6514 10920
rect 6276 10736 6328 10742
rect 6276 10678 6328 10684
rect 6366 10704 6422 10713
rect 6366 10639 6422 10648
rect 6196 10560 6316 10588
rect 6092 10542 6144 10548
rect 6184 10464 6236 10470
rect 5920 10390 6132 10418
rect 6184 10406 6236 10412
rect 6288 10418 6316 10560
rect 6380 10538 6408 10639
rect 6368 10532 6420 10538
rect 6368 10474 6420 10480
rect 6472 10441 6500 10911
rect 6564 10606 6592 11834
rect 6656 11393 6684 14010
rect 7484 13569 7512 14200
rect 7840 14136 7892 14142
rect 7840 14078 7892 14084
rect 7470 13560 7526 13569
rect 7470 13495 7526 13504
rect 7656 13456 7708 13462
rect 7484 13404 7656 13410
rect 7484 13398 7708 13404
rect 7484 13382 7696 13398
rect 7104 13320 7156 13326
rect 7104 13262 7156 13268
rect 7194 13288 7250 13297
rect 7116 12918 7144 13262
rect 7194 13223 7250 13232
rect 7104 12912 7156 12918
rect 7104 12854 7156 12860
rect 7012 12776 7064 12782
rect 7012 12718 7064 12724
rect 7024 12442 7052 12718
rect 7208 12646 7236 13223
rect 7288 13184 7340 13190
rect 7288 13126 7340 13132
rect 7300 12918 7328 13126
rect 7484 12986 7512 13382
rect 7656 13320 7708 13326
rect 7656 13262 7708 13268
rect 7668 13190 7696 13262
rect 7656 13184 7708 13190
rect 7656 13126 7708 13132
rect 7472 12980 7524 12986
rect 7472 12922 7524 12928
rect 7288 12912 7340 12918
rect 7288 12854 7340 12860
rect 7104 12640 7156 12646
rect 7104 12582 7156 12588
rect 7196 12640 7248 12646
rect 7196 12582 7248 12588
rect 7012 12436 7064 12442
rect 7012 12378 7064 12384
rect 7116 12238 7144 12582
rect 7300 12374 7328 12854
rect 7656 12844 7708 12850
rect 7656 12786 7708 12792
rect 7288 12368 7340 12374
rect 7288 12310 7340 12316
rect 7380 12368 7432 12374
rect 7380 12310 7432 12316
rect 7472 12368 7524 12374
rect 7472 12310 7524 12316
rect 7104 12232 7156 12238
rect 6826 12200 6882 12209
rect 7104 12174 7156 12180
rect 6826 12135 6882 12144
rect 7012 12164 7064 12170
rect 6734 11792 6790 11801
rect 6840 11762 6868 12135
rect 7012 12106 7064 12112
rect 6734 11727 6790 11736
rect 6828 11756 6880 11762
rect 6642 11384 6698 11393
rect 6642 11319 6698 11328
rect 6644 11280 6696 11286
rect 6644 11222 6696 11228
rect 6656 10810 6684 11222
rect 6748 11014 6776 11727
rect 7024 11744 7052 12106
rect 7392 11898 7420 12310
rect 7484 12238 7512 12310
rect 7472 12232 7524 12238
rect 7472 12174 7524 12180
rect 7668 12170 7696 12786
rect 7656 12164 7708 12170
rect 7656 12106 7708 12112
rect 7562 12064 7618 12073
rect 7562 11999 7618 12008
rect 7380 11892 7432 11898
rect 7380 11834 7432 11840
rect 7472 11892 7524 11898
rect 7472 11834 7524 11840
rect 7104 11756 7156 11762
rect 7024 11716 7104 11744
rect 6828 11698 6880 11704
rect 7104 11698 7156 11704
rect 6840 11268 6868 11698
rect 6920 11688 6972 11694
rect 6920 11630 6972 11636
rect 7194 11656 7250 11665
rect 6932 11529 6960 11630
rect 7104 11620 7156 11626
rect 7194 11591 7250 11600
rect 7104 11562 7156 11568
rect 7012 11552 7064 11558
rect 6918 11520 6974 11529
rect 7012 11494 7064 11500
rect 6918 11455 6974 11464
rect 6840 11240 6960 11268
rect 6828 11144 6880 11150
rect 6828 11086 6880 11092
rect 6736 11008 6788 11014
rect 6736 10950 6788 10956
rect 6644 10804 6696 10810
rect 6644 10746 6696 10752
rect 6656 10656 6684 10746
rect 6736 10668 6788 10674
rect 6656 10628 6736 10656
rect 6736 10610 6788 10616
rect 6552 10600 6604 10606
rect 6604 10560 6684 10588
rect 6552 10542 6604 10548
rect 6552 10464 6604 10470
rect 6458 10432 6514 10441
rect 6104 10198 6132 10390
rect 6092 10192 6144 10198
rect 6092 10134 6144 10140
rect 5816 10124 5868 10130
rect 5816 10066 5868 10072
rect 5828 9625 5856 10066
rect 6092 10056 6144 10062
rect 6092 9998 6144 10004
rect 5814 9616 5870 9625
rect 5814 9551 5870 9560
rect 5908 9580 5960 9586
rect 5724 9444 5776 9450
rect 5724 9386 5776 9392
rect 5828 9178 5856 9551
rect 5908 9522 5960 9528
rect 5816 9172 5868 9178
rect 5816 9114 5868 9120
rect 5540 8968 5592 8974
rect 5540 8910 5592 8916
rect 5632 8968 5684 8974
rect 5632 8910 5684 8916
rect 5448 8900 5500 8906
rect 5448 8842 5500 8848
rect 5460 8378 5488 8842
rect 5552 8498 5580 8910
rect 5644 8566 5672 8910
rect 5632 8560 5684 8566
rect 5632 8502 5684 8508
rect 5828 8498 5856 9114
rect 5920 8974 5948 9522
rect 5908 8968 5960 8974
rect 5908 8910 5960 8916
rect 5540 8492 5592 8498
rect 5540 8434 5592 8440
rect 5816 8492 5868 8498
rect 5816 8434 5868 8440
rect 5460 8350 5580 8378
rect 5552 7478 5580 8350
rect 5816 8356 5868 8362
rect 5816 8298 5868 8304
rect 5828 8090 5856 8298
rect 5816 8084 5868 8090
rect 5816 8026 5868 8032
rect 5920 7886 5948 8910
rect 6104 8498 6132 9998
rect 6092 8492 6144 8498
rect 6092 8434 6144 8440
rect 5908 7880 5960 7886
rect 5908 7822 5960 7828
rect 5920 7546 5948 7822
rect 5908 7540 5960 7546
rect 5908 7482 5960 7488
rect 5540 7472 5592 7478
rect 5540 7414 5592 7420
rect 5540 7200 5592 7206
rect 5540 7142 5592 7148
rect 5552 6866 5580 7142
rect 5540 6860 5592 6866
rect 5540 6802 5592 6808
rect 5632 6792 5684 6798
rect 5632 6734 5684 6740
rect 5540 6656 5592 6662
rect 5540 6598 5592 6604
rect 5552 6322 5580 6598
rect 5540 6316 5592 6322
rect 5540 6258 5592 6264
rect 5448 5908 5500 5914
rect 5448 5850 5500 5856
rect 5460 5710 5488 5850
rect 5552 5794 5580 6258
rect 5644 5930 5672 6734
rect 6196 6474 6224 10406
rect 6288 10390 6408 10418
rect 6274 10160 6330 10169
rect 6274 10095 6330 10104
rect 6288 9994 6316 10095
rect 6276 9988 6328 9994
rect 6276 9930 6328 9936
rect 6288 9722 6316 9930
rect 6276 9716 6328 9722
rect 6276 9658 6328 9664
rect 6274 9208 6330 9217
rect 6274 9143 6330 9152
rect 6288 8974 6316 9143
rect 6276 8968 6328 8974
rect 6276 8910 6328 8916
rect 6276 8628 6328 8634
rect 6276 8570 6328 8576
rect 6288 7274 6316 8570
rect 6276 7268 6328 7274
rect 6276 7210 6328 7216
rect 6380 6934 6408 10390
rect 6552 10406 6604 10412
rect 6458 10367 6514 10376
rect 6472 10033 6500 10367
rect 6564 10266 6592 10406
rect 6552 10260 6604 10266
rect 6552 10202 6604 10208
rect 6550 10160 6606 10169
rect 6550 10095 6606 10104
rect 6458 10024 6514 10033
rect 6458 9959 6514 9968
rect 6564 9926 6592 10095
rect 6552 9920 6604 9926
rect 6458 9888 6514 9897
rect 6552 9862 6604 9868
rect 6458 9823 6514 9832
rect 6472 9586 6500 9823
rect 6460 9580 6512 9586
rect 6460 9522 6512 9528
rect 6472 7886 6500 9522
rect 6564 8634 6592 9862
rect 6552 8628 6604 8634
rect 6552 8570 6604 8576
rect 6656 8566 6684 10560
rect 6736 10532 6788 10538
rect 6736 10474 6788 10480
rect 6748 10198 6776 10474
rect 6736 10192 6788 10198
rect 6736 10134 6788 10140
rect 6736 10034 6788 10040
rect 6734 10024 6736 10033
rect 6788 10024 6790 10033
rect 6734 9959 6790 9968
rect 6736 9920 6788 9926
rect 6736 9862 6788 9868
rect 6748 9489 6776 9862
rect 6734 9480 6790 9489
rect 6734 9415 6790 9424
rect 6748 8974 6776 9415
rect 6840 9178 6868 11086
rect 6932 10198 6960 11240
rect 7024 11014 7052 11494
rect 7116 11218 7144 11562
rect 7104 11212 7156 11218
rect 7104 11154 7156 11160
rect 7208 11082 7236 11591
rect 7288 11552 7340 11558
rect 7288 11494 7340 11500
rect 7300 11218 7328 11494
rect 7288 11212 7340 11218
rect 7288 11154 7340 11160
rect 7196 11076 7248 11082
rect 7196 11018 7248 11024
rect 7012 11008 7064 11014
rect 7300 10962 7328 11154
rect 7012 10950 7064 10956
rect 7208 10934 7328 10962
rect 7012 10804 7064 10810
rect 7012 10746 7064 10752
rect 7024 10713 7052 10746
rect 7010 10704 7066 10713
rect 7010 10639 7066 10648
rect 7104 10668 7156 10674
rect 6920 10192 6972 10198
rect 6920 10134 6972 10140
rect 7024 10130 7052 10639
rect 7104 10610 7156 10616
rect 7012 10124 7064 10130
rect 7012 10066 7064 10072
rect 7012 9988 7064 9994
rect 7012 9930 7064 9936
rect 6920 9920 6972 9926
rect 7024 9897 7052 9930
rect 6920 9862 6972 9868
rect 7010 9888 7066 9897
rect 6932 9568 6960 9862
rect 7010 9823 7066 9832
rect 7012 9580 7064 9586
rect 6932 9540 7012 9568
rect 7012 9522 7064 9528
rect 7116 9500 7144 10610
rect 7208 10577 7236 10934
rect 7288 10668 7340 10674
rect 7288 10610 7340 10616
rect 7194 10568 7250 10577
rect 7194 10503 7250 10512
rect 7196 10124 7248 10130
rect 7196 10066 7248 10072
rect 7208 9761 7236 10066
rect 7300 9926 7328 10610
rect 7392 10538 7420 11834
rect 7484 11665 7512 11834
rect 7470 11656 7526 11665
rect 7470 11591 7526 11600
rect 7470 11520 7526 11529
rect 7470 11455 7526 11464
rect 7484 11286 7512 11455
rect 7472 11280 7524 11286
rect 7472 11222 7524 11228
rect 7472 10668 7524 10674
rect 7472 10610 7524 10616
rect 7380 10532 7432 10538
rect 7380 10474 7432 10480
rect 7378 10296 7434 10305
rect 7378 10231 7434 10240
rect 7288 9920 7340 9926
rect 7288 9862 7340 9868
rect 7194 9752 7250 9761
rect 7194 9687 7196 9696
rect 7248 9687 7250 9696
rect 7196 9658 7248 9664
rect 7288 9512 7340 9518
rect 7116 9472 7288 9500
rect 7288 9454 7340 9460
rect 7012 9444 7064 9450
rect 7012 9386 7064 9392
rect 7024 9178 7052 9386
rect 7116 9382 7144 9413
rect 7104 9376 7156 9382
rect 7102 9344 7104 9353
rect 7156 9344 7158 9353
rect 7102 9279 7158 9288
rect 6828 9172 6880 9178
rect 6828 9114 6880 9120
rect 7012 9172 7064 9178
rect 7012 9114 7064 9120
rect 7116 9042 7144 9279
rect 7104 9036 7156 9042
rect 7104 8978 7156 8984
rect 6736 8968 6788 8974
rect 6736 8910 6788 8916
rect 6918 8936 6974 8945
rect 6918 8871 6974 8880
rect 6644 8560 6696 8566
rect 6644 8502 6696 8508
rect 6736 8492 6788 8498
rect 6736 8434 6788 8440
rect 6550 8256 6606 8265
rect 6550 8191 6606 8200
rect 6460 7880 6512 7886
rect 6460 7822 6512 7828
rect 6564 7206 6592 8191
rect 6748 7954 6776 8434
rect 6736 7948 6788 7954
rect 6736 7890 6788 7896
rect 6644 7812 6696 7818
rect 6644 7754 6696 7760
rect 6552 7200 6604 7206
rect 6552 7142 6604 7148
rect 6368 6928 6420 6934
rect 6368 6870 6420 6876
rect 6196 6446 6316 6474
rect 6184 6384 6236 6390
rect 6288 6361 6316 6446
rect 6184 6326 6236 6332
rect 6274 6352 6330 6361
rect 5998 6216 6054 6225
rect 5998 6151 6054 6160
rect 5816 6112 5868 6118
rect 5816 6054 5868 6060
rect 5644 5902 5764 5930
rect 5736 5846 5764 5902
rect 5724 5840 5776 5846
rect 5552 5766 5672 5794
rect 5724 5782 5776 5788
rect 5184 5630 5304 5658
rect 5448 5704 5500 5710
rect 5448 5646 5500 5652
rect 5540 5704 5592 5710
rect 5540 5646 5592 5652
rect 5184 4554 5212 5630
rect 5552 5556 5580 5646
rect 5262 5536 5318 5545
rect 5262 5471 5318 5480
rect 5368 5528 5580 5556
rect 5276 5166 5304 5471
rect 5264 5160 5316 5166
rect 5264 5102 5316 5108
rect 5172 4548 5224 4554
rect 5172 4490 5224 4496
rect 5172 4208 5224 4214
rect 5172 4150 5224 4156
rect 5080 3732 5132 3738
rect 5080 3674 5132 3680
rect 5184 3670 5212 4150
rect 5172 3664 5224 3670
rect 5172 3606 5224 3612
rect 4988 3460 5040 3466
rect 4908 3420 4988 3448
rect 4988 3402 5040 3408
rect 4712 3052 4764 3058
rect 4712 2994 4764 3000
rect 4620 2984 4672 2990
rect 4080 2910 4200 2938
rect 4620 2926 4672 2932
rect 4172 2854 4200 2910
rect 4160 2848 4212 2854
rect 4160 2790 4212 2796
rect 3804 2746 3924 2774
rect 3700 2508 3752 2514
rect 3700 2450 3752 2456
rect 3712 1873 3740 2450
rect 3698 1864 3754 1873
rect 3698 1799 3754 1808
rect 3516 1488 3568 1494
rect 3516 1430 3568 1436
rect 3424 1352 3476 1358
rect 3252 1312 3424 1340
rect 3424 1294 3476 1300
rect 3608 1352 3660 1358
rect 3896 1329 3924 2746
rect 4214 2748 4522 2757
rect 4214 2746 4220 2748
rect 4276 2746 4300 2748
rect 4356 2746 4380 2748
rect 4436 2746 4460 2748
rect 4516 2746 4522 2748
rect 4276 2694 4278 2746
rect 4458 2694 4460 2746
rect 4214 2692 4220 2694
rect 4276 2692 4300 2694
rect 4356 2692 4380 2694
rect 4436 2692 4460 2694
rect 4516 2692 4522 2694
rect 4214 2683 4522 2692
rect 4068 2644 4120 2650
rect 4068 2586 4120 2592
rect 4080 2417 4108 2586
rect 4066 2408 4122 2417
rect 4066 2343 4122 2352
rect 4160 2372 4212 2378
rect 3976 1556 4028 1562
rect 3976 1498 4028 1504
rect 3988 1426 4016 1498
rect 3976 1420 4028 1426
rect 3976 1362 4028 1368
rect 4080 1340 4108 2343
rect 4160 2314 4212 2320
rect 4172 2009 4200 2314
rect 4436 2304 4488 2310
rect 4436 2246 4488 2252
rect 4158 2000 4214 2009
rect 4158 1935 4214 1944
rect 4448 1766 4476 2246
rect 4620 2100 4672 2106
rect 4724 2088 4752 2994
rect 4896 2440 4948 2446
rect 5000 2428 5028 3402
rect 5172 3120 5224 3126
rect 5172 3062 5224 3068
rect 5080 2984 5132 2990
rect 5080 2926 5132 2932
rect 5092 2689 5120 2926
rect 5184 2854 5212 3062
rect 5276 2854 5304 5102
rect 5368 4690 5396 5528
rect 5644 5234 5672 5766
rect 5632 5228 5684 5234
rect 5632 5170 5684 5176
rect 5540 5024 5592 5030
rect 5540 4966 5592 4972
rect 5736 4978 5764 5782
rect 5828 5574 5856 6054
rect 5816 5568 5868 5574
rect 5816 5510 5868 5516
rect 5356 4684 5408 4690
rect 5356 4626 5408 4632
rect 5368 4060 5396 4626
rect 5552 4554 5580 4966
rect 5736 4950 5856 4978
rect 5540 4548 5592 4554
rect 5540 4490 5592 4496
rect 5724 4276 5776 4282
rect 5724 4218 5776 4224
rect 5448 4072 5500 4078
rect 5368 4032 5448 4060
rect 5172 2848 5224 2854
rect 5172 2790 5224 2796
rect 5264 2848 5316 2854
rect 5264 2790 5316 2796
rect 5078 2680 5134 2689
rect 5078 2615 5134 2624
rect 5092 2514 5120 2615
rect 5080 2508 5132 2514
rect 5080 2450 5132 2456
rect 5276 2446 5304 2790
rect 5368 2514 5396 4032
rect 5448 4014 5500 4020
rect 5448 3936 5500 3942
rect 5448 3878 5500 3884
rect 5460 3602 5488 3878
rect 5448 3596 5500 3602
rect 5448 3538 5500 3544
rect 5460 3058 5488 3538
rect 5540 3460 5592 3466
rect 5540 3402 5592 3408
rect 5448 3052 5500 3058
rect 5448 2994 5500 3000
rect 5552 2972 5580 3402
rect 5736 2990 5764 4218
rect 5828 3618 5856 4950
rect 5908 3936 5960 3942
rect 5908 3878 5960 3884
rect 5920 3738 5948 3878
rect 6012 3738 6040 6151
rect 6196 5234 6224 6326
rect 6274 6287 6330 6296
rect 6656 6254 6684 7754
rect 6748 7478 6776 7890
rect 6828 7812 6880 7818
rect 6828 7754 6880 7760
rect 6736 7472 6788 7478
rect 6736 7414 6788 7420
rect 6736 7200 6788 7206
rect 6736 7142 6788 7148
rect 6748 6644 6776 7142
rect 6840 6798 6868 7754
rect 6828 6792 6880 6798
rect 6828 6734 6880 6740
rect 6932 6746 6960 8871
rect 7116 8838 7144 8978
rect 7196 8900 7248 8906
rect 7196 8842 7248 8848
rect 7104 8832 7156 8838
rect 7104 8774 7156 8780
rect 7012 8628 7064 8634
rect 7012 8570 7064 8576
rect 7024 8430 7052 8570
rect 7116 8498 7144 8774
rect 7104 8492 7156 8498
rect 7104 8434 7156 8440
rect 7012 8424 7064 8430
rect 7208 8401 7236 8842
rect 7012 8366 7064 8372
rect 7194 8392 7250 8401
rect 7024 8090 7052 8366
rect 7104 8356 7156 8362
rect 7194 8327 7250 8336
rect 7104 8298 7156 8304
rect 7012 8084 7064 8090
rect 7012 8026 7064 8032
rect 7012 7744 7064 7750
rect 7012 7686 7064 7692
rect 7024 7410 7052 7686
rect 7012 7404 7064 7410
rect 7012 7346 7064 7352
rect 7024 6866 7052 7346
rect 7116 7342 7144 8298
rect 7194 8120 7250 8129
rect 7194 8055 7250 8064
rect 7208 7410 7236 8055
rect 7300 7886 7328 9454
rect 7392 9178 7420 10231
rect 7484 10198 7512 10610
rect 7472 10192 7524 10198
rect 7472 10134 7524 10140
rect 7484 9722 7512 10134
rect 7472 9716 7524 9722
rect 7472 9658 7524 9664
rect 7576 9466 7604 11999
rect 7668 11200 7696 12106
rect 7748 12096 7800 12102
rect 7748 12038 7800 12044
rect 7760 11558 7788 12038
rect 7852 11898 7880 14078
rect 7932 13932 7984 13938
rect 7932 13874 7984 13880
rect 7944 12434 7972 13874
rect 8588 13734 8616 14200
rect 9772 14136 9824 14142
rect 9772 14078 9824 14084
rect 9784 13841 9812 14078
rect 9770 13832 9826 13841
rect 9680 13796 9732 13802
rect 9770 13767 9826 13776
rect 9680 13738 9732 13744
rect 8024 13728 8076 13734
rect 8024 13670 8076 13676
rect 8576 13728 8628 13734
rect 8576 13670 8628 13676
rect 8036 13326 8064 13670
rect 8298 13424 8354 13433
rect 8298 13359 8354 13368
rect 8850 13424 8906 13433
rect 8850 13359 8906 13368
rect 8312 13326 8340 13359
rect 8024 13320 8076 13326
rect 8024 13262 8076 13268
rect 8300 13320 8352 13326
rect 8484 13320 8536 13326
rect 8300 13262 8352 13268
rect 8482 13288 8484 13297
rect 8760 13320 8812 13326
rect 8536 13288 8538 13297
rect 8208 13252 8260 13258
rect 8128 13212 8208 13240
rect 8128 12832 8156 13212
rect 8760 13262 8812 13268
rect 8482 13223 8538 13232
rect 8208 13194 8260 13200
rect 8214 13084 8522 13093
rect 8214 13082 8220 13084
rect 8276 13082 8300 13084
rect 8356 13082 8380 13084
rect 8436 13082 8460 13084
rect 8516 13082 8522 13084
rect 8276 13030 8278 13082
rect 8458 13030 8460 13082
rect 8214 13028 8220 13030
rect 8276 13028 8300 13030
rect 8356 13028 8380 13030
rect 8436 13028 8460 13030
rect 8516 13028 8522 13030
rect 8214 13019 8522 13028
rect 8772 12850 8800 13262
rect 8392 12844 8444 12850
rect 8128 12804 8392 12832
rect 7944 12406 8064 12434
rect 7932 12232 7984 12238
rect 7932 12174 7984 12180
rect 7944 11937 7972 12174
rect 7930 11928 7986 11937
rect 7840 11892 7892 11898
rect 7930 11863 7986 11872
rect 7840 11834 7892 11840
rect 7932 11824 7984 11830
rect 7930 11792 7932 11801
rect 7984 11792 7986 11801
rect 7930 11727 7986 11736
rect 7932 11688 7984 11694
rect 7932 11630 7984 11636
rect 7748 11552 7800 11558
rect 7748 11494 7800 11500
rect 7840 11552 7892 11558
rect 7840 11494 7892 11500
rect 7668 11172 7788 11200
rect 7760 10962 7788 11172
rect 7852 11082 7880 11494
rect 7840 11076 7892 11082
rect 7840 11018 7892 11024
rect 7944 10985 7972 11630
rect 7930 10976 7986 10985
rect 7760 10934 7880 10962
rect 7746 10840 7802 10849
rect 7656 10804 7708 10810
rect 7746 10775 7802 10784
rect 7656 10746 7708 10752
rect 7668 9489 7696 10746
rect 7484 9438 7604 9466
rect 7654 9480 7710 9489
rect 7380 9172 7432 9178
rect 7380 9114 7432 9120
rect 7380 8900 7432 8906
rect 7380 8842 7432 8848
rect 7288 7880 7340 7886
rect 7288 7822 7340 7828
rect 7196 7404 7248 7410
rect 7196 7346 7248 7352
rect 7104 7336 7156 7342
rect 7104 7278 7156 7284
rect 7012 6860 7064 6866
rect 7012 6802 7064 6808
rect 6932 6718 7052 6746
rect 6920 6656 6972 6662
rect 6748 6616 6868 6644
rect 6644 6248 6696 6254
rect 6644 6190 6696 6196
rect 6368 6112 6420 6118
rect 6368 6054 6420 6060
rect 6184 5228 6236 5234
rect 6184 5170 6236 5176
rect 6196 4740 6224 5170
rect 6380 5098 6408 6054
rect 6656 5148 6684 6190
rect 6736 5160 6788 5166
rect 6656 5120 6736 5148
rect 6736 5102 6788 5108
rect 6368 5092 6420 5098
rect 6368 5034 6420 5040
rect 6460 5024 6512 5030
rect 6460 4966 6512 4972
rect 6276 4752 6328 4758
rect 6196 4712 6276 4740
rect 6276 4694 6328 4700
rect 6368 4208 6420 4214
rect 6368 4150 6420 4156
rect 6092 3936 6144 3942
rect 6092 3878 6144 3884
rect 5908 3732 5960 3738
rect 5908 3674 5960 3680
rect 6000 3732 6052 3738
rect 6000 3674 6052 3680
rect 5828 3602 5948 3618
rect 5828 3596 5960 3602
rect 5828 3590 5908 3596
rect 5908 3538 5960 3544
rect 5816 3528 5868 3534
rect 5816 3470 5868 3476
rect 5828 3194 5856 3470
rect 5816 3188 5868 3194
rect 5816 3130 5868 3136
rect 5908 3052 5960 3058
rect 6012 3040 6040 3674
rect 6104 3126 6132 3878
rect 6380 3738 6408 4150
rect 6368 3732 6420 3738
rect 6368 3674 6420 3680
rect 6472 3534 6500 4966
rect 6840 4214 6868 6616
rect 6920 6598 6972 6604
rect 6932 6322 6960 6598
rect 7024 6390 7052 6718
rect 7012 6384 7064 6390
rect 7012 6326 7064 6332
rect 6920 6316 6972 6322
rect 6920 6258 6972 6264
rect 6932 5234 6960 6258
rect 7392 6254 7420 8842
rect 7484 6780 7512 9438
rect 7654 9415 7710 9424
rect 7656 9376 7708 9382
rect 7656 9318 7708 9324
rect 7668 9178 7696 9318
rect 7656 9172 7708 9178
rect 7656 9114 7708 9120
rect 7564 8424 7616 8430
rect 7564 8366 7616 8372
rect 7576 7886 7604 8366
rect 7760 8294 7788 10775
rect 7852 10742 7880 10934
rect 7930 10911 7986 10920
rect 7932 10804 7984 10810
rect 7932 10746 7984 10752
rect 7840 10736 7892 10742
rect 7840 10678 7892 10684
rect 7840 10600 7892 10606
rect 7944 10588 7972 10746
rect 7892 10560 7972 10588
rect 7840 10542 7892 10548
rect 7932 9920 7984 9926
rect 7932 9862 7984 9868
rect 7838 9480 7894 9489
rect 7838 9415 7840 9424
rect 7892 9415 7894 9424
rect 7840 9386 7892 9392
rect 7840 8968 7892 8974
rect 7838 8936 7840 8945
rect 7892 8936 7894 8945
rect 7838 8871 7894 8880
rect 7838 8664 7894 8673
rect 7838 8599 7840 8608
rect 7892 8599 7894 8608
rect 7840 8570 7892 8576
rect 7944 8566 7972 9862
rect 7932 8560 7984 8566
rect 7932 8502 7984 8508
rect 7932 8356 7984 8362
rect 7932 8298 7984 8304
rect 7668 8266 7788 8294
rect 7564 7880 7616 7886
rect 7564 7822 7616 7828
rect 7576 7750 7604 7822
rect 7564 7744 7616 7750
rect 7564 7686 7616 7692
rect 7668 7546 7696 8266
rect 7840 8084 7892 8090
rect 7840 8026 7892 8032
rect 7656 7540 7708 7546
rect 7656 7482 7708 7488
rect 7748 7336 7800 7342
rect 7748 7278 7800 7284
rect 7564 6792 7616 6798
rect 7484 6752 7564 6780
rect 7564 6734 7616 6740
rect 7656 6724 7708 6730
rect 7656 6666 7708 6672
rect 7380 6248 7432 6254
rect 7380 6190 7432 6196
rect 7012 5636 7064 5642
rect 7012 5578 7064 5584
rect 6920 5228 6972 5234
rect 6920 5170 6972 5176
rect 6920 4548 6972 4554
rect 6920 4490 6972 4496
rect 6828 4208 6880 4214
rect 6828 4150 6880 4156
rect 6644 3936 6696 3942
rect 6644 3878 6696 3884
rect 6656 3602 6684 3878
rect 6644 3596 6696 3602
rect 6644 3538 6696 3544
rect 6460 3528 6512 3534
rect 6512 3488 6592 3516
rect 6460 3470 6512 3476
rect 6276 3392 6328 3398
rect 6276 3334 6328 3340
rect 6092 3120 6144 3126
rect 6092 3062 6144 3068
rect 6288 3058 6316 3334
rect 5960 3012 6040 3040
rect 6276 3052 6328 3058
rect 5908 2994 5960 3000
rect 6276 2994 6328 3000
rect 5724 2984 5776 2990
rect 5552 2944 5672 2972
rect 5356 2508 5408 2514
rect 5356 2450 5408 2456
rect 5540 2508 5592 2514
rect 5540 2450 5592 2456
rect 4948 2400 5028 2428
rect 5264 2440 5316 2446
rect 4896 2382 4948 2388
rect 5264 2382 5316 2388
rect 4896 2304 4948 2310
rect 4896 2246 4948 2252
rect 4988 2304 5040 2310
rect 4988 2246 5040 2252
rect 4908 2106 4936 2246
rect 4672 2060 4752 2088
rect 4620 2042 4672 2048
rect 4436 1760 4488 1766
rect 4436 1702 4488 1708
rect 4620 1760 4672 1766
rect 4620 1702 4672 1708
rect 4214 1660 4522 1669
rect 4214 1658 4220 1660
rect 4276 1658 4300 1660
rect 4356 1658 4380 1660
rect 4436 1658 4460 1660
rect 4516 1658 4522 1660
rect 4276 1606 4278 1658
rect 4458 1606 4460 1658
rect 4214 1604 4220 1606
rect 4276 1604 4300 1606
rect 4356 1604 4380 1606
rect 4436 1604 4460 1606
rect 4516 1604 4522 1606
rect 4214 1595 4522 1604
rect 4160 1352 4212 1358
rect 3608 1294 3660 1300
rect 3882 1320 3938 1329
rect 2964 1012 3016 1018
rect 2964 954 3016 960
rect 3436 950 3464 1294
rect 3424 944 3476 950
rect 3424 886 3476 892
rect 3620 898 3648 1294
rect 4080 1312 4160 1340
rect 4160 1294 4212 1300
rect 4632 1290 4660 1702
rect 4724 1358 4752 2060
rect 4896 2100 4948 2106
rect 4896 2042 4948 2048
rect 5000 1426 5028 2246
rect 5448 2032 5500 2038
rect 5552 2020 5580 2450
rect 5644 2446 5672 2944
rect 5724 2926 5776 2932
rect 5632 2440 5684 2446
rect 5632 2382 5684 2388
rect 5736 2310 5764 2926
rect 5724 2304 5776 2310
rect 5724 2246 5776 2252
rect 5632 2032 5684 2038
rect 5552 1992 5632 2020
rect 5448 1974 5500 1980
rect 5632 1974 5684 1980
rect 4988 1420 5040 1426
rect 4988 1362 5040 1368
rect 4712 1352 4764 1358
rect 4712 1294 4764 1300
rect 5460 1290 5488 1974
rect 5736 1340 5764 2246
rect 6564 1970 6592 3488
rect 6828 3392 6880 3398
rect 6828 3334 6880 3340
rect 6840 3194 6868 3334
rect 6828 3188 6880 3194
rect 6828 3130 6880 3136
rect 6932 3126 6960 4490
rect 7024 4282 7052 5578
rect 7392 4758 7420 6190
rect 7668 5778 7696 6666
rect 7760 6458 7788 7278
rect 7852 6730 7880 8026
rect 7944 7818 7972 8298
rect 7932 7812 7984 7818
rect 7932 7754 7984 7760
rect 7840 6724 7892 6730
rect 7840 6666 7892 6672
rect 8036 6662 8064 12406
rect 8220 12374 8248 12804
rect 8312 12646 8340 12804
rect 8576 12844 8628 12850
rect 8392 12786 8444 12792
rect 8496 12804 8576 12832
rect 8300 12640 8352 12646
rect 8300 12582 8352 12588
rect 8208 12368 8260 12374
rect 8208 12310 8260 12316
rect 8496 12306 8524 12804
rect 8576 12786 8628 12792
rect 8760 12844 8812 12850
rect 8760 12786 8812 12792
rect 8576 12708 8628 12714
rect 8576 12650 8628 12656
rect 8484 12300 8536 12306
rect 8484 12242 8536 12248
rect 8208 12232 8260 12238
rect 8128 12192 8208 12220
rect 8128 11150 8156 12192
rect 8208 12174 8260 12180
rect 8214 11996 8522 12005
rect 8214 11994 8220 11996
rect 8276 11994 8300 11996
rect 8356 11994 8380 11996
rect 8436 11994 8460 11996
rect 8516 11994 8522 11996
rect 8276 11942 8278 11994
rect 8458 11942 8460 11994
rect 8214 11940 8220 11942
rect 8276 11940 8300 11942
rect 8356 11940 8380 11942
rect 8436 11940 8460 11942
rect 8516 11940 8522 11942
rect 8214 11931 8522 11940
rect 8588 11762 8616 12650
rect 8668 12232 8720 12238
rect 8666 12200 8668 12209
rect 8720 12200 8722 12209
rect 8666 12135 8722 12144
rect 8666 12064 8722 12073
rect 8666 11999 8722 12008
rect 8576 11756 8628 11762
rect 8576 11698 8628 11704
rect 8484 11688 8536 11694
rect 8484 11630 8536 11636
rect 8300 11620 8352 11626
rect 8300 11562 8352 11568
rect 8312 11370 8340 11562
rect 8496 11529 8524 11630
rect 8482 11520 8538 11529
rect 8482 11455 8538 11464
rect 8220 11342 8340 11370
rect 8390 11384 8446 11393
rect 8220 11286 8248 11342
rect 8390 11319 8446 11328
rect 8208 11280 8260 11286
rect 8208 11222 8260 11228
rect 8116 11144 8168 11150
rect 8114 11112 8116 11121
rect 8168 11112 8170 11121
rect 8114 11047 8170 11056
rect 8404 11014 8432 11319
rect 8496 11218 8524 11455
rect 8588 11286 8616 11698
rect 8680 11529 8708 11999
rect 8666 11520 8722 11529
rect 8666 11455 8722 11464
rect 8576 11280 8628 11286
rect 8576 11222 8628 11228
rect 8484 11212 8536 11218
rect 8484 11154 8536 11160
rect 8576 11144 8628 11150
rect 8576 11086 8628 11092
rect 8392 11008 8444 11014
rect 8392 10950 8444 10956
rect 8214 10908 8522 10917
rect 8214 10906 8220 10908
rect 8276 10906 8300 10908
rect 8356 10906 8380 10908
rect 8436 10906 8460 10908
rect 8516 10906 8522 10908
rect 8276 10854 8278 10906
rect 8458 10854 8460 10906
rect 8214 10852 8220 10854
rect 8276 10852 8300 10854
rect 8356 10852 8380 10854
rect 8436 10852 8460 10854
rect 8516 10852 8522 10854
rect 8214 10843 8522 10852
rect 8588 10810 8616 11086
rect 8668 11076 8720 11082
rect 8668 11018 8720 11024
rect 8576 10804 8628 10810
rect 8576 10746 8628 10752
rect 8298 10704 8354 10713
rect 8116 10668 8168 10674
rect 8680 10674 8708 11018
rect 8298 10639 8300 10648
rect 8116 10610 8168 10616
rect 8352 10639 8354 10648
rect 8668 10668 8720 10674
rect 8300 10610 8352 10616
rect 8668 10610 8720 10616
rect 8128 10538 8156 10610
rect 8392 10600 8444 10606
rect 8390 10568 8392 10577
rect 8444 10568 8446 10577
rect 8116 10532 8168 10538
rect 8390 10503 8446 10512
rect 8116 10474 8168 10480
rect 8574 10296 8630 10305
rect 8300 10260 8352 10266
rect 8772 10266 8800 12786
rect 8864 12374 8892 13359
rect 9220 13184 9272 13190
rect 9220 13126 9272 13132
rect 9232 12986 9260 13126
rect 9220 12980 9272 12986
rect 9220 12922 9272 12928
rect 8944 12912 8996 12918
rect 8944 12854 8996 12860
rect 8852 12368 8904 12374
rect 8852 12310 8904 12316
rect 8864 12238 8892 12310
rect 8852 12232 8904 12238
rect 8852 12174 8904 12180
rect 8852 12096 8904 12102
rect 8956 12073 8984 12854
rect 9692 12850 9720 13738
rect 9968 13734 9996 14334
rect 10784 14340 10930 14346
rect 10836 14334 10930 14340
rect 10784 14282 10836 14288
rect 10416 14000 10468 14006
rect 10416 13942 10468 13948
rect 9956 13728 10008 13734
rect 9956 13670 10008 13676
rect 9864 13388 9916 13394
rect 9864 13330 9916 13336
rect 9772 13252 9824 13258
rect 9772 13194 9824 13200
rect 9680 12844 9732 12850
rect 9680 12786 9732 12792
rect 9784 12714 9812 13194
rect 9876 12850 9904 13330
rect 9864 12844 9916 12850
rect 9864 12786 9916 12792
rect 9772 12708 9824 12714
rect 9772 12650 9824 12656
rect 9588 12640 9640 12646
rect 9588 12582 9640 12588
rect 9036 12368 9088 12374
rect 9036 12310 9088 12316
rect 8852 12038 8904 12044
rect 8942 12064 8998 12073
rect 8864 11898 8892 12038
rect 8942 11999 8998 12008
rect 8942 11928 8998 11937
rect 8852 11892 8904 11898
rect 8942 11863 8998 11872
rect 8852 11834 8904 11840
rect 8852 11756 8904 11762
rect 8852 11698 8904 11704
rect 8864 11354 8892 11698
rect 8852 11348 8904 11354
rect 8852 11290 8904 11296
rect 8956 11082 8984 11863
rect 9048 11762 9076 12310
rect 9128 12300 9180 12306
rect 9180 12260 9260 12288
rect 9128 12242 9180 12248
rect 9128 12096 9180 12102
rect 9128 12038 9180 12044
rect 9140 11898 9168 12038
rect 9128 11892 9180 11898
rect 9128 11834 9180 11840
rect 9232 11801 9260 12260
rect 9404 12232 9456 12238
rect 9404 12174 9456 12180
rect 9310 11928 9366 11937
rect 9310 11863 9366 11872
rect 9218 11792 9274 11801
rect 9036 11756 9088 11762
rect 9036 11698 9088 11704
rect 9128 11756 9180 11762
rect 9324 11762 9352 11863
rect 9416 11762 9444 12174
rect 9600 12170 9628 12582
rect 9876 12442 9904 12786
rect 9864 12436 9916 12442
rect 9864 12378 9916 12384
rect 9968 12238 9996 13670
rect 10048 13524 10100 13530
rect 10048 13466 10100 13472
rect 10060 12306 10088 13466
rect 10140 13252 10192 13258
rect 10140 13194 10192 13200
rect 10232 13252 10284 13258
rect 10232 13194 10284 13200
rect 10152 12442 10180 13194
rect 10244 12918 10272 13194
rect 10232 12912 10284 12918
rect 10232 12854 10284 12860
rect 10140 12436 10192 12442
rect 10140 12378 10192 12384
rect 10048 12300 10100 12306
rect 10048 12242 10100 12248
rect 10140 12300 10192 12306
rect 10140 12242 10192 12248
rect 9956 12232 10008 12238
rect 9956 12174 10008 12180
rect 9588 12164 9640 12170
rect 9588 12106 9640 12112
rect 10048 12164 10100 12170
rect 10048 12106 10100 12112
rect 9218 11727 9274 11736
rect 9312 11756 9364 11762
rect 9128 11698 9180 11704
rect 9312 11698 9364 11704
rect 9404 11756 9456 11762
rect 9404 11698 9456 11704
rect 9140 11626 9168 11698
rect 9128 11620 9180 11626
rect 9128 11562 9180 11568
rect 9140 11393 9168 11562
rect 9310 11520 9366 11529
rect 9310 11455 9366 11464
rect 9126 11384 9182 11393
rect 9036 11348 9088 11354
rect 9126 11319 9182 11328
rect 9036 11290 9088 11296
rect 9048 11218 9076 11290
rect 9036 11212 9088 11218
rect 9036 11154 9088 11160
rect 9220 11144 9272 11150
rect 9324 11132 9352 11455
rect 9416 11393 9444 11698
rect 9600 11626 9628 12106
rect 10060 11762 10088 12106
rect 10152 11830 10180 12242
rect 10244 12238 10272 12854
rect 10428 12442 10456 13942
rect 10692 13320 10744 13326
rect 10692 13262 10744 13268
rect 10416 12436 10468 12442
rect 10416 12378 10468 12384
rect 10232 12232 10284 12238
rect 10232 12174 10284 12180
rect 10600 12232 10652 12238
rect 10600 12174 10652 12180
rect 10508 12096 10560 12102
rect 10230 12064 10286 12073
rect 10508 12038 10560 12044
rect 10230 11999 10286 12008
rect 10244 11830 10272 11999
rect 10140 11824 10192 11830
rect 10140 11766 10192 11772
rect 10232 11824 10284 11830
rect 10232 11766 10284 11772
rect 10416 11824 10468 11830
rect 10416 11766 10468 11772
rect 10048 11756 10100 11762
rect 10048 11698 10100 11704
rect 9588 11620 9640 11626
rect 9588 11562 9640 11568
rect 9402 11384 9458 11393
rect 9402 11319 9458 11328
rect 9772 11212 9824 11218
rect 9772 11154 9824 11160
rect 9496 11144 9548 11150
rect 9324 11104 9496 11132
rect 9220 11086 9272 11092
rect 9496 11086 9548 11092
rect 8944 11076 8996 11082
rect 8944 11018 8996 11024
rect 9232 11014 9260 11086
rect 9036 11008 9088 11014
rect 8942 10976 8998 10985
rect 9036 10950 9088 10956
rect 9220 11008 9272 11014
rect 9220 10950 9272 10956
rect 9678 10976 9734 10985
rect 8942 10911 8998 10920
rect 8956 10742 8984 10911
rect 9048 10826 9076 10950
rect 9678 10911 9734 10920
rect 9310 10840 9366 10849
rect 9048 10798 9260 10826
rect 8944 10736 8996 10742
rect 8944 10678 8996 10684
rect 8852 10668 8904 10674
rect 8852 10610 8904 10616
rect 9036 10668 9088 10674
rect 9036 10610 9088 10616
rect 8574 10231 8576 10240
rect 8300 10202 8352 10208
rect 8628 10231 8630 10240
rect 8760 10260 8812 10266
rect 8576 10202 8628 10208
rect 8760 10202 8812 10208
rect 8312 10130 8340 10202
rect 8392 10192 8444 10198
rect 8444 10152 8524 10180
rect 8392 10134 8444 10140
rect 8300 10124 8352 10130
rect 8300 10066 8352 10072
rect 8496 9926 8524 10152
rect 8864 10112 8892 10610
rect 8944 10124 8996 10130
rect 8864 10084 8944 10112
rect 8768 10056 8820 10062
rect 8864 10044 8892 10084
rect 9048 10112 9076 10610
rect 9126 10568 9182 10577
rect 9126 10503 9128 10512
rect 9180 10503 9182 10512
rect 9128 10474 9180 10480
rect 9232 10198 9260 10798
rect 9310 10775 9366 10784
rect 9220 10192 9272 10198
rect 9220 10134 9272 10140
rect 9048 10084 9168 10112
rect 8944 10066 8996 10072
rect 8820 10016 8892 10044
rect 8768 9998 8820 10004
rect 8484 9920 8536 9926
rect 8484 9862 8536 9868
rect 8214 9820 8522 9829
rect 8214 9818 8220 9820
rect 8276 9818 8300 9820
rect 8356 9818 8380 9820
rect 8436 9818 8460 9820
rect 8516 9818 8522 9820
rect 8276 9766 8278 9818
rect 8458 9766 8460 9818
rect 8214 9764 8220 9766
rect 8276 9764 8300 9766
rect 8356 9764 8380 9766
rect 8436 9764 8460 9766
rect 8516 9764 8522 9766
rect 8214 9755 8522 9764
rect 8208 9716 8260 9722
rect 8208 9658 8260 9664
rect 8220 9586 8248 9658
rect 8208 9580 8260 9586
rect 8208 9522 8260 9528
rect 8392 9580 8444 9586
rect 8392 9522 8444 9528
rect 8576 9580 8628 9586
rect 8576 9522 8628 9528
rect 8404 9042 8432 9522
rect 8392 9036 8444 9042
rect 8392 8978 8444 8984
rect 8298 8936 8354 8945
rect 8298 8871 8354 8880
rect 8312 8838 8340 8871
rect 8588 8838 8616 9522
rect 8760 9512 8812 9518
rect 8760 9454 8812 9460
rect 8772 9217 8800 9454
rect 8758 9208 8814 9217
rect 8680 9166 8758 9194
rect 8116 8832 8168 8838
rect 8116 8774 8168 8780
rect 8300 8832 8352 8838
rect 8300 8774 8352 8780
rect 8576 8832 8628 8838
rect 8576 8774 8628 8780
rect 8128 8634 8156 8774
rect 8214 8732 8522 8741
rect 8214 8730 8220 8732
rect 8276 8730 8300 8732
rect 8356 8730 8380 8732
rect 8436 8730 8460 8732
rect 8516 8730 8522 8732
rect 8276 8678 8278 8730
rect 8458 8678 8460 8730
rect 8214 8676 8220 8678
rect 8276 8676 8300 8678
rect 8356 8676 8380 8678
rect 8436 8676 8460 8678
rect 8516 8676 8522 8678
rect 8214 8667 8522 8676
rect 8588 8634 8616 8774
rect 8116 8628 8168 8634
rect 8116 8570 8168 8576
rect 8576 8628 8628 8634
rect 8576 8570 8628 8576
rect 8206 8528 8262 8537
rect 8206 8463 8262 8472
rect 8220 8362 8248 8463
rect 8680 8430 8708 9166
rect 8758 9143 8814 9152
rect 8758 9072 8814 9081
rect 8758 9007 8814 9016
rect 8668 8424 8720 8430
rect 8588 8384 8668 8412
rect 8208 8356 8260 8362
rect 8208 8298 8260 8304
rect 8116 8288 8168 8294
rect 8116 8230 8168 8236
rect 8128 7002 8156 8230
rect 8588 8090 8616 8384
rect 8668 8366 8720 8372
rect 8772 8276 8800 9007
rect 8864 8974 8892 10016
rect 9034 10024 9090 10033
rect 9034 9959 9090 9968
rect 9048 9382 9076 9959
rect 9140 9654 9168 10084
rect 9220 9920 9272 9926
rect 9220 9862 9272 9868
rect 9128 9648 9180 9654
rect 9128 9590 9180 9596
rect 9036 9376 9088 9382
rect 9036 9318 9088 9324
rect 8944 9172 8996 9178
rect 8944 9114 8996 9120
rect 8956 8974 8984 9114
rect 8852 8968 8904 8974
rect 8852 8910 8904 8916
rect 8944 8968 8996 8974
rect 8944 8910 8996 8916
rect 9048 8498 9076 9318
rect 9128 8968 9180 8974
rect 9232 8956 9260 9862
rect 9180 8928 9260 8956
rect 9128 8910 9180 8916
rect 9036 8492 9088 8498
rect 9036 8434 9088 8440
rect 8944 8424 8996 8430
rect 8944 8366 8996 8372
rect 8680 8248 8800 8276
rect 8576 8084 8628 8090
rect 8576 8026 8628 8032
rect 8208 7948 8260 7954
rect 8208 7890 8260 7896
rect 8576 7948 8628 7954
rect 8576 7890 8628 7896
rect 8220 7750 8248 7890
rect 8208 7744 8260 7750
rect 8208 7686 8260 7692
rect 8214 7644 8522 7653
rect 8214 7642 8220 7644
rect 8276 7642 8300 7644
rect 8356 7642 8380 7644
rect 8436 7642 8460 7644
rect 8516 7642 8522 7644
rect 8276 7590 8278 7642
rect 8458 7590 8460 7642
rect 8214 7588 8220 7590
rect 8276 7588 8300 7590
rect 8356 7588 8380 7590
rect 8436 7588 8460 7590
rect 8516 7588 8522 7590
rect 8214 7579 8522 7588
rect 8392 7472 8444 7478
rect 8390 7440 8392 7449
rect 8444 7440 8446 7449
rect 8390 7375 8446 7384
rect 8116 6996 8168 7002
rect 8116 6938 8168 6944
rect 8024 6656 8076 6662
rect 8024 6598 8076 6604
rect 8214 6556 8522 6565
rect 8214 6554 8220 6556
rect 8276 6554 8300 6556
rect 8356 6554 8380 6556
rect 8436 6554 8460 6556
rect 8516 6554 8522 6556
rect 8276 6502 8278 6554
rect 8458 6502 8460 6554
rect 8214 6500 8220 6502
rect 8276 6500 8300 6502
rect 8356 6500 8380 6502
rect 8436 6500 8460 6502
rect 8516 6500 8522 6502
rect 8214 6491 8522 6500
rect 7748 6452 7800 6458
rect 7748 6394 7800 6400
rect 8588 6390 8616 7890
rect 8680 6866 8708 8248
rect 8852 8016 8904 8022
rect 8852 7958 8904 7964
rect 8760 7812 8812 7818
rect 8760 7754 8812 7760
rect 8668 6860 8720 6866
rect 8668 6802 8720 6808
rect 8772 6458 8800 7754
rect 8864 7721 8892 7958
rect 8850 7712 8906 7721
rect 8850 7647 8906 7656
rect 8956 7410 8984 8366
rect 9140 8294 9168 8910
rect 9324 8616 9352 10775
rect 9692 10742 9720 10911
rect 9680 10736 9732 10742
rect 9402 10704 9458 10713
rect 9680 10678 9732 10684
rect 9784 10674 9812 11154
rect 9864 11144 9916 11150
rect 9864 11086 9916 11092
rect 9954 11112 10010 11121
rect 9402 10639 9458 10648
rect 9772 10668 9824 10674
rect 9416 9654 9444 10639
rect 9772 10610 9824 10616
rect 9680 10600 9732 10606
rect 9494 10568 9550 10577
rect 9876 10554 9904 11086
rect 9954 11047 10010 11056
rect 9732 10548 9904 10554
rect 9680 10542 9904 10548
rect 9692 10526 9904 10542
rect 9494 10503 9550 10512
rect 9404 9648 9456 9654
rect 9404 9590 9456 9596
rect 9404 9512 9456 9518
rect 9404 9454 9456 9460
rect 9416 9110 9444 9454
rect 9508 9450 9536 10503
rect 9772 10464 9824 10470
rect 9586 10432 9642 10441
rect 9772 10406 9824 10412
rect 9586 10367 9642 10376
rect 9600 10198 9628 10367
rect 9588 10192 9640 10198
rect 9640 10152 9720 10180
rect 9588 10134 9640 10140
rect 9588 10056 9640 10062
rect 9588 9998 9640 10004
rect 9600 9586 9628 9998
rect 9588 9580 9640 9586
rect 9588 9522 9640 9528
rect 9496 9444 9548 9450
rect 9496 9386 9548 9392
rect 9692 9110 9720 10152
rect 9404 9104 9456 9110
rect 9680 9104 9732 9110
rect 9404 9046 9456 9052
rect 9494 9072 9550 9081
rect 9680 9046 9732 9052
rect 9494 9007 9550 9016
rect 9508 8974 9536 9007
rect 9496 8968 9548 8974
rect 9496 8910 9548 8916
rect 9784 8906 9812 10406
rect 9876 10198 9904 10526
rect 9864 10192 9916 10198
rect 9864 10134 9916 10140
rect 9968 10130 9996 11047
rect 10060 10169 10088 11698
rect 10152 10282 10180 11766
rect 10428 11354 10456 11766
rect 10520 11558 10548 12038
rect 10612 11558 10640 12174
rect 10704 11937 10732 13262
rect 10796 12238 10824 14282
rect 10874 14200 10930 14334
rect 11808 14334 12126 14362
rect 11704 13864 11756 13870
rect 11704 13806 11756 13812
rect 11244 13796 11296 13802
rect 11244 13738 11296 13744
rect 10968 13728 11020 13734
rect 10968 13670 11020 13676
rect 10980 13530 11008 13670
rect 10968 13524 11020 13530
rect 10968 13466 11020 13472
rect 11256 13326 11284 13738
rect 11716 13326 11744 13806
rect 10968 13320 11020 13326
rect 10968 13262 11020 13268
rect 11244 13320 11296 13326
rect 11244 13262 11296 13268
rect 11520 13320 11572 13326
rect 11520 13262 11572 13268
rect 11704 13320 11756 13326
rect 11704 13262 11756 13268
rect 10784 12232 10836 12238
rect 10784 12174 10836 12180
rect 10690 11928 10746 11937
rect 10690 11863 10746 11872
rect 10690 11792 10746 11801
rect 10690 11727 10746 11736
rect 10704 11626 10732 11727
rect 10782 11656 10838 11665
rect 10692 11620 10744 11626
rect 10782 11591 10838 11600
rect 10692 11562 10744 11568
rect 10508 11552 10560 11558
rect 10508 11494 10560 11500
rect 10600 11552 10652 11558
rect 10600 11494 10652 11500
rect 10416 11348 10468 11354
rect 10520 11336 10548 11494
rect 10600 11348 10652 11354
rect 10520 11308 10600 11336
rect 10416 11290 10468 11296
rect 10600 11290 10652 11296
rect 10230 11248 10286 11257
rect 10230 11183 10286 11192
rect 10244 11150 10272 11183
rect 10232 11144 10284 11150
rect 10232 11086 10284 11092
rect 10232 10736 10284 10742
rect 10232 10678 10284 10684
rect 10244 10577 10272 10678
rect 10230 10568 10286 10577
rect 10230 10503 10286 10512
rect 10232 10464 10284 10470
rect 10428 10452 10456 11290
rect 10506 10704 10562 10713
rect 10612 10674 10640 11290
rect 10692 11144 10744 11150
rect 10692 11086 10744 11092
rect 10506 10639 10508 10648
rect 10560 10639 10562 10648
rect 10600 10668 10652 10674
rect 10508 10610 10560 10616
rect 10600 10610 10652 10616
rect 10704 10606 10732 11086
rect 10692 10600 10744 10606
rect 10598 10568 10654 10577
rect 10692 10542 10744 10548
rect 10598 10503 10654 10512
rect 10284 10424 10456 10452
rect 10232 10406 10284 10412
rect 10152 10254 10272 10282
rect 10046 10160 10102 10169
rect 9956 10124 10008 10130
rect 10046 10095 10102 10104
rect 9956 10066 10008 10072
rect 9864 9580 9916 9586
rect 9864 9522 9916 9528
rect 9876 9353 9904 9522
rect 9862 9344 9918 9353
rect 9862 9279 9918 9288
rect 9876 9178 9904 9279
rect 9864 9172 9916 9178
rect 9864 9114 9916 9120
rect 9772 8900 9824 8906
rect 9772 8842 9824 8848
rect 9404 8832 9456 8838
rect 9404 8774 9456 8780
rect 9232 8588 9352 8616
rect 9128 8288 9180 8294
rect 9128 8230 9180 8236
rect 9128 7880 9180 7886
rect 9128 7822 9180 7828
rect 9036 7744 9088 7750
rect 9036 7686 9088 7692
rect 9048 7410 9076 7686
rect 8944 7404 8996 7410
rect 8944 7346 8996 7352
rect 9036 7404 9088 7410
rect 9036 7346 9088 7352
rect 9140 7342 9168 7822
rect 9128 7336 9180 7342
rect 9128 7278 9180 7284
rect 8852 7200 8904 7206
rect 8852 7142 8904 7148
rect 8760 6452 8812 6458
rect 8760 6394 8812 6400
rect 8576 6384 8628 6390
rect 8576 6326 8628 6332
rect 7748 6316 7800 6322
rect 7748 6258 7800 6264
rect 7760 5914 7788 6258
rect 7932 6180 7984 6186
rect 7932 6122 7984 6128
rect 7840 6112 7892 6118
rect 7840 6054 7892 6060
rect 7852 5914 7880 6054
rect 7748 5908 7800 5914
rect 7748 5850 7800 5856
rect 7840 5908 7892 5914
rect 7840 5850 7892 5856
rect 7656 5772 7708 5778
rect 7656 5714 7708 5720
rect 7840 5772 7892 5778
rect 7840 5714 7892 5720
rect 7852 5370 7880 5714
rect 7944 5710 7972 6122
rect 8392 6112 8444 6118
rect 8392 6054 8444 6060
rect 8116 5840 8168 5846
rect 8116 5782 8168 5788
rect 7932 5704 7984 5710
rect 7932 5646 7984 5652
rect 8024 5568 8076 5574
rect 8024 5510 8076 5516
rect 7840 5364 7892 5370
rect 7840 5306 7892 5312
rect 8036 5302 8064 5510
rect 8024 5296 8076 5302
rect 8024 5238 8076 5244
rect 7748 5160 7800 5166
rect 7748 5102 7800 5108
rect 7380 4752 7432 4758
rect 7380 4694 7432 4700
rect 7760 4690 7788 5102
rect 7748 4684 7800 4690
rect 7748 4626 7800 4632
rect 7012 4276 7064 4282
rect 7012 4218 7064 4224
rect 7104 4276 7156 4282
rect 7104 4218 7156 4224
rect 7012 4140 7064 4146
rect 7012 4082 7064 4088
rect 6920 3120 6972 3126
rect 6920 3062 6972 3068
rect 7024 3058 7052 4082
rect 7116 3738 7144 4218
rect 7196 4140 7248 4146
rect 7196 4082 7248 4088
rect 7104 3732 7156 3738
rect 7104 3674 7156 3680
rect 7208 3058 7236 4082
rect 7760 4078 7788 4626
rect 7932 4548 7984 4554
rect 7932 4490 7984 4496
rect 7748 4072 7800 4078
rect 7748 4014 7800 4020
rect 7760 3602 7788 4014
rect 7748 3596 7800 3602
rect 7748 3538 7800 3544
rect 7564 3460 7616 3466
rect 7564 3402 7616 3408
rect 7380 3120 7432 3126
rect 7300 3080 7380 3108
rect 7012 3052 7064 3058
rect 7012 2994 7064 3000
rect 7196 3052 7248 3058
rect 7196 2994 7248 3000
rect 6736 2984 6788 2990
rect 6736 2926 6788 2932
rect 6644 2100 6696 2106
rect 6644 2042 6696 2048
rect 6656 1970 6684 2042
rect 6552 1964 6604 1970
rect 6552 1906 6604 1912
rect 6644 1964 6696 1970
rect 6644 1906 6696 1912
rect 6460 1896 6512 1902
rect 6460 1838 6512 1844
rect 6472 1426 6500 1838
rect 6460 1420 6512 1426
rect 6460 1362 6512 1368
rect 6656 1358 6684 1906
rect 6748 1902 6776 2926
rect 7104 2576 7156 2582
rect 7102 2544 7104 2553
rect 7156 2544 7158 2553
rect 7300 2514 7328 3080
rect 7380 3062 7432 3068
rect 7380 2984 7432 2990
rect 7380 2926 7432 2932
rect 7102 2479 7158 2488
rect 7288 2508 7340 2514
rect 7288 2450 7340 2456
rect 7288 2372 7340 2378
rect 7288 2314 7340 2320
rect 7300 2106 7328 2314
rect 7288 2100 7340 2106
rect 7288 2042 7340 2048
rect 6736 1896 6788 1902
rect 6736 1838 6788 1844
rect 7196 1896 7248 1902
rect 7196 1838 7248 1844
rect 7208 1562 7236 1838
rect 7196 1556 7248 1562
rect 7196 1498 7248 1504
rect 5816 1352 5868 1358
rect 5736 1312 5816 1340
rect 5816 1294 5868 1300
rect 6644 1352 6696 1358
rect 6644 1294 6696 1300
rect 7392 1290 7420 2926
rect 7576 2514 7604 3402
rect 7944 3194 7972 4490
rect 8128 4078 8156 5782
rect 8404 5710 8432 6054
rect 8392 5704 8444 5710
rect 8392 5646 8444 5652
rect 8576 5568 8628 5574
rect 8576 5510 8628 5516
rect 8214 5468 8522 5477
rect 8214 5466 8220 5468
rect 8276 5466 8300 5468
rect 8356 5466 8380 5468
rect 8436 5466 8460 5468
rect 8516 5466 8522 5468
rect 8276 5414 8278 5466
rect 8458 5414 8460 5466
rect 8214 5412 8220 5414
rect 8276 5412 8300 5414
rect 8356 5412 8380 5414
rect 8436 5412 8460 5414
rect 8516 5412 8522 5414
rect 8214 5403 8522 5412
rect 8588 4554 8616 5510
rect 8668 5296 8720 5302
rect 8668 5238 8720 5244
rect 8576 4548 8628 4554
rect 8576 4490 8628 4496
rect 8214 4380 8522 4389
rect 8214 4378 8220 4380
rect 8276 4378 8300 4380
rect 8356 4378 8380 4380
rect 8436 4378 8460 4380
rect 8516 4378 8522 4380
rect 8276 4326 8278 4378
rect 8458 4326 8460 4378
rect 8214 4324 8220 4326
rect 8276 4324 8300 4326
rect 8356 4324 8380 4326
rect 8436 4324 8460 4326
rect 8516 4324 8522 4326
rect 8214 4315 8522 4324
rect 8300 4208 8352 4214
rect 8352 4168 8432 4196
rect 8300 4150 8352 4156
rect 8404 4078 8432 4168
rect 8116 4072 8168 4078
rect 8116 4014 8168 4020
rect 8392 4072 8444 4078
rect 8392 4014 8444 4020
rect 8116 3936 8168 3942
rect 8116 3878 8168 3884
rect 8128 3516 8156 3878
rect 8680 3670 8708 5238
rect 8760 4820 8812 4826
rect 8760 4762 8812 4768
rect 8668 3664 8720 3670
rect 8668 3606 8720 3612
rect 8772 3602 8800 4762
rect 8864 4622 8892 7142
rect 9232 6458 9260 8588
rect 9312 8492 9364 8498
rect 9312 8434 9364 8440
rect 9324 6458 9352 8434
rect 9416 7886 9444 8774
rect 9784 8498 9812 8842
rect 9496 8492 9548 8498
rect 9496 8434 9548 8440
rect 9772 8492 9824 8498
rect 9772 8434 9824 8440
rect 9508 7954 9536 8434
rect 9864 8424 9916 8430
rect 9864 8366 9916 8372
rect 9588 8288 9640 8294
rect 9588 8230 9640 8236
rect 9772 8288 9824 8294
rect 9772 8230 9824 8236
rect 9496 7948 9548 7954
rect 9496 7890 9548 7896
rect 9404 7880 9456 7886
rect 9404 7822 9456 7828
rect 9496 7812 9548 7818
rect 9496 7754 9548 7760
rect 9404 7540 9456 7546
rect 9404 7482 9456 7488
rect 9416 6798 9444 7482
rect 9508 7206 9536 7754
rect 9496 7200 9548 7206
rect 9496 7142 9548 7148
rect 9404 6792 9456 6798
rect 9404 6734 9456 6740
rect 9220 6452 9272 6458
rect 9220 6394 9272 6400
rect 9312 6452 9364 6458
rect 9312 6394 9364 6400
rect 9128 5092 9180 5098
rect 9128 5034 9180 5040
rect 8852 4616 8904 4622
rect 8852 4558 8904 4564
rect 9036 4208 9088 4214
rect 9036 4150 9088 4156
rect 9048 3670 9076 4150
rect 9036 3664 9088 3670
rect 9036 3606 9088 3612
rect 9140 3602 9168 5034
rect 9220 4480 9272 4486
rect 9220 4422 9272 4428
rect 8760 3596 8812 3602
rect 8760 3538 8812 3544
rect 9128 3596 9180 3602
rect 9128 3538 9180 3544
rect 8208 3528 8260 3534
rect 8128 3488 8208 3516
rect 7932 3188 7984 3194
rect 7932 3130 7984 3136
rect 8128 3126 8156 3488
rect 8208 3470 8260 3476
rect 8576 3528 8628 3534
rect 8576 3470 8628 3476
rect 9036 3528 9088 3534
rect 9036 3470 9088 3476
rect 8214 3292 8522 3301
rect 8214 3290 8220 3292
rect 8276 3290 8300 3292
rect 8356 3290 8380 3292
rect 8436 3290 8460 3292
rect 8516 3290 8522 3292
rect 8276 3238 8278 3290
rect 8458 3238 8460 3290
rect 8214 3236 8220 3238
rect 8276 3236 8300 3238
rect 8356 3236 8380 3238
rect 8436 3236 8460 3238
rect 8516 3236 8522 3238
rect 8214 3227 8522 3236
rect 8588 3194 8616 3470
rect 8760 3392 8812 3398
rect 8760 3334 8812 3340
rect 8772 3194 8800 3334
rect 8576 3188 8628 3194
rect 8576 3130 8628 3136
rect 8760 3188 8812 3194
rect 8760 3130 8812 3136
rect 8116 3120 8168 3126
rect 8116 3062 8168 3068
rect 8300 2984 8352 2990
rect 8300 2926 8352 2932
rect 8024 2916 8076 2922
rect 8024 2858 8076 2864
rect 8036 2802 8064 2858
rect 8208 2848 8260 2854
rect 8036 2796 8208 2802
rect 8036 2790 8260 2796
rect 8036 2774 8248 2790
rect 7748 2644 7800 2650
rect 7748 2586 7800 2592
rect 7564 2508 7616 2514
rect 7564 2450 7616 2456
rect 7472 2440 7524 2446
rect 7472 2382 7524 2388
rect 7484 1970 7512 2382
rect 7656 2372 7708 2378
rect 7656 2314 7708 2320
rect 7668 1970 7696 2314
rect 7760 2106 7788 2586
rect 8036 2446 8064 2774
rect 8312 2666 8340 2926
rect 8128 2638 8340 2666
rect 8024 2440 8076 2446
rect 8024 2382 8076 2388
rect 7748 2100 7800 2106
rect 7748 2042 7800 2048
rect 7472 1964 7524 1970
rect 7472 1906 7524 1912
rect 7656 1964 7708 1970
rect 7656 1906 7708 1912
rect 7668 1426 7696 1906
rect 7760 1562 7788 2042
rect 8128 2038 8156 2638
rect 8482 2544 8538 2553
rect 8588 2530 8616 3130
rect 9048 2922 9076 3470
rect 9128 3392 9180 3398
rect 9128 3334 9180 3340
rect 9036 2916 9088 2922
rect 9036 2858 9088 2864
rect 9140 2650 9168 3334
rect 9232 3058 9260 4422
rect 9600 4078 9628 8230
rect 9784 8129 9812 8230
rect 9770 8120 9826 8129
rect 9692 8078 9770 8106
rect 9692 7410 9720 8078
rect 9770 8055 9826 8064
rect 9770 7848 9826 7857
rect 9770 7783 9826 7792
rect 9680 7404 9732 7410
rect 9784 7392 9812 7783
rect 9876 7750 9904 8366
rect 9864 7744 9916 7750
rect 9864 7686 9916 7692
rect 9968 7546 9996 10066
rect 10048 10056 10100 10062
rect 10046 10024 10048 10033
rect 10100 10024 10102 10033
rect 10046 9959 10102 9968
rect 10138 9752 10194 9761
rect 10138 9687 10194 9696
rect 10152 9450 10180 9687
rect 10140 9444 10192 9450
rect 10140 9386 10192 9392
rect 10244 9178 10272 10254
rect 10324 10260 10376 10266
rect 10324 10202 10376 10208
rect 10336 9722 10364 10202
rect 10612 10198 10640 10503
rect 10600 10192 10652 10198
rect 10600 10134 10652 10140
rect 10704 10130 10732 10542
rect 10692 10124 10744 10130
rect 10692 10066 10744 10072
rect 10416 10056 10468 10062
rect 10416 9998 10468 10004
rect 10324 9716 10376 9722
rect 10324 9658 10376 9664
rect 10324 9580 10376 9586
rect 10428 9568 10456 9998
rect 10508 9920 10560 9926
rect 10508 9862 10560 9868
rect 10376 9540 10456 9568
rect 10324 9522 10376 9528
rect 10140 9172 10192 9178
rect 10140 9114 10192 9120
rect 10232 9172 10284 9178
rect 10232 9114 10284 9120
rect 10046 8392 10102 8401
rect 10046 8327 10102 8336
rect 10060 8294 10088 8327
rect 10048 8288 10100 8294
rect 10048 8230 10100 8236
rect 10152 8090 10180 9114
rect 10232 8968 10284 8974
rect 10232 8910 10284 8916
rect 10244 8265 10272 8910
rect 10336 8634 10364 9522
rect 10416 9444 10468 9450
rect 10416 9386 10468 9392
rect 10428 8974 10456 9386
rect 10416 8968 10468 8974
rect 10416 8910 10468 8916
rect 10520 8838 10548 9862
rect 10704 9654 10732 10066
rect 10796 9761 10824 11591
rect 10876 11552 10928 11558
rect 10876 11494 10928 11500
rect 10782 9752 10838 9761
rect 10782 9687 10838 9696
rect 10692 9648 10744 9654
rect 10692 9590 10744 9596
rect 10600 9580 10652 9586
rect 10600 9522 10652 9528
rect 10612 8906 10640 9522
rect 10704 9466 10732 9590
rect 10704 9438 10824 9466
rect 10692 9376 10744 9382
rect 10690 9344 10692 9353
rect 10744 9344 10746 9353
rect 10690 9279 10746 9288
rect 10600 8900 10652 8906
rect 10600 8842 10652 8848
rect 10508 8832 10560 8838
rect 10508 8774 10560 8780
rect 10520 8634 10548 8774
rect 10324 8628 10376 8634
rect 10324 8570 10376 8576
rect 10508 8628 10560 8634
rect 10508 8570 10560 8576
rect 10336 8378 10364 8570
rect 10416 8560 10468 8566
rect 10468 8508 10548 8514
rect 10416 8502 10548 8508
rect 10428 8486 10548 8502
rect 10704 8498 10732 9279
rect 10796 9110 10824 9438
rect 10784 9104 10836 9110
rect 10784 9046 10836 9052
rect 10888 8974 10916 11494
rect 10980 11286 11008 13262
rect 11256 12918 11284 13262
rect 11244 12912 11296 12918
rect 11244 12854 11296 12860
rect 11532 12850 11560 13262
rect 11612 12980 11664 12986
rect 11612 12922 11664 12928
rect 11520 12844 11572 12850
rect 11520 12786 11572 12792
rect 11532 12374 11560 12786
rect 11520 12368 11572 12374
rect 11520 12310 11572 12316
rect 11624 12238 11652 12922
rect 11520 12232 11572 12238
rect 11520 12174 11572 12180
rect 11612 12232 11664 12238
rect 11612 12174 11664 12180
rect 11336 12164 11388 12170
rect 11336 12106 11388 12112
rect 11060 11756 11112 11762
rect 11060 11698 11112 11704
rect 11072 11286 11100 11698
rect 11348 11694 11376 12106
rect 11428 11824 11480 11830
rect 11428 11766 11480 11772
rect 11336 11688 11388 11694
rect 11336 11630 11388 11636
rect 11440 11506 11468 11766
rect 11532 11762 11560 12174
rect 11520 11756 11572 11762
rect 11520 11698 11572 11704
rect 11348 11478 11468 11506
rect 10968 11280 11020 11286
rect 10968 11222 11020 11228
rect 11060 11280 11112 11286
rect 11060 11222 11112 11228
rect 10980 10470 11008 11222
rect 11072 11150 11100 11222
rect 11060 11144 11112 11150
rect 11060 11086 11112 11092
rect 11072 10742 11100 11086
rect 11150 10976 11206 10985
rect 11150 10911 11206 10920
rect 11164 10826 11192 10911
rect 11164 10810 11284 10826
rect 11164 10804 11296 10810
rect 11164 10798 11244 10804
rect 11244 10746 11296 10752
rect 11060 10736 11112 10742
rect 11060 10678 11112 10684
rect 11244 10668 11296 10674
rect 11164 10628 11244 10656
rect 11060 10600 11112 10606
rect 11060 10542 11112 10548
rect 10968 10464 11020 10470
rect 11072 10441 11100 10542
rect 10968 10406 11020 10412
rect 11058 10432 11114 10441
rect 11058 10367 11114 10376
rect 10968 10056 11020 10062
rect 10966 10024 10968 10033
rect 11020 10024 11022 10033
rect 10966 9959 11022 9968
rect 10980 9722 11008 9959
rect 10968 9716 11020 9722
rect 10968 9658 11020 9664
rect 11058 9616 11114 9625
rect 11058 9551 11114 9560
rect 10968 9444 11020 9450
rect 10968 9386 11020 9392
rect 10784 8968 10836 8974
rect 10784 8910 10836 8916
rect 10876 8968 10928 8974
rect 10876 8910 10928 8916
rect 10336 8350 10456 8378
rect 10324 8288 10376 8294
rect 10230 8256 10286 8265
rect 10324 8230 10376 8236
rect 10230 8191 10286 8200
rect 10048 8084 10100 8090
rect 10048 8026 10100 8032
rect 10140 8084 10192 8090
rect 10140 8026 10192 8032
rect 10232 8084 10284 8090
rect 10336 8072 10364 8230
rect 10284 8044 10364 8072
rect 10232 8026 10284 8032
rect 10060 7936 10088 8026
rect 10428 8022 10456 8350
rect 10416 8016 10468 8022
rect 10230 7984 10286 7993
rect 10060 7908 10180 7936
rect 10230 7919 10286 7928
rect 10414 7984 10416 7993
rect 10468 7984 10470 7993
rect 10414 7919 10470 7928
rect 9956 7540 10008 7546
rect 9956 7482 10008 7488
rect 9864 7404 9916 7410
rect 9784 7364 9864 7392
rect 9680 7346 9732 7352
rect 9864 7346 9916 7352
rect 9692 6798 9720 7346
rect 10046 7032 10102 7041
rect 10046 6967 10102 6976
rect 9680 6792 9732 6798
rect 9680 6734 9732 6740
rect 9956 6656 10008 6662
rect 9956 6598 10008 6604
rect 9968 6458 9996 6598
rect 9956 6452 10008 6458
rect 9956 6394 10008 6400
rect 9680 6180 9732 6186
rect 9680 6122 9732 6128
rect 9692 5710 9720 6122
rect 9772 6112 9824 6118
rect 9772 6054 9824 6060
rect 9680 5704 9732 5710
rect 9680 5646 9732 5652
rect 9784 4554 9812 6054
rect 9956 5908 10008 5914
rect 9956 5850 10008 5856
rect 9968 4690 9996 5850
rect 9956 4684 10008 4690
rect 9956 4626 10008 4632
rect 9772 4548 9824 4554
rect 9772 4490 9824 4496
rect 9588 4072 9640 4078
rect 9588 4014 9640 4020
rect 9680 3936 9732 3942
rect 9680 3878 9732 3884
rect 9692 3670 9720 3878
rect 9680 3664 9732 3670
rect 9680 3606 9732 3612
rect 9496 3528 9548 3534
rect 9496 3470 9548 3476
rect 9220 3052 9272 3058
rect 9220 2994 9272 3000
rect 9508 2990 9536 3470
rect 10060 3466 10088 6967
rect 10152 6934 10180 7908
rect 10140 6928 10192 6934
rect 10140 6870 10192 6876
rect 10244 5370 10272 7919
rect 10520 7410 10548 8486
rect 10692 8492 10744 8498
rect 10692 8434 10744 8440
rect 10690 8120 10746 8129
rect 10690 8055 10746 8064
rect 10598 7984 10654 7993
rect 10704 7954 10732 8055
rect 10796 7993 10824 8910
rect 10888 8566 10916 8910
rect 10876 8560 10928 8566
rect 10876 8502 10928 8508
rect 10876 8016 10928 8022
rect 10782 7984 10838 7993
rect 10598 7919 10654 7928
rect 10692 7948 10744 7954
rect 10508 7404 10560 7410
rect 10508 7346 10560 7352
rect 10416 7336 10468 7342
rect 10416 7278 10468 7284
rect 10428 6934 10456 7278
rect 10416 6928 10468 6934
rect 10416 6870 10468 6876
rect 10612 6798 10640 7919
rect 10876 7958 10928 7964
rect 10782 7919 10838 7928
rect 10692 7890 10744 7896
rect 10782 7848 10838 7857
rect 10692 7812 10744 7818
rect 10782 7783 10838 7792
rect 10692 7754 10744 7760
rect 10704 7721 10732 7754
rect 10690 7712 10746 7721
rect 10690 7647 10746 7656
rect 10796 6798 10824 7783
rect 10888 6934 10916 7958
rect 10876 6928 10928 6934
rect 10876 6870 10928 6876
rect 10324 6792 10376 6798
rect 10324 6734 10376 6740
rect 10600 6792 10652 6798
rect 10600 6734 10652 6740
rect 10784 6792 10836 6798
rect 10784 6734 10836 6740
rect 10336 6186 10364 6734
rect 10416 6656 10468 6662
rect 10416 6598 10468 6604
rect 10428 6254 10456 6598
rect 10508 6316 10560 6322
rect 10508 6258 10560 6264
rect 10416 6248 10468 6254
rect 10416 6190 10468 6196
rect 10324 6180 10376 6186
rect 10324 6122 10376 6128
rect 10232 5364 10284 5370
rect 10232 5306 10284 5312
rect 10140 5228 10192 5234
rect 10140 5170 10192 5176
rect 10152 4146 10180 5170
rect 10428 4826 10456 6190
rect 10520 5370 10548 6258
rect 10508 5364 10560 5370
rect 10508 5306 10560 5312
rect 10796 5234 10824 6734
rect 10980 6225 11008 9386
rect 11072 8974 11100 9551
rect 11164 9489 11192 10628
rect 11244 10610 11296 10616
rect 11244 9920 11296 9926
rect 11244 9862 11296 9868
rect 11150 9480 11206 9489
rect 11150 9415 11206 9424
rect 11152 9104 11204 9110
rect 11152 9046 11204 9052
rect 11060 8968 11112 8974
rect 11060 8910 11112 8916
rect 11072 8838 11100 8910
rect 11164 8906 11192 9046
rect 11152 8900 11204 8906
rect 11152 8842 11204 8848
rect 11060 8832 11112 8838
rect 11060 8774 11112 8780
rect 11072 8498 11100 8774
rect 11060 8492 11112 8498
rect 11060 8434 11112 8440
rect 11152 8492 11204 8498
rect 11152 8434 11204 8440
rect 11060 7880 11112 7886
rect 11058 7848 11060 7857
rect 11112 7848 11114 7857
rect 11058 7783 11114 7792
rect 11060 7404 11112 7410
rect 11060 7346 11112 7352
rect 11072 6390 11100 7346
rect 11164 7342 11192 8434
rect 11256 8362 11284 9862
rect 11348 8974 11376 11478
rect 11532 11354 11560 11698
rect 11624 11694 11652 12174
rect 11612 11688 11664 11694
rect 11612 11630 11664 11636
rect 11520 11348 11572 11354
rect 11520 11290 11572 11296
rect 11702 11248 11758 11257
rect 11702 11183 11758 11192
rect 11428 11144 11480 11150
rect 11428 11086 11480 11092
rect 11612 11144 11664 11150
rect 11612 11086 11664 11092
rect 11440 9994 11468 11086
rect 11520 10192 11572 10198
rect 11520 10134 11572 10140
rect 11428 9988 11480 9994
rect 11428 9930 11480 9936
rect 11428 9580 11480 9586
rect 11428 9522 11480 9528
rect 11440 9353 11468 9522
rect 11426 9344 11482 9353
rect 11426 9279 11482 9288
rect 11336 8968 11388 8974
rect 11336 8910 11388 8916
rect 11244 8356 11296 8362
rect 11244 8298 11296 8304
rect 11244 7880 11296 7886
rect 11244 7822 11296 7828
rect 11152 7336 11204 7342
rect 11152 7278 11204 7284
rect 11164 6662 11192 7278
rect 11256 7274 11284 7822
rect 11244 7268 11296 7274
rect 11244 7210 11296 7216
rect 11244 6792 11296 6798
rect 11244 6734 11296 6740
rect 11152 6656 11204 6662
rect 11152 6598 11204 6604
rect 11256 6390 11284 6734
rect 11060 6384 11112 6390
rect 11060 6326 11112 6332
rect 11244 6384 11296 6390
rect 11244 6326 11296 6332
rect 11152 6248 11204 6254
rect 10966 6216 11022 6225
rect 11348 6202 11376 8910
rect 11428 8900 11480 8906
rect 11428 8842 11480 8848
rect 11440 8430 11468 8842
rect 11532 8498 11560 10134
rect 11624 9178 11652 11086
rect 11716 11082 11744 11183
rect 11704 11076 11756 11082
rect 11704 11018 11756 11024
rect 11716 9874 11744 11018
rect 11808 10674 11836 14334
rect 12070 14200 12126 14334
rect 13174 14200 13230 15000
rect 14370 14200 14426 15000
rect 12214 13628 12522 13637
rect 12214 13626 12220 13628
rect 12276 13626 12300 13628
rect 12356 13626 12380 13628
rect 12436 13626 12460 13628
rect 12516 13626 12522 13628
rect 12276 13574 12278 13626
rect 12458 13574 12460 13626
rect 12214 13572 12220 13574
rect 12276 13572 12300 13574
rect 12356 13572 12380 13574
rect 12436 13572 12460 13574
rect 12516 13572 12522 13574
rect 12214 13563 12522 13572
rect 11980 13456 12032 13462
rect 11980 13398 12032 13404
rect 11888 13184 11940 13190
rect 11888 13126 11940 13132
rect 11900 12850 11928 13126
rect 11888 12844 11940 12850
rect 11888 12786 11940 12792
rect 11900 12238 11928 12786
rect 11888 12232 11940 12238
rect 11888 12174 11940 12180
rect 11888 12096 11940 12102
rect 11888 12038 11940 12044
rect 11900 10996 11928 12038
rect 11992 11830 12020 13398
rect 12072 13252 12124 13258
rect 12072 13194 12124 13200
rect 12084 12918 12112 13194
rect 13084 13184 13136 13190
rect 13084 13126 13136 13132
rect 12072 12912 12124 12918
rect 12072 12854 12124 12860
rect 12214 12540 12522 12549
rect 12214 12538 12220 12540
rect 12276 12538 12300 12540
rect 12356 12538 12380 12540
rect 12436 12538 12460 12540
rect 12516 12538 12522 12540
rect 12276 12486 12278 12538
rect 12458 12486 12460 12538
rect 12214 12484 12220 12486
rect 12276 12484 12300 12486
rect 12356 12484 12380 12486
rect 12436 12484 12460 12486
rect 12516 12484 12522 12486
rect 12214 12475 12522 12484
rect 13096 11830 13124 13126
rect 13188 12306 13216 14200
rect 13452 13320 13504 13326
rect 13452 13262 13504 13268
rect 13268 13252 13320 13258
rect 13268 13194 13320 13200
rect 13280 12646 13308 13194
rect 13360 13184 13412 13190
rect 13360 13126 13412 13132
rect 13268 12640 13320 12646
rect 13268 12582 13320 12588
rect 13176 12300 13228 12306
rect 13176 12242 13228 12248
rect 13280 12238 13308 12582
rect 13268 12232 13320 12238
rect 13268 12174 13320 12180
rect 11980 11824 12032 11830
rect 11980 11766 12032 11772
rect 13084 11824 13136 11830
rect 13084 11766 13136 11772
rect 12624 11688 12676 11694
rect 12624 11630 12676 11636
rect 12214 11452 12522 11461
rect 12214 11450 12220 11452
rect 12276 11450 12300 11452
rect 12356 11450 12380 11452
rect 12436 11450 12460 11452
rect 12516 11450 12522 11452
rect 12276 11398 12278 11450
rect 12458 11398 12460 11450
rect 12214 11396 12220 11398
rect 12276 11396 12300 11398
rect 12356 11396 12380 11398
rect 12436 11396 12460 11398
rect 12516 11396 12522 11398
rect 12214 11387 12522 11396
rect 12636 11150 12664 11630
rect 12992 11620 13044 11626
rect 12992 11562 13044 11568
rect 12716 11552 12768 11558
rect 12716 11494 12768 11500
rect 12624 11144 12676 11150
rect 12624 11086 12676 11092
rect 11980 11008 12032 11014
rect 11900 10968 11980 10996
rect 11980 10950 12032 10956
rect 12254 10976 12310 10985
rect 11796 10668 11848 10674
rect 11796 10610 11848 10616
rect 11808 9994 11836 10610
rect 11888 10532 11940 10538
rect 11888 10474 11940 10480
rect 11900 10266 11928 10474
rect 11888 10260 11940 10266
rect 11888 10202 11940 10208
rect 11796 9988 11848 9994
rect 11796 9930 11848 9936
rect 11716 9846 11836 9874
rect 11702 9752 11758 9761
rect 11702 9687 11758 9696
rect 11612 9172 11664 9178
rect 11612 9114 11664 9120
rect 11610 8528 11666 8537
rect 11520 8492 11572 8498
rect 11610 8463 11612 8472
rect 11520 8434 11572 8440
rect 11664 8463 11666 8472
rect 11612 8434 11664 8440
rect 11428 8424 11480 8430
rect 11428 8366 11480 8372
rect 11440 7886 11468 8366
rect 11716 7970 11744 9687
rect 11532 7942 11744 7970
rect 11428 7880 11480 7886
rect 11428 7822 11480 7828
rect 11428 7540 11480 7546
rect 11428 7482 11480 7488
rect 11440 7041 11468 7482
rect 11426 7032 11482 7041
rect 11426 6967 11482 6976
rect 11532 6882 11560 7942
rect 11612 7880 11664 7886
rect 11612 7822 11664 7828
rect 11624 7410 11652 7822
rect 11704 7812 11756 7818
rect 11704 7754 11756 7760
rect 11716 7410 11744 7754
rect 11612 7404 11664 7410
rect 11612 7346 11664 7352
rect 11704 7404 11756 7410
rect 11704 7346 11756 7352
rect 11440 6854 11560 6882
rect 11440 6254 11468 6854
rect 11520 6724 11572 6730
rect 11520 6666 11572 6672
rect 11532 6458 11560 6666
rect 11520 6452 11572 6458
rect 11520 6394 11572 6400
rect 11152 6190 11204 6196
rect 10966 6151 11022 6160
rect 11164 5914 11192 6190
rect 11256 6174 11376 6202
rect 11428 6248 11480 6254
rect 11428 6190 11480 6196
rect 11152 5908 11204 5914
rect 11152 5850 11204 5856
rect 11164 5658 11192 5850
rect 11072 5630 11192 5658
rect 11072 5234 11100 5630
rect 10784 5228 10836 5234
rect 10784 5170 10836 5176
rect 11060 5228 11112 5234
rect 11060 5170 11112 5176
rect 11152 5092 11204 5098
rect 11152 5034 11204 5040
rect 10416 4820 10468 4826
rect 10416 4762 10468 4768
rect 11164 4554 11192 5034
rect 10600 4548 10652 4554
rect 10600 4490 10652 4496
rect 11152 4548 11204 4554
rect 11152 4490 11204 4496
rect 10612 4282 10640 4490
rect 10600 4276 10652 4282
rect 10600 4218 10652 4224
rect 10140 4140 10192 4146
rect 10140 4082 10192 4088
rect 10508 4004 10560 4010
rect 10508 3946 10560 3952
rect 10048 3460 10100 3466
rect 10048 3402 10100 3408
rect 9496 2984 9548 2990
rect 9496 2926 9548 2932
rect 9220 2916 9272 2922
rect 9220 2858 9272 2864
rect 9128 2644 9180 2650
rect 9128 2586 9180 2592
rect 8588 2502 8708 2530
rect 8482 2479 8484 2488
rect 8536 2479 8538 2488
rect 8484 2450 8536 2456
rect 8576 2440 8628 2446
rect 8576 2382 8628 2388
rect 8214 2204 8522 2213
rect 8214 2202 8220 2204
rect 8276 2202 8300 2204
rect 8356 2202 8380 2204
rect 8436 2202 8460 2204
rect 8516 2202 8522 2204
rect 8276 2150 8278 2202
rect 8458 2150 8460 2202
rect 8214 2148 8220 2150
rect 8276 2148 8300 2150
rect 8356 2148 8380 2150
rect 8436 2148 8460 2150
rect 8516 2148 8522 2150
rect 8214 2139 8522 2148
rect 8116 2032 8168 2038
rect 8116 1974 8168 1980
rect 7748 1556 7800 1562
rect 7748 1498 7800 1504
rect 7656 1420 7708 1426
rect 7656 1362 7708 1368
rect 8128 1290 8156 1974
rect 8588 1766 8616 2382
rect 8680 1902 8708 2502
rect 9128 2440 9180 2446
rect 9232 2428 9260 2858
rect 10520 2854 10548 3946
rect 11256 3670 11284 6174
rect 11336 5772 11388 5778
rect 11336 5714 11388 5720
rect 11348 5234 11376 5714
rect 11428 5636 11480 5642
rect 11428 5578 11480 5584
rect 11336 5228 11388 5234
rect 11336 5170 11388 5176
rect 11440 4758 11468 5578
rect 11624 5370 11652 7346
rect 11808 6866 11836 9846
rect 11888 9580 11940 9586
rect 11992 9568 12020 10950
rect 12254 10911 12310 10920
rect 12164 10736 12216 10742
rect 12162 10704 12164 10713
rect 12216 10704 12218 10713
rect 12268 10674 12296 10911
rect 12440 10804 12492 10810
rect 12728 10792 12756 11494
rect 13004 11082 13032 11562
rect 13280 11150 13308 12174
rect 13084 11144 13136 11150
rect 13084 11086 13136 11092
rect 13268 11144 13320 11150
rect 13268 11086 13320 11092
rect 12992 11076 13044 11082
rect 12992 11018 13044 11024
rect 12492 10764 12756 10792
rect 12440 10746 12492 10752
rect 12162 10639 12218 10648
rect 12256 10668 12308 10674
rect 12256 10610 12308 10616
rect 12072 10532 12124 10538
rect 12072 10474 12124 10480
rect 12084 10266 12112 10474
rect 12214 10364 12522 10373
rect 12214 10362 12220 10364
rect 12276 10362 12300 10364
rect 12356 10362 12380 10364
rect 12436 10362 12460 10364
rect 12516 10362 12522 10364
rect 12276 10310 12278 10362
rect 12458 10310 12460 10362
rect 12214 10308 12220 10310
rect 12276 10308 12300 10310
rect 12356 10308 12380 10310
rect 12436 10308 12460 10310
rect 12516 10308 12522 10310
rect 12214 10299 12522 10308
rect 12072 10260 12124 10266
rect 12072 10202 12124 10208
rect 12728 10112 12756 10764
rect 13096 10742 13124 11086
rect 13176 11008 13228 11014
rect 13176 10950 13228 10956
rect 13084 10736 13136 10742
rect 13084 10678 13136 10684
rect 12900 10668 12952 10674
rect 12900 10610 12952 10616
rect 12992 10668 13044 10674
rect 12992 10610 13044 10616
rect 12912 10577 12940 10610
rect 12898 10568 12954 10577
rect 12898 10503 12954 10512
rect 12636 10084 12756 10112
rect 12072 10056 12124 10062
rect 12072 9998 12124 10004
rect 12440 10056 12492 10062
rect 12636 10044 12664 10084
rect 12492 10016 12664 10044
rect 12808 10056 12860 10062
rect 12440 9998 12492 10004
rect 12808 9998 12860 10004
rect 11940 9540 12020 9568
rect 11888 9522 11940 9528
rect 11900 9178 11928 9522
rect 11980 9376 12032 9382
rect 11980 9318 12032 9324
rect 11888 9172 11940 9178
rect 11888 9114 11940 9120
rect 11992 8022 12020 9318
rect 12084 9217 12112 9998
rect 12452 9382 12480 9998
rect 12820 9586 12848 9998
rect 13004 9625 13032 10610
rect 13188 10198 13216 10950
rect 13176 10192 13228 10198
rect 13176 10134 13228 10140
rect 13188 9654 13216 10134
rect 13372 10130 13400 13126
rect 13464 11830 13492 13262
rect 14384 12714 14412 14200
rect 14372 12708 14424 12714
rect 14372 12650 14424 12656
rect 13452 11824 13504 11830
rect 13452 11766 13504 11772
rect 13360 10124 13412 10130
rect 13360 10066 13412 10072
rect 13464 9654 13492 11766
rect 13544 11076 13596 11082
rect 13544 11018 13596 11024
rect 13176 9648 13228 9654
rect 12990 9616 13046 9625
rect 12808 9580 12860 9586
rect 13176 9590 13228 9596
rect 13268 9648 13320 9654
rect 13268 9590 13320 9596
rect 13452 9648 13504 9654
rect 13452 9590 13504 9596
rect 12990 9551 13046 9560
rect 12808 9522 12860 9528
rect 12440 9376 12492 9382
rect 12440 9318 12492 9324
rect 12214 9276 12522 9285
rect 12214 9274 12220 9276
rect 12276 9274 12300 9276
rect 12356 9274 12380 9276
rect 12436 9274 12460 9276
rect 12516 9274 12522 9276
rect 12276 9222 12278 9274
rect 12458 9222 12460 9274
rect 12214 9220 12220 9222
rect 12276 9220 12300 9222
rect 12356 9220 12380 9222
rect 12436 9220 12460 9222
rect 12516 9220 12522 9222
rect 12070 9208 12126 9217
rect 12214 9211 12522 9220
rect 12070 9143 12126 9152
rect 12164 9172 12216 9178
rect 12084 8838 12112 9143
rect 12164 9114 12216 9120
rect 12072 8832 12124 8838
rect 12072 8774 12124 8780
rect 12072 8356 12124 8362
rect 12072 8298 12124 8304
rect 11980 8016 12032 8022
rect 11980 7958 12032 7964
rect 11980 7880 12032 7886
rect 11900 7840 11980 7868
rect 11704 6860 11756 6866
rect 11704 6802 11756 6808
rect 11796 6860 11848 6866
rect 11796 6802 11848 6808
rect 11716 6322 11744 6802
rect 11796 6656 11848 6662
rect 11796 6598 11848 6604
rect 11704 6316 11756 6322
rect 11704 6258 11756 6264
rect 11716 5710 11744 6258
rect 11704 5704 11756 5710
rect 11704 5646 11756 5652
rect 11716 5370 11744 5646
rect 11612 5364 11664 5370
rect 11612 5306 11664 5312
rect 11704 5364 11756 5370
rect 11704 5306 11756 5312
rect 11808 5302 11836 6598
rect 11900 5914 11928 7840
rect 11980 7822 12032 7828
rect 11980 7744 12032 7750
rect 11980 7686 12032 7692
rect 11992 6798 12020 7686
rect 11980 6792 12032 6798
rect 11980 6734 12032 6740
rect 11980 6656 12032 6662
rect 11980 6598 12032 6604
rect 11992 6322 12020 6598
rect 11980 6316 12032 6322
rect 11980 6258 12032 6264
rect 11888 5908 11940 5914
rect 11888 5850 11940 5856
rect 12084 5710 12112 8298
rect 12176 8294 12204 9114
rect 13280 8974 13308 9590
rect 13452 9376 13504 9382
rect 13452 9318 13504 9324
rect 12992 8968 13044 8974
rect 12992 8910 13044 8916
rect 13268 8968 13320 8974
rect 13268 8910 13320 8916
rect 12348 8832 12400 8838
rect 12348 8774 12400 8780
rect 12360 8430 12388 8774
rect 12716 8492 12768 8498
rect 12716 8434 12768 8440
rect 12348 8424 12400 8430
rect 12348 8366 12400 8372
rect 12164 8288 12216 8294
rect 12624 8288 12676 8294
rect 12164 8230 12216 8236
rect 12622 8256 12624 8265
rect 12676 8256 12678 8265
rect 12214 8188 12522 8197
rect 12622 8191 12678 8200
rect 12214 8186 12220 8188
rect 12276 8186 12300 8188
rect 12356 8186 12380 8188
rect 12436 8186 12460 8188
rect 12516 8186 12522 8188
rect 12276 8134 12278 8186
rect 12458 8134 12460 8186
rect 12214 8132 12220 8134
rect 12276 8132 12300 8134
rect 12356 8132 12380 8134
rect 12436 8132 12460 8134
rect 12516 8132 12522 8134
rect 12214 8123 12522 8132
rect 12624 8084 12676 8090
rect 12624 8026 12676 8032
rect 12164 7948 12216 7954
rect 12164 7890 12216 7896
rect 12256 7948 12308 7954
rect 12256 7890 12308 7896
rect 12176 7546 12204 7890
rect 12164 7540 12216 7546
rect 12164 7482 12216 7488
rect 12268 7410 12296 7890
rect 12256 7404 12308 7410
rect 12256 7346 12308 7352
rect 12214 7100 12522 7109
rect 12214 7098 12220 7100
rect 12276 7098 12300 7100
rect 12356 7098 12380 7100
rect 12436 7098 12460 7100
rect 12516 7098 12522 7100
rect 12276 7046 12278 7098
rect 12458 7046 12460 7098
rect 12214 7044 12220 7046
rect 12276 7044 12300 7046
rect 12356 7044 12380 7046
rect 12436 7044 12460 7046
rect 12516 7044 12522 7046
rect 12214 7035 12522 7044
rect 12256 6996 12308 7002
rect 12256 6938 12308 6944
rect 12268 6866 12296 6938
rect 12256 6860 12308 6866
rect 12256 6802 12308 6808
rect 12214 6012 12522 6021
rect 12214 6010 12220 6012
rect 12276 6010 12300 6012
rect 12356 6010 12380 6012
rect 12436 6010 12460 6012
rect 12516 6010 12522 6012
rect 12276 5958 12278 6010
rect 12458 5958 12460 6010
rect 12214 5956 12220 5958
rect 12276 5956 12300 5958
rect 12356 5956 12380 5958
rect 12436 5956 12460 5958
rect 12516 5956 12522 5958
rect 12214 5947 12522 5956
rect 12072 5704 12124 5710
rect 12072 5646 12124 5652
rect 11796 5296 11848 5302
rect 11796 5238 11848 5244
rect 11888 5296 11940 5302
rect 11888 5238 11940 5244
rect 11520 5228 11572 5234
rect 11520 5170 11572 5176
rect 11428 4752 11480 4758
rect 11428 4694 11480 4700
rect 11532 4690 11560 5170
rect 11520 4684 11572 4690
rect 11520 4626 11572 4632
rect 11612 4616 11664 4622
rect 11612 4558 11664 4564
rect 11428 4548 11480 4554
rect 11428 4490 11480 4496
rect 11520 4548 11572 4554
rect 11520 4490 11572 4496
rect 11336 4140 11388 4146
rect 11336 4082 11388 4088
rect 11244 3664 11296 3670
rect 11244 3606 11296 3612
rect 11348 3210 11376 4082
rect 11440 4078 11468 4490
rect 11428 4072 11480 4078
rect 11428 4014 11480 4020
rect 11532 4010 11560 4490
rect 11624 4214 11652 4558
rect 11796 4480 11848 4486
rect 11796 4422 11848 4428
rect 11612 4208 11664 4214
rect 11612 4150 11664 4156
rect 11520 4004 11572 4010
rect 11520 3946 11572 3952
rect 11532 3670 11560 3946
rect 11520 3664 11572 3670
rect 11520 3606 11572 3612
rect 11624 3534 11652 4150
rect 11808 4146 11836 4422
rect 11900 4282 11928 5238
rect 11980 4616 12032 4622
rect 11980 4558 12032 4564
rect 11888 4276 11940 4282
rect 11888 4218 11940 4224
rect 11796 4140 11848 4146
rect 11796 4082 11848 4088
rect 11704 3936 11756 3942
rect 11704 3878 11756 3884
rect 11716 3738 11744 3878
rect 11992 3738 12020 4558
rect 12084 4146 12112 5646
rect 12214 4924 12522 4933
rect 12214 4922 12220 4924
rect 12276 4922 12300 4924
rect 12356 4922 12380 4924
rect 12436 4922 12460 4924
rect 12516 4922 12522 4924
rect 12276 4870 12278 4922
rect 12458 4870 12460 4922
rect 12214 4868 12220 4870
rect 12276 4868 12300 4870
rect 12356 4868 12380 4870
rect 12436 4868 12460 4870
rect 12516 4868 12522 4870
rect 12214 4859 12522 4868
rect 12072 4140 12124 4146
rect 12072 4082 12124 4088
rect 12072 4004 12124 4010
rect 12072 3946 12124 3952
rect 11704 3732 11756 3738
rect 11704 3674 11756 3680
rect 11980 3732 12032 3738
rect 11980 3674 12032 3680
rect 11612 3528 11664 3534
rect 11612 3470 11664 3476
rect 11980 3528 12032 3534
rect 11980 3470 12032 3476
rect 11796 3392 11848 3398
rect 11796 3334 11848 3340
rect 11072 3194 11376 3210
rect 11808 3194 11836 3334
rect 11060 3188 11376 3194
rect 11112 3182 11376 3188
rect 11796 3188 11848 3194
rect 11060 3130 11112 3136
rect 11796 3130 11848 3136
rect 11888 3188 11940 3194
rect 11888 3130 11940 3136
rect 11244 3120 11296 3126
rect 11244 3062 11296 3068
rect 11060 3052 11112 3058
rect 11060 2994 11112 3000
rect 10508 2848 10560 2854
rect 10508 2790 10560 2796
rect 10140 2644 10192 2650
rect 10140 2586 10192 2592
rect 9180 2400 9260 2428
rect 9128 2382 9180 2388
rect 9140 2281 9168 2382
rect 9680 2304 9732 2310
rect 9126 2272 9182 2281
rect 9732 2252 9812 2258
rect 9680 2246 9812 2252
rect 9692 2230 9812 2246
rect 9126 2207 9182 2216
rect 9680 2100 9732 2106
rect 9680 2042 9732 2048
rect 9220 1964 9272 1970
rect 9220 1906 9272 1912
rect 8668 1896 8720 1902
rect 8668 1838 8720 1844
rect 8576 1760 8628 1766
rect 8576 1702 8628 1708
rect 8680 1340 8708 1838
rect 8760 1352 8812 1358
rect 8680 1312 8760 1340
rect 8760 1294 8812 1300
rect 3882 1255 3938 1264
rect 4620 1284 4672 1290
rect 4620 1226 4672 1232
rect 5448 1284 5500 1290
rect 5448 1226 5500 1232
rect 7380 1284 7432 1290
rect 7380 1226 7432 1232
rect 8116 1284 8168 1290
rect 8116 1226 8168 1232
rect 9232 1222 9260 1906
rect 9310 1864 9366 1873
rect 9310 1799 9312 1808
rect 9364 1799 9366 1808
rect 9312 1770 9364 1776
rect 9324 1358 9352 1770
rect 9692 1426 9720 2042
rect 9784 1562 9812 2230
rect 10152 2038 10180 2586
rect 10140 2032 10192 2038
rect 10140 1974 10192 1980
rect 10520 1970 10548 2790
rect 11072 2553 11100 2994
rect 11256 2689 11284 3062
rect 11900 3058 11928 3130
rect 11888 3052 11940 3058
rect 11888 2994 11940 3000
rect 11992 2990 12020 3470
rect 12084 3466 12112 3946
rect 12214 3836 12522 3845
rect 12214 3834 12220 3836
rect 12276 3834 12300 3836
rect 12356 3834 12380 3836
rect 12436 3834 12460 3836
rect 12516 3834 12522 3836
rect 12276 3782 12278 3834
rect 12458 3782 12460 3834
rect 12214 3780 12220 3782
rect 12276 3780 12300 3782
rect 12356 3780 12380 3782
rect 12436 3780 12460 3782
rect 12516 3780 12522 3782
rect 12214 3771 12522 3780
rect 12072 3460 12124 3466
rect 12072 3402 12124 3408
rect 11520 2984 11572 2990
rect 11520 2926 11572 2932
rect 11980 2984 12032 2990
rect 12164 2984 12216 2990
rect 11980 2926 12032 2932
rect 12084 2944 12164 2972
rect 11242 2680 11298 2689
rect 11242 2615 11298 2624
rect 11058 2544 11114 2553
rect 11058 2479 11114 2488
rect 11072 1970 11100 2479
rect 11256 1970 11284 2615
rect 11428 2440 11480 2446
rect 11428 2382 11480 2388
rect 10232 1964 10284 1970
rect 10232 1906 10284 1912
rect 10508 1964 10560 1970
rect 10508 1906 10560 1912
rect 11060 1964 11112 1970
rect 11060 1906 11112 1912
rect 11244 1964 11296 1970
rect 11244 1906 11296 1912
rect 10140 1828 10192 1834
rect 10140 1770 10192 1776
rect 9772 1556 9824 1562
rect 9772 1498 9824 1504
rect 9680 1420 9732 1426
rect 9680 1362 9732 1368
rect 9312 1352 9364 1358
rect 9312 1294 9364 1300
rect 10152 1290 10180 1770
rect 10140 1284 10192 1290
rect 10140 1226 10192 1232
rect 5908 1216 5960 1222
rect 5908 1158 5960 1164
rect 6092 1216 6144 1222
rect 6092 1158 6144 1164
rect 9220 1216 9272 1222
rect 9220 1158 9272 1164
rect 5920 1018 5948 1158
rect 5908 1012 5960 1018
rect 5908 954 5960 960
rect 3620 882 3740 898
rect 6104 882 6132 1158
rect 8214 1116 8522 1125
rect 8214 1114 8220 1116
rect 8276 1114 8300 1116
rect 8356 1114 8380 1116
rect 8436 1114 8460 1116
rect 8516 1114 8522 1116
rect 8276 1062 8278 1114
rect 8458 1062 8460 1114
rect 8214 1060 8220 1062
rect 8276 1060 8300 1062
rect 8356 1060 8380 1062
rect 8436 1060 8460 1062
rect 8516 1060 8522 1062
rect 8214 1051 8522 1060
rect 10244 1018 10272 1906
rect 10980 1562 11192 1578
rect 10968 1556 11192 1562
rect 11020 1550 11192 1556
rect 10968 1498 11020 1504
rect 10232 1012 10284 1018
rect 10232 954 10284 960
rect 3608 876 3740 882
rect 3660 870 3740 876
rect 3608 818 3660 824
rect 3712 800 3740 870
rect 6092 876 6144 882
rect 6092 818 6144 824
rect 11164 800 11192 1550
rect 11256 1426 11284 1906
rect 11440 1562 11468 2382
rect 11532 2378 11560 2926
rect 11888 2916 11940 2922
rect 11888 2858 11940 2864
rect 11900 2514 11928 2858
rect 11888 2508 11940 2514
rect 11888 2450 11940 2456
rect 11612 2440 11664 2446
rect 11612 2382 11664 2388
rect 11520 2372 11572 2378
rect 11520 2314 11572 2320
rect 11518 2272 11574 2281
rect 11518 2207 11574 2216
rect 11532 1970 11560 2207
rect 11624 2106 11652 2382
rect 11612 2100 11664 2106
rect 11612 2042 11664 2048
rect 11520 1964 11572 1970
rect 11520 1906 11572 1912
rect 11428 1556 11480 1562
rect 11428 1498 11480 1504
rect 11900 1494 11928 2450
rect 12084 2378 12112 2944
rect 12164 2926 12216 2932
rect 12214 2748 12522 2757
rect 12214 2746 12220 2748
rect 12276 2746 12300 2748
rect 12356 2746 12380 2748
rect 12436 2746 12460 2748
rect 12516 2746 12522 2748
rect 12276 2694 12278 2746
rect 12458 2694 12460 2746
rect 12214 2692 12220 2694
rect 12276 2692 12300 2694
rect 12356 2692 12380 2694
rect 12436 2692 12460 2694
rect 12516 2692 12522 2694
rect 12214 2683 12522 2692
rect 12636 2650 12664 8026
rect 12728 3777 12756 8434
rect 13004 8430 13032 8910
rect 13360 8900 13412 8906
rect 13360 8842 13412 8848
rect 12992 8424 13044 8430
rect 12992 8366 13044 8372
rect 13372 8362 13400 8842
rect 13464 8498 13492 9318
rect 13556 8566 13584 11018
rect 13728 10668 13780 10674
rect 13728 10610 13780 10616
rect 13636 10600 13688 10606
rect 13636 10542 13688 10548
rect 13648 8809 13676 10542
rect 13634 8800 13690 8809
rect 13634 8735 13690 8744
rect 13544 8560 13596 8566
rect 13544 8502 13596 8508
rect 13452 8492 13504 8498
rect 13452 8434 13504 8440
rect 13268 8356 13320 8362
rect 13268 8298 13320 8304
rect 13360 8356 13412 8362
rect 13360 8298 13412 8304
rect 12808 8288 12860 8294
rect 12808 8230 12860 8236
rect 12898 8256 12954 8265
rect 12820 7886 12848 8230
rect 12898 8191 12954 8200
rect 12808 7880 12860 7886
rect 12808 7822 12860 7828
rect 12820 7410 12848 7822
rect 12808 7404 12860 7410
rect 12808 7346 12860 7352
rect 12806 6352 12862 6361
rect 12806 6287 12862 6296
rect 12820 4078 12848 6287
rect 12808 4072 12860 4078
rect 12808 4014 12860 4020
rect 12714 3768 12770 3777
rect 12714 3703 12770 3712
rect 12912 3602 12940 8191
rect 13280 8090 13308 8298
rect 13268 8084 13320 8090
rect 13268 8026 13320 8032
rect 13176 7812 13228 7818
rect 13176 7754 13228 7760
rect 13188 7478 13216 7754
rect 13176 7472 13228 7478
rect 13174 7440 13176 7449
rect 13228 7440 13230 7449
rect 13174 7375 13230 7384
rect 13268 7336 13320 7342
rect 13268 7278 13320 7284
rect 13176 7268 13228 7274
rect 13176 7210 13228 7216
rect 13188 6866 13216 7210
rect 13176 6860 13228 6866
rect 13176 6802 13228 6808
rect 13176 6724 13228 6730
rect 13176 6666 13228 6672
rect 13188 6186 13216 6666
rect 13176 6180 13228 6186
rect 13176 6122 13228 6128
rect 13188 5794 13216 6122
rect 13280 5914 13308 7278
rect 13268 5908 13320 5914
rect 13268 5850 13320 5856
rect 13188 5766 13308 5794
rect 13280 5642 13308 5766
rect 12992 5636 13044 5642
rect 12992 5578 13044 5584
rect 13268 5636 13320 5642
rect 13268 5578 13320 5584
rect 13004 5030 13032 5578
rect 12992 5024 13044 5030
rect 12992 4966 13044 4972
rect 13004 4146 13032 4966
rect 13280 4622 13308 5578
rect 13268 4616 13320 4622
rect 13268 4558 13320 4564
rect 13084 4480 13136 4486
rect 13084 4422 13136 4428
rect 12992 4140 13044 4146
rect 12992 4082 13044 4088
rect 13096 3738 13124 4422
rect 13176 4072 13228 4078
rect 13176 4014 13228 4020
rect 13084 3732 13136 3738
rect 13084 3674 13136 3680
rect 12900 3596 12952 3602
rect 12900 3538 12952 3544
rect 12912 3194 12940 3538
rect 13188 3194 13216 4014
rect 12900 3188 12952 3194
rect 12900 3130 12952 3136
rect 13176 3188 13228 3194
rect 13176 3130 13228 3136
rect 13280 3058 13308 4558
rect 13372 4214 13400 8298
rect 13544 8084 13596 8090
rect 13544 8026 13596 8032
rect 13452 7880 13504 7886
rect 13452 7822 13504 7828
rect 13464 6322 13492 7822
rect 13452 6316 13504 6322
rect 13452 6258 13504 6264
rect 13464 5710 13492 6258
rect 13452 5704 13504 5710
rect 13452 5646 13504 5652
rect 13360 4208 13412 4214
rect 13360 4150 13412 4156
rect 13464 3942 13492 5646
rect 13452 3936 13504 3942
rect 13452 3878 13504 3884
rect 13360 3528 13412 3534
rect 13360 3470 13412 3476
rect 13268 3052 13320 3058
rect 13268 2994 13320 3000
rect 12624 2644 12676 2650
rect 12624 2586 12676 2592
rect 13372 2514 13400 3470
rect 13360 2508 13412 2514
rect 13360 2450 13412 2456
rect 13176 2440 13228 2446
rect 13176 2382 13228 2388
rect 12072 2372 12124 2378
rect 12072 2314 12124 2320
rect 11980 2304 12032 2310
rect 11980 2246 12032 2252
rect 11992 1766 12020 2246
rect 12992 1896 13044 1902
rect 12992 1838 13044 1844
rect 11980 1760 12032 1766
rect 11980 1702 12032 1708
rect 11888 1488 11940 1494
rect 11888 1430 11940 1436
rect 11244 1420 11296 1426
rect 11244 1362 11296 1368
rect 11992 1222 12020 1702
rect 12214 1660 12522 1669
rect 12214 1658 12220 1660
rect 12276 1658 12300 1660
rect 12356 1658 12380 1660
rect 12436 1658 12460 1660
rect 12516 1658 12522 1660
rect 12276 1606 12278 1658
rect 12458 1606 12460 1658
rect 12214 1604 12220 1606
rect 12276 1604 12300 1606
rect 12356 1604 12380 1606
rect 12436 1604 12460 1606
rect 12516 1604 12522 1606
rect 12214 1595 12522 1604
rect 13004 1562 13032 1838
rect 12992 1556 13044 1562
rect 12992 1498 13044 1504
rect 13188 1358 13216 2382
rect 13176 1352 13228 1358
rect 13556 1329 13584 8026
rect 13648 5370 13676 8735
rect 13740 7410 13768 10610
rect 13728 7404 13780 7410
rect 13728 7346 13780 7352
rect 13636 5364 13688 5370
rect 13636 5306 13688 5312
rect 13176 1294 13228 1300
rect 13542 1320 13598 1329
rect 13542 1255 13598 1264
rect 11520 1216 11572 1222
rect 11520 1158 11572 1164
rect 11980 1216 12032 1222
rect 11980 1158 12032 1164
rect 11532 950 11560 1158
rect 11520 944 11572 950
rect 11520 886 11572 892
rect 1398 504 1454 513
rect 1398 439 1454 448
rect 3698 0 3754 800
rect 11150 0 11206 800
<< via2 >>
rect 3238 14456 3294 14512
rect 1674 13368 1730 13424
rect 1398 12552 1454 12608
rect 1950 13504 2006 13560
rect 2870 13268 2872 13288
rect 2872 13268 2924 13288
rect 2924 13268 2926 13288
rect 2870 13232 2926 13268
rect 1950 12824 2006 12880
rect 1490 8880 1546 8936
rect 2410 11756 2466 11792
rect 2410 11736 2412 11756
rect 2412 11736 2464 11756
rect 2464 11736 2466 11756
rect 3054 11600 3110 11656
rect 4220 13626 4276 13628
rect 4300 13626 4356 13628
rect 4380 13626 4436 13628
rect 4460 13626 4516 13628
rect 4220 13574 4266 13626
rect 4266 13574 4276 13626
rect 4300 13574 4330 13626
rect 4330 13574 4342 13626
rect 4342 13574 4356 13626
rect 4380 13574 4394 13626
rect 4394 13574 4406 13626
rect 4406 13574 4436 13626
rect 4460 13574 4470 13626
rect 4470 13574 4516 13626
rect 4220 13572 4276 13574
rect 4300 13572 4356 13574
rect 4380 13572 4436 13574
rect 4460 13572 4516 13574
rect 3146 10784 3202 10840
rect 1398 5072 1454 5128
rect 2962 7928 3018 7984
rect 2594 6160 2650 6216
rect 2870 6976 2926 7032
rect 2962 6024 3018 6080
rect 1674 2388 1676 2408
rect 1676 2388 1728 2408
rect 1728 2388 1730 2408
rect 1674 2352 1730 2388
rect 1674 1964 1730 2000
rect 1674 1944 1676 1964
rect 1676 1944 1728 1964
rect 1728 1944 1730 1964
rect 2318 2508 2374 2544
rect 2318 2488 2320 2508
rect 2320 2488 2372 2508
rect 2372 2488 2374 2508
rect 2870 5208 2926 5264
rect 4220 12538 4276 12540
rect 4300 12538 4356 12540
rect 4380 12538 4436 12540
rect 4460 12538 4516 12540
rect 4220 12486 4266 12538
rect 4266 12486 4276 12538
rect 4300 12486 4330 12538
rect 4330 12486 4342 12538
rect 4342 12486 4356 12538
rect 4380 12486 4394 12538
rect 4394 12486 4406 12538
rect 4406 12486 4436 12538
rect 4460 12486 4470 12538
rect 4470 12486 4516 12538
rect 4220 12484 4276 12486
rect 4300 12484 4356 12486
rect 4380 12484 4436 12486
rect 4460 12484 4516 12486
rect 3974 12008 4030 12064
rect 3974 9696 4030 9752
rect 3790 9152 3846 9208
rect 3606 7928 3662 7984
rect 3882 8744 3938 8800
rect 3054 3168 3110 3224
rect 2778 2216 2834 2272
rect 4526 11600 4582 11656
rect 4220 11450 4276 11452
rect 4300 11450 4356 11452
rect 4380 11450 4436 11452
rect 4460 11450 4516 11452
rect 4220 11398 4266 11450
rect 4266 11398 4276 11450
rect 4300 11398 4330 11450
rect 4330 11398 4342 11450
rect 4342 11398 4356 11450
rect 4380 11398 4394 11450
rect 4394 11398 4406 11450
rect 4406 11398 4436 11450
rect 4460 11398 4470 11450
rect 4470 11398 4516 11450
rect 4220 11396 4276 11398
rect 4300 11396 4356 11398
rect 4380 11396 4436 11398
rect 4460 11396 4516 11398
rect 4220 10362 4276 10364
rect 4300 10362 4356 10364
rect 4380 10362 4436 10364
rect 4460 10362 4516 10364
rect 4220 10310 4266 10362
rect 4266 10310 4276 10362
rect 4300 10310 4330 10362
rect 4330 10310 4342 10362
rect 4342 10310 4356 10362
rect 4380 10310 4394 10362
rect 4394 10310 4406 10362
rect 4406 10310 4436 10362
rect 4460 10310 4470 10362
rect 4470 10310 4516 10362
rect 4220 10308 4276 10310
rect 4300 10308 4356 10310
rect 4380 10308 4436 10310
rect 4460 10308 4516 10310
rect 4802 11192 4858 11248
rect 4710 9968 4766 10024
rect 4220 9274 4276 9276
rect 4300 9274 4356 9276
rect 4380 9274 4436 9276
rect 4460 9274 4516 9276
rect 4220 9222 4266 9274
rect 4266 9222 4276 9274
rect 4300 9222 4330 9274
rect 4330 9222 4342 9274
rect 4342 9222 4356 9274
rect 4380 9222 4394 9274
rect 4394 9222 4406 9274
rect 4406 9222 4436 9274
rect 4460 9222 4470 9274
rect 4470 9222 4516 9274
rect 4220 9220 4276 9222
rect 4300 9220 4356 9222
rect 4380 9220 4436 9222
rect 4460 9220 4516 9222
rect 4220 8186 4276 8188
rect 4300 8186 4356 8188
rect 4380 8186 4436 8188
rect 4460 8186 4516 8188
rect 4220 8134 4266 8186
rect 4266 8134 4276 8186
rect 4300 8134 4330 8186
rect 4330 8134 4342 8186
rect 4342 8134 4356 8186
rect 4380 8134 4394 8186
rect 4394 8134 4406 8186
rect 4406 8134 4436 8186
rect 4460 8134 4470 8186
rect 4470 8134 4516 8186
rect 4220 8132 4276 8134
rect 4300 8132 4356 8134
rect 4380 8132 4436 8134
rect 4460 8132 4516 8134
rect 5078 8608 5134 8664
rect 5170 8064 5226 8120
rect 4220 7098 4276 7100
rect 4300 7098 4356 7100
rect 4380 7098 4436 7100
rect 4460 7098 4516 7100
rect 4220 7046 4266 7098
rect 4266 7046 4276 7098
rect 4300 7046 4330 7098
rect 4330 7046 4342 7098
rect 4342 7046 4356 7098
rect 4380 7046 4394 7098
rect 4394 7046 4406 7098
rect 4406 7046 4436 7098
rect 4460 7046 4470 7098
rect 4470 7046 4516 7098
rect 4220 7044 4276 7046
rect 4300 7044 4356 7046
rect 4380 7044 4436 7046
rect 4460 7044 4516 7046
rect 4250 6160 4306 6216
rect 3974 6024 4030 6080
rect 4220 6010 4276 6012
rect 4300 6010 4356 6012
rect 4380 6010 4436 6012
rect 4460 6010 4516 6012
rect 4220 5958 4266 6010
rect 4266 5958 4276 6010
rect 4300 5958 4330 6010
rect 4330 5958 4342 6010
rect 4342 5958 4356 6010
rect 4380 5958 4394 6010
rect 4394 5958 4406 6010
rect 4406 5958 4436 6010
rect 4460 5958 4470 6010
rect 4470 5958 4516 6010
rect 4220 5956 4276 5958
rect 4300 5956 4356 5958
rect 4380 5956 4436 5958
rect 4460 5956 4516 5958
rect 4618 5208 4674 5264
rect 4066 5072 4122 5128
rect 4220 4922 4276 4924
rect 4300 4922 4356 4924
rect 4380 4922 4436 4924
rect 4460 4922 4516 4924
rect 4220 4870 4266 4922
rect 4266 4870 4276 4922
rect 4300 4870 4330 4922
rect 4330 4870 4342 4922
rect 4342 4870 4356 4922
rect 4380 4870 4394 4922
rect 4394 4870 4406 4922
rect 4406 4870 4436 4922
rect 4460 4870 4470 4922
rect 4470 4870 4516 4922
rect 4220 4868 4276 4870
rect 4300 4868 4356 4870
rect 4380 4868 4436 4870
rect 4460 4868 4516 4870
rect 4066 4120 4122 4176
rect 4986 5630 4988 5672
rect 4988 5630 5040 5672
rect 5040 5630 5042 5672
rect 4986 5616 5042 5630
rect 4220 3834 4276 3836
rect 4300 3834 4356 3836
rect 4380 3834 4436 3836
rect 4460 3834 4516 3836
rect 4220 3782 4266 3834
rect 4266 3782 4276 3834
rect 4300 3782 4330 3834
rect 4330 3782 4342 3834
rect 4342 3782 4356 3834
rect 4380 3782 4394 3834
rect 4394 3782 4406 3834
rect 4406 3782 4436 3834
rect 4460 3782 4470 3834
rect 4470 3782 4516 3834
rect 4220 3780 4276 3782
rect 4300 3780 4356 3782
rect 4380 3780 4436 3782
rect 4460 3780 4516 3782
rect 4066 3168 4122 3224
rect 5906 11736 5962 11792
rect 6458 11192 6514 11248
rect 6458 10956 6460 10976
rect 6460 10956 6512 10976
rect 6512 10956 6514 10976
rect 6458 10920 6514 10956
rect 6366 10648 6422 10704
rect 7470 13504 7526 13560
rect 7194 13232 7250 13288
rect 6826 12144 6882 12200
rect 6734 11736 6790 11792
rect 6642 11328 6698 11384
rect 7562 12008 7618 12064
rect 7194 11600 7250 11656
rect 6918 11464 6974 11520
rect 5814 9560 5870 9616
rect 6274 10104 6330 10160
rect 6274 9152 6330 9208
rect 6458 10376 6514 10432
rect 6550 10104 6606 10160
rect 6458 9968 6514 10024
rect 6458 9832 6514 9888
rect 6734 9982 6736 10024
rect 6736 9982 6788 10024
rect 6788 9982 6790 10024
rect 6734 9968 6790 9982
rect 6734 9424 6790 9480
rect 7010 10648 7066 10704
rect 7010 9832 7066 9888
rect 7194 10512 7250 10568
rect 7470 11600 7526 11656
rect 7470 11464 7526 11520
rect 7378 10240 7434 10296
rect 7194 9716 7250 9752
rect 7194 9696 7196 9716
rect 7196 9696 7248 9716
rect 7248 9696 7250 9716
rect 7102 9324 7104 9344
rect 7104 9324 7156 9344
rect 7156 9324 7158 9344
rect 7102 9288 7158 9324
rect 6918 8880 6974 8936
rect 6550 8200 6606 8256
rect 5998 6160 6054 6216
rect 5262 5480 5318 5536
rect 3698 1808 3754 1864
rect 4220 2746 4276 2748
rect 4300 2746 4356 2748
rect 4380 2746 4436 2748
rect 4460 2746 4516 2748
rect 4220 2694 4266 2746
rect 4266 2694 4276 2746
rect 4300 2694 4330 2746
rect 4330 2694 4342 2746
rect 4342 2694 4356 2746
rect 4380 2694 4394 2746
rect 4394 2694 4406 2746
rect 4406 2694 4436 2746
rect 4460 2694 4470 2746
rect 4470 2694 4516 2746
rect 4220 2692 4276 2694
rect 4300 2692 4356 2694
rect 4380 2692 4436 2694
rect 4460 2692 4516 2694
rect 4066 2352 4122 2408
rect 4158 1944 4214 2000
rect 5078 2624 5134 2680
rect 6274 6296 6330 6352
rect 7194 8336 7250 8392
rect 7194 8064 7250 8120
rect 9770 13776 9826 13832
rect 8298 13368 8354 13424
rect 8850 13368 8906 13424
rect 8482 13268 8484 13288
rect 8484 13268 8536 13288
rect 8536 13268 8538 13288
rect 8482 13232 8538 13268
rect 8220 13082 8276 13084
rect 8300 13082 8356 13084
rect 8380 13082 8436 13084
rect 8460 13082 8516 13084
rect 8220 13030 8266 13082
rect 8266 13030 8276 13082
rect 8300 13030 8330 13082
rect 8330 13030 8342 13082
rect 8342 13030 8356 13082
rect 8380 13030 8394 13082
rect 8394 13030 8406 13082
rect 8406 13030 8436 13082
rect 8460 13030 8470 13082
rect 8470 13030 8516 13082
rect 8220 13028 8276 13030
rect 8300 13028 8356 13030
rect 8380 13028 8436 13030
rect 8460 13028 8516 13030
rect 7930 11872 7986 11928
rect 7930 11772 7932 11792
rect 7932 11772 7984 11792
rect 7984 11772 7986 11792
rect 7930 11736 7986 11772
rect 7746 10784 7802 10840
rect 7654 9424 7710 9480
rect 7930 10920 7986 10976
rect 7838 9444 7894 9480
rect 7838 9424 7840 9444
rect 7840 9424 7892 9444
rect 7892 9424 7894 9444
rect 7838 8916 7840 8936
rect 7840 8916 7892 8936
rect 7892 8916 7894 8936
rect 7838 8880 7894 8916
rect 7838 8628 7894 8664
rect 7838 8608 7840 8628
rect 7840 8608 7892 8628
rect 7892 8608 7894 8628
rect 4220 1658 4276 1660
rect 4300 1658 4356 1660
rect 4380 1658 4436 1660
rect 4460 1658 4516 1660
rect 4220 1606 4266 1658
rect 4266 1606 4276 1658
rect 4300 1606 4330 1658
rect 4330 1606 4342 1658
rect 4342 1606 4356 1658
rect 4380 1606 4394 1658
rect 4394 1606 4406 1658
rect 4406 1606 4436 1658
rect 4460 1606 4470 1658
rect 4470 1606 4516 1658
rect 4220 1604 4276 1606
rect 4300 1604 4356 1606
rect 4380 1604 4436 1606
rect 4460 1604 4516 1606
rect 3882 1264 3938 1320
rect 8220 11994 8276 11996
rect 8300 11994 8356 11996
rect 8380 11994 8436 11996
rect 8460 11994 8516 11996
rect 8220 11942 8266 11994
rect 8266 11942 8276 11994
rect 8300 11942 8330 11994
rect 8330 11942 8342 11994
rect 8342 11942 8356 11994
rect 8380 11942 8394 11994
rect 8394 11942 8406 11994
rect 8406 11942 8436 11994
rect 8460 11942 8470 11994
rect 8470 11942 8516 11994
rect 8220 11940 8276 11942
rect 8300 11940 8356 11942
rect 8380 11940 8436 11942
rect 8460 11940 8516 11942
rect 8666 12180 8668 12200
rect 8668 12180 8720 12200
rect 8720 12180 8722 12200
rect 8666 12144 8722 12180
rect 8666 12008 8722 12064
rect 8482 11464 8538 11520
rect 8390 11328 8446 11384
rect 8114 11092 8116 11112
rect 8116 11092 8168 11112
rect 8168 11092 8170 11112
rect 8114 11056 8170 11092
rect 8666 11464 8722 11520
rect 8220 10906 8276 10908
rect 8300 10906 8356 10908
rect 8380 10906 8436 10908
rect 8460 10906 8516 10908
rect 8220 10854 8266 10906
rect 8266 10854 8276 10906
rect 8300 10854 8330 10906
rect 8330 10854 8342 10906
rect 8342 10854 8356 10906
rect 8380 10854 8394 10906
rect 8394 10854 8406 10906
rect 8406 10854 8436 10906
rect 8460 10854 8470 10906
rect 8470 10854 8516 10906
rect 8220 10852 8276 10854
rect 8300 10852 8356 10854
rect 8380 10852 8436 10854
rect 8460 10852 8516 10854
rect 8298 10668 8354 10704
rect 8298 10648 8300 10668
rect 8300 10648 8352 10668
rect 8352 10648 8354 10668
rect 8390 10548 8392 10568
rect 8392 10548 8444 10568
rect 8444 10548 8446 10568
rect 8390 10512 8446 10548
rect 8574 10260 8630 10296
rect 8942 12008 8998 12064
rect 8942 11872 8998 11928
rect 9310 11872 9366 11928
rect 9218 11736 9274 11792
rect 9310 11464 9366 11520
rect 9126 11328 9182 11384
rect 10230 12008 10286 12064
rect 9402 11328 9458 11384
rect 8942 10920 8998 10976
rect 9678 10920 9734 10976
rect 8574 10240 8576 10260
rect 8576 10240 8628 10260
rect 8628 10240 8630 10260
rect 9126 10532 9182 10568
rect 9126 10512 9128 10532
rect 9128 10512 9180 10532
rect 9180 10512 9182 10532
rect 9310 10784 9366 10840
rect 8220 9818 8276 9820
rect 8300 9818 8356 9820
rect 8380 9818 8436 9820
rect 8460 9818 8516 9820
rect 8220 9766 8266 9818
rect 8266 9766 8276 9818
rect 8300 9766 8330 9818
rect 8330 9766 8342 9818
rect 8342 9766 8356 9818
rect 8380 9766 8394 9818
rect 8394 9766 8406 9818
rect 8406 9766 8436 9818
rect 8460 9766 8470 9818
rect 8470 9766 8516 9818
rect 8220 9764 8276 9766
rect 8300 9764 8356 9766
rect 8380 9764 8436 9766
rect 8460 9764 8516 9766
rect 8298 8880 8354 8936
rect 8220 8730 8276 8732
rect 8300 8730 8356 8732
rect 8380 8730 8436 8732
rect 8460 8730 8516 8732
rect 8220 8678 8266 8730
rect 8266 8678 8276 8730
rect 8300 8678 8330 8730
rect 8330 8678 8342 8730
rect 8342 8678 8356 8730
rect 8380 8678 8394 8730
rect 8394 8678 8406 8730
rect 8406 8678 8436 8730
rect 8460 8678 8470 8730
rect 8470 8678 8516 8730
rect 8220 8676 8276 8678
rect 8300 8676 8356 8678
rect 8380 8676 8436 8678
rect 8460 8676 8516 8678
rect 8206 8472 8262 8528
rect 8758 9152 8814 9208
rect 8758 9016 8814 9072
rect 9034 9968 9090 10024
rect 8220 7642 8276 7644
rect 8300 7642 8356 7644
rect 8380 7642 8436 7644
rect 8460 7642 8516 7644
rect 8220 7590 8266 7642
rect 8266 7590 8276 7642
rect 8300 7590 8330 7642
rect 8330 7590 8342 7642
rect 8342 7590 8356 7642
rect 8380 7590 8394 7642
rect 8394 7590 8406 7642
rect 8406 7590 8436 7642
rect 8460 7590 8470 7642
rect 8470 7590 8516 7642
rect 8220 7588 8276 7590
rect 8300 7588 8356 7590
rect 8380 7588 8436 7590
rect 8460 7588 8516 7590
rect 8390 7420 8392 7440
rect 8392 7420 8444 7440
rect 8444 7420 8446 7440
rect 8390 7384 8446 7420
rect 8220 6554 8276 6556
rect 8300 6554 8356 6556
rect 8380 6554 8436 6556
rect 8460 6554 8516 6556
rect 8220 6502 8266 6554
rect 8266 6502 8276 6554
rect 8300 6502 8330 6554
rect 8330 6502 8342 6554
rect 8342 6502 8356 6554
rect 8380 6502 8394 6554
rect 8394 6502 8406 6554
rect 8406 6502 8436 6554
rect 8460 6502 8470 6554
rect 8470 6502 8516 6554
rect 8220 6500 8276 6502
rect 8300 6500 8356 6502
rect 8380 6500 8436 6502
rect 8460 6500 8516 6502
rect 8850 7656 8906 7712
rect 9402 10648 9458 10704
rect 9494 10512 9550 10568
rect 9954 11056 10010 11112
rect 9586 10376 9642 10432
rect 9494 9016 9550 9072
rect 10690 11872 10746 11928
rect 10690 11736 10746 11792
rect 10782 11600 10838 11656
rect 10230 11192 10286 11248
rect 10230 10512 10286 10568
rect 10506 10668 10562 10704
rect 10506 10648 10508 10668
rect 10508 10648 10560 10668
rect 10560 10648 10562 10668
rect 10598 10512 10654 10568
rect 10046 10104 10102 10160
rect 9862 9288 9918 9344
rect 7102 2524 7104 2544
rect 7104 2524 7156 2544
rect 7156 2524 7158 2544
rect 7102 2488 7158 2524
rect 8220 5466 8276 5468
rect 8300 5466 8356 5468
rect 8380 5466 8436 5468
rect 8460 5466 8516 5468
rect 8220 5414 8266 5466
rect 8266 5414 8276 5466
rect 8300 5414 8330 5466
rect 8330 5414 8342 5466
rect 8342 5414 8356 5466
rect 8380 5414 8394 5466
rect 8394 5414 8406 5466
rect 8406 5414 8436 5466
rect 8460 5414 8470 5466
rect 8470 5414 8516 5466
rect 8220 5412 8276 5414
rect 8300 5412 8356 5414
rect 8380 5412 8436 5414
rect 8460 5412 8516 5414
rect 8220 4378 8276 4380
rect 8300 4378 8356 4380
rect 8380 4378 8436 4380
rect 8460 4378 8516 4380
rect 8220 4326 8266 4378
rect 8266 4326 8276 4378
rect 8300 4326 8330 4378
rect 8330 4326 8342 4378
rect 8342 4326 8356 4378
rect 8380 4326 8394 4378
rect 8394 4326 8406 4378
rect 8406 4326 8436 4378
rect 8460 4326 8470 4378
rect 8470 4326 8516 4378
rect 8220 4324 8276 4326
rect 8300 4324 8356 4326
rect 8380 4324 8436 4326
rect 8460 4324 8516 4326
rect 8220 3290 8276 3292
rect 8300 3290 8356 3292
rect 8380 3290 8436 3292
rect 8460 3290 8516 3292
rect 8220 3238 8266 3290
rect 8266 3238 8276 3290
rect 8300 3238 8330 3290
rect 8330 3238 8342 3290
rect 8342 3238 8356 3290
rect 8380 3238 8394 3290
rect 8394 3238 8406 3290
rect 8406 3238 8436 3290
rect 8460 3238 8470 3290
rect 8470 3238 8516 3290
rect 8220 3236 8276 3238
rect 8300 3236 8356 3238
rect 8380 3236 8436 3238
rect 8460 3236 8516 3238
rect 8482 2508 8538 2544
rect 8482 2488 8484 2508
rect 8484 2488 8536 2508
rect 8536 2488 8538 2508
rect 9770 8064 9826 8120
rect 9770 7792 9826 7848
rect 10046 10004 10048 10024
rect 10048 10004 10100 10024
rect 10100 10004 10102 10024
rect 10046 9968 10102 10004
rect 10138 9696 10194 9752
rect 10046 8336 10102 8392
rect 10782 9696 10838 9752
rect 10690 9324 10692 9344
rect 10692 9324 10744 9344
rect 10744 9324 10746 9344
rect 10690 9288 10746 9324
rect 11150 10920 11206 10976
rect 11058 10376 11114 10432
rect 10966 10004 10968 10024
rect 10968 10004 11020 10024
rect 11020 10004 11022 10024
rect 10966 9968 11022 10004
rect 11058 9560 11114 9616
rect 10230 8200 10286 8256
rect 10230 7928 10286 7984
rect 10414 7964 10416 7984
rect 10416 7964 10468 7984
rect 10468 7964 10470 7984
rect 10414 7928 10470 7964
rect 10046 6976 10102 7032
rect 10690 8064 10746 8120
rect 10598 7928 10654 7984
rect 10782 7928 10838 7984
rect 10782 7792 10838 7848
rect 10690 7656 10746 7712
rect 11150 9424 11206 9480
rect 11058 7828 11060 7848
rect 11060 7828 11112 7848
rect 11112 7828 11114 7848
rect 11058 7792 11114 7828
rect 11702 11192 11758 11248
rect 11426 9288 11482 9344
rect 10966 6160 11022 6216
rect 12220 13626 12276 13628
rect 12300 13626 12356 13628
rect 12380 13626 12436 13628
rect 12460 13626 12516 13628
rect 12220 13574 12266 13626
rect 12266 13574 12276 13626
rect 12300 13574 12330 13626
rect 12330 13574 12342 13626
rect 12342 13574 12356 13626
rect 12380 13574 12394 13626
rect 12394 13574 12406 13626
rect 12406 13574 12436 13626
rect 12460 13574 12470 13626
rect 12470 13574 12516 13626
rect 12220 13572 12276 13574
rect 12300 13572 12356 13574
rect 12380 13572 12436 13574
rect 12460 13572 12516 13574
rect 12220 12538 12276 12540
rect 12300 12538 12356 12540
rect 12380 12538 12436 12540
rect 12460 12538 12516 12540
rect 12220 12486 12266 12538
rect 12266 12486 12276 12538
rect 12300 12486 12330 12538
rect 12330 12486 12342 12538
rect 12342 12486 12356 12538
rect 12380 12486 12394 12538
rect 12394 12486 12406 12538
rect 12406 12486 12436 12538
rect 12460 12486 12470 12538
rect 12470 12486 12516 12538
rect 12220 12484 12276 12486
rect 12300 12484 12356 12486
rect 12380 12484 12436 12486
rect 12460 12484 12516 12486
rect 12220 11450 12276 11452
rect 12300 11450 12356 11452
rect 12380 11450 12436 11452
rect 12460 11450 12516 11452
rect 12220 11398 12266 11450
rect 12266 11398 12276 11450
rect 12300 11398 12330 11450
rect 12330 11398 12342 11450
rect 12342 11398 12356 11450
rect 12380 11398 12394 11450
rect 12394 11398 12406 11450
rect 12406 11398 12436 11450
rect 12460 11398 12470 11450
rect 12470 11398 12516 11450
rect 12220 11396 12276 11398
rect 12300 11396 12356 11398
rect 12380 11396 12436 11398
rect 12460 11396 12516 11398
rect 11702 9696 11758 9752
rect 11610 8492 11666 8528
rect 11610 8472 11612 8492
rect 11612 8472 11664 8492
rect 11664 8472 11666 8492
rect 11426 6976 11482 7032
rect 8220 2202 8276 2204
rect 8300 2202 8356 2204
rect 8380 2202 8436 2204
rect 8460 2202 8516 2204
rect 8220 2150 8266 2202
rect 8266 2150 8276 2202
rect 8300 2150 8330 2202
rect 8330 2150 8342 2202
rect 8342 2150 8356 2202
rect 8380 2150 8394 2202
rect 8394 2150 8406 2202
rect 8406 2150 8436 2202
rect 8460 2150 8470 2202
rect 8470 2150 8516 2202
rect 8220 2148 8276 2150
rect 8300 2148 8356 2150
rect 8380 2148 8436 2150
rect 8460 2148 8516 2150
rect 12254 10920 12310 10976
rect 12162 10684 12164 10704
rect 12164 10684 12216 10704
rect 12216 10684 12218 10704
rect 12162 10648 12218 10684
rect 12220 10362 12276 10364
rect 12300 10362 12356 10364
rect 12380 10362 12436 10364
rect 12460 10362 12516 10364
rect 12220 10310 12266 10362
rect 12266 10310 12276 10362
rect 12300 10310 12330 10362
rect 12330 10310 12342 10362
rect 12342 10310 12356 10362
rect 12380 10310 12394 10362
rect 12394 10310 12406 10362
rect 12406 10310 12436 10362
rect 12460 10310 12470 10362
rect 12470 10310 12516 10362
rect 12220 10308 12276 10310
rect 12300 10308 12356 10310
rect 12380 10308 12436 10310
rect 12460 10308 12516 10310
rect 12898 10512 12954 10568
rect 12990 9560 13046 9616
rect 12220 9274 12276 9276
rect 12300 9274 12356 9276
rect 12380 9274 12436 9276
rect 12460 9274 12516 9276
rect 12220 9222 12266 9274
rect 12266 9222 12276 9274
rect 12300 9222 12330 9274
rect 12330 9222 12342 9274
rect 12342 9222 12356 9274
rect 12380 9222 12394 9274
rect 12394 9222 12406 9274
rect 12406 9222 12436 9274
rect 12460 9222 12470 9274
rect 12470 9222 12516 9274
rect 12220 9220 12276 9222
rect 12300 9220 12356 9222
rect 12380 9220 12436 9222
rect 12460 9220 12516 9222
rect 12070 9152 12126 9208
rect 12622 8236 12624 8256
rect 12624 8236 12676 8256
rect 12676 8236 12678 8256
rect 12622 8200 12678 8236
rect 12220 8186 12276 8188
rect 12300 8186 12356 8188
rect 12380 8186 12436 8188
rect 12460 8186 12516 8188
rect 12220 8134 12266 8186
rect 12266 8134 12276 8186
rect 12300 8134 12330 8186
rect 12330 8134 12342 8186
rect 12342 8134 12356 8186
rect 12380 8134 12394 8186
rect 12394 8134 12406 8186
rect 12406 8134 12436 8186
rect 12460 8134 12470 8186
rect 12470 8134 12516 8186
rect 12220 8132 12276 8134
rect 12300 8132 12356 8134
rect 12380 8132 12436 8134
rect 12460 8132 12516 8134
rect 12220 7098 12276 7100
rect 12300 7098 12356 7100
rect 12380 7098 12436 7100
rect 12460 7098 12516 7100
rect 12220 7046 12266 7098
rect 12266 7046 12276 7098
rect 12300 7046 12330 7098
rect 12330 7046 12342 7098
rect 12342 7046 12356 7098
rect 12380 7046 12394 7098
rect 12394 7046 12406 7098
rect 12406 7046 12436 7098
rect 12460 7046 12470 7098
rect 12470 7046 12516 7098
rect 12220 7044 12276 7046
rect 12300 7044 12356 7046
rect 12380 7044 12436 7046
rect 12460 7044 12516 7046
rect 12220 6010 12276 6012
rect 12300 6010 12356 6012
rect 12380 6010 12436 6012
rect 12460 6010 12516 6012
rect 12220 5958 12266 6010
rect 12266 5958 12276 6010
rect 12300 5958 12330 6010
rect 12330 5958 12342 6010
rect 12342 5958 12356 6010
rect 12380 5958 12394 6010
rect 12394 5958 12406 6010
rect 12406 5958 12436 6010
rect 12460 5958 12470 6010
rect 12470 5958 12516 6010
rect 12220 5956 12276 5958
rect 12300 5956 12356 5958
rect 12380 5956 12436 5958
rect 12460 5956 12516 5958
rect 12220 4922 12276 4924
rect 12300 4922 12356 4924
rect 12380 4922 12436 4924
rect 12460 4922 12516 4924
rect 12220 4870 12266 4922
rect 12266 4870 12276 4922
rect 12300 4870 12330 4922
rect 12330 4870 12342 4922
rect 12342 4870 12356 4922
rect 12380 4870 12394 4922
rect 12394 4870 12406 4922
rect 12406 4870 12436 4922
rect 12460 4870 12470 4922
rect 12470 4870 12516 4922
rect 12220 4868 12276 4870
rect 12300 4868 12356 4870
rect 12380 4868 12436 4870
rect 12460 4868 12516 4870
rect 9126 2216 9182 2272
rect 9310 1828 9366 1864
rect 9310 1808 9312 1828
rect 9312 1808 9364 1828
rect 9364 1808 9366 1828
rect 12220 3834 12276 3836
rect 12300 3834 12356 3836
rect 12380 3834 12436 3836
rect 12460 3834 12516 3836
rect 12220 3782 12266 3834
rect 12266 3782 12276 3834
rect 12300 3782 12330 3834
rect 12330 3782 12342 3834
rect 12342 3782 12356 3834
rect 12380 3782 12394 3834
rect 12394 3782 12406 3834
rect 12406 3782 12436 3834
rect 12460 3782 12470 3834
rect 12470 3782 12516 3834
rect 12220 3780 12276 3782
rect 12300 3780 12356 3782
rect 12380 3780 12436 3782
rect 12460 3780 12516 3782
rect 11242 2624 11298 2680
rect 11058 2488 11114 2544
rect 8220 1114 8276 1116
rect 8300 1114 8356 1116
rect 8380 1114 8436 1116
rect 8460 1114 8516 1116
rect 8220 1062 8266 1114
rect 8266 1062 8276 1114
rect 8300 1062 8330 1114
rect 8330 1062 8342 1114
rect 8342 1062 8356 1114
rect 8380 1062 8394 1114
rect 8394 1062 8406 1114
rect 8406 1062 8436 1114
rect 8460 1062 8470 1114
rect 8470 1062 8516 1114
rect 8220 1060 8276 1062
rect 8300 1060 8356 1062
rect 8380 1060 8436 1062
rect 8460 1060 8516 1062
rect 11518 2216 11574 2272
rect 12220 2746 12276 2748
rect 12300 2746 12356 2748
rect 12380 2746 12436 2748
rect 12460 2746 12516 2748
rect 12220 2694 12266 2746
rect 12266 2694 12276 2746
rect 12300 2694 12330 2746
rect 12330 2694 12342 2746
rect 12342 2694 12356 2746
rect 12380 2694 12394 2746
rect 12394 2694 12406 2746
rect 12406 2694 12436 2746
rect 12460 2694 12470 2746
rect 12470 2694 12516 2746
rect 12220 2692 12276 2694
rect 12300 2692 12356 2694
rect 12380 2692 12436 2694
rect 12460 2692 12516 2694
rect 13634 8744 13690 8800
rect 12898 8200 12954 8256
rect 12806 6296 12862 6352
rect 12714 3712 12770 3768
rect 13174 7420 13176 7440
rect 13176 7420 13228 7440
rect 13228 7420 13230 7440
rect 13174 7384 13230 7420
rect 12220 1658 12276 1660
rect 12300 1658 12356 1660
rect 12380 1658 12436 1660
rect 12460 1658 12516 1660
rect 12220 1606 12266 1658
rect 12266 1606 12276 1658
rect 12300 1606 12330 1658
rect 12330 1606 12342 1658
rect 12342 1606 12356 1658
rect 12380 1606 12394 1658
rect 12394 1606 12406 1658
rect 12406 1606 12436 1658
rect 12460 1606 12470 1658
rect 12470 1606 12516 1658
rect 12220 1604 12276 1606
rect 12300 1604 12356 1606
rect 12380 1604 12436 1606
rect 12460 1604 12516 1606
rect 13542 1264 13598 1320
rect 1398 448 1454 504
<< metal3 >>
rect 0 14514 800 14544
rect 3233 14514 3299 14517
rect 0 14512 3299 14514
rect 0 14456 3238 14512
rect 3294 14456 3299 14512
rect 0 14454 3299 14456
rect 0 14424 800 14454
rect 3233 14451 3299 14454
rect 9765 13834 9831 13837
rect 9765 13832 12818 13834
rect 9765 13776 9770 13832
rect 9826 13776 12818 13832
rect 9765 13774 12818 13776
rect 9765 13771 9831 13774
rect 12758 13698 12818 13774
rect 14200 13698 15000 13728
rect 12758 13638 15000 13698
rect 4210 13632 4526 13633
rect 0 13562 800 13592
rect 4210 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4526 13632
rect 4210 13567 4526 13568
rect 12210 13632 12526 13633
rect 12210 13568 12216 13632
rect 12280 13568 12296 13632
rect 12360 13568 12376 13632
rect 12440 13568 12456 13632
rect 12520 13568 12526 13632
rect 14200 13608 15000 13638
rect 12210 13567 12526 13568
rect 1945 13562 2011 13565
rect 0 13560 2011 13562
rect 0 13504 1950 13560
rect 2006 13504 2011 13560
rect 0 13502 2011 13504
rect 0 13472 800 13502
rect 1945 13499 2011 13502
rect 6310 13500 6316 13564
rect 6380 13562 6386 13564
rect 7465 13562 7531 13565
rect 6380 13560 7531 13562
rect 6380 13504 7470 13560
rect 7526 13504 7531 13560
rect 6380 13502 7531 13504
rect 6380 13500 6386 13502
rect 7465 13499 7531 13502
rect 1669 13426 1735 13429
rect 8293 13426 8359 13429
rect 8845 13426 8911 13429
rect 1669 13424 8911 13426
rect 1669 13368 1674 13424
rect 1730 13368 8298 13424
rect 8354 13368 8850 13424
rect 8906 13368 8911 13424
rect 1669 13366 8911 13368
rect 1669 13363 1735 13366
rect 8293 13363 8359 13366
rect 8845 13363 8911 13366
rect 2865 13290 2931 13293
rect 7189 13290 7255 13293
rect 2865 13288 7255 13290
rect 2865 13232 2870 13288
rect 2926 13232 7194 13288
rect 7250 13232 7255 13288
rect 2865 13230 7255 13232
rect 2865 13227 2931 13230
rect 7189 13227 7255 13230
rect 8477 13290 8543 13293
rect 9438 13290 9444 13292
rect 8477 13288 9444 13290
rect 8477 13232 8482 13288
rect 8538 13232 9444 13288
rect 8477 13230 9444 13232
rect 8477 13227 8543 13230
rect 9438 13228 9444 13230
rect 9508 13228 9514 13292
rect 8210 13088 8526 13089
rect 8210 13024 8216 13088
rect 8280 13024 8296 13088
rect 8360 13024 8376 13088
rect 8440 13024 8456 13088
rect 8520 13024 8526 13088
rect 8210 13023 8526 13024
rect 1945 12882 2011 12885
rect 8702 12882 8708 12884
rect 1945 12880 8708 12882
rect 1945 12824 1950 12880
rect 2006 12824 8708 12880
rect 1945 12822 8708 12824
rect 1945 12819 2011 12822
rect 8702 12820 8708 12822
rect 8772 12820 8778 12884
rect 0 12610 800 12640
rect 1393 12610 1459 12613
rect 0 12608 1459 12610
rect 0 12552 1398 12608
rect 1454 12552 1459 12608
rect 0 12550 1459 12552
rect 0 12520 800 12550
rect 1393 12547 1459 12550
rect 4210 12544 4526 12545
rect 4210 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4526 12544
rect 4210 12479 4526 12480
rect 12210 12544 12526 12545
rect 12210 12480 12216 12544
rect 12280 12480 12296 12544
rect 12360 12480 12376 12544
rect 12440 12480 12456 12544
rect 12520 12480 12526 12544
rect 12210 12479 12526 12480
rect 6821 12202 6887 12205
rect 8661 12202 8727 12205
rect 6821 12200 8727 12202
rect 6821 12144 6826 12200
rect 6882 12144 8666 12200
rect 8722 12144 8727 12200
rect 6821 12142 8727 12144
rect 6821 12139 6887 12142
rect 8661 12139 8727 12142
rect 8664 12069 8724 12139
rect 3969 12066 4035 12069
rect 7557 12066 7623 12069
rect 3969 12064 7623 12066
rect 3969 12008 3974 12064
rect 4030 12008 7562 12064
rect 7618 12008 7623 12064
rect 3969 12006 7623 12008
rect 3969 12003 4035 12006
rect 7557 12003 7623 12006
rect 8661 12064 8727 12069
rect 8661 12008 8666 12064
rect 8722 12008 8727 12064
rect 8661 12003 8727 12008
rect 8937 12066 9003 12069
rect 10225 12066 10291 12069
rect 8937 12064 10291 12066
rect 8937 12008 8942 12064
rect 8998 12008 10230 12064
rect 10286 12008 10291 12064
rect 8937 12006 10291 12008
rect 8937 12003 9003 12006
rect 10225 12003 10291 12006
rect 8210 12000 8526 12001
rect 8210 11936 8216 12000
rect 8280 11936 8296 12000
rect 8360 11936 8376 12000
rect 8440 11936 8456 12000
rect 8520 11936 8526 12000
rect 8210 11935 8526 11936
rect 7925 11930 7991 11933
rect 7790 11928 7991 11930
rect 7790 11872 7930 11928
rect 7986 11872 7991 11928
rect 7790 11870 7991 11872
rect 2405 11794 2471 11797
rect 5901 11794 5967 11797
rect 6729 11794 6795 11797
rect 2405 11792 6795 11794
rect 2405 11736 2410 11792
rect 2466 11736 5906 11792
rect 5962 11736 6734 11792
rect 6790 11736 6795 11792
rect 2405 11734 6795 11736
rect 2405 11731 2471 11734
rect 5901 11731 5967 11734
rect 6729 11731 6795 11734
rect 0 11658 800 11688
rect 3049 11658 3115 11661
rect 0 11656 3115 11658
rect 0 11600 3054 11656
rect 3110 11600 3115 11656
rect 0 11598 3115 11600
rect 0 11568 800 11598
rect 3049 11595 3115 11598
rect 4521 11658 4587 11661
rect 7189 11658 7255 11661
rect 7465 11658 7531 11661
rect 4521 11656 4722 11658
rect 4521 11600 4526 11656
rect 4582 11600 4722 11656
rect 4521 11598 4722 11600
rect 4521 11595 4587 11598
rect 4210 11456 4526 11457
rect 4210 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4526 11456
rect 4210 11391 4526 11392
rect 4662 11250 4722 11598
rect 7189 11656 7531 11658
rect 7189 11600 7194 11656
rect 7250 11600 7470 11656
rect 7526 11600 7531 11656
rect 7189 11598 7531 11600
rect 7189 11595 7255 11598
rect 7465 11595 7531 11598
rect 6913 11522 6979 11525
rect 7465 11522 7531 11525
rect 6913 11520 7531 11522
rect 6913 11464 6918 11520
rect 6974 11464 7470 11520
rect 7526 11464 7531 11520
rect 6913 11462 7531 11464
rect 7790 11522 7850 11870
rect 7925 11867 7991 11870
rect 8937 11930 9003 11933
rect 9305 11930 9371 11933
rect 8937 11928 9371 11930
rect 8937 11872 8942 11928
rect 8998 11872 9310 11928
rect 9366 11872 9371 11928
rect 8937 11870 9371 11872
rect 8937 11867 9003 11870
rect 9305 11867 9371 11870
rect 10174 11868 10180 11932
rect 10244 11930 10250 11932
rect 10685 11930 10751 11933
rect 10244 11928 10751 11930
rect 10244 11872 10690 11928
rect 10746 11872 10751 11928
rect 10244 11870 10751 11872
rect 10244 11868 10250 11870
rect 10685 11867 10751 11870
rect 7925 11794 7991 11797
rect 9213 11794 9279 11797
rect 10685 11794 10751 11797
rect 7925 11792 8540 11794
rect 7925 11736 7930 11792
rect 7986 11736 8540 11792
rect 7925 11734 8540 11736
rect 7925 11731 7991 11734
rect 8480 11658 8540 11734
rect 9213 11792 10751 11794
rect 9213 11736 9218 11792
rect 9274 11736 10690 11792
rect 10746 11736 10751 11792
rect 9213 11734 10751 11736
rect 9213 11731 9279 11734
rect 10685 11731 10751 11734
rect 10777 11658 10843 11661
rect 8480 11656 10843 11658
rect 8480 11600 10782 11656
rect 10838 11600 10843 11656
rect 8480 11598 10843 11600
rect 10777 11595 10843 11598
rect 8477 11522 8543 11525
rect 7790 11520 8543 11522
rect 7790 11464 8482 11520
rect 8538 11464 8543 11520
rect 7790 11462 8543 11464
rect 6913 11459 6979 11462
rect 7465 11459 7531 11462
rect 8477 11459 8543 11462
rect 8661 11522 8727 11525
rect 9305 11522 9371 11525
rect 8661 11520 9371 11522
rect 8661 11464 8666 11520
rect 8722 11464 9310 11520
rect 9366 11464 9371 11520
rect 8661 11462 9371 11464
rect 8661 11459 8727 11462
rect 9305 11459 9371 11462
rect 12210 11456 12526 11457
rect 12210 11392 12216 11456
rect 12280 11392 12296 11456
rect 12360 11392 12376 11456
rect 12440 11392 12456 11456
rect 12520 11392 12526 11456
rect 12210 11391 12526 11392
rect 6637 11386 6703 11389
rect 8385 11386 8451 11389
rect 9121 11388 9187 11389
rect 9070 11386 9076 11388
rect 6637 11384 8451 11386
rect 6637 11328 6642 11384
rect 6698 11328 8390 11384
rect 8446 11328 8451 11384
rect 6637 11326 8451 11328
rect 9030 11326 9076 11386
rect 9140 11384 9187 11388
rect 9182 11328 9187 11384
rect 6637 11323 6703 11326
rect 8385 11323 8451 11326
rect 9070 11324 9076 11326
rect 9140 11324 9187 11328
rect 9254 11324 9260 11388
rect 9324 11386 9330 11388
rect 9397 11386 9463 11389
rect 9324 11384 9463 11386
rect 9324 11328 9402 11384
rect 9458 11328 9463 11384
rect 9324 11326 9463 11328
rect 9324 11324 9330 11326
rect 9121 11323 9187 11324
rect 9397 11323 9463 11326
rect 4797 11250 4863 11253
rect 4662 11248 4863 11250
rect 4662 11192 4802 11248
rect 4858 11192 4863 11248
rect 4662 11190 4863 11192
rect 4797 11187 4863 11190
rect 6453 11250 6519 11253
rect 7966 11250 7972 11252
rect 6453 11248 7972 11250
rect 6453 11192 6458 11248
rect 6514 11192 7972 11248
rect 6453 11190 7972 11192
rect 6453 11187 6519 11190
rect 7966 11188 7972 11190
rect 8036 11250 8042 11252
rect 9990 11250 9996 11252
rect 8036 11190 9996 11250
rect 8036 11188 8042 11190
rect 9990 11188 9996 11190
rect 10060 11250 10066 11252
rect 10225 11250 10291 11253
rect 10060 11248 10291 11250
rect 10060 11192 10230 11248
rect 10286 11192 10291 11248
rect 10060 11190 10291 11192
rect 10060 11188 10066 11190
rect 10225 11187 10291 11190
rect 11697 11250 11763 11253
rect 14200 11250 15000 11280
rect 11697 11248 15000 11250
rect 11697 11192 11702 11248
rect 11758 11192 15000 11248
rect 11697 11190 15000 11192
rect 11697 11187 11763 11190
rect 14200 11160 15000 11190
rect 8109 11114 8175 11117
rect 9949 11114 10015 11117
rect 8109 11112 10015 11114
rect 8109 11056 8114 11112
rect 8170 11056 9954 11112
rect 10010 11056 10015 11112
rect 8109 11054 10015 11056
rect 8109 11051 8175 11054
rect 9949 11051 10015 11054
rect 6453 10978 6519 10981
rect 7925 10978 7991 10981
rect 6453 10976 7991 10978
rect 6453 10920 6458 10976
rect 6514 10920 7930 10976
rect 7986 10920 7991 10976
rect 6453 10918 7991 10920
rect 6453 10915 6519 10918
rect 7925 10915 7991 10918
rect 8937 10978 9003 10981
rect 9673 10978 9739 10981
rect 8937 10976 9739 10978
rect 8937 10920 8942 10976
rect 8998 10920 9678 10976
rect 9734 10920 9739 10976
rect 8937 10918 9739 10920
rect 8937 10915 9003 10918
rect 9673 10915 9739 10918
rect 11145 10978 11211 10981
rect 12249 10978 12315 10981
rect 11145 10976 12315 10978
rect 11145 10920 11150 10976
rect 11206 10920 12254 10976
rect 12310 10920 12315 10976
rect 11145 10918 12315 10920
rect 11145 10915 11211 10918
rect 12249 10915 12315 10918
rect 8210 10912 8526 10913
rect 8210 10848 8216 10912
rect 8280 10848 8296 10912
rect 8360 10848 8376 10912
rect 8440 10848 8456 10912
rect 8520 10848 8526 10912
rect 8210 10847 8526 10848
rect 3141 10842 3207 10845
rect 7741 10842 7807 10845
rect 3141 10840 7807 10842
rect 3141 10784 3146 10840
rect 3202 10784 7746 10840
rect 7802 10784 7807 10840
rect 3141 10782 7807 10784
rect 3141 10779 3207 10782
rect 7741 10779 7807 10782
rect 8702 10780 8708 10844
rect 8772 10842 8778 10844
rect 9305 10842 9371 10845
rect 8772 10840 9371 10842
rect 8772 10784 9310 10840
rect 9366 10784 9371 10840
rect 8772 10782 9371 10784
rect 8772 10780 8778 10782
rect 9305 10779 9371 10782
rect 0 10706 800 10736
rect 6361 10706 6427 10709
rect 0 10704 6427 10706
rect 0 10648 6366 10704
rect 6422 10648 6427 10704
rect 0 10646 6427 10648
rect 0 10616 800 10646
rect 6361 10643 6427 10646
rect 7005 10706 7071 10709
rect 8293 10706 8359 10709
rect 7005 10704 8359 10706
rect 7005 10648 7010 10704
rect 7066 10648 8298 10704
rect 8354 10648 8359 10704
rect 7005 10646 8359 10648
rect 7005 10643 7071 10646
rect 8293 10643 8359 10646
rect 9254 10644 9260 10708
rect 9324 10706 9330 10708
rect 9397 10706 9463 10709
rect 9324 10704 9463 10706
rect 9324 10648 9402 10704
rect 9458 10648 9463 10704
rect 9324 10646 9463 10648
rect 9324 10644 9330 10646
rect 9397 10643 9463 10646
rect 10501 10706 10567 10709
rect 12157 10706 12223 10709
rect 10501 10704 12223 10706
rect 10501 10648 10506 10704
rect 10562 10648 12162 10704
rect 12218 10648 12223 10704
rect 10501 10646 12223 10648
rect 10501 10643 10567 10646
rect 12157 10643 12223 10646
rect 7189 10570 7255 10573
rect 8385 10570 8451 10573
rect 9121 10570 9187 10573
rect 9489 10572 9555 10573
rect 7189 10568 9187 10570
rect 7189 10512 7194 10568
rect 7250 10512 8390 10568
rect 8446 10512 9126 10568
rect 9182 10512 9187 10568
rect 7189 10510 9187 10512
rect 7189 10507 7255 10510
rect 8385 10507 8451 10510
rect 9121 10507 9187 10510
rect 9438 10508 9444 10572
rect 9508 10570 9555 10572
rect 10225 10570 10291 10573
rect 10593 10570 10659 10573
rect 12893 10570 12959 10573
rect 9508 10568 9600 10570
rect 9550 10512 9600 10568
rect 9508 10510 9600 10512
rect 10225 10568 10659 10570
rect 10225 10512 10230 10568
rect 10286 10512 10598 10568
rect 10654 10512 10659 10568
rect 10225 10510 10659 10512
rect 9508 10508 9555 10510
rect 9489 10507 9555 10508
rect 10225 10507 10291 10510
rect 10593 10507 10659 10510
rect 11056 10568 12959 10570
rect 11056 10512 12898 10568
rect 12954 10512 12959 10568
rect 11056 10510 12959 10512
rect 11056 10437 11116 10510
rect 12893 10507 12959 10510
rect 6453 10434 6519 10437
rect 9581 10434 9647 10437
rect 11053 10434 11119 10437
rect 6453 10432 11119 10434
rect 6453 10376 6458 10432
rect 6514 10376 9586 10432
rect 9642 10376 11058 10432
rect 11114 10376 11119 10432
rect 6453 10374 11119 10376
rect 6453 10371 6519 10374
rect 9581 10371 9647 10374
rect 11053 10371 11119 10374
rect 4210 10368 4526 10369
rect 4210 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4526 10368
rect 4210 10303 4526 10304
rect 12210 10368 12526 10369
rect 12210 10304 12216 10368
rect 12280 10304 12296 10368
rect 12360 10304 12376 10368
rect 12440 10304 12456 10368
rect 12520 10304 12526 10368
rect 12210 10303 12526 10304
rect 7373 10298 7439 10301
rect 8569 10298 8635 10301
rect 10174 10298 10180 10300
rect 7373 10296 10180 10298
rect 7373 10240 7378 10296
rect 7434 10240 8574 10296
rect 8630 10240 10180 10296
rect 7373 10238 10180 10240
rect 7373 10235 7439 10238
rect 8569 10235 8635 10238
rect 10174 10236 10180 10238
rect 10244 10236 10250 10300
rect 6269 10164 6335 10165
rect 6269 10162 6316 10164
rect 6224 10160 6316 10162
rect 6224 10104 6274 10160
rect 6224 10102 6316 10104
rect 6269 10100 6316 10102
rect 6380 10100 6386 10164
rect 6545 10162 6611 10165
rect 10041 10162 10107 10165
rect 6545 10160 10107 10162
rect 6545 10104 6550 10160
rect 6606 10104 10046 10160
rect 10102 10104 10107 10160
rect 6545 10102 10107 10104
rect 6269 10099 6335 10100
rect 6545 10099 6611 10102
rect 10041 10099 10107 10102
rect 4705 10026 4771 10029
rect 6453 10026 6519 10029
rect 4705 10024 6519 10026
rect 4705 9968 4710 10024
rect 4766 9968 6458 10024
rect 6514 9968 6519 10024
rect 4705 9966 6519 9968
rect 4705 9963 4771 9966
rect 6453 9963 6519 9966
rect 6729 10026 6795 10029
rect 9029 10026 9095 10029
rect 10041 10028 10107 10029
rect 9990 10026 9996 10028
rect 6729 10024 9095 10026
rect 6729 9968 6734 10024
rect 6790 9968 9034 10024
rect 9090 9968 9095 10024
rect 6729 9966 9095 9968
rect 9950 9966 9996 10026
rect 10060 10026 10107 10028
rect 10961 10026 11027 10029
rect 10060 10024 11027 10026
rect 10102 9968 10966 10024
rect 11022 9968 11027 10024
rect 6729 9963 6795 9966
rect 9029 9963 9095 9966
rect 9990 9964 9996 9966
rect 10060 9966 11027 9968
rect 10060 9964 10107 9966
rect 10041 9963 10107 9964
rect 10961 9963 11027 9966
rect 6453 9890 6519 9893
rect 7005 9890 7071 9893
rect 6453 9888 7071 9890
rect 6453 9832 6458 9888
rect 6514 9832 7010 9888
rect 7066 9832 7071 9888
rect 6453 9830 7071 9832
rect 6453 9827 6519 9830
rect 7005 9827 7071 9830
rect 8210 9824 8526 9825
rect 0 9754 800 9784
rect 8210 9760 8216 9824
rect 8280 9760 8296 9824
rect 8360 9760 8376 9824
rect 8440 9760 8456 9824
rect 8520 9760 8526 9824
rect 8210 9759 8526 9760
rect 3969 9754 4035 9757
rect 0 9752 4035 9754
rect 0 9696 3974 9752
rect 4030 9696 4035 9752
rect 0 9694 4035 9696
rect 0 9664 800 9694
rect 3969 9691 4035 9694
rect 7189 9752 7255 9757
rect 10133 9756 10199 9757
rect 10133 9754 10180 9756
rect 7189 9696 7194 9752
rect 7250 9696 7255 9752
rect 7189 9691 7255 9696
rect 10088 9752 10180 9754
rect 10088 9696 10138 9752
rect 10088 9694 10180 9696
rect 10133 9692 10180 9694
rect 10244 9692 10250 9756
rect 10777 9754 10843 9757
rect 11697 9754 11763 9757
rect 10777 9752 11763 9754
rect 10777 9696 10782 9752
rect 10838 9696 11702 9752
rect 11758 9696 11763 9752
rect 10777 9694 11763 9696
rect 10133 9691 10199 9692
rect 10777 9691 10843 9694
rect 11697 9691 11763 9694
rect 5809 9618 5875 9621
rect 7192 9618 7252 9691
rect 11053 9618 11119 9621
rect 12985 9618 13051 9621
rect 5809 9616 7252 9618
rect 5809 9560 5814 9616
rect 5870 9560 7252 9616
rect 5809 9558 7252 9560
rect 7468 9616 13051 9618
rect 7468 9560 11058 9616
rect 11114 9560 12990 9616
rect 13046 9560 13051 9616
rect 7468 9558 13051 9560
rect 5809 9555 5875 9558
rect 6729 9482 6795 9485
rect 7468 9482 7528 9558
rect 11053 9555 11119 9558
rect 12985 9555 13051 9558
rect 6729 9480 7528 9482
rect 6729 9424 6734 9480
rect 6790 9424 7528 9480
rect 6729 9422 7528 9424
rect 7649 9480 7715 9485
rect 7649 9424 7654 9480
rect 7710 9424 7715 9480
rect 6729 9419 6795 9422
rect 7649 9419 7715 9424
rect 7833 9482 7899 9485
rect 11145 9482 11211 9485
rect 7833 9480 11211 9482
rect 7833 9424 7838 9480
rect 7894 9424 11150 9480
rect 11206 9424 11211 9480
rect 7833 9422 11211 9424
rect 7833 9419 7899 9422
rect 11145 9419 11211 9422
rect 7097 9346 7163 9349
rect 7652 9346 7712 9419
rect 9857 9346 9923 9349
rect 7097 9344 9923 9346
rect 7097 9288 7102 9344
rect 7158 9288 9862 9344
rect 9918 9288 9923 9344
rect 7097 9286 9923 9288
rect 7097 9283 7163 9286
rect 9857 9283 9923 9286
rect 10685 9346 10751 9349
rect 11421 9346 11487 9349
rect 10685 9344 11487 9346
rect 10685 9288 10690 9344
rect 10746 9288 11426 9344
rect 11482 9288 11487 9344
rect 10685 9286 11487 9288
rect 10685 9283 10751 9286
rect 11421 9283 11487 9286
rect 4210 9280 4526 9281
rect 4210 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4526 9280
rect 4210 9215 4526 9216
rect 12210 9280 12526 9281
rect 12210 9216 12216 9280
rect 12280 9216 12296 9280
rect 12360 9216 12376 9280
rect 12440 9216 12456 9280
rect 12520 9216 12526 9280
rect 12210 9215 12526 9216
rect 3785 9210 3851 9213
rect 6269 9210 6335 9213
rect 8753 9210 8819 9213
rect 12065 9210 12131 9213
rect 3785 9208 3986 9210
rect 3785 9152 3790 9208
rect 3846 9152 3986 9208
rect 3785 9150 3986 9152
rect 3785 9147 3851 9150
rect 3926 9074 3986 9150
rect 6269 9208 12131 9210
rect 6269 9152 6274 9208
rect 6330 9152 8758 9208
rect 8814 9152 12070 9208
rect 12126 9152 12131 9208
rect 6269 9150 12131 9152
rect 6269 9147 6335 9150
rect 8753 9147 8819 9150
rect 12065 9147 12131 9150
rect 8753 9074 8819 9077
rect 9489 9074 9555 9077
rect 3926 9072 8819 9074
rect 3926 9016 8758 9072
rect 8814 9016 8819 9072
rect 3926 9014 8819 9016
rect 8753 9011 8819 9014
rect 8894 9072 9555 9074
rect 8894 9016 9494 9072
rect 9550 9016 9555 9072
rect 8894 9014 9555 9016
rect 1485 8938 1551 8941
rect 6913 8938 6979 8941
rect 1485 8936 6979 8938
rect 1485 8880 1490 8936
rect 1546 8880 6918 8936
rect 6974 8880 6979 8936
rect 1485 8878 6979 8880
rect 1485 8875 1551 8878
rect 6913 8875 6979 8878
rect 7833 8938 7899 8941
rect 7966 8938 7972 8940
rect 7833 8936 7972 8938
rect 7833 8880 7838 8936
rect 7894 8880 7972 8936
rect 7833 8878 7972 8880
rect 7833 8875 7899 8878
rect 7966 8876 7972 8878
rect 8036 8876 8042 8940
rect 8293 8938 8359 8941
rect 8894 8938 8954 9014
rect 9489 9011 9555 9014
rect 8293 8936 8954 8938
rect 8293 8880 8298 8936
rect 8354 8880 8954 8936
rect 8293 8878 8954 8880
rect 8293 8875 8359 8878
rect 0 8802 800 8832
rect 3877 8802 3943 8805
rect 0 8800 3943 8802
rect 0 8744 3882 8800
rect 3938 8744 3943 8800
rect 0 8742 3943 8744
rect 0 8712 800 8742
rect 3877 8739 3943 8742
rect 13629 8802 13695 8805
rect 14200 8802 15000 8832
rect 13629 8800 15000 8802
rect 13629 8744 13634 8800
rect 13690 8744 15000 8800
rect 13629 8742 15000 8744
rect 13629 8739 13695 8742
rect 8210 8736 8526 8737
rect 8210 8672 8216 8736
rect 8280 8672 8296 8736
rect 8360 8672 8376 8736
rect 8440 8672 8456 8736
rect 8520 8672 8526 8736
rect 14200 8712 15000 8742
rect 8210 8671 8526 8672
rect 5073 8666 5139 8669
rect 7833 8666 7899 8669
rect 5073 8664 7899 8666
rect 5073 8608 5078 8664
rect 5134 8608 7838 8664
rect 7894 8608 7899 8664
rect 5073 8606 7899 8608
rect 5073 8603 5139 8606
rect 7833 8603 7899 8606
rect 8201 8530 8267 8533
rect 9070 8530 9076 8532
rect 8201 8528 9076 8530
rect 8201 8472 8206 8528
rect 8262 8472 9076 8528
rect 8201 8470 9076 8472
rect 8201 8467 8267 8470
rect 9070 8468 9076 8470
rect 9140 8530 9146 8532
rect 11605 8530 11671 8533
rect 9140 8528 11671 8530
rect 9140 8472 11610 8528
rect 11666 8472 11671 8528
rect 9140 8470 11671 8472
rect 9140 8468 9146 8470
rect 11605 8467 11671 8470
rect 7189 8394 7255 8397
rect 10041 8394 10107 8397
rect 7189 8392 10107 8394
rect 7189 8336 7194 8392
rect 7250 8336 10046 8392
rect 10102 8336 10107 8392
rect 7189 8334 10107 8336
rect 7189 8331 7255 8334
rect 10041 8331 10107 8334
rect 6545 8258 6611 8261
rect 10225 8258 10291 8261
rect 6545 8256 10291 8258
rect 6545 8200 6550 8256
rect 6606 8200 10230 8256
rect 10286 8200 10291 8256
rect 6545 8198 10291 8200
rect 6545 8195 6611 8198
rect 10225 8195 10291 8198
rect 12617 8258 12683 8261
rect 12893 8258 12959 8261
rect 12617 8256 12959 8258
rect 12617 8200 12622 8256
rect 12678 8200 12898 8256
rect 12954 8200 12959 8256
rect 12617 8198 12959 8200
rect 12617 8195 12683 8198
rect 12893 8195 12959 8198
rect 4210 8192 4526 8193
rect 4210 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4526 8192
rect 4210 8127 4526 8128
rect 12210 8192 12526 8193
rect 12210 8128 12216 8192
rect 12280 8128 12296 8192
rect 12360 8128 12376 8192
rect 12440 8128 12456 8192
rect 12520 8128 12526 8192
rect 12210 8127 12526 8128
rect 5165 8122 5231 8125
rect 7189 8122 7255 8125
rect 5165 8120 7255 8122
rect 5165 8064 5170 8120
rect 5226 8064 7194 8120
rect 7250 8064 7255 8120
rect 5165 8062 7255 8064
rect 5165 8059 5231 8062
rect 7189 8059 7255 8062
rect 9765 8122 9831 8125
rect 10685 8122 10751 8125
rect 9765 8120 10751 8122
rect 9765 8064 9770 8120
rect 9826 8064 10690 8120
rect 10746 8064 10751 8120
rect 9765 8062 10751 8064
rect 9765 8059 9831 8062
rect 10685 8059 10751 8062
rect 0 7986 800 8016
rect 2957 7986 3023 7989
rect 3601 7986 3667 7989
rect 0 7984 3667 7986
rect 0 7928 2962 7984
rect 3018 7928 3606 7984
rect 3662 7928 3667 7984
rect 0 7926 3667 7928
rect 0 7896 800 7926
rect 2957 7923 3023 7926
rect 3601 7923 3667 7926
rect 10225 7986 10291 7989
rect 10409 7986 10475 7989
rect 10225 7984 10475 7986
rect 10225 7928 10230 7984
rect 10286 7928 10414 7984
rect 10470 7928 10475 7984
rect 10225 7926 10475 7928
rect 10225 7923 10291 7926
rect 10409 7923 10475 7926
rect 10593 7986 10659 7989
rect 10777 7986 10843 7989
rect 10593 7984 10843 7986
rect 10593 7928 10598 7984
rect 10654 7928 10782 7984
rect 10838 7928 10843 7984
rect 10593 7926 10843 7928
rect 10593 7923 10659 7926
rect 10777 7923 10843 7926
rect 7966 7788 7972 7852
rect 8036 7850 8042 7852
rect 9765 7850 9831 7853
rect 8036 7848 9831 7850
rect 8036 7792 9770 7848
rect 9826 7792 9831 7848
rect 8036 7790 9831 7792
rect 8036 7788 8042 7790
rect 9765 7787 9831 7790
rect 10777 7850 10843 7853
rect 11053 7850 11119 7853
rect 10777 7848 11119 7850
rect 10777 7792 10782 7848
rect 10838 7792 11058 7848
rect 11114 7792 11119 7848
rect 10777 7790 11119 7792
rect 10777 7787 10843 7790
rect 11053 7787 11119 7790
rect 8845 7714 8911 7717
rect 10685 7714 10751 7717
rect 8845 7712 10751 7714
rect 8845 7656 8850 7712
rect 8906 7656 10690 7712
rect 10746 7656 10751 7712
rect 8845 7654 10751 7656
rect 8845 7651 8911 7654
rect 10685 7651 10751 7654
rect 8210 7648 8526 7649
rect 8210 7584 8216 7648
rect 8280 7584 8296 7648
rect 8360 7584 8376 7648
rect 8440 7584 8456 7648
rect 8520 7584 8526 7648
rect 8210 7583 8526 7584
rect 8385 7442 8451 7445
rect 13169 7442 13235 7445
rect 8385 7440 13235 7442
rect 8385 7384 8390 7440
rect 8446 7384 13174 7440
rect 13230 7384 13235 7440
rect 8385 7382 13235 7384
rect 8385 7379 8451 7382
rect 13169 7379 13235 7382
rect 4210 7104 4526 7105
rect 0 7034 800 7064
rect 4210 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4526 7104
rect 4210 7039 4526 7040
rect 12210 7104 12526 7105
rect 12210 7040 12216 7104
rect 12280 7040 12296 7104
rect 12360 7040 12376 7104
rect 12440 7040 12456 7104
rect 12520 7040 12526 7104
rect 12210 7039 12526 7040
rect 2865 7034 2931 7037
rect 0 7032 2931 7034
rect 0 6976 2870 7032
rect 2926 6976 2931 7032
rect 0 6974 2931 6976
rect 0 6944 800 6974
rect 2865 6971 2931 6974
rect 10041 7034 10107 7037
rect 11421 7034 11487 7037
rect 10041 7032 11487 7034
rect 10041 6976 10046 7032
rect 10102 6976 11426 7032
rect 11482 6976 11487 7032
rect 10041 6974 11487 6976
rect 10041 6971 10107 6974
rect 11421 6971 11487 6974
rect 8210 6560 8526 6561
rect 8210 6496 8216 6560
rect 8280 6496 8296 6560
rect 8360 6496 8376 6560
rect 8440 6496 8456 6560
rect 8520 6496 8526 6560
rect 8210 6495 8526 6496
rect 6269 6354 6335 6357
rect 12801 6354 12867 6357
rect 6269 6352 12867 6354
rect 6269 6296 6274 6352
rect 6330 6296 12806 6352
rect 12862 6296 12867 6352
rect 6269 6294 12867 6296
rect 6269 6291 6335 6294
rect 12801 6291 12867 6294
rect 2589 6218 2655 6221
rect 4245 6218 4311 6221
rect 5993 6218 6059 6221
rect 2589 6216 6059 6218
rect 2589 6160 2594 6216
rect 2650 6160 4250 6216
rect 4306 6160 5998 6216
rect 6054 6160 6059 6216
rect 2589 6158 6059 6160
rect 2589 6155 2655 6158
rect 4245 6155 4311 6158
rect 5993 6155 6059 6158
rect 10961 6218 11027 6221
rect 14200 6218 15000 6248
rect 10961 6216 15000 6218
rect 10961 6160 10966 6216
rect 11022 6160 15000 6216
rect 10961 6158 15000 6160
rect 10961 6155 11027 6158
rect 14200 6128 15000 6158
rect 0 6082 800 6112
rect 2957 6082 3023 6085
rect 3969 6082 4035 6085
rect 0 6080 4035 6082
rect 0 6024 2962 6080
rect 3018 6024 3974 6080
rect 4030 6024 4035 6080
rect 0 6022 4035 6024
rect 0 5992 800 6022
rect 2957 6019 3023 6022
rect 3969 6019 4035 6022
rect 4210 6016 4526 6017
rect 4210 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4526 6016
rect 4210 5951 4526 5952
rect 12210 6016 12526 6017
rect 12210 5952 12216 6016
rect 12280 5952 12296 6016
rect 12360 5952 12376 6016
rect 12440 5952 12456 6016
rect 12520 5952 12526 6016
rect 12210 5951 12526 5952
rect 4981 5674 5047 5677
rect 4981 5672 5090 5674
rect 4981 5616 4986 5672
rect 5042 5616 5090 5672
rect 4981 5611 5090 5616
rect 5030 5538 5090 5611
rect 5257 5538 5323 5541
rect 5030 5536 5323 5538
rect 5030 5480 5262 5536
rect 5318 5480 5323 5536
rect 5030 5478 5323 5480
rect 5257 5475 5323 5478
rect 8210 5472 8526 5473
rect 8210 5408 8216 5472
rect 8280 5408 8296 5472
rect 8360 5408 8376 5472
rect 8440 5408 8456 5472
rect 8520 5408 8526 5472
rect 8210 5407 8526 5408
rect 2865 5266 2931 5269
rect 4613 5266 4679 5269
rect 2865 5264 4679 5266
rect 2865 5208 2870 5264
rect 2926 5208 4618 5264
rect 4674 5208 4679 5264
rect 2865 5206 4679 5208
rect 2865 5203 2931 5206
rect 4613 5203 4679 5206
rect 0 5130 800 5160
rect 1393 5130 1459 5133
rect 4061 5130 4127 5133
rect 0 5128 4127 5130
rect 0 5072 1398 5128
rect 1454 5072 4066 5128
rect 4122 5072 4127 5128
rect 0 5070 4127 5072
rect 0 5040 800 5070
rect 1393 5067 1459 5070
rect 4061 5067 4127 5070
rect 4210 4928 4526 4929
rect 4210 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4526 4928
rect 4210 4863 4526 4864
rect 12210 4928 12526 4929
rect 12210 4864 12216 4928
rect 12280 4864 12296 4928
rect 12360 4864 12376 4928
rect 12440 4864 12456 4928
rect 12520 4864 12526 4928
rect 12210 4863 12526 4864
rect 8210 4384 8526 4385
rect 8210 4320 8216 4384
rect 8280 4320 8296 4384
rect 8360 4320 8376 4384
rect 8440 4320 8456 4384
rect 8520 4320 8526 4384
rect 8210 4319 8526 4320
rect 0 4178 800 4208
rect 4061 4178 4127 4181
rect 0 4176 4127 4178
rect 0 4120 4066 4176
rect 4122 4120 4127 4176
rect 0 4118 4127 4120
rect 0 4088 800 4118
rect 4061 4115 4127 4118
rect 4210 3840 4526 3841
rect 4210 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4526 3840
rect 4210 3775 4526 3776
rect 12210 3840 12526 3841
rect 12210 3776 12216 3840
rect 12280 3776 12296 3840
rect 12360 3776 12376 3840
rect 12440 3776 12456 3840
rect 12520 3776 12526 3840
rect 12210 3775 12526 3776
rect 12709 3770 12775 3773
rect 14200 3770 15000 3800
rect 12709 3768 15000 3770
rect 12709 3712 12714 3768
rect 12770 3712 15000 3768
rect 12709 3710 15000 3712
rect 12709 3707 12775 3710
rect 14200 3680 15000 3710
rect 8210 3296 8526 3297
rect 0 3226 800 3256
rect 8210 3232 8216 3296
rect 8280 3232 8296 3296
rect 8360 3232 8376 3296
rect 8440 3232 8456 3296
rect 8520 3232 8526 3296
rect 8210 3231 8526 3232
rect 3049 3226 3115 3229
rect 4061 3226 4127 3229
rect 0 3224 4127 3226
rect 0 3168 3054 3224
rect 3110 3168 4066 3224
rect 4122 3168 4127 3224
rect 0 3166 4127 3168
rect 0 3136 800 3166
rect 3049 3163 3115 3166
rect 4061 3163 4127 3166
rect 4210 2752 4526 2753
rect 4210 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4526 2752
rect 4210 2687 4526 2688
rect 12210 2752 12526 2753
rect 12210 2688 12216 2752
rect 12280 2688 12296 2752
rect 12360 2688 12376 2752
rect 12440 2688 12456 2752
rect 12520 2688 12526 2752
rect 12210 2687 12526 2688
rect 5073 2682 5139 2685
rect 11237 2682 11303 2685
rect 5073 2680 11303 2682
rect 5073 2624 5078 2680
rect 5134 2624 11242 2680
rect 11298 2624 11303 2680
rect 5073 2622 11303 2624
rect 5073 2619 5139 2622
rect 11237 2619 11303 2622
rect 2313 2546 2379 2549
rect 7097 2546 7163 2549
rect 2313 2544 7163 2546
rect 2313 2488 2318 2544
rect 2374 2488 7102 2544
rect 7158 2488 7163 2544
rect 2313 2486 7163 2488
rect 2313 2483 2379 2486
rect 7097 2483 7163 2486
rect 8477 2546 8543 2549
rect 11053 2546 11119 2549
rect 8477 2544 11119 2546
rect 8477 2488 8482 2544
rect 8538 2488 11058 2544
rect 11114 2488 11119 2544
rect 8477 2486 11119 2488
rect 8477 2483 8543 2486
rect 11053 2483 11119 2486
rect 1669 2410 1735 2413
rect 4061 2410 4127 2413
rect 1669 2408 4127 2410
rect 1669 2352 1674 2408
rect 1730 2352 4066 2408
rect 4122 2352 4127 2408
rect 1669 2350 4127 2352
rect 1669 2347 1735 2350
rect 4061 2347 4127 2350
rect 0 2274 800 2304
rect 2773 2274 2839 2277
rect 0 2272 2839 2274
rect 0 2216 2778 2272
rect 2834 2216 2839 2272
rect 0 2214 2839 2216
rect 0 2184 800 2214
rect 2773 2211 2839 2214
rect 9121 2274 9187 2277
rect 11513 2274 11579 2277
rect 9121 2272 11579 2274
rect 9121 2216 9126 2272
rect 9182 2216 11518 2272
rect 11574 2216 11579 2272
rect 9121 2214 11579 2216
rect 9121 2211 9187 2214
rect 11513 2211 11579 2214
rect 8210 2208 8526 2209
rect 8210 2144 8216 2208
rect 8280 2144 8296 2208
rect 8360 2144 8376 2208
rect 8440 2144 8456 2208
rect 8520 2144 8526 2208
rect 8210 2143 8526 2144
rect 1669 2002 1735 2005
rect 4153 2002 4219 2005
rect 1669 2000 4219 2002
rect 1669 1944 1674 2000
rect 1730 1944 4158 2000
rect 4214 1944 4219 2000
rect 1669 1942 4219 1944
rect 1669 1939 1735 1942
rect 4153 1939 4219 1942
rect 3693 1866 3759 1869
rect 9305 1866 9371 1869
rect 3693 1864 9371 1866
rect 3693 1808 3698 1864
rect 3754 1808 9310 1864
rect 9366 1808 9371 1864
rect 3693 1806 9371 1808
rect 3693 1803 3759 1806
rect 9305 1803 9371 1806
rect 4210 1664 4526 1665
rect 4210 1600 4216 1664
rect 4280 1600 4296 1664
rect 4360 1600 4376 1664
rect 4440 1600 4456 1664
rect 4520 1600 4526 1664
rect 4210 1599 4526 1600
rect 12210 1664 12526 1665
rect 12210 1600 12216 1664
rect 12280 1600 12296 1664
rect 12360 1600 12376 1664
rect 12440 1600 12456 1664
rect 12520 1600 12526 1664
rect 12210 1599 12526 1600
rect 0 1322 800 1352
rect 3877 1322 3943 1325
rect 0 1320 3943 1322
rect 0 1264 3882 1320
rect 3938 1264 3943 1320
rect 0 1262 3943 1264
rect 0 1232 800 1262
rect 3877 1259 3943 1262
rect 13537 1322 13603 1325
rect 14200 1322 15000 1352
rect 13537 1320 15000 1322
rect 13537 1264 13542 1320
rect 13598 1264 15000 1320
rect 13537 1262 15000 1264
rect 13537 1259 13603 1262
rect 14200 1232 15000 1262
rect 8210 1120 8526 1121
rect 8210 1056 8216 1120
rect 8280 1056 8296 1120
rect 8360 1056 8376 1120
rect 8440 1056 8456 1120
rect 8520 1056 8526 1120
rect 8210 1055 8526 1056
rect 0 506 800 536
rect 1393 506 1459 509
rect 0 504 1459 506
rect 0 448 1398 504
rect 1454 448 1459 504
rect 0 446 1459 448
rect 0 416 800 446
rect 1393 443 1459 446
<< via3 >>
rect 4216 13628 4280 13632
rect 4216 13572 4220 13628
rect 4220 13572 4276 13628
rect 4276 13572 4280 13628
rect 4216 13568 4280 13572
rect 4296 13628 4360 13632
rect 4296 13572 4300 13628
rect 4300 13572 4356 13628
rect 4356 13572 4360 13628
rect 4296 13568 4360 13572
rect 4376 13628 4440 13632
rect 4376 13572 4380 13628
rect 4380 13572 4436 13628
rect 4436 13572 4440 13628
rect 4376 13568 4440 13572
rect 4456 13628 4520 13632
rect 4456 13572 4460 13628
rect 4460 13572 4516 13628
rect 4516 13572 4520 13628
rect 4456 13568 4520 13572
rect 12216 13628 12280 13632
rect 12216 13572 12220 13628
rect 12220 13572 12276 13628
rect 12276 13572 12280 13628
rect 12216 13568 12280 13572
rect 12296 13628 12360 13632
rect 12296 13572 12300 13628
rect 12300 13572 12356 13628
rect 12356 13572 12360 13628
rect 12296 13568 12360 13572
rect 12376 13628 12440 13632
rect 12376 13572 12380 13628
rect 12380 13572 12436 13628
rect 12436 13572 12440 13628
rect 12376 13568 12440 13572
rect 12456 13628 12520 13632
rect 12456 13572 12460 13628
rect 12460 13572 12516 13628
rect 12516 13572 12520 13628
rect 12456 13568 12520 13572
rect 6316 13500 6380 13564
rect 9444 13228 9508 13292
rect 8216 13084 8280 13088
rect 8216 13028 8220 13084
rect 8220 13028 8276 13084
rect 8276 13028 8280 13084
rect 8216 13024 8280 13028
rect 8296 13084 8360 13088
rect 8296 13028 8300 13084
rect 8300 13028 8356 13084
rect 8356 13028 8360 13084
rect 8296 13024 8360 13028
rect 8376 13084 8440 13088
rect 8376 13028 8380 13084
rect 8380 13028 8436 13084
rect 8436 13028 8440 13084
rect 8376 13024 8440 13028
rect 8456 13084 8520 13088
rect 8456 13028 8460 13084
rect 8460 13028 8516 13084
rect 8516 13028 8520 13084
rect 8456 13024 8520 13028
rect 8708 12820 8772 12884
rect 4216 12540 4280 12544
rect 4216 12484 4220 12540
rect 4220 12484 4276 12540
rect 4276 12484 4280 12540
rect 4216 12480 4280 12484
rect 4296 12540 4360 12544
rect 4296 12484 4300 12540
rect 4300 12484 4356 12540
rect 4356 12484 4360 12540
rect 4296 12480 4360 12484
rect 4376 12540 4440 12544
rect 4376 12484 4380 12540
rect 4380 12484 4436 12540
rect 4436 12484 4440 12540
rect 4376 12480 4440 12484
rect 4456 12540 4520 12544
rect 4456 12484 4460 12540
rect 4460 12484 4516 12540
rect 4516 12484 4520 12540
rect 4456 12480 4520 12484
rect 12216 12540 12280 12544
rect 12216 12484 12220 12540
rect 12220 12484 12276 12540
rect 12276 12484 12280 12540
rect 12216 12480 12280 12484
rect 12296 12540 12360 12544
rect 12296 12484 12300 12540
rect 12300 12484 12356 12540
rect 12356 12484 12360 12540
rect 12296 12480 12360 12484
rect 12376 12540 12440 12544
rect 12376 12484 12380 12540
rect 12380 12484 12436 12540
rect 12436 12484 12440 12540
rect 12376 12480 12440 12484
rect 12456 12540 12520 12544
rect 12456 12484 12460 12540
rect 12460 12484 12516 12540
rect 12516 12484 12520 12540
rect 12456 12480 12520 12484
rect 8216 11996 8280 12000
rect 8216 11940 8220 11996
rect 8220 11940 8276 11996
rect 8276 11940 8280 11996
rect 8216 11936 8280 11940
rect 8296 11996 8360 12000
rect 8296 11940 8300 11996
rect 8300 11940 8356 11996
rect 8356 11940 8360 11996
rect 8296 11936 8360 11940
rect 8376 11996 8440 12000
rect 8376 11940 8380 11996
rect 8380 11940 8436 11996
rect 8436 11940 8440 11996
rect 8376 11936 8440 11940
rect 8456 11996 8520 12000
rect 8456 11940 8460 11996
rect 8460 11940 8516 11996
rect 8516 11940 8520 11996
rect 8456 11936 8520 11940
rect 4216 11452 4280 11456
rect 4216 11396 4220 11452
rect 4220 11396 4276 11452
rect 4276 11396 4280 11452
rect 4216 11392 4280 11396
rect 4296 11452 4360 11456
rect 4296 11396 4300 11452
rect 4300 11396 4356 11452
rect 4356 11396 4360 11452
rect 4296 11392 4360 11396
rect 4376 11452 4440 11456
rect 4376 11396 4380 11452
rect 4380 11396 4436 11452
rect 4436 11396 4440 11452
rect 4376 11392 4440 11396
rect 4456 11452 4520 11456
rect 4456 11396 4460 11452
rect 4460 11396 4516 11452
rect 4516 11396 4520 11452
rect 4456 11392 4520 11396
rect 10180 11868 10244 11932
rect 12216 11452 12280 11456
rect 12216 11396 12220 11452
rect 12220 11396 12276 11452
rect 12276 11396 12280 11452
rect 12216 11392 12280 11396
rect 12296 11452 12360 11456
rect 12296 11396 12300 11452
rect 12300 11396 12356 11452
rect 12356 11396 12360 11452
rect 12296 11392 12360 11396
rect 12376 11452 12440 11456
rect 12376 11396 12380 11452
rect 12380 11396 12436 11452
rect 12436 11396 12440 11452
rect 12376 11392 12440 11396
rect 12456 11452 12520 11456
rect 12456 11396 12460 11452
rect 12460 11396 12516 11452
rect 12516 11396 12520 11452
rect 12456 11392 12520 11396
rect 9076 11384 9140 11388
rect 9076 11328 9126 11384
rect 9126 11328 9140 11384
rect 9076 11324 9140 11328
rect 9260 11324 9324 11388
rect 7972 11188 8036 11252
rect 9996 11188 10060 11252
rect 8216 10908 8280 10912
rect 8216 10852 8220 10908
rect 8220 10852 8276 10908
rect 8276 10852 8280 10908
rect 8216 10848 8280 10852
rect 8296 10908 8360 10912
rect 8296 10852 8300 10908
rect 8300 10852 8356 10908
rect 8356 10852 8360 10908
rect 8296 10848 8360 10852
rect 8376 10908 8440 10912
rect 8376 10852 8380 10908
rect 8380 10852 8436 10908
rect 8436 10852 8440 10908
rect 8376 10848 8440 10852
rect 8456 10908 8520 10912
rect 8456 10852 8460 10908
rect 8460 10852 8516 10908
rect 8516 10852 8520 10908
rect 8456 10848 8520 10852
rect 8708 10780 8772 10844
rect 9260 10644 9324 10708
rect 9444 10568 9508 10572
rect 9444 10512 9494 10568
rect 9494 10512 9508 10568
rect 9444 10508 9508 10512
rect 4216 10364 4280 10368
rect 4216 10308 4220 10364
rect 4220 10308 4276 10364
rect 4276 10308 4280 10364
rect 4216 10304 4280 10308
rect 4296 10364 4360 10368
rect 4296 10308 4300 10364
rect 4300 10308 4356 10364
rect 4356 10308 4360 10364
rect 4296 10304 4360 10308
rect 4376 10364 4440 10368
rect 4376 10308 4380 10364
rect 4380 10308 4436 10364
rect 4436 10308 4440 10364
rect 4376 10304 4440 10308
rect 4456 10364 4520 10368
rect 4456 10308 4460 10364
rect 4460 10308 4516 10364
rect 4516 10308 4520 10364
rect 4456 10304 4520 10308
rect 12216 10364 12280 10368
rect 12216 10308 12220 10364
rect 12220 10308 12276 10364
rect 12276 10308 12280 10364
rect 12216 10304 12280 10308
rect 12296 10364 12360 10368
rect 12296 10308 12300 10364
rect 12300 10308 12356 10364
rect 12356 10308 12360 10364
rect 12296 10304 12360 10308
rect 12376 10364 12440 10368
rect 12376 10308 12380 10364
rect 12380 10308 12436 10364
rect 12436 10308 12440 10364
rect 12376 10304 12440 10308
rect 12456 10364 12520 10368
rect 12456 10308 12460 10364
rect 12460 10308 12516 10364
rect 12516 10308 12520 10364
rect 12456 10304 12520 10308
rect 10180 10236 10244 10300
rect 6316 10160 6380 10164
rect 6316 10104 6330 10160
rect 6330 10104 6380 10160
rect 6316 10100 6380 10104
rect 9996 10024 10060 10028
rect 9996 9968 10046 10024
rect 10046 9968 10060 10024
rect 9996 9964 10060 9968
rect 8216 9820 8280 9824
rect 8216 9764 8220 9820
rect 8220 9764 8276 9820
rect 8276 9764 8280 9820
rect 8216 9760 8280 9764
rect 8296 9820 8360 9824
rect 8296 9764 8300 9820
rect 8300 9764 8356 9820
rect 8356 9764 8360 9820
rect 8296 9760 8360 9764
rect 8376 9820 8440 9824
rect 8376 9764 8380 9820
rect 8380 9764 8436 9820
rect 8436 9764 8440 9820
rect 8376 9760 8440 9764
rect 8456 9820 8520 9824
rect 8456 9764 8460 9820
rect 8460 9764 8516 9820
rect 8516 9764 8520 9820
rect 8456 9760 8520 9764
rect 10180 9752 10244 9756
rect 10180 9696 10194 9752
rect 10194 9696 10244 9752
rect 10180 9692 10244 9696
rect 4216 9276 4280 9280
rect 4216 9220 4220 9276
rect 4220 9220 4276 9276
rect 4276 9220 4280 9276
rect 4216 9216 4280 9220
rect 4296 9276 4360 9280
rect 4296 9220 4300 9276
rect 4300 9220 4356 9276
rect 4356 9220 4360 9276
rect 4296 9216 4360 9220
rect 4376 9276 4440 9280
rect 4376 9220 4380 9276
rect 4380 9220 4436 9276
rect 4436 9220 4440 9276
rect 4376 9216 4440 9220
rect 4456 9276 4520 9280
rect 4456 9220 4460 9276
rect 4460 9220 4516 9276
rect 4516 9220 4520 9276
rect 4456 9216 4520 9220
rect 12216 9276 12280 9280
rect 12216 9220 12220 9276
rect 12220 9220 12276 9276
rect 12276 9220 12280 9276
rect 12216 9216 12280 9220
rect 12296 9276 12360 9280
rect 12296 9220 12300 9276
rect 12300 9220 12356 9276
rect 12356 9220 12360 9276
rect 12296 9216 12360 9220
rect 12376 9276 12440 9280
rect 12376 9220 12380 9276
rect 12380 9220 12436 9276
rect 12436 9220 12440 9276
rect 12376 9216 12440 9220
rect 12456 9276 12520 9280
rect 12456 9220 12460 9276
rect 12460 9220 12516 9276
rect 12516 9220 12520 9276
rect 12456 9216 12520 9220
rect 7972 8876 8036 8940
rect 8216 8732 8280 8736
rect 8216 8676 8220 8732
rect 8220 8676 8276 8732
rect 8276 8676 8280 8732
rect 8216 8672 8280 8676
rect 8296 8732 8360 8736
rect 8296 8676 8300 8732
rect 8300 8676 8356 8732
rect 8356 8676 8360 8732
rect 8296 8672 8360 8676
rect 8376 8732 8440 8736
rect 8376 8676 8380 8732
rect 8380 8676 8436 8732
rect 8436 8676 8440 8732
rect 8376 8672 8440 8676
rect 8456 8732 8520 8736
rect 8456 8676 8460 8732
rect 8460 8676 8516 8732
rect 8516 8676 8520 8732
rect 8456 8672 8520 8676
rect 9076 8468 9140 8532
rect 4216 8188 4280 8192
rect 4216 8132 4220 8188
rect 4220 8132 4276 8188
rect 4276 8132 4280 8188
rect 4216 8128 4280 8132
rect 4296 8188 4360 8192
rect 4296 8132 4300 8188
rect 4300 8132 4356 8188
rect 4356 8132 4360 8188
rect 4296 8128 4360 8132
rect 4376 8188 4440 8192
rect 4376 8132 4380 8188
rect 4380 8132 4436 8188
rect 4436 8132 4440 8188
rect 4376 8128 4440 8132
rect 4456 8188 4520 8192
rect 4456 8132 4460 8188
rect 4460 8132 4516 8188
rect 4516 8132 4520 8188
rect 4456 8128 4520 8132
rect 12216 8188 12280 8192
rect 12216 8132 12220 8188
rect 12220 8132 12276 8188
rect 12276 8132 12280 8188
rect 12216 8128 12280 8132
rect 12296 8188 12360 8192
rect 12296 8132 12300 8188
rect 12300 8132 12356 8188
rect 12356 8132 12360 8188
rect 12296 8128 12360 8132
rect 12376 8188 12440 8192
rect 12376 8132 12380 8188
rect 12380 8132 12436 8188
rect 12436 8132 12440 8188
rect 12376 8128 12440 8132
rect 12456 8188 12520 8192
rect 12456 8132 12460 8188
rect 12460 8132 12516 8188
rect 12516 8132 12520 8188
rect 12456 8128 12520 8132
rect 7972 7788 8036 7852
rect 8216 7644 8280 7648
rect 8216 7588 8220 7644
rect 8220 7588 8276 7644
rect 8276 7588 8280 7644
rect 8216 7584 8280 7588
rect 8296 7644 8360 7648
rect 8296 7588 8300 7644
rect 8300 7588 8356 7644
rect 8356 7588 8360 7644
rect 8296 7584 8360 7588
rect 8376 7644 8440 7648
rect 8376 7588 8380 7644
rect 8380 7588 8436 7644
rect 8436 7588 8440 7644
rect 8376 7584 8440 7588
rect 8456 7644 8520 7648
rect 8456 7588 8460 7644
rect 8460 7588 8516 7644
rect 8516 7588 8520 7644
rect 8456 7584 8520 7588
rect 4216 7100 4280 7104
rect 4216 7044 4220 7100
rect 4220 7044 4276 7100
rect 4276 7044 4280 7100
rect 4216 7040 4280 7044
rect 4296 7100 4360 7104
rect 4296 7044 4300 7100
rect 4300 7044 4356 7100
rect 4356 7044 4360 7100
rect 4296 7040 4360 7044
rect 4376 7100 4440 7104
rect 4376 7044 4380 7100
rect 4380 7044 4436 7100
rect 4436 7044 4440 7100
rect 4376 7040 4440 7044
rect 4456 7100 4520 7104
rect 4456 7044 4460 7100
rect 4460 7044 4516 7100
rect 4516 7044 4520 7100
rect 4456 7040 4520 7044
rect 12216 7100 12280 7104
rect 12216 7044 12220 7100
rect 12220 7044 12276 7100
rect 12276 7044 12280 7100
rect 12216 7040 12280 7044
rect 12296 7100 12360 7104
rect 12296 7044 12300 7100
rect 12300 7044 12356 7100
rect 12356 7044 12360 7100
rect 12296 7040 12360 7044
rect 12376 7100 12440 7104
rect 12376 7044 12380 7100
rect 12380 7044 12436 7100
rect 12436 7044 12440 7100
rect 12376 7040 12440 7044
rect 12456 7100 12520 7104
rect 12456 7044 12460 7100
rect 12460 7044 12516 7100
rect 12516 7044 12520 7100
rect 12456 7040 12520 7044
rect 8216 6556 8280 6560
rect 8216 6500 8220 6556
rect 8220 6500 8276 6556
rect 8276 6500 8280 6556
rect 8216 6496 8280 6500
rect 8296 6556 8360 6560
rect 8296 6500 8300 6556
rect 8300 6500 8356 6556
rect 8356 6500 8360 6556
rect 8296 6496 8360 6500
rect 8376 6556 8440 6560
rect 8376 6500 8380 6556
rect 8380 6500 8436 6556
rect 8436 6500 8440 6556
rect 8376 6496 8440 6500
rect 8456 6556 8520 6560
rect 8456 6500 8460 6556
rect 8460 6500 8516 6556
rect 8516 6500 8520 6556
rect 8456 6496 8520 6500
rect 4216 6012 4280 6016
rect 4216 5956 4220 6012
rect 4220 5956 4276 6012
rect 4276 5956 4280 6012
rect 4216 5952 4280 5956
rect 4296 6012 4360 6016
rect 4296 5956 4300 6012
rect 4300 5956 4356 6012
rect 4356 5956 4360 6012
rect 4296 5952 4360 5956
rect 4376 6012 4440 6016
rect 4376 5956 4380 6012
rect 4380 5956 4436 6012
rect 4436 5956 4440 6012
rect 4376 5952 4440 5956
rect 4456 6012 4520 6016
rect 4456 5956 4460 6012
rect 4460 5956 4516 6012
rect 4516 5956 4520 6012
rect 4456 5952 4520 5956
rect 12216 6012 12280 6016
rect 12216 5956 12220 6012
rect 12220 5956 12276 6012
rect 12276 5956 12280 6012
rect 12216 5952 12280 5956
rect 12296 6012 12360 6016
rect 12296 5956 12300 6012
rect 12300 5956 12356 6012
rect 12356 5956 12360 6012
rect 12296 5952 12360 5956
rect 12376 6012 12440 6016
rect 12376 5956 12380 6012
rect 12380 5956 12436 6012
rect 12436 5956 12440 6012
rect 12376 5952 12440 5956
rect 12456 6012 12520 6016
rect 12456 5956 12460 6012
rect 12460 5956 12516 6012
rect 12516 5956 12520 6012
rect 12456 5952 12520 5956
rect 8216 5468 8280 5472
rect 8216 5412 8220 5468
rect 8220 5412 8276 5468
rect 8276 5412 8280 5468
rect 8216 5408 8280 5412
rect 8296 5468 8360 5472
rect 8296 5412 8300 5468
rect 8300 5412 8356 5468
rect 8356 5412 8360 5468
rect 8296 5408 8360 5412
rect 8376 5468 8440 5472
rect 8376 5412 8380 5468
rect 8380 5412 8436 5468
rect 8436 5412 8440 5468
rect 8376 5408 8440 5412
rect 8456 5468 8520 5472
rect 8456 5412 8460 5468
rect 8460 5412 8516 5468
rect 8516 5412 8520 5468
rect 8456 5408 8520 5412
rect 4216 4924 4280 4928
rect 4216 4868 4220 4924
rect 4220 4868 4276 4924
rect 4276 4868 4280 4924
rect 4216 4864 4280 4868
rect 4296 4924 4360 4928
rect 4296 4868 4300 4924
rect 4300 4868 4356 4924
rect 4356 4868 4360 4924
rect 4296 4864 4360 4868
rect 4376 4924 4440 4928
rect 4376 4868 4380 4924
rect 4380 4868 4436 4924
rect 4436 4868 4440 4924
rect 4376 4864 4440 4868
rect 4456 4924 4520 4928
rect 4456 4868 4460 4924
rect 4460 4868 4516 4924
rect 4516 4868 4520 4924
rect 4456 4864 4520 4868
rect 12216 4924 12280 4928
rect 12216 4868 12220 4924
rect 12220 4868 12276 4924
rect 12276 4868 12280 4924
rect 12216 4864 12280 4868
rect 12296 4924 12360 4928
rect 12296 4868 12300 4924
rect 12300 4868 12356 4924
rect 12356 4868 12360 4924
rect 12296 4864 12360 4868
rect 12376 4924 12440 4928
rect 12376 4868 12380 4924
rect 12380 4868 12436 4924
rect 12436 4868 12440 4924
rect 12376 4864 12440 4868
rect 12456 4924 12520 4928
rect 12456 4868 12460 4924
rect 12460 4868 12516 4924
rect 12516 4868 12520 4924
rect 12456 4864 12520 4868
rect 8216 4380 8280 4384
rect 8216 4324 8220 4380
rect 8220 4324 8276 4380
rect 8276 4324 8280 4380
rect 8216 4320 8280 4324
rect 8296 4380 8360 4384
rect 8296 4324 8300 4380
rect 8300 4324 8356 4380
rect 8356 4324 8360 4380
rect 8296 4320 8360 4324
rect 8376 4380 8440 4384
rect 8376 4324 8380 4380
rect 8380 4324 8436 4380
rect 8436 4324 8440 4380
rect 8376 4320 8440 4324
rect 8456 4380 8520 4384
rect 8456 4324 8460 4380
rect 8460 4324 8516 4380
rect 8516 4324 8520 4380
rect 8456 4320 8520 4324
rect 4216 3836 4280 3840
rect 4216 3780 4220 3836
rect 4220 3780 4276 3836
rect 4276 3780 4280 3836
rect 4216 3776 4280 3780
rect 4296 3836 4360 3840
rect 4296 3780 4300 3836
rect 4300 3780 4356 3836
rect 4356 3780 4360 3836
rect 4296 3776 4360 3780
rect 4376 3836 4440 3840
rect 4376 3780 4380 3836
rect 4380 3780 4436 3836
rect 4436 3780 4440 3836
rect 4376 3776 4440 3780
rect 4456 3836 4520 3840
rect 4456 3780 4460 3836
rect 4460 3780 4516 3836
rect 4516 3780 4520 3836
rect 4456 3776 4520 3780
rect 12216 3836 12280 3840
rect 12216 3780 12220 3836
rect 12220 3780 12276 3836
rect 12276 3780 12280 3836
rect 12216 3776 12280 3780
rect 12296 3836 12360 3840
rect 12296 3780 12300 3836
rect 12300 3780 12356 3836
rect 12356 3780 12360 3836
rect 12296 3776 12360 3780
rect 12376 3836 12440 3840
rect 12376 3780 12380 3836
rect 12380 3780 12436 3836
rect 12436 3780 12440 3836
rect 12376 3776 12440 3780
rect 12456 3836 12520 3840
rect 12456 3780 12460 3836
rect 12460 3780 12516 3836
rect 12516 3780 12520 3836
rect 12456 3776 12520 3780
rect 8216 3292 8280 3296
rect 8216 3236 8220 3292
rect 8220 3236 8276 3292
rect 8276 3236 8280 3292
rect 8216 3232 8280 3236
rect 8296 3292 8360 3296
rect 8296 3236 8300 3292
rect 8300 3236 8356 3292
rect 8356 3236 8360 3292
rect 8296 3232 8360 3236
rect 8376 3292 8440 3296
rect 8376 3236 8380 3292
rect 8380 3236 8436 3292
rect 8436 3236 8440 3292
rect 8376 3232 8440 3236
rect 8456 3292 8520 3296
rect 8456 3236 8460 3292
rect 8460 3236 8516 3292
rect 8516 3236 8520 3292
rect 8456 3232 8520 3236
rect 4216 2748 4280 2752
rect 4216 2692 4220 2748
rect 4220 2692 4276 2748
rect 4276 2692 4280 2748
rect 4216 2688 4280 2692
rect 4296 2748 4360 2752
rect 4296 2692 4300 2748
rect 4300 2692 4356 2748
rect 4356 2692 4360 2748
rect 4296 2688 4360 2692
rect 4376 2748 4440 2752
rect 4376 2692 4380 2748
rect 4380 2692 4436 2748
rect 4436 2692 4440 2748
rect 4376 2688 4440 2692
rect 4456 2748 4520 2752
rect 4456 2692 4460 2748
rect 4460 2692 4516 2748
rect 4516 2692 4520 2748
rect 4456 2688 4520 2692
rect 12216 2748 12280 2752
rect 12216 2692 12220 2748
rect 12220 2692 12276 2748
rect 12276 2692 12280 2748
rect 12216 2688 12280 2692
rect 12296 2748 12360 2752
rect 12296 2692 12300 2748
rect 12300 2692 12356 2748
rect 12356 2692 12360 2748
rect 12296 2688 12360 2692
rect 12376 2748 12440 2752
rect 12376 2692 12380 2748
rect 12380 2692 12436 2748
rect 12436 2692 12440 2748
rect 12376 2688 12440 2692
rect 12456 2748 12520 2752
rect 12456 2692 12460 2748
rect 12460 2692 12516 2748
rect 12516 2692 12520 2748
rect 12456 2688 12520 2692
rect 8216 2204 8280 2208
rect 8216 2148 8220 2204
rect 8220 2148 8276 2204
rect 8276 2148 8280 2204
rect 8216 2144 8280 2148
rect 8296 2204 8360 2208
rect 8296 2148 8300 2204
rect 8300 2148 8356 2204
rect 8356 2148 8360 2204
rect 8296 2144 8360 2148
rect 8376 2204 8440 2208
rect 8376 2148 8380 2204
rect 8380 2148 8436 2204
rect 8436 2148 8440 2204
rect 8376 2144 8440 2148
rect 8456 2204 8520 2208
rect 8456 2148 8460 2204
rect 8460 2148 8516 2204
rect 8516 2148 8520 2204
rect 8456 2144 8520 2148
rect 4216 1660 4280 1664
rect 4216 1604 4220 1660
rect 4220 1604 4276 1660
rect 4276 1604 4280 1660
rect 4216 1600 4280 1604
rect 4296 1660 4360 1664
rect 4296 1604 4300 1660
rect 4300 1604 4356 1660
rect 4356 1604 4360 1660
rect 4296 1600 4360 1604
rect 4376 1660 4440 1664
rect 4376 1604 4380 1660
rect 4380 1604 4436 1660
rect 4436 1604 4440 1660
rect 4376 1600 4440 1604
rect 4456 1660 4520 1664
rect 4456 1604 4460 1660
rect 4460 1604 4516 1660
rect 4516 1604 4520 1660
rect 4456 1600 4520 1604
rect 12216 1660 12280 1664
rect 12216 1604 12220 1660
rect 12220 1604 12276 1660
rect 12276 1604 12280 1660
rect 12216 1600 12280 1604
rect 12296 1660 12360 1664
rect 12296 1604 12300 1660
rect 12300 1604 12356 1660
rect 12356 1604 12360 1660
rect 12296 1600 12360 1604
rect 12376 1660 12440 1664
rect 12376 1604 12380 1660
rect 12380 1604 12436 1660
rect 12436 1604 12440 1660
rect 12376 1600 12440 1604
rect 12456 1660 12520 1664
rect 12456 1604 12460 1660
rect 12460 1604 12516 1660
rect 12516 1604 12520 1660
rect 12456 1600 12520 1604
rect 8216 1116 8280 1120
rect 8216 1060 8220 1116
rect 8220 1060 8276 1116
rect 8276 1060 8280 1116
rect 8216 1056 8280 1060
rect 8296 1116 8360 1120
rect 8296 1060 8300 1116
rect 8300 1060 8356 1116
rect 8356 1060 8360 1116
rect 8296 1056 8360 1060
rect 8376 1116 8440 1120
rect 8376 1060 8380 1116
rect 8380 1060 8436 1116
rect 8436 1060 8440 1116
rect 8376 1056 8440 1060
rect 8456 1116 8520 1120
rect 8456 1060 8460 1116
rect 8460 1060 8516 1116
rect 8516 1060 8520 1116
rect 8456 1056 8520 1060
<< metal4 >>
rect 4208 13632 4528 13648
rect 4208 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4528 13632
rect 4208 12544 4528 13568
rect 6315 13564 6381 13565
rect 6315 13500 6316 13564
rect 6380 13500 6381 13564
rect 6315 13499 6381 13500
rect 4208 12480 4216 12544
rect 4280 12488 4296 12544
rect 4360 12488 4376 12544
rect 4440 12488 4456 12544
rect 4520 12480 4528 12544
rect 4208 12252 4250 12480
rect 4486 12252 4528 12480
rect 4208 11456 4528 12252
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 4208 10368 4528 11392
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 4208 9280 4528 10304
rect 6318 10165 6378 13499
rect 8208 13088 8528 13648
rect 12208 13632 12528 13648
rect 12208 13568 12216 13632
rect 12280 13568 12296 13632
rect 12360 13568 12376 13632
rect 12440 13568 12456 13632
rect 12520 13568 12528 13632
rect 9443 13292 9509 13293
rect 9443 13228 9444 13292
rect 9508 13228 9509 13292
rect 9443 13227 9509 13228
rect 8208 13024 8216 13088
rect 8280 13024 8296 13088
rect 8360 13024 8376 13088
rect 8440 13024 8456 13088
rect 8520 13024 8528 13088
rect 8208 12000 8528 13024
rect 8707 12884 8773 12885
rect 8707 12820 8708 12884
rect 8772 12820 8773 12884
rect 8707 12819 8773 12820
rect 8208 11936 8216 12000
rect 8280 11936 8296 12000
rect 8360 11936 8376 12000
rect 8440 11936 8456 12000
rect 8520 11936 8528 12000
rect 7971 11252 8037 11253
rect 7971 11188 7972 11252
rect 8036 11188 8037 11252
rect 7971 11187 8037 11188
rect 6315 10164 6381 10165
rect 6315 10100 6316 10164
rect 6380 10100 6381 10164
rect 6315 10099 6381 10100
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 8192 4528 9216
rect 7974 8941 8034 11187
rect 8208 10912 8528 11936
rect 8208 10848 8216 10912
rect 8280 10848 8296 10912
rect 8360 10848 8376 10912
rect 8440 10848 8456 10912
rect 8520 10848 8528 10912
rect 8208 9824 8528 10848
rect 8710 10845 8770 12819
rect 9075 11388 9141 11389
rect 9075 11324 9076 11388
rect 9140 11324 9141 11388
rect 9075 11323 9141 11324
rect 9259 11388 9325 11389
rect 9259 11324 9260 11388
rect 9324 11324 9325 11388
rect 9259 11323 9325 11324
rect 8707 10844 8773 10845
rect 8707 10780 8708 10844
rect 8772 10780 8773 10844
rect 8707 10779 8773 10780
rect 8208 9760 8216 9824
rect 8280 9760 8296 9824
rect 8360 9760 8376 9824
rect 8440 9760 8456 9824
rect 8520 9760 8528 9824
rect 7971 8940 8037 8941
rect 7971 8876 7972 8940
rect 8036 8876 8037 8940
rect 7971 8875 8037 8876
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 7104 4528 8128
rect 7974 7853 8034 8875
rect 8208 8736 8528 9760
rect 8208 8672 8216 8736
rect 8280 8672 8296 8736
rect 8360 8672 8376 8736
rect 8440 8672 8456 8736
rect 8520 8672 8528 8736
rect 8208 8488 8528 8672
rect 9078 8533 9138 11323
rect 9262 10709 9322 11323
rect 9259 10708 9325 10709
rect 9259 10644 9260 10708
rect 9324 10644 9325 10708
rect 9259 10643 9325 10644
rect 9446 10573 9506 13227
rect 12208 12544 12528 13568
rect 12208 12480 12216 12544
rect 12280 12488 12296 12544
rect 12360 12488 12376 12544
rect 12440 12488 12456 12544
rect 12520 12480 12528 12544
rect 12208 12252 12250 12480
rect 12486 12252 12528 12480
rect 10179 11932 10245 11933
rect 10179 11868 10180 11932
rect 10244 11868 10245 11932
rect 10179 11867 10245 11868
rect 9995 11252 10061 11253
rect 9995 11188 9996 11252
rect 10060 11188 10061 11252
rect 9995 11187 10061 11188
rect 9443 10572 9509 10573
rect 9443 10508 9444 10572
rect 9508 10508 9509 10572
rect 9443 10507 9509 10508
rect 9998 10029 10058 11187
rect 10182 10301 10242 11867
rect 12208 11456 12528 12252
rect 12208 11392 12216 11456
rect 12280 11392 12296 11456
rect 12360 11392 12376 11456
rect 12440 11392 12456 11456
rect 12520 11392 12528 11456
rect 12208 10368 12528 11392
rect 12208 10304 12216 10368
rect 12280 10304 12296 10368
rect 12360 10304 12376 10368
rect 12440 10304 12456 10368
rect 12520 10304 12528 10368
rect 10179 10300 10245 10301
rect 10179 10236 10180 10300
rect 10244 10236 10245 10300
rect 10179 10235 10245 10236
rect 9995 10028 10061 10029
rect 9995 9964 9996 10028
rect 10060 9964 10061 10028
rect 9995 9963 10061 9964
rect 10182 9757 10242 10235
rect 10179 9756 10245 9757
rect 10179 9692 10180 9756
rect 10244 9692 10245 9756
rect 10179 9691 10245 9692
rect 12208 9280 12528 10304
rect 12208 9216 12216 9280
rect 12280 9216 12296 9280
rect 12360 9216 12376 9280
rect 12440 9216 12456 9280
rect 12520 9216 12528 9280
rect 8208 8252 8250 8488
rect 8486 8252 8528 8488
rect 9075 8532 9141 8533
rect 9075 8468 9076 8532
rect 9140 8468 9141 8532
rect 9075 8467 9141 8468
rect 7971 7852 8037 7853
rect 7971 7788 7972 7852
rect 8036 7788 8037 7852
rect 7971 7787 8037 7788
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 6016 4528 7040
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 4928 4528 5952
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 4488 4528 4864
rect 4208 4252 4250 4488
rect 4486 4252 4528 4488
rect 4208 3840 4528 4252
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 2752 4528 3776
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 1664 4528 2688
rect 4208 1600 4216 1664
rect 4280 1600 4296 1664
rect 4360 1600 4376 1664
rect 4440 1600 4456 1664
rect 4520 1600 4528 1664
rect 4208 1040 4528 1600
rect 8208 7648 8528 8252
rect 8208 7584 8216 7648
rect 8280 7584 8296 7648
rect 8360 7584 8376 7648
rect 8440 7584 8456 7648
rect 8520 7584 8528 7648
rect 8208 6560 8528 7584
rect 8208 6496 8216 6560
rect 8280 6496 8296 6560
rect 8360 6496 8376 6560
rect 8440 6496 8456 6560
rect 8520 6496 8528 6560
rect 8208 5472 8528 6496
rect 8208 5408 8216 5472
rect 8280 5408 8296 5472
rect 8360 5408 8376 5472
rect 8440 5408 8456 5472
rect 8520 5408 8528 5472
rect 8208 4384 8528 5408
rect 8208 4320 8216 4384
rect 8280 4320 8296 4384
rect 8360 4320 8376 4384
rect 8440 4320 8456 4384
rect 8520 4320 8528 4384
rect 8208 3296 8528 4320
rect 8208 3232 8216 3296
rect 8280 3232 8296 3296
rect 8360 3232 8376 3296
rect 8440 3232 8456 3296
rect 8520 3232 8528 3296
rect 8208 2208 8528 3232
rect 8208 2144 8216 2208
rect 8280 2144 8296 2208
rect 8360 2144 8376 2208
rect 8440 2144 8456 2208
rect 8520 2144 8528 2208
rect 8208 1120 8528 2144
rect 8208 1056 8216 1120
rect 8280 1056 8296 1120
rect 8360 1056 8376 1120
rect 8440 1056 8456 1120
rect 8520 1056 8528 1120
rect 8208 1040 8528 1056
rect 12208 8192 12528 9216
rect 12208 8128 12216 8192
rect 12280 8128 12296 8192
rect 12360 8128 12376 8192
rect 12440 8128 12456 8192
rect 12520 8128 12528 8192
rect 12208 7104 12528 8128
rect 12208 7040 12216 7104
rect 12280 7040 12296 7104
rect 12360 7040 12376 7104
rect 12440 7040 12456 7104
rect 12520 7040 12528 7104
rect 12208 6016 12528 7040
rect 12208 5952 12216 6016
rect 12280 5952 12296 6016
rect 12360 5952 12376 6016
rect 12440 5952 12456 6016
rect 12520 5952 12528 6016
rect 12208 4928 12528 5952
rect 12208 4864 12216 4928
rect 12280 4864 12296 4928
rect 12360 4864 12376 4928
rect 12440 4864 12456 4928
rect 12520 4864 12528 4928
rect 12208 4488 12528 4864
rect 12208 4252 12250 4488
rect 12486 4252 12528 4488
rect 12208 3840 12528 4252
rect 12208 3776 12216 3840
rect 12280 3776 12296 3840
rect 12360 3776 12376 3840
rect 12440 3776 12456 3840
rect 12520 3776 12528 3840
rect 12208 2752 12528 3776
rect 12208 2688 12216 2752
rect 12280 2688 12296 2752
rect 12360 2688 12376 2752
rect 12440 2688 12456 2752
rect 12520 2688 12528 2752
rect 12208 1664 12528 2688
rect 12208 1600 12216 1664
rect 12280 1600 12296 1664
rect 12360 1600 12376 1664
rect 12440 1600 12456 1664
rect 12520 1600 12528 1664
rect 12208 1040 12528 1600
<< via4 >>
rect 4250 12480 4280 12488
rect 4280 12480 4296 12488
rect 4296 12480 4360 12488
rect 4360 12480 4376 12488
rect 4376 12480 4440 12488
rect 4440 12480 4456 12488
rect 4456 12480 4486 12488
rect 4250 12252 4486 12480
rect 12250 12480 12280 12488
rect 12280 12480 12296 12488
rect 12296 12480 12360 12488
rect 12360 12480 12376 12488
rect 12376 12480 12440 12488
rect 12440 12480 12456 12488
rect 12456 12480 12486 12488
rect 12250 12252 12486 12480
rect 8250 8252 8486 8488
rect 4250 4252 4486 4488
rect 12250 4252 12486 4488
<< metal5 >>
rect 1056 12488 13940 12530
rect 1056 12252 4250 12488
rect 4486 12252 12250 12488
rect 12486 12252 13940 12488
rect 1056 12210 13940 12252
rect 1056 8488 13940 8530
rect 1056 8252 8250 8488
rect 8486 8252 13940 8488
rect 1056 8210 13940 8252
rect 1056 4488 13940 4530
rect 1056 4252 4250 4488
rect 4486 4252 12250 4488
rect 12486 4252 13940 4488
rect 1056 4210 13940 4252
use sky130_fd_sc_hd__diode_2  ANTENNA__243__A $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform -1 0 6992 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__244__A
timestamp 1665323087
transform -1 0 8372 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__252__A
timestamp 1665323087
transform -1 0 5336 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__257__A_N
timestamp 1665323087
transform -1 0 9568 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__258__A
timestamp 1665323087
transform -1 0 6256 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__260__A1
timestamp 1665323087
transform -1 0 1564 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__266__A
timestamp 1665323087
transform -1 0 5060 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__267__A1
timestamp 1665323087
transform 1 0 6348 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__270__A1
timestamp 1665323087
transform -1 0 3956 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__287__B1
timestamp 1665323087
transform -1 0 7820 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__289__A1
timestamp 1665323087
transform 1 0 5428 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__348__A
timestamp 1665323087
transform -1 0 8648 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__349__A
timestamp 1665323087
transform -1 0 1564 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__350__A
timestamp 1665323087
transform -1 0 4048 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__358__A
timestamp 1665323087
transform 1 0 6072 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__360__A2
timestamp 1665323087
transform -1 0 4968 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__361__B
timestamp 1665323087
transform 1 0 7176 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__363__A2
timestamp 1665323087
transform 1 0 7636 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__364__A2
timestamp 1665323087
transform -1 0 8464 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__369__A2
timestamp 1665323087
transform -1 0 8188 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__373__A2
timestamp 1665323087
transform -1 0 9200 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__374__B1
timestamp 1665323087
transform 1 0 5428 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__375__A2
timestamp 1665323087
transform -1 0 8832 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__378__A2
timestamp 1665323087
transform -1 0 3680 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__379__A
timestamp 1665323087
transform 1 0 6348 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__380__A2
timestamp 1665323087
transform 1 0 3496 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__383__A2
timestamp 1665323087
transform -1 0 8832 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__384__A_N
timestamp 1665323087
transform -1 0 2208 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__387__B1
timestamp 1665323087
transform 1 0 5152 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__389__A2
timestamp 1665323087
transform -1 0 3956 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__392__A2
timestamp 1665323087
transform -1 0 6256 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__396__A2
timestamp 1665323087
transform -1 0 4324 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__399__A2
timestamp 1665323087
transform -1 0 13616 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__404__A2
timestamp 1665323087
transform -1 0 3680 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__409__B1
timestamp 1665323087
transform -1 0 13616 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__410__A2
timestamp 1665323087
transform -1 0 10856 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__411__A2
timestamp 1665323087
transform -1 0 5520 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__417__B1
timestamp 1665323087
transform 1 0 7728 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__419__A2
timestamp 1665323087
transform -1 0 13616 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__421__B1
timestamp 1665323087
transform -1 0 13616 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__422__A2
timestamp 1665323087
transform -1 0 11684 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__423__A2
timestamp 1665323087
transform -1 0 13616 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__424__A2
timestamp 1665323087
transform 1 0 13432 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__425__A
timestamp 1665323087
transform -1 0 11684 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__425__B
timestamp 1665323087
transform -1 0 6256 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__447__A
timestamp 1665323087
transform -1 0 3956 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__470__D
timestamp 1665323087
transform -1 0 9108 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform 1 0 4324 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_83
timestamp 1665323087
transform 1 0 8740 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_111
timestamp 1665323087
transform 1 0 11316 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_115 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform 1 0 11684 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_135
timestamp 1665323087
transform 1 0 13524 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_3
timestamp 1665323087
transform 1 0 1380 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_111
timestamp 1665323087
transform 1 0 11316 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_134 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform 1 0 13432 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_2_76
timestamp 1665323087
transform 1 0 8096 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_2_108
timestamp 1665323087
transform 1 0 11040 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_3_3
timestamp 1665323087
transform 1 0 1380 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_134
timestamp 1665323087
transform 1 0 13432 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_4_12
timestamp 1665323087
transform 1 0 2208 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_29
timestamp 1665323087
transform 1 0 3772 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_55
timestamp 1665323087
transform 1 0 6164 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_92
timestamp 1665323087
transform 1 0 9568 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_134
timestamp 1665323087
transform 1 0 13432 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_5_101
timestamp 1665323087
transform 1 0 10396 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_5_135
timestamp 1665323087
transform 1 0 13524 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_3
timestamp 1665323087
transform 1 0 1380 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_85
timestamp 1665323087
transform 1 0 8924 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_90
timestamp 1665323087
transform 1 0 9384 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_7_3
timestamp 1665323087
transform 1 0 1380 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_21
timestamp 1665323087
transform 1 0 3036 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_64
timestamp 1665323087
transform 1 0 6992 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_71
timestamp 1665323087
transform 1 0 7636 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_97
timestamp 1665323087
transform 1 0 10028 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_105
timestamp 1665323087
transform 1 0 10764 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_8_41
timestamp 1665323087
transform 1 0 4876 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_8_83
timestamp 1665323087
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_89
timestamp 1665323087
transform 1 0 9292 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_9_45
timestamp 1665323087
transform 1 0 5244 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_88
timestamp 1665323087
transform 1 0 9200 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_9_102
timestamp 1665323087
transform 1 0 10488 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_27
timestamp 1665323087
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_126
timestamp 1665323087
transform 1 0 12696 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_11_3
timestamp 1665323087
transform 1 0 1380 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_11_102
timestamp 1665323087
transform 1 0 10488 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_37
timestamp 1665323087
transform 1 0 4508 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_69
timestamp 1665323087
transform 1 0 7452 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_83
timestamp 1665323087
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_85
timestamp 1665323087
transform 1 0 8924 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_116
timestamp 1665323087
transform 1 0 11776 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_122
timestamp 1665323087
transform 1 0 12328 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_23
timestamp 1665323087
transform 1 0 3220 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_90
timestamp 1665323087
transform 1 0 9384 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_15_122
timestamp 1665323087
transform 1 0 12328 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_39
timestamp 1665323087
transform 1 0 4692 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_85
timestamp 1665323087
transform 1 0 8924 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_17_28
timestamp 1665323087
transform 1 0 3680 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_17_87
timestamp 1665323087
transform 1 0 9108 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_17_96
timestamp 1665323087
transform 1 0 9936 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_18_65
timestamp 1665323087
transform 1 0 7084 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_18_95
timestamp 1665323087
transform 1 0 9844 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_19_48
timestamp 1665323087
transform 1 0 5520 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_19_57
timestamp 1665323087
transform 1 0 6348 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_19_123
timestamp 1665323087
transform 1 0 12420 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_19_135
timestamp 1665323087
transform 1 0 13524 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_20_64
timestamp 1665323087
transform 1 0 6992 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_20_85
timestamp 1665323087
transform 1 0 8924 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_21_3
timestamp 1665323087
transform 1 0 1380 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_21_55
timestamp 1665323087
transform 1 0 6164 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_21_68
timestamp 1665323087
transform 1 0 7360 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_21_135
timestamp 1665323087
transform 1 0 13524 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_22_57
timestamp 1665323087
transform 1 0 6348 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_22_65
timestamp 1665323087
transform 1 0 7084 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_22_85
timestamp 1665323087
transform 1 0 8924 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_22_111
timestamp 1665323087
transform 1 0 11316 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_22_113
timestamp 1665323087
transform 1 0 11500 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1665323087
transform 1 0 1104 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1665323087
transform -1 0 13892 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1665323087
transform 1 0 1104 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1665323087
transform -1 0 13892 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1665323087
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1665323087
transform -1 0 13892 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1665323087
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1665323087
transform -1 0 13892 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1665323087
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1665323087
transform -1 0 13892 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1665323087
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1665323087
transform -1 0 13892 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1665323087
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1665323087
transform -1 0 13892 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1665323087
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1665323087
transform -1 0 13892 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1665323087
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1665323087
transform -1 0 13892 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1665323087
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1665323087
transform -1 0 13892 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1665323087
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1665323087
transform -1 0 13892 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1665323087
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1665323087
transform -1 0 13892 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1665323087
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1665323087
transform -1 0 13892 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1665323087
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1665323087
transform -1 0 13892 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1665323087
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1665323087
transform -1 0 13892 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1665323087
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1665323087
transform -1 0 13892 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1665323087
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1665323087
transform -1 0 13892 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1665323087
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1665323087
transform -1 0 13892 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1665323087
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1665323087
transform -1 0 13892 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1665323087
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1665323087
transform -1 0 13892 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1665323087
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1665323087
transform -1 0 13892 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1665323087
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1665323087
transform -1 0 13892 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1665323087
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1665323087
transform -1 0 13892 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_46 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform 1 0 3680 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_47
timestamp 1665323087
transform 1 0 6256 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_48
timestamp 1665323087
transform 1 0 8832 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_49
timestamp 1665323087
transform 1 0 11408 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_50
timestamp 1665323087
transform 1 0 6256 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_51
timestamp 1665323087
transform 1 0 11408 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_52
timestamp 1665323087
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_53
timestamp 1665323087
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_54
timestamp 1665323087
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_55
timestamp 1665323087
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_56
timestamp 1665323087
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_57
timestamp 1665323087
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_58
timestamp 1665323087
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_59
timestamp 1665323087
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_60
timestamp 1665323087
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_61
timestamp 1665323087
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_62
timestamp 1665323087
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_63
timestamp 1665323087
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_64
timestamp 1665323087
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_65
timestamp 1665323087
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_66
timestamp 1665323087
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_67
timestamp 1665323087
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_68
timestamp 1665323087
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_69
timestamp 1665323087
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_70
timestamp 1665323087
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_71
timestamp 1665323087
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_72
timestamp 1665323087
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_73
timestamp 1665323087
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_74
timestamp 1665323087
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_75
timestamp 1665323087
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_76
timestamp 1665323087
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_77
timestamp 1665323087
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_78
timestamp 1665323087
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_79
timestamp 1665323087
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_80
timestamp 1665323087
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_81
timestamp 1665323087
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_82
timestamp 1665323087
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_83
timestamp 1665323087
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_84
timestamp 1665323087
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_85
timestamp 1665323087
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_86
timestamp 1665323087
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_87
timestamp 1665323087
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_88
timestamp 1665323087
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_89
timestamp 1665323087
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_90
timestamp 1665323087
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_91
timestamp 1665323087
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_92
timestamp 1665323087
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_93
timestamp 1665323087
transform 1 0 6256 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_94
timestamp 1665323087
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_95
timestamp 1665323087
transform 1 0 11408 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__xnor2_2  _214_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform 1 0 11316 0 1 2176
box -38 -48 1234 592
use sky130_fd_sc_hd__buf_2  _215_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform 1 0 13156 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _216_
timestamp 1665323087
transform -1 0 11316 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_2  _217_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform 1 0 4416 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _218_
timestamp 1665323087
transform -1 0 3496 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_2  _219_
timestamp 1665323087
transform 1 0 3956 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _220_
timestamp 1665323087
transform -1 0 2208 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_2  _221_
timestamp 1665323087
transform 1 0 2208 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _222_
timestamp 1665323087
transform -1 0 1840 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_2  _223_
timestamp 1665323087
transform 1 0 4324 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _224_
timestamp 1665323087
transform -1 0 1748 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _225_
timestamp 1665323087
transform -1 0 1748 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_2  _226_
timestamp 1665323087
transform 1 0 3772 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _227_
timestamp 1665323087
transform -1 0 2024 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _228_
timestamp 1665323087
transform 1 0 8464 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _229_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform -1 0 7636 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _230_
timestamp 1665323087
transform 1 0 3404 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__nand2b_2  _231_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform -1 0 4416 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__and2_2  _232_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform -1 0 4324 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_2  _233_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform -1 0 5060 0 1 3264
box -38 -48 1234 592
use sky130_fd_sc_hd__and2_2  _234_
timestamp 1665323087
transform 1 0 2484 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__and2_2  _235_
timestamp 1665323087
transform -1 0 4140 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__a211o_2  _236_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform 1 0 3036 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_2  _237_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform -1 0 4876 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _238_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform 1 0 5428 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_2  _239_
timestamp 1665323087
transform 1 0 4416 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__and3_2  _240_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform -1 0 3220 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_2  _241_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform -1 0 3588 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_2  _242_
timestamp 1665323087
transform -1 0 2944 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _243_
timestamp 1665323087
transform 1 0 1380 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _244_
timestamp 1665323087
transform -1 0 2392 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_2  _245_
timestamp 1665323087
transform 1 0 3036 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_2  _246_
timestamp 1665323087
transform -1 0 2484 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _247_
timestamp 1665323087
transform 1 0 2576 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_2  _248_
timestamp 1665323087
transform -1 0 2576 0 -1 6528
box -38 -48 1234 592
use sky130_fd_sc_hd__o32a_2  _249_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform 1 0 1656 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_2  _250_
timestamp 1665323087
transform -1 0 1932 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_2  _251_
timestamp 1665323087
transform -1 0 3496 0 1 3264
box -38 -48 1234 592
use sky130_fd_sc_hd__inv_2  _252_
timestamp 1665323087
transform 1 0 5980 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__nand2b_2  _253_
timestamp 1665323087
transform -1 0 2116 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_2  _254_
timestamp 1665323087
transform -1 0 1932 0 -1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _255_
timestamp 1665323087
transform -1 0 6072 0 1 1088
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _256_
timestamp 1665323087
transform 1 0 10212 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__nand3b_2  _257_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform -1 0 2576 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__and2_2  _258_
timestamp 1665323087
transform -1 0 3128 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_2  _259_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform 1 0 1564 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__o2111a_2  _260_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform 1 0 1380 0 1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__xor2_2  _261_
timestamp 1665323087
transform -1 0 5796 0 1 7616
box -38 -48 1234 592
use sky130_fd_sc_hd__inv_2  _262_
timestamp 1665323087
transform 1 0 5980 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__and2_2  _263_
timestamp 1665323087
transform -1 0 4968 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_2  _264_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform 1 0 3772 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_2  _265_
timestamp 1665323087
transform 1 0 3220 0 -1 7616
box -38 -48 1234 592
use sky130_fd_sc_hd__and2_2  _266_
timestamp 1665323087
transform -1 0 4692 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_2  _267_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform 1 0 2760 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_2  _268_
timestamp 1665323087
transform 1 0 4968 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _269_
timestamp 1665323087
transform -1 0 5152 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_2  _270_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform -1 0 4508 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__o31a_2  _271_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform 1 0 1932 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _272_
timestamp 1665323087
transform -1 0 9384 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _273_
timestamp 1665323087
transform -1 0 6716 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__and2_2  _274_
timestamp 1665323087
transform 1 0 11776 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _275_
timestamp 1665323087
transform 1 0 12144 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _276_
timestamp 1665323087
transform 1 0 13340 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _277_
timestamp 1665323087
transform 1 0 8832 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__nand4_2  _278_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform 1 0 9384 0 1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__nand2_2  _279_
timestamp 1665323087
transform 1 0 10580 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _280_
timestamp 1665323087
transform 1 0 10212 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _281_
timestamp 1665323087
transform 1 0 8924 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _282_
timestamp 1665323087
transform 1 0 8372 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _283_
timestamp 1665323087
transform -1 0 10948 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _284_
timestamp 1665323087
transform 1 0 10948 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__and3_2  _285_
timestamp 1665323087
transform 1 0 9936 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__and4b_2  _286_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform -1 0 13340 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__o21ai_2  _287_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform -1 0 3220 0 1 2176
box -38 -48 682 592
use sky130_fd_sc_hd__and4b_2  _288_
timestamp 1665323087
transform 1 0 1748 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__o211a_2  _289_
timestamp 1665323087
transform 1 0 2024 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__nand4b_2  _290_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform -1 0 3404 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__and3b_2  _291_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform 1 0 10304 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__o31a_2  _292_
timestamp 1665323087
transform -1 0 10856 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _293_
timestamp 1665323087
transform -1 0 10764 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_2  _294_
timestamp 1665323087
transform 1 0 5612 0 1 6528
box -38 -48 1234 592
use sky130_fd_sc_hd__nor2_2  _295_
timestamp 1665323087
transform 1 0 6532 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and2_2  _296_
timestamp 1665323087
transform -1 0 6624 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_2  _297_
timestamp 1665323087
transform 1 0 7636 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _298_
timestamp 1665323087
transform 1 0 11040 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _299_
timestamp 1665323087
transform 1 0 11592 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_2  _300_
timestamp 1665323087
transform -1 0 11408 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _301_
timestamp 1665323087
transform 1 0 9752 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_2  _302_
timestamp 1665323087
transform 1 0 8464 0 -1 7616
box -38 -48 1234 592
use sky130_fd_sc_hd__inv_2  _303_
timestamp 1665323087
transform -1 0 9660 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_2  _304_
timestamp 1665323087
transform -1 0 9936 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__a32o_2  _305_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform -1 0 10488 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _306_
timestamp 1665323087
transform -1 0 8372 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_2  _307_
timestamp 1665323087
transform 1 0 6624 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__xnor2_2  _308_
timestamp 1665323087
transform -1 0 8004 0 1 6528
box -38 -48 1234 592
use sky130_fd_sc_hd__and2_2  _309_
timestamp 1665323087
transform 1 0 7084 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_2  _310_
timestamp 1665323087
transform 1 0 6532 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_2  _311_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform -1 0 8372 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_2  _312_
timestamp 1665323087
transform -1 0 7636 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_2  _313_
timestamp 1665323087
transform 1 0 6716 0 -1 7616
box -38 -48 1234 592
use sky130_fd_sc_hd__mux2_2  _314_
timestamp 1665323087
transform -1 0 8004 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _315_
timestamp 1665323087
transform 1 0 8924 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__xor2_2  _316_
timestamp 1665323087
transform 1 0 7544 0 1 7616
box -38 -48 1234 592
use sky130_fd_sc_hd__mux2_2  _317_
timestamp 1665323087
transform 1 0 8188 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _318_
timestamp 1665323087
transform 1 0 8372 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_2  _319_
timestamp 1665323087
transform -1 0 11408 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__o211a_2  _320_
timestamp 1665323087
transform 1 0 11040 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_2  _321_
timestamp 1665323087
transform -1 0 12696 0 -1 7616
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_2  _322_
timestamp 1665323087
transform 1 0 8924 0 1 6528
box -38 -48 1234 592
use sky130_fd_sc_hd__o2bb2a_2  _323_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform 1 0 9660 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_2  _324_
timestamp 1665323087
transform 1 0 11868 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_2  _325_
timestamp 1665323087
transform -1 0 12696 0 1 6528
box -38 -48 1234 592
use sky130_fd_sc_hd__mux2_2  _326_
timestamp 1665323087
transform 1 0 10580 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _327_
timestamp 1665323087
transform -1 0 9844 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_2  _328_
timestamp 1665323087
transform 1 0 11500 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_2  _329_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform -1 0 11500 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__and3_2  _330_
timestamp 1665323087
transform 1 0 6348 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__and2_2  _331_
timestamp 1665323087
transform 1 0 5060 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_2  _332_
timestamp 1665323087
transform 1 0 5612 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__nand2b_2  _333_
timestamp 1665323087
transform -1 0 5980 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_2  _334_
timestamp 1665323087
transform 1 0 4968 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_2  _335_
timestamp 1665323087
transform 1 0 5336 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_2  _336_
timestamp 1665323087
transform 1 0 6348 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_2  _337_
timestamp 1665323087
transform 1 0 5520 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__and2_2  _338_
timestamp 1665323087
transform 1 0 6348 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _339_
timestamp 1665323087
transform 1 0 11500 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_2  _340_
timestamp 1665323087
transform 1 0 4416 0 1 1088
box -38 -48 1234 592
use sky130_fd_sc_hd__a21boi_2  _341_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform -1 0 7176 0 -1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__nand3_2  _342_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform 1 0 4968 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_2  _343_
timestamp 1665323087
transform -1 0 12788 0 1 1088
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _344_
timestamp 1665323087
transform 1 0 12788 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_2  _345_
timestamp 1665323087
transform -1 0 12788 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _346_
timestamp 1665323087
transform 1 0 12788 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__nand2b_2  _347_
timestamp 1665323087
transform -1 0 8832 0 1 2176
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _348_
timestamp 1665323087
transform 1 0 1656 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _349_
timestamp 1665323087
transform 1 0 4048 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_2  _350_
timestamp 1665323087
transform -1 0 4232 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_2  _351_
timestamp 1665323087
transform -1 0 4876 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _352_
timestamp 1665323087
transform -1 0 5152 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_2  _353_
timestamp 1665323087
transform -1 0 7176 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__and2b_2  _354_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform -1 0 7636 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__and3_2  _355_
timestamp 1665323087
transform 1 0 8280 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_2  _356_
timestamp 1665323087
transform 1 0 9384 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _357_
timestamp 1665323087
transform -1 0 7452 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _358_
timestamp 1665323087
transform 1 0 5796 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and2_2  _359_
timestamp 1665323087
transform -1 0 8004 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_2  _360_
timestamp 1665323087
transform 1 0 3772 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_2  _361_
timestamp 1665323087
transform -1 0 8280 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _362_
timestamp 1665323087
transform -1 0 10672 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__a211o_2  _363_
timestamp 1665323087
transform 1 0 9016 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_2  _364_
timestamp 1665323087
transform 1 0 5520 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _365_
timestamp 1665323087
transform -1 0 8832 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__and2_2  _366_
timestamp 1665323087
transform -1 0 10120 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_2  _367_
timestamp 1665323087
transform -1 0 9108 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_2  _368_
timestamp 1665323087
transform 1 0 7912 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_2  _369_
timestamp 1665323087
transform -1 0 2024 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_2  _370_
timestamp 1665323087
transform 1 0 13156 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _371_
timestamp 1665323087
transform -1 0 9384 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_2  _372_
timestamp 1665323087
transform 1 0 7820 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_2  _373_
timestamp 1665323087
transform 1 0 1380 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_2  _374_
timestamp 1665323087
transform -1 0 6992 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_2  _375_
timestamp 1665323087
transform 1 0 2208 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_2  _376_
timestamp 1665323087
transform 1 0 7452 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_2  _377_
timestamp 1665323087
transform 1 0 5612 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_2  _378_
timestamp 1665323087
transform -1 0 3864 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _379_
timestamp 1665323087
transform -1 0 8464 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_2  _380_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform -1 0 7820 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _381_
timestamp 1665323087
transform 1 0 11960 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_2  _382_
timestamp 1665323087
transform -1 0 7912 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _383_
timestamp 1665323087
transform 1 0 8832 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__nand2b_2  _384_
timestamp 1665323087
transform 1 0 4048 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__o31a_2  _385_
timestamp 1665323087
transform -1 0 10212 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_2  _386_
timestamp 1665323087
transform -1 0 6900 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_2  _387_
timestamp 1665323087
transform -1 0 7728 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__o21a_2  _388_
timestamp 1665323087
transform 1 0 6348 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_2  _389_
timestamp 1665323087
transform -1 0 6256 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _390_
timestamp 1665323087
transform 1 0 5888 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_2  _391_
timestamp 1665323087
transform 1 0 5612 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_2  _392_
timestamp 1665323087
transform 1 0 5704 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_2  _393_
timestamp 1665323087
transform 1 0 7636 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_2  _394_
timestamp 1665323087
transform 1 0 8372 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_2  _395_
timestamp 1665323087
transform 1 0 7360 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _396_
timestamp 1665323087
transform -1 0 8556 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_2  _397_
timestamp 1665323087
transform -1 0 11040 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__and2_2  _398_
timestamp 1665323087
transform 1 0 9016 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_2  _399_
timestamp 1665323087
transform 1 0 9292 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__nand2b_2  _400_
timestamp 1665323087
transform 1 0 10672 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_2  _401_
timestamp 1665323087
transform 1 0 10120 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__o22a_2  _402_
timestamp 1665323087
transform -1 0 10672 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__and3_2  _403_
timestamp 1665323087
transform 1 0 10212 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_2  _404_
timestamp 1665323087
transform 1 0 10304 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__nand3_2  _405_
timestamp 1665323087
transform -1 0 12052 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__nand3b_2  _406_
timestamp 1665323087
transform -1 0 11316 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__and3_2  _407_
timestamp 1665323087
transform 1 0 10028 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_2  _408_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform 1 0 10580 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__a32o_2  _409_
timestamp 1665323087
transform 1 0 11500 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_2  _410_
timestamp 1665323087
transform 1 0 9568 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_2  _411_
timestamp 1665323087
transform -1 0 8740 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__o22a_2  _412_
timestamp 1665323087
transform 1 0 9200 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_2  _413_
timestamp 1665323087
transform -1 0 8648 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__o2111a_2  _414_
timestamp 1665323087
transform 1 0 7912 0 -1 11968
box -38 -48 958 592
use sky130_fd_sc_hd__o21ai_2  _415_
timestamp 1665323087
transform 1 0 6716 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_2  _416_
timestamp 1665323087
transform -1 0 6716 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_2  _417_
timestamp 1665323087
transform 1 0 6256 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__o31a_2  _418_
timestamp 1665323087
transform -1 0 11592 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_2  _419_
timestamp 1665323087
transform 1 0 11316 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__nand3_2  _420_
timestamp 1665323087
transform 1 0 12052 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__a32o_2  _421_
timestamp 1665323087
transform -1 0 13156 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_2  _422_
timestamp 1665323087
transform -1 0 12328 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_2  _423_
timestamp 1665323087
transform 1 0 12236 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _424_
timestamp 1665323087
transform 1 0 11500 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_2  _425_
timestamp 1665323087
transform -1 0 3680 0 1 1088
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _426_
timestamp 1665323087
transform 1 0 4600 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_2  _427_
timestamp 1665323087
transform -1 0 11960 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _428_
timestamp 1665323087
transform 1 0 12512 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _429_
timestamp 1665323087
transform -1 0 10028 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_2  _430_
timestamp 1665323087
transform 1 0 10488 0 -1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _431_
timestamp 1665323087
transform -1 0 7636 0 -1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _432_
timestamp 1665323087
transform -1 0 6808 0 1 1088
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _433_
timestamp 1665323087
transform -1 0 8096 0 1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _434_
timestamp 1665323087
transform 1 0 10028 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_2  _435_
timestamp 1665323087
transform -1 0 7360 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _436_
timestamp 1665323087
transform -1 0 7360 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _437_
timestamp 1665323087
transform 1 0 10948 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _438_
timestamp 1665323087
transform -1 0 7728 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_2  _439_
timestamp 1665323087
transform 1 0 11500 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _440_
timestamp 1665323087
transform 1 0 10488 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _441_
timestamp 1665323087
transform 1 0 11592 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _442_
timestamp 1665323087
transform -1 0 9384 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _443_
timestamp 1665323087
transform -1 0 10028 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_2  _444_
timestamp 1665323087
transform -1 0 8280 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _445_
timestamp 1665323087
transform 1 0 8372 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _446_
timestamp 1665323087
transform -1 0 7820 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _447_
timestamp 1665323087
transform -1 0 3680 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_2  _448_
timestamp 1665323087
transform -1 0 9384 0 1 1088
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _449_
timestamp 1665323087
transform 1 0 9752 0 -1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _450_
timestamp 1665323087
transform -1 0 2392 0 -1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _451_
timestamp 1665323087
transform 1 0 3220 0 1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _452_
timestamp 1665323087
transform -1 0 3588 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _453_
timestamp 1665323087
transform 1 0 3956 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _454_
timestamp 1665323087
transform 1 0 5060 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__dfrtp_2  _455_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform 1 0 9108 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _456_
timestamp 1665323087
transform 1 0 9476 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _457_
timestamp 1665323087
transform 1 0 11500 0 -1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _458_
timestamp 1665323087
transform 1 0 5704 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _459_
timestamp 1665323087
transform -1 0 6256 0 -1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _460_
timestamp 1665323087
transform -1 0 8188 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _461_
timestamp 1665323087
transform 1 0 5704 0 1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _462_
timestamp 1665323087
transform 1 0 4968 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _463_
timestamp 1665323087
transform 1 0 11500 0 -1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _464_
timestamp 1665323087
transform 1 0 9844 0 1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _465_
timestamp 1665323087
transform 1 0 9568 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _466_
timestamp 1665323087
transform 1 0 9660 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _467_
timestamp 1665323087
transform 1 0 7728 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _468_
timestamp 1665323087
transform -1 0 8832 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _469_
timestamp 1665323087
transform 1 0 7728 0 -1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _470_
timestamp 1665323087
transform -1 0 8740 0 1 1088
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _471_
timestamp 1665323087
transform 1 0 7820 0 -1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _472_
timestamp 1665323087
transform 1 0 9384 0 1 1088
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _473_
timestamp 1665323087
transform 1 0 2392 0 -1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _474_
timestamp 1665323087
transform 1 0 2392 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _475_
timestamp 1665323087
transform 1 0 1472 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _476_
timestamp 1665323087
transform 1 0 3496 0 -1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _477_
timestamp 1665323087
transform 1 0 4140 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__clkbuf_16  clockp_buffer_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform -1 0 3220 0 1 1088
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clockp_buffer_1
timestamp 1665323087
transform 1 0 1380 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[0\].id.delaybuf0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform -1 0 6716 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[0\].id.delaybuf1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform 1 0 5796 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[0\].id.delayen0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform 1 0 4784 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[0\].id.delayen1
timestamp 1665323087
transform 1 0 5152 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__einvn_8  ringosc.dstage\[0\].id.delayenb0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform 1 0 4416 0 -1 9792
box -38 -48 1694 592
use sky130_fd_sc_hd__einvn_4  ringosc.dstage\[0\].id.delayenb1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform 1 0 5060 0 1 8704
box -38 -48 1050 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[0\].id.delayint0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform -1 0 5704 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[1\].id.delaybuf0
timestamp 1665323087
transform -1 0 5520 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[1\].id.delaybuf1
timestamp 1665323087
transform -1 0 4048 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[1\].id.delayen0
timestamp 1665323087
transform 1 0 3864 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[1\].id.delayen1
timestamp 1665323087
transform -1 0 5152 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__einvn_8  ringosc.dstage\[1\].id.delayenb0
timestamp 1665323087
transform 1 0 3956 0 1 10880
box -38 -48 1694 592
use sky130_fd_sc_hd__einvn_4  ringosc.dstage\[1\].id.delayenb1
timestamp 1665323087
transform 1 0 4416 0 -1 10880
box -38 -48 1050 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[1\].id.delayint0
timestamp 1665323087
transform 1 0 4968 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[2\].id.delaybuf0
timestamp 1665323087
transform 1 0 5244 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[2\].id.delaybuf1
timestamp 1665323087
transform 1 0 11040 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[2\].id.delayen0
timestamp 1665323087
transform 1 0 9292 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[2\].id.delayen1
timestamp 1665323087
transform 1 0 9936 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__einvn_8  ringosc.dstage\[2\].id.delayenb0
timestamp 1665323087
transform 1 0 8740 0 -1 13056
box -38 -48 1694 592
use sky130_fd_sc_hd__einvn_4  ringosc.dstage\[2\].id.delayenb1
timestamp 1665323087
transform 1 0 10396 0 -1 13056
box -38 -48 1050 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[2\].id.delayint0
timestamp 1665323087
transform -1 0 10304 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[3\].id.delaybuf0
timestamp 1665323087
transform -1 0 7544 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[3\].id.delaybuf1
timestamp 1665323087
transform 1 0 7544 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[3\].id.delayen0
timestamp 1665323087
transform 1 0 5612 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[3\].id.delayen1
timestamp 1665323087
transform 1 0 6440 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__einvn_8  ringosc.dstage\[3\].id.delayenb0
timestamp 1665323087
transform 1 0 5336 0 1 11968
box -38 -48 1694 592
use sky130_fd_sc_hd__einvn_4  ringosc.dstage\[3\].id.delayenb1
timestamp 1665323087
transform 1 0 6348 0 -1 13056
box -38 -48 1050 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[3\].id.delayint0
timestamp 1665323087
transform 1 0 8556 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[4\].id.delaybuf0
timestamp 1665323087
transform -1 0 3220 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[4\].id.delaybuf1
timestamp 1665323087
transform -1 0 2852 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[4\].id.delayen0
timestamp 1665323087
transform 1 0 2024 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[4\].id.delayen1
timestamp 1665323087
transform -1 0 4140 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__einvn_8  ringosc.dstage\[4\].id.delayenb0
timestamp 1665323087
transform 1 0 2024 0 1 9792
box -38 -48 1694 592
use sky130_fd_sc_hd__einvn_4  ringosc.dstage\[4\].id.delayenb1
timestamp 1665323087
transform -1 0 3864 0 -1 9792
box -38 -48 1050 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[4\].id.delayint0
timestamp 1665323087
transform -1 0 1656 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[5\].id.delaybuf0
timestamp 1665323087
transform 1 0 1380 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[5\].id.delaybuf1
timestamp 1665323087
transform -1 0 3036 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[5\].id.delayen0
timestamp 1665323087
transform 1 0 1564 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[5\].id.delayen1
timestamp 1665323087
transform -1 0 3680 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__einvn_8  ringosc.dstage\[5\].id.delayenb0
timestamp 1665323087
transform 1 0 1380 0 1 10880
box -38 -48 1694 592
use sky130_fd_sc_hd__einvn_4  ringosc.dstage\[5\].id.delayenb1
timestamp 1665323087
transform -1 0 3680 0 -1 10880
box -38 -48 1050 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[5\].id.delayint0
timestamp 1665323087
transform -1 0 1656 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[6\].id.delaybuf0
timestamp 1665323087
transform 1 0 1472 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[6\].id.delaybuf1
timestamp 1665323087
transform 1 0 8004 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[6\].id.delayen0
timestamp 1665323087
transform 1 0 2208 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[6\].id.delayen1
timestamp 1665323087
transform 1 0 2852 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__einvn_8  ringosc.dstage\[6\].id.delayenb0
timestamp 1665323087
transform 1 0 1840 0 -1 13056
box -38 -48 1694 592
use sky130_fd_sc_hd__einvn_4  ringosc.dstage\[6\].id.delayenb1
timestamp 1665323087
transform -1 0 2760 0 1 11968
box -38 -48 1050 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[6\].id.delayint0
timestamp 1665323087
transform 1 0 7912 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[7\].id.delaybuf0
timestamp 1665323087
transform 1 0 3772 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[7\].id.delaybuf1
timestamp 1665323087
transform -1 0 1656 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[7\].id.delayen0
timestamp 1665323087
transform 1 0 4324 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[7\].id.delayen1
timestamp 1665323087
transform -1 0 3680 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__einvn_8  ringosc.dstage\[7\].id.delayenb0
timestamp 1665323087
transform 1 0 3680 0 -1 13056
box -38 -48 1694 592
use sky130_fd_sc_hd__einvn_4  ringosc.dstage\[7\].id.delayenb1
timestamp 1665323087
transform -1 0 4784 0 1 11968
box -38 -48 1050 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[7\].id.delayint0
timestamp 1665323087
transform -1 0 3680 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[8\].id.delaybuf0
timestamp 1665323087
transform 1 0 12236 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[8\].id.delaybuf1
timestamp 1665323087
transform 1 0 12604 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[8\].id.delayen0
timestamp 1665323087
transform 1 0 11592 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[8\].id.delayen1
timestamp 1665323087
transform 1 0 11500 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__einvn_8  ringosc.dstage\[8\].id.delayenb0
timestamp 1665323087
transform 1 0 11500 0 -1 13056
box -38 -48 1694 592
use sky130_fd_sc_hd__einvn_4  ringosc.dstage\[8\].id.delayenb1
timestamp 1665323087
transform 1 0 10948 0 1 11968
box -38 -48 1050 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[8\].id.delayint0
timestamp 1665323087
transform -1 0 9292 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[9\].id.delaybuf0
timestamp 1665323087
transform -1 0 13524 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[9\].id.delaybuf1
timestamp 1665323087
transform -1 0 13156 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[9\].id.delayen0
timestamp 1665323087
transform -1 0 11408 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[9\].id.delayen1
timestamp 1665323087
transform 1 0 12512 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__einvn_8  ringosc.dstage\[9\].id.delayenb0
timestamp 1665323087
transform 1 0 11960 0 1 11968
box -38 -48 1694 592
use sky130_fd_sc_hd__einvn_4  ringosc.dstage\[9\].id.delayenb1
timestamp 1665323087
transform 1 0 12328 0 1 10880
box -38 -48 1050 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[9\].id.delayint0
timestamp 1665323087
transform -1 0 9292 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[10\].id.delaybuf0
timestamp 1665323087
transform 1 0 13156 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[10\].id.delaybuf1
timestamp 1665323087
transform -1 0 13432 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[10\].id.delayen0
timestamp 1665323087
transform 1 0 12972 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[10\].id.delayen1
timestamp 1665323087
transform 1 0 12788 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__einvn_8  ringosc.dstage\[10\].id.delayenb0
timestamp 1665323087
transform 1 0 11960 0 1 8704
box -38 -48 1694 592
use sky130_fd_sc_hd__einvn_4  ringosc.dstage\[10\].id.delayenb1
timestamp 1665323087
transform 1 0 12420 0 -1 9792
box -38 -48 1050 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[10\].id.delayint0
timestamp 1665323087
transform 1 0 13340 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[11\].id.delaybuf0
timestamp 1665323087
transform -1 0 13524 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[11\].id.delaybuf1
timestamp 1665323087
transform 1 0 13340 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[11\].id.delayen0
timestamp 1665323087
transform 1 0 12788 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[11\].id.delayen1
timestamp 1665323087
transform 1 0 12696 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__einvn_8  ringosc.dstage\[11\].id.delayenb0
timestamp 1665323087
transform 1 0 11960 0 -1 6528
box -38 -48 1694 592
use sky130_fd_sc_hd__einvn_4  ringosc.dstage\[11\].id.delayenb1
timestamp 1665323087
transform 1 0 12420 0 1 7616
box -38 -48 1050 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[11\].id.delayint0
timestamp 1665323087
transform -1 0 8464 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  ringosc.ibufp00 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform -1 0 9384 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_8  ringosc.ibufp01 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform -1 0 9476 0 -1 3264
box -38 -48 1234 592
use sky130_fd_sc_hd__clkinv_2  ringosc.ibufp10
timestamp 1665323087
transform 1 0 1656 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_8  ringosc.ibufp11
timestamp 1665323087
transform 1 0 1380 0 -1 9792
box -38 -48 1234 592
use sky130_fd_sc_hd__conb_1  ringosc.iss.const1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform 1 0 13340 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__or2_2  ringosc.iss.ctrlen0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform 1 0 12052 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.iss.delaybuf0
timestamp 1665323087
transform 1 0 13156 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_2  ringosc.iss.delayen0
timestamp 1665323087
transform -1 0 12512 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__einvp_2  ringosc.iss.delayen1
timestamp 1665323087
transform 1 0 12512 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__einvn_8  ringosc.iss.delayenb0
timestamp 1665323087
transform 1 0 11960 0 1 4352
box -38 -48 1694 592
use sky130_fd_sc_hd__einvn_4  ringosc.iss.delayenb1
timestamp 1665323087
transform 1 0 12328 0 1 5440
box -38 -48 1050 592
use sky130_fd_sc_hd__clkinv_1  ringosc.iss.delayint0
timestamp 1665323087
transform -1 0 10396 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_1  ringosc.iss.reseten0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform 1 0 12972 0 1 3264
box -38 -48 498 592
<< labels >>
flabel metal4 s 8208 1040 8528 13648 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal5 s 1056 8210 13940 8530 0 FreeSans 2560 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 4208 1040 4528 13648 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 12208 1040 12528 13648 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal5 s 1056 4210 13940 4530 0 FreeSans 2560 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal5 s 1056 12210 13940 12530 0 FreeSans 2560 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal3 s 0 416 800 536 0 FreeSans 480 0 0 0 clockp[0]
port 2 nsew signal tristate
flabel metal3 s 0 1232 800 1352 0 FreeSans 480 0 0 0 clockp[1]
port 3 nsew signal tristate
flabel metal3 s 0 7896 800 8016 0 FreeSans 480 0 0 0 dco
port 4 nsew signal input
flabel metal3 s 0 2184 800 2304 0 FreeSans 480 0 0 0 div[0]
port 5 nsew signal input
flabel metal3 s 0 3136 800 3256 0 FreeSans 480 0 0 0 div[1]
port 6 nsew signal input
flabel metal3 s 0 4088 800 4208 0 FreeSans 480 0 0 0 div[2]
port 7 nsew signal input
flabel metal3 s 0 5040 800 5160 0 FreeSans 480 0 0 0 div[3]
port 8 nsew signal input
flabel metal3 s 0 5992 800 6112 0 FreeSans 480 0 0 0 div[4]
port 9 nsew signal input
flabel metal3 s 0 6944 800 7064 0 FreeSans 480 0 0 0 enable
port 10 nsew signal input
flabel metal3 s 0 8712 800 8832 0 FreeSans 480 0 0 0 ext_trim[0]
port 11 nsew signal input
flabel metal2 s 3974 14200 4030 15000 0 FreeSans 224 90 0 0 ext_trim[10]
port 12 nsew signal input
flabel metal2 s 5170 14200 5226 15000 0 FreeSans 224 90 0 0 ext_trim[11]
port 13 nsew signal input
flabel metal2 s 6274 14200 6330 15000 0 FreeSans 224 90 0 0 ext_trim[12]
port 14 nsew signal input
flabel metal2 s 7470 14200 7526 15000 0 FreeSans 224 90 0 0 ext_trim[13]
port 15 nsew signal input
flabel metal2 s 8574 14200 8630 15000 0 FreeSans 224 90 0 0 ext_trim[14]
port 16 nsew signal input
flabel metal2 s 9770 14200 9826 15000 0 FreeSans 224 90 0 0 ext_trim[15]
port 17 nsew signal input
flabel metal2 s 10874 14200 10930 15000 0 FreeSans 224 90 0 0 ext_trim[16]
port 18 nsew signal input
flabel metal2 s 12070 14200 12126 15000 0 FreeSans 224 90 0 0 ext_trim[17]
port 19 nsew signal input
flabel metal2 s 13174 14200 13230 15000 0 FreeSans 224 90 0 0 ext_trim[18]
port 20 nsew signal input
flabel metal2 s 14370 14200 14426 15000 0 FreeSans 224 90 0 0 ext_trim[19]
port 21 nsew signal input
flabel metal3 s 0 9664 800 9784 0 FreeSans 480 0 0 0 ext_trim[1]
port 22 nsew signal input
flabel metal3 s 14200 13608 15000 13728 0 FreeSans 480 0 0 0 ext_trim[20]
port 23 nsew signal input
flabel metal3 s 14200 11160 15000 11280 0 FreeSans 480 0 0 0 ext_trim[21]
port 24 nsew signal input
flabel metal3 s 14200 8712 15000 8832 0 FreeSans 480 0 0 0 ext_trim[22]
port 25 nsew signal input
flabel metal3 s 14200 6128 15000 6248 0 FreeSans 480 0 0 0 ext_trim[23]
port 26 nsew signal input
flabel metal3 s 14200 3680 15000 3800 0 FreeSans 480 0 0 0 ext_trim[24]
port 27 nsew signal input
flabel metal3 s 14200 1232 15000 1352 0 FreeSans 480 0 0 0 ext_trim[25]
port 28 nsew signal input
flabel metal3 s 0 10616 800 10736 0 FreeSans 480 0 0 0 ext_trim[2]
port 29 nsew signal input
flabel metal3 s 0 11568 800 11688 0 FreeSans 480 0 0 0 ext_trim[3]
port 30 nsew signal input
flabel metal3 s 0 12520 800 12640 0 FreeSans 480 0 0 0 ext_trim[4]
port 31 nsew signal input
flabel metal3 s 0 13472 800 13592 0 FreeSans 480 0 0 0 ext_trim[5]
port 32 nsew signal input
flabel metal3 s 0 14424 800 14544 0 FreeSans 480 0 0 0 ext_trim[6]
port 33 nsew signal input
flabel metal2 s 570 14200 626 15000 0 FreeSans 224 90 0 0 ext_trim[7]
port 34 nsew signal input
flabel metal2 s 1674 14200 1730 15000 0 FreeSans 224 90 0 0 ext_trim[8]
port 35 nsew signal input
flabel metal2 s 2870 14200 2926 15000 0 FreeSans 224 90 0 0 ext_trim[9]
port 36 nsew signal input
flabel metal2 s 11150 0 11206 800 0 FreeSans 224 90 0 0 osc
port 37 nsew signal input
flabel metal2 s 3698 0 3754 800 0 FreeSans 224 90 0 0 resetb
port 38 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 15000 15000
<< end >>
