magic
tech sky130A
magscale 1 2
timestamp 1636983106
<< locali >>
rect 8769 13175 8803 13277
rect 14933 12223 14967 14977
rect 14933 9027 14967 10557
rect 15025 9571 15059 10965
rect 14933 8483 14967 8993
rect 14933 7531 14967 8449
rect 15025 7871 15059 8993
rect 14933 5627 14967 6613
rect 15025 6443 15059 7837
rect 15117 8007 15151 10081
rect 15117 7327 15151 7973
rect 15209 7395 15243 10829
rect 15301 8959 15335 11781
rect 15209 6375 15243 7361
rect 15393 7259 15427 11169
rect 3065 3587 3099 3689
rect 14933 1071 14967 3417
rect 15025 2635 15059 6273
<< viali >>
rect 14933 14977 14967 15011
rect 2881 13481 2915 13515
rect 4537 13481 4571 13515
rect 7573 13481 7607 13515
rect 8953 13481 8987 13515
rect 14289 13481 14323 13515
rect 3985 13413 4019 13447
rect 5181 13413 5215 13447
rect 8309 13413 8343 13447
rect 3801 13345 3835 13379
rect 5733 13345 5767 13379
rect 9505 13345 9539 13379
rect 12081 13345 12115 13379
rect 2789 13277 2823 13311
rect 3065 13277 3099 13311
rect 4077 13277 4111 13311
rect 4353 13287 4387 13321
rect 4445 13287 4479 13321
rect 4629 13277 4663 13311
rect 7481 13277 7515 13311
rect 8217 13277 8251 13311
rect 8493 13277 8527 13311
rect 8769 13277 8803 13311
rect 9137 13277 9171 13311
rect 9413 13277 9447 13311
rect 9873 13277 9907 13311
rect 11805 13277 11839 13311
rect 12449 13277 12483 13311
rect 14105 13277 14139 13311
rect 11621 13209 11655 13243
rect 2697 13141 2731 13175
rect 3801 13141 3835 13175
rect 4261 13141 4295 13175
rect 4721 13141 4755 13175
rect 5549 13141 5583 13175
rect 5641 13141 5675 13175
rect 7941 13141 7975 13175
rect 8677 13141 8711 13175
rect 8769 13141 8803 13175
rect 11299 13141 11333 13175
rect 11989 13141 12023 13175
rect 13875 13141 13909 13175
rect 5457 12937 5491 12971
rect 5825 12937 5859 12971
rect 6377 12937 6411 12971
rect 13323 12937 13357 12971
rect 14197 12937 14231 12971
rect 5089 12869 5123 12903
rect 8769 12869 8803 12903
rect 10701 12869 10735 12903
rect 2513 12801 2547 12835
rect 2881 12801 2915 12835
rect 4629 12801 4663 12835
rect 4813 12801 4847 12835
rect 5365 12801 5399 12835
rect 6745 12801 6779 12835
rect 7021 12801 7055 12835
rect 7288 12801 7322 12835
rect 11161 12801 11195 12835
rect 11529 12801 11563 12835
rect 13829 12801 13863 12835
rect 14105 12801 14139 12835
rect 14289 12801 14323 12835
rect 5917 12733 5951 12767
rect 6009 12733 6043 12767
rect 6653 12733 6687 12767
rect 8493 12733 8527 12767
rect 10517 12733 10551 12767
rect 11897 12733 11931 12767
rect 13737 12733 13771 12767
rect 4307 12665 4341 12699
rect 13461 12665 13495 12699
rect 8401 12597 8435 12631
rect 10885 12597 10919 12631
rect 10977 12597 11011 12631
rect 11253 12597 11287 12631
rect 7573 12393 7607 12427
rect 8033 12393 8067 12427
rect 8309 12393 8343 12427
rect 11621 12393 11655 12427
rect 14289 12393 14323 12427
rect 4077 12325 4111 12359
rect 3525 12257 3559 12291
rect 4813 12257 4847 12291
rect 5089 12257 5123 12291
rect 5733 12257 5767 12291
rect 10149 12257 10183 12291
rect 13921 12257 13955 12291
rect 1777 12189 1811 12223
rect 3985 12189 4019 12223
rect 4077 12189 4111 12223
rect 4261 12189 4295 12223
rect 4353 12189 4387 12223
rect 4721 12189 4755 12223
rect 6193 12189 6227 12223
rect 7757 12189 7791 12223
rect 8309 12189 8343 12223
rect 8585 12189 8619 12223
rect 9873 12189 9907 12223
rect 14197 12189 14231 12223
rect 14473 12189 14507 12223
rect 14933 12189 14967 12223
rect 2053 12121 2087 12155
rect 3801 12121 3835 12155
rect 6460 12121 6494 12155
rect 8401 12121 8435 12155
rect 11897 12121 11931 12155
rect 13645 12121 13679 12155
rect 5181 12053 5215 12087
rect 5549 12053 5583 12087
rect 5641 12053 5675 12087
rect 8217 12053 8251 12087
rect 8769 12053 8803 12087
rect 9321 12053 9355 12087
rect 9689 12053 9723 12087
rect 11713 12053 11747 12087
rect 3249 11849 3283 11883
rect 3801 11849 3835 11883
rect 4997 11849 5031 11883
rect 5457 11849 5491 11883
rect 8309 11849 8343 11883
rect 10149 11849 10183 11883
rect 10333 11849 10367 11883
rect 10977 11849 11011 11883
rect 11345 11849 11379 11883
rect 14289 11849 14323 11883
rect 5825 11781 5859 11815
rect 9413 11781 9447 11815
rect 10241 11781 10275 11815
rect 11621 11781 11655 11815
rect 12817 11781 12851 11815
rect 15301 11781 15335 11815
rect 3525 11713 3559 11747
rect 3801 11713 3835 11747
rect 3985 11713 4019 11747
rect 4537 11713 4571 11747
rect 4629 11713 4663 11747
rect 4813 11713 4847 11747
rect 4905 11713 4939 11747
rect 5089 11713 5123 11747
rect 6377 11713 6411 11747
rect 6633 11713 6667 11747
rect 8033 11713 8067 11747
rect 8585 11713 8619 11747
rect 9045 11713 9079 11747
rect 9321 11713 9355 11747
rect 9505 11713 9539 11747
rect 9597 11713 9631 11747
rect 9965 11713 9999 11747
rect 10057 11713 10091 11747
rect 11069 11713 11103 11747
rect 11253 11713 11287 11747
rect 11345 11713 11379 11747
rect 12081 11713 12115 11747
rect 3249 11645 3283 11679
rect 5917 11645 5951 11679
rect 6009 11645 6043 11679
rect 7849 11645 7883 11679
rect 8309 11645 8343 11679
rect 8769 11645 8803 11679
rect 10701 11645 10735 11679
rect 10793 11645 10827 11679
rect 12173 11645 12207 11679
rect 12265 11645 12299 11679
rect 12541 11645 12575 11679
rect 3433 11577 3467 11611
rect 7757 11577 7791 11611
rect 8217 11577 8251 11611
rect 8493 11577 8527 11611
rect 9229 11577 9263 11611
rect 3617 11509 3651 11543
rect 4077 11509 4111 11543
rect 4445 11509 4479 11543
rect 4721 11509 4755 11543
rect 8861 11509 8895 11543
rect 9689 11509 9723 11543
rect 11713 11509 11747 11543
rect 3617 11305 3651 11339
rect 3985 11305 4019 11339
rect 4399 11305 4433 11339
rect 8723 11305 8757 11339
rect 9505 11305 9539 11339
rect 11161 11305 11195 11339
rect 14197 11305 14231 11339
rect 3893 11237 3927 11271
rect 6009 11237 6043 11271
rect 6377 11237 6411 11271
rect 11069 11237 11103 11271
rect 2145 11169 2179 11203
rect 3801 11169 3835 11203
rect 5733 11169 5767 11203
rect 6929 11169 6963 11203
rect 7297 11169 7331 11203
rect 10609 11169 10643 11203
rect 11713 11169 11747 11203
rect 12449 11169 12483 11203
rect 1869 11101 1903 11135
rect 4077 11101 4111 11135
rect 4169 11101 4203 11135
rect 6193 11101 6227 11135
rect 6837 11101 6871 11135
rect 9141 11101 9175 11135
rect 9229 11079 9263 11113
rect 9321 11101 9355 11135
rect 9781 11101 9815 11135
rect 9965 11101 9999 11135
rect 10425 11101 10459 11135
rect 10701 11101 10735 11135
rect 11529 11101 11563 11135
rect 12081 11101 12115 11135
rect 14105 11101 14139 11135
rect 5457 11033 5491 11067
rect 5549 11033 5583 11067
rect 6285 11033 6319 11067
rect 6469 11033 6503 11067
rect 10149 11033 10183 11067
rect 10333 11033 10367 11067
rect 5089 10965 5123 10999
rect 6745 10965 6779 10999
rect 8953 10965 8987 10999
rect 9689 10965 9723 10999
rect 10425 10965 10459 10999
rect 11621 10965 11655 10999
rect 13875 10965 13909 10999
rect 14473 10965 14507 10999
rect 15025 10965 15059 10999
rect 4261 10761 4295 10795
rect 4353 10761 4387 10795
rect 4721 10761 4755 10795
rect 5641 10761 5675 10795
rect 6009 10761 6043 10795
rect 8953 10761 8987 10795
rect 11299 10761 11333 10795
rect 3341 10693 3375 10727
rect 4813 10693 4847 10727
rect 5365 10693 5399 10727
rect 6377 10693 6411 10727
rect 9229 10693 9263 10727
rect 12357 10693 12391 10727
rect 1685 10625 1719 10659
rect 3525 10625 3559 10659
rect 3709 10625 3743 10659
rect 3801 10625 3835 10659
rect 3985 10625 4019 10659
rect 4077 10625 4111 10659
rect 4261 10625 4295 10659
rect 5549 10625 5583 10659
rect 5641 10625 5675 10659
rect 5779 10625 5813 10659
rect 5917 10625 5951 10659
rect 6561 10625 6595 10659
rect 6929 10625 6963 10659
rect 8585 10625 8619 10659
rect 8953 10625 8987 10659
rect 9045 10625 9079 10659
rect 9505 10625 9539 10659
rect 11897 10625 11931 10659
rect 14105 10625 14139 10659
rect 4905 10557 4939 10591
rect 8769 10557 8803 10591
rect 9873 10557 9907 10591
rect 11989 10557 12023 10591
rect 12081 10557 12115 10591
rect 14473 10557 14507 10591
rect 14933 10557 14967 10591
rect 3157 10489 3191 10523
rect 3985 10489 4019 10523
rect 1593 10421 1627 10455
rect 3617 10421 3651 10455
rect 6193 10421 6227 10455
rect 8355 10421 8389 10455
rect 9321 10421 9355 10455
rect 11529 10421 11563 10455
rect 3157 10217 3191 10251
rect 3341 10217 3375 10251
rect 7021 10217 7055 10251
rect 10977 10217 11011 10251
rect 12173 10217 12207 10251
rect 13001 10217 13035 10251
rect 13829 10217 13863 10251
rect 4721 10149 4755 10183
rect 5181 10149 5215 10183
rect 5273 10149 5307 10183
rect 7573 10149 7607 10183
rect 9505 10149 9539 10183
rect 11069 10149 11103 10183
rect 1409 10081 1443 10115
rect 8585 10081 8619 10115
rect 9045 10081 9079 10115
rect 10333 10081 10367 10115
rect 10701 10081 10735 10115
rect 11897 10081 11931 10115
rect 12633 10081 12667 10115
rect 12817 10081 12851 10115
rect 13645 10081 13679 10115
rect 3249 10013 3283 10047
rect 3801 10013 3835 10047
rect 4169 10013 4203 10047
rect 4353 10013 4387 10047
rect 4445 10013 4479 10047
rect 4629 10013 4663 10047
rect 4997 10013 5031 10047
rect 5089 10013 5123 10047
rect 5365 10013 5399 10047
rect 5457 10013 5491 10047
rect 5733 10013 5767 10047
rect 7573 10013 7607 10047
rect 7757 10013 7791 10047
rect 8033 10013 8067 10047
rect 8677 10013 8711 10047
rect 9137 10013 9171 10047
rect 9965 10013 9999 10047
rect 10057 10013 10091 10047
rect 10793 10013 10827 10047
rect 11069 10013 11103 10047
rect 11253 10013 11287 10047
rect 12541 10013 12575 10047
rect 1685 9945 1719 9979
rect 13369 9945 13403 9979
rect 14381 9945 14415 9979
rect 3525 9877 3559 9911
rect 3893 9877 3927 9911
rect 4077 9877 4111 9911
rect 4537 9877 4571 9911
rect 5549 9877 5583 9911
rect 7941 9877 7975 9911
rect 9597 9877 9631 9911
rect 10241 9877 10275 9911
rect 11345 9877 11379 9911
rect 11713 9877 11747 9911
rect 11805 9877 11839 9911
rect 13461 9877 13495 9911
rect 14289 9877 14323 9911
rect 4997 9673 5031 9707
rect 7205 9673 7239 9707
rect 11529 9673 11563 9707
rect 11897 9673 11931 9707
rect 5825 9605 5859 9639
rect 8217 9605 8251 9639
rect 10333 9605 10367 9639
rect 10977 9605 11011 9639
rect 1409 9537 1443 9571
rect 4261 9537 4295 9571
rect 4445 9537 4479 9571
rect 4629 9537 4663 9571
rect 4721 9537 4755 9571
rect 4813 9537 4847 9571
rect 5733 9537 5767 9571
rect 6377 9537 6411 9571
rect 6653 9537 6687 9571
rect 6929 9537 6963 9571
rect 7573 9537 7607 9571
rect 8125 9537 8159 9571
rect 8493 9537 8527 9571
rect 8861 9537 8895 9571
rect 9045 9537 9079 9571
rect 9354 9537 9388 9571
rect 9965 9537 9999 9571
rect 10149 9537 10183 9571
rect 10517 9537 10551 9571
rect 11529 9537 11563 9571
rect 11621 9537 11655 9571
rect 11805 9537 11839 9571
rect 12265 9537 12299 9571
rect 12725 9537 12759 9571
rect 1777 9469 1811 9503
rect 3893 9469 3927 9503
rect 5917 9469 5951 9503
rect 7665 9469 7699 9503
rect 7849 9469 7883 9503
rect 8309 9469 8343 9503
rect 9137 9469 9171 9503
rect 10793 9469 10827 9503
rect 10885 9469 10919 9503
rect 12357 9469 12391 9503
rect 12541 9469 12575 9503
rect 3433 9401 3467 9435
rect 3617 9401 3651 9435
rect 5365 9401 5399 9435
rect 6469 9401 6503 9435
rect 7113 9401 7147 9435
rect 9045 9401 9079 9435
rect 9873 9401 9907 9435
rect 11345 9401 11379 9435
rect 3203 9333 3237 9367
rect 3985 9333 4019 9367
rect 4261 9333 4295 9367
rect 14013 9333 14047 9367
rect 2789 9129 2823 9163
rect 3249 9129 3283 9163
rect 8125 9129 8159 9163
rect 8677 9129 8711 9163
rect 9137 9129 9171 9163
rect 11713 9129 11747 9163
rect 14197 9129 14231 9163
rect 2881 9061 2915 9095
rect 3525 9061 3559 9095
rect 15209 10829 15243 10863
rect 15025 9537 15059 9571
rect 15117 10081 15151 10115
rect 2697 8963 2731 8997
rect 6377 8993 6411 9027
rect 6929 8993 6963 9027
rect 7113 8993 7147 9027
rect 7849 8993 7883 9027
rect 9597 8993 9631 9027
rect 9781 8993 9815 9027
rect 10241 8993 10275 9027
rect 13921 8993 13955 9027
rect 14933 8993 14967 9027
rect 2973 8925 3007 8959
rect 3341 8925 3375 8959
rect 3985 8925 4019 8959
rect 4077 8925 4111 8959
rect 4629 8925 4663 8959
rect 7665 8925 7699 8959
rect 8217 8925 8251 8959
rect 8585 8925 8619 8959
rect 9965 8925 9999 8959
rect 14105 8925 14139 8959
rect 4445 8857 4479 8891
rect 4905 8857 4939 8891
rect 6837 8857 6871 8891
rect 11897 8857 11931 8891
rect 13645 8857 13679 8891
rect 3801 8789 3835 8823
rect 6469 8789 6503 8823
rect 7297 8789 7331 8823
rect 7757 8789 7791 8823
rect 8953 8789 8987 8823
rect 9505 8789 9539 8823
rect 14381 8789 14415 8823
rect 2881 8585 2915 8619
rect 4813 8585 4847 8619
rect 5089 8585 5123 8619
rect 6745 8585 6779 8619
rect 7757 8585 7791 8619
rect 4353 8517 4387 8551
rect 8585 8517 8619 8551
rect 11161 8517 11195 8551
rect 11345 8517 11379 8551
rect 12081 8517 12115 8551
rect 12357 8517 12391 8551
rect 4905 8449 4939 8483
rect 5273 8449 5307 8483
rect 6101 8449 6135 8483
rect 7389 8449 7423 8483
rect 8033 8449 8067 8483
rect 8493 8449 8527 8483
rect 8769 8449 8803 8483
rect 8861 8449 8895 8483
rect 10977 8449 11011 8483
rect 11897 8449 11931 8483
rect 12449 8449 12483 8483
rect 14473 8449 14507 8483
rect 14933 8449 14967 8483
rect 4629 8381 4663 8415
rect 6837 8381 6871 8415
rect 6929 8381 6963 8415
rect 7297 8381 7331 8415
rect 7941 8381 7975 8415
rect 9229 8381 9263 8415
rect 12173 8381 12207 8415
rect 12725 8381 12759 8415
rect 14197 8381 14231 8415
rect 6377 8313 6411 8347
rect 8677 8313 8711 8347
rect 11621 8313 11655 8347
rect 5365 8245 5399 8279
rect 5733 8245 5767 8279
rect 5917 8245 5951 8279
rect 8401 8245 8435 8279
rect 10655 8245 10689 8279
rect 10793 8245 10827 8279
rect 9597 8041 9631 8075
rect 14289 8041 14323 8075
rect 11713 7973 11747 8007
rect 13921 7973 13955 8007
rect 2513 7905 2547 7939
rect 5457 7905 5491 7939
rect 5825 7905 5859 7939
rect 7251 7905 7285 7939
rect 9873 7905 9907 7939
rect 12449 7905 12483 7939
rect 2237 7837 2271 7871
rect 2697 7837 2731 7871
rect 2789 7837 2823 7871
rect 7389 7837 7423 7871
rect 7757 7837 7791 7871
rect 8217 7837 8251 7871
rect 8953 7837 8987 7871
rect 9229 7837 9263 7871
rect 9413 7837 9447 7871
rect 9505 7837 9539 7871
rect 9689 7837 9723 7871
rect 9965 7837 9999 7871
rect 10333 7837 10367 7871
rect 12173 7837 12207 7871
rect 14473 7837 14507 7871
rect 7941 7769 7975 7803
rect 9045 7769 9079 7803
rect 10600 7769 10634 7803
rect 2145 7701 2179 7735
rect 2513 7701 2547 7735
rect 3341 7701 3375 7735
rect 3985 7701 4019 7735
rect 5365 7701 5399 7735
rect 8677 7701 8711 7735
rect 10149 7701 10183 7735
rect 11897 7701 11931 7735
rect 11989 7701 12023 7735
rect 14105 7701 14139 7735
rect 7113 7497 7147 7531
rect 7665 7497 7699 7531
rect 11529 7497 11563 7531
rect 13369 7497 13403 7531
rect 13737 7497 13771 7531
rect 13829 7497 13863 7531
rect 14933 7497 14967 7531
rect 15025 8993 15059 9027
rect 15025 7837 15059 7871
rect 6837 7429 6871 7463
rect 9137 7429 9171 7463
rect 1961 7361 1995 7395
rect 2329 7361 2363 7395
rect 3755 7361 3789 7395
rect 4169 7361 4203 7395
rect 4629 7361 4663 7395
rect 4813 7361 4847 7395
rect 7113 7361 7147 7395
rect 7205 7361 7239 7395
rect 9413 7361 9447 7395
rect 9597 7361 9631 7395
rect 10149 7361 10183 7395
rect 11345 7361 11379 7395
rect 13277 7361 13311 7395
rect 14473 7361 14507 7395
rect 4077 7293 4111 7327
rect 7021 7293 7055 7327
rect 7481 7293 7515 7327
rect 10057 7293 10091 7327
rect 10701 7293 10735 7327
rect 13001 7293 13035 7327
rect 14013 7293 14047 7327
rect 14289 7225 14323 7259
rect 4445 7157 4479 7191
rect 4629 7157 4663 7191
rect 6745 7157 6779 7191
rect 7297 7157 7331 7191
rect 7389 7157 7423 7191
rect 9873 7157 9907 7191
rect 10425 7157 10459 7191
rect 10609 7157 10643 7191
rect 2145 6953 2179 6987
rect 8125 6953 8159 6987
rect 10609 6953 10643 6987
rect 7481 6885 7515 6919
rect 11069 6885 11103 6919
rect 2329 6817 2363 6851
rect 3341 6817 3375 6851
rect 3617 6817 3651 6851
rect 5641 6817 5675 6851
rect 8217 6817 8251 6851
rect 13921 6817 13955 6851
rect 2053 6749 2087 6783
rect 2237 6749 2271 6783
rect 2513 6749 2547 6783
rect 2605 6749 2639 6783
rect 2973 6749 3007 6783
rect 3249 6749 3283 6783
rect 3801 6749 3835 6783
rect 4169 6749 4203 6783
rect 4629 6749 4663 6783
rect 4721 6749 4755 6783
rect 6009 6749 6043 6783
rect 7481 6749 7515 6783
rect 7665 6749 7699 6783
rect 7941 6749 7975 6783
rect 8401 6749 8435 6783
rect 9229 6749 9263 6783
rect 11437 6749 11471 6783
rect 14473 6749 14507 6783
rect 5457 6681 5491 6715
rect 6276 6681 6310 6715
rect 8769 6681 8803 6715
rect 9496 6681 9530 6715
rect 11345 6681 11379 6715
rect 11529 6681 11563 6715
rect 11713 6681 11747 6715
rect 11897 6681 11931 6715
rect 13645 6681 13679 6715
rect 2329 6613 2363 6647
rect 2881 6613 2915 6647
rect 3893 6613 3927 6647
rect 4813 6613 4847 6647
rect 5089 6613 5123 6647
rect 5549 6613 5583 6647
rect 7389 6613 7423 6647
rect 7757 6613 7791 6647
rect 8493 6613 8527 6647
rect 9045 6613 9079 6647
rect 10885 6613 10919 6647
rect 11437 6613 11471 6647
rect 14105 6613 14139 6647
rect 14289 6613 14323 6647
rect 14933 6613 14967 6647
rect 3157 6409 3191 6443
rect 5089 6409 5123 6443
rect 6745 6409 6779 6443
rect 6837 6409 6871 6443
rect 11345 6409 11379 6443
rect 11989 6409 12023 6443
rect 14473 6409 14507 6443
rect 4537 6341 4571 6375
rect 5641 6341 5675 6375
rect 7849 6341 7883 6375
rect 13461 6341 13495 6375
rect 14289 6341 14323 6375
rect 1409 6273 1443 6307
rect 3249 6273 3283 6307
rect 3341 6273 3375 6307
rect 3525 6273 3559 6307
rect 3985 6273 4019 6307
rect 4445 6273 4479 6307
rect 4629 6273 4663 6307
rect 5549 6273 5583 6307
rect 5825 6273 5859 6307
rect 5917 6273 5951 6307
rect 7205 6273 7239 6307
rect 7389 6273 7423 6307
rect 7481 6273 7515 6307
rect 9873 6273 9907 6307
rect 10232 6273 10266 6307
rect 11713 6273 11747 6307
rect 11897 6273 11931 6307
rect 1685 6205 1719 6239
rect 4077 6205 4111 6239
rect 4261 6205 4295 6239
rect 5181 6205 5215 6239
rect 5273 6205 5307 6239
rect 6929 6205 6963 6239
rect 7573 6205 7607 6239
rect 9597 6205 9631 6239
rect 9965 6205 9999 6239
rect 13737 6205 13771 6239
rect 3617 6137 3651 6171
rect 5733 6137 5767 6171
rect 11897 6137 11931 6171
rect 14105 6137 14139 6171
rect 3433 6069 3467 6103
rect 4721 6069 4755 6103
rect 6009 6069 6043 6103
rect 6377 6069 6411 6103
rect 7481 6069 7515 6103
rect 9781 6069 9815 6103
rect 11529 6069 11563 6103
rect 13829 6069 13863 6103
rect 4813 5865 4847 5899
rect 7619 5865 7653 5899
rect 12173 5865 12207 5899
rect 3433 5797 3467 5831
rect 11989 5797 12023 5831
rect 1409 5729 1443 5763
rect 3249 5729 3283 5763
rect 4353 5729 4387 5763
rect 5457 5729 5491 5763
rect 5733 5729 5767 5763
rect 8309 5729 8343 5763
rect 8677 5729 8711 5763
rect 8999 5729 9033 5763
rect 10793 5729 10827 5763
rect 11437 5729 11471 5763
rect 13921 5729 13955 5763
rect 3525 5661 3559 5695
rect 4629 5661 4663 5695
rect 5814 5661 5848 5695
rect 6193 5661 6227 5695
rect 7849 5661 7883 5695
rect 7941 5661 7975 5695
rect 8033 5661 8067 5695
rect 8493 5661 8527 5695
rect 8769 5661 8803 5695
rect 10425 5661 10459 5695
rect 10885 5661 10919 5695
rect 11069 5661 11103 5695
rect 11621 5661 11655 5695
rect 14473 5661 14507 5695
rect 15117 7973 15151 8007
rect 15117 7293 15151 7327
rect 15301 8925 15335 8959
rect 15393 11169 15427 11203
rect 15209 7361 15243 7395
rect 15025 6409 15059 6443
rect 15393 7225 15427 7259
rect 15209 6341 15243 6375
rect 1685 5593 1719 5627
rect 3249 5593 3283 5627
rect 5181 5593 5215 5627
rect 8217 5593 8251 5627
rect 11805 5593 11839 5627
rect 13645 5593 13679 5627
rect 14933 5593 14967 5627
rect 15025 6273 15059 6307
rect 3157 5525 3191 5559
rect 5273 5525 5307 5559
rect 14105 5525 14139 5559
rect 14289 5525 14323 5559
rect 2513 5321 2547 5355
rect 3341 5321 3375 5355
rect 3801 5321 3835 5355
rect 4169 5321 4203 5355
rect 5365 5321 5399 5355
rect 7021 5321 7055 5355
rect 10517 5321 10551 5355
rect 11529 5321 11563 5355
rect 11989 5321 12023 5355
rect 4905 5253 4939 5287
rect 6101 5253 6135 5287
rect 1685 5185 1719 5219
rect 2329 5185 2363 5219
rect 2513 5185 2547 5219
rect 2789 5185 2823 5219
rect 2881 5185 2915 5219
rect 3065 5185 3099 5219
rect 3157 5185 3191 5219
rect 3341 5185 3375 5219
rect 3525 5185 3559 5219
rect 3709 5185 3743 5219
rect 4261 5185 4295 5219
rect 4721 5185 4755 5219
rect 4997 5185 5031 5219
rect 5089 5185 5123 5219
rect 5273 5185 5307 5219
rect 5641 5185 5675 5219
rect 5825 5185 5859 5219
rect 5917 5185 5951 5219
rect 6193 5185 6227 5219
rect 6561 5185 6595 5219
rect 6837 5185 6871 5219
rect 7113 5185 7147 5219
rect 8953 5185 8987 5219
rect 9137 5185 9171 5219
rect 9505 5185 9539 5219
rect 9965 5185 9999 5219
rect 10425 5185 10459 5219
rect 10517 5185 10551 5219
rect 10701 5185 10735 5219
rect 10977 5185 11011 5219
rect 11897 5185 11931 5219
rect 12349 5185 12383 5219
rect 12541 5185 12575 5219
rect 12633 5185 12667 5219
rect 14427 5185 14461 5219
rect 2697 5117 2731 5151
rect 4445 5117 4479 5151
rect 5549 5117 5583 5151
rect 6469 5117 6503 5151
rect 6653 5117 6687 5151
rect 10057 5117 10091 5151
rect 10885 5117 10919 5151
rect 12173 5117 12207 5151
rect 13001 5117 13035 5151
rect 4997 5049 5031 5083
rect 1593 4981 1627 5015
rect 2237 4981 2271 5015
rect 3065 4981 3099 5015
rect 3525 4981 3559 5015
rect 5733 4981 5767 5015
rect 6193 4981 6227 5015
rect 8401 4981 8435 5015
rect 9137 4981 9171 5015
rect 9413 4981 9447 5015
rect 9689 4981 9723 5015
rect 10241 4981 10275 5015
rect 11253 4981 11287 5015
rect 12449 4981 12483 5015
rect 3341 4777 3375 4811
rect 4813 4777 4847 4811
rect 6745 4777 6779 4811
rect 11667 4777 11701 4811
rect 14105 4777 14139 4811
rect 3525 4709 3559 4743
rect 8953 4709 8987 4743
rect 1409 4641 1443 4675
rect 4629 4641 4663 4675
rect 4905 4641 4939 4675
rect 5641 4641 5675 4675
rect 5917 4641 5951 4675
rect 7573 4641 7607 4675
rect 7757 4641 7791 4675
rect 8217 4641 8251 4675
rect 8677 4641 8711 4675
rect 9505 4641 9539 4675
rect 10241 4641 10275 4675
rect 13921 4641 13955 4675
rect 3249 4573 3283 4607
rect 3985 4573 4019 4607
rect 4353 4573 4387 4607
rect 4721 4573 4755 4607
rect 4997 4573 5031 4607
rect 5273 4573 5307 4607
rect 5365 4573 5399 4607
rect 5549 4573 5583 4607
rect 7481 4573 7515 4607
rect 8125 4573 8159 4607
rect 8585 4573 8619 4607
rect 9321 4573 9355 4607
rect 9873 4573 9907 4607
rect 13553 4573 13587 4607
rect 14473 4573 14507 4607
rect 1685 4505 1719 4539
rect 6653 4505 6687 4539
rect 3157 4437 3191 4471
rect 3893 4437 3927 4471
rect 4261 4437 4295 4471
rect 6929 4437 6963 4471
rect 7113 4437 7147 4471
rect 8493 4437 8527 4471
rect 9413 4437 9447 4471
rect 11805 4437 11839 4471
rect 14289 4437 14323 4471
rect 3617 4233 3651 4267
rect 4813 4233 4847 4267
rect 5641 4233 5675 4267
rect 6377 4233 6411 4267
rect 7573 4233 7607 4267
rect 8677 4233 8711 4267
rect 9137 4233 9171 4267
rect 9505 4233 9539 4267
rect 10149 4233 10183 4267
rect 10793 4233 10827 4267
rect 11529 4233 11563 4267
rect 11897 4233 11931 4267
rect 12587 4233 12621 4267
rect 3203 4165 3237 4199
rect 5181 4165 5215 4199
rect 7205 4165 7239 4199
rect 7389 4165 7423 4199
rect 1409 4097 1443 4131
rect 3341 4097 3375 4131
rect 3433 4097 3467 4131
rect 3709 4097 3743 4131
rect 3893 4097 3927 4131
rect 4721 4097 4755 4131
rect 5273 4097 5307 4131
rect 5917 4097 5951 4131
rect 6745 4097 6779 4131
rect 7113 4097 7147 4131
rect 8033 4097 8067 4131
rect 9965 4097 9999 4131
rect 10885 4097 10919 4131
rect 14013 4097 14047 4131
rect 14381 4097 14415 4131
rect 1777 4029 1811 4063
rect 4445 4029 4479 4063
rect 5365 4029 5399 4063
rect 5641 4029 5675 4063
rect 5825 4029 5859 4063
rect 6837 4029 6871 4063
rect 7941 4029 7975 4063
rect 8769 4029 8803 4063
rect 8953 4029 8987 4063
rect 9597 4029 9631 4063
rect 9689 4029 9723 4063
rect 10977 4029 11011 4063
rect 11989 4029 12023 4063
rect 12173 4029 12207 4063
rect 4169 3961 4203 3995
rect 8309 3961 8343 3995
rect 10425 3961 10459 3995
rect 3985 3893 4019 3927
rect 4629 3893 4663 3927
rect 6101 3893 6135 3927
rect 7021 3893 7055 3927
rect 7113 3893 7147 3927
rect 8217 3893 8251 3927
rect 11345 3893 11379 3927
rect 12357 3893 12391 3927
rect 2789 3689 2823 3723
rect 3065 3689 3099 3723
rect 3433 3689 3467 3723
rect 4537 3689 4571 3723
rect 5181 3689 5215 3723
rect 8401 3689 8435 3723
rect 10057 3689 10091 3723
rect 2881 3621 2915 3655
rect 8953 3621 8987 3655
rect 10793 3621 10827 3655
rect 10885 3621 10919 3655
rect 2697 3553 2731 3587
rect 3065 3553 3099 3587
rect 3157 3553 3191 3587
rect 4077 3553 4111 3587
rect 5641 3553 5675 3587
rect 6009 3553 6043 3587
rect 8217 3553 8251 3587
rect 9505 3553 9539 3587
rect 10517 3553 10551 3587
rect 11345 3553 11379 3587
rect 11529 3553 11563 3587
rect 13921 3553 13955 3587
rect 2973 3485 3007 3519
rect 3433 3485 3467 3519
rect 3617 3485 3651 3519
rect 3985 3485 4019 3519
rect 4445 3485 4479 3519
rect 4709 3485 4743 3519
rect 4813 3463 4847 3497
rect 4923 3485 4957 3519
rect 5089 3485 5123 3519
rect 5365 3485 5399 3519
rect 5549 3485 5583 3519
rect 7435 3485 7469 3519
rect 7941 3485 7975 3519
rect 8401 3485 8435 3519
rect 8493 3485 8527 3519
rect 10057 3485 10091 3519
rect 10425 3485 10459 3519
rect 5457 3417 5491 3451
rect 8677 3417 8711 3451
rect 11897 3417 11931 3451
rect 13645 3417 13679 3451
rect 14933 3417 14967 3451
rect 2605 3349 2639 3383
rect 3801 3349 3835 3383
rect 7573 3349 7607 3383
rect 8033 3349 8067 3383
rect 9321 3349 9355 3383
rect 9413 3349 9447 3383
rect 11253 3349 11287 3383
rect 11713 3349 11747 3383
rect 14105 3349 14139 3383
rect 14473 3349 14507 3383
rect 4353 3145 4387 3179
rect 7021 3145 7055 3179
rect 10517 3145 10551 3179
rect 11621 3145 11655 3179
rect 12633 3145 12667 3179
rect 2881 3077 2915 3111
rect 7757 3077 7791 3111
rect 10057 3077 10091 3111
rect 11069 3077 11103 3111
rect 12081 3077 12115 3111
rect 14105 3077 14139 3111
rect 6653 3009 6687 3043
rect 7205 3009 7239 3043
rect 7481 3009 7515 3043
rect 9413 3009 9447 3043
rect 9689 3009 9723 3043
rect 9781 3031 9815 3065
rect 9869 3009 9903 3043
rect 11345 3009 11379 3043
rect 11529 3009 11563 3043
rect 12449 3009 12483 3043
rect 14381 3009 14415 3043
rect 2605 2941 2639 2975
rect 4445 2941 4479 2975
rect 4721 2941 4755 2975
rect 6377 2941 6411 2975
rect 6561 2941 6595 2975
rect 7297 2941 7331 2975
rect 10609 2941 10643 2975
rect 10701 2941 10735 2975
rect 6193 2873 6227 2907
rect 10149 2873 10183 2907
rect 11253 2873 11287 2907
rect 11345 2873 11379 2907
rect 9229 2805 9263 2839
rect 8585 2601 8619 2635
rect 11345 2601 11379 2635
rect 14197 2601 14231 2635
rect 7849 2465 7883 2499
rect 8125 2465 8159 2499
rect 9597 2465 9631 2499
rect 11805 2465 11839 2499
rect 12081 2465 12115 2499
rect 12173 2465 12207 2499
rect 14381 2465 14415 2499
rect 3617 2397 3651 2431
rect 4077 2397 4111 2431
rect 7757 2397 7791 2431
rect 7941 2397 7975 2431
rect 8217 2397 8251 2431
rect 9045 2397 9079 2431
rect 9229 2397 9263 2431
rect 9321 2397 9355 2431
rect 11713 2397 11747 2431
rect 14105 2397 14139 2431
rect 5273 2329 5307 2363
rect 9873 2329 9907 2363
rect 12449 2329 12483 2363
rect 3985 2261 4019 2295
rect 6469 2261 6503 2295
rect 7297 2261 7331 2295
rect 9137 2261 9171 2295
rect 9505 2261 9539 2295
rect 13921 2261 13955 2295
rect 15025 2601 15059 2635
rect 14933 1037 14967 1071
<< metal1 >>
rect 14918 15008 14924 15020
rect 14879 14980 14924 15008
rect 14918 14968 14924 14980
rect 14976 14968 14982 15020
rect 1104 13626 14812 13648
rect 1104 13574 3248 13626
rect 3300 13574 3312 13626
rect 3364 13574 3376 13626
rect 3428 13574 3440 13626
rect 3492 13574 3504 13626
rect 3556 13574 7846 13626
rect 7898 13574 7910 13626
rect 7962 13574 7974 13626
rect 8026 13574 8038 13626
rect 8090 13574 8102 13626
rect 8154 13574 12443 13626
rect 12495 13574 12507 13626
rect 12559 13574 12571 13626
rect 12623 13574 12635 13626
rect 12687 13574 12699 13626
rect 12751 13574 14812 13626
rect 1104 13552 14812 13574
rect 2774 13472 2780 13524
rect 2832 13512 2838 13524
rect 2869 13515 2927 13521
rect 2869 13512 2881 13515
rect 2832 13484 2881 13512
rect 2832 13472 2838 13484
rect 2869 13481 2881 13484
rect 2915 13481 2927 13515
rect 4525 13515 4583 13521
rect 4525 13512 4537 13515
rect 2869 13475 2927 13481
rect 3804 13484 4537 13512
rect 3804 13385 3832 13484
rect 4525 13481 4537 13484
rect 4571 13481 4583 13515
rect 7558 13512 7564 13524
rect 7519 13484 7564 13512
rect 4525 13475 4583 13481
rect 7558 13472 7564 13484
rect 7616 13472 7622 13524
rect 8202 13472 8208 13524
rect 8260 13512 8266 13524
rect 8941 13515 8999 13521
rect 8941 13512 8953 13515
rect 8260 13484 8953 13512
rect 8260 13472 8266 13484
rect 8941 13481 8953 13484
rect 8987 13481 8999 13515
rect 13262 13512 13268 13524
rect 8941 13475 8999 13481
rect 9140 13484 13268 13512
rect 3973 13447 4031 13453
rect 3973 13413 3985 13447
rect 4019 13444 4031 13447
rect 5169 13447 5227 13453
rect 4019 13416 4476 13444
rect 4019 13413 4031 13416
rect 3973 13407 4031 13413
rect 3789 13379 3847 13385
rect 3789 13345 3801 13379
rect 3835 13345 3847 13379
rect 3789 13339 3847 13345
rect 2774 13268 2780 13320
rect 2832 13308 2838 13320
rect 3053 13311 3111 13317
rect 2832 13280 2877 13308
rect 2832 13268 2838 13280
rect 3053 13277 3065 13311
rect 3099 13277 3111 13311
rect 3053 13271 3111 13277
rect 3068 13240 3096 13271
rect 3970 13268 3976 13320
rect 4028 13308 4034 13320
rect 4065 13311 4123 13317
rect 4065 13308 4077 13311
rect 4028 13280 4077 13308
rect 4028 13268 4034 13280
rect 4065 13277 4077 13280
rect 4111 13308 4123 13311
rect 4154 13308 4160 13320
rect 4111 13280 4160 13308
rect 4111 13277 4123 13280
rect 4065 13271 4123 13277
rect 4154 13268 4160 13280
rect 4212 13268 4218 13320
rect 4338 13318 4344 13330
rect 4299 13290 4344 13318
rect 4338 13278 4344 13290
rect 4396 13278 4402 13330
rect 4448 13327 4476 13416
rect 5169 13413 5181 13447
rect 5215 13413 5227 13447
rect 5169 13407 5227 13413
rect 8297 13447 8355 13453
rect 8297 13413 8309 13447
rect 8343 13444 8355 13447
rect 8478 13444 8484 13456
rect 8343 13416 8484 13444
rect 8343 13413 8355 13416
rect 8297 13407 8355 13413
rect 4433 13321 4491 13327
rect 4433 13287 4445 13321
rect 4479 13308 4491 13321
rect 4522 13308 4528 13320
rect 4479 13287 4528 13308
rect 4433 13281 4528 13287
rect 4448 13280 4528 13281
rect 4522 13268 4528 13280
rect 4580 13268 4586 13320
rect 4617 13311 4675 13317
rect 4617 13277 4629 13311
rect 4663 13308 4675 13311
rect 5184 13308 5212 13407
rect 8478 13404 8484 13416
rect 8536 13404 8542 13456
rect 5258 13336 5264 13388
rect 5316 13376 5322 13388
rect 5721 13379 5779 13385
rect 5721 13376 5733 13379
rect 5316 13348 5733 13376
rect 5316 13336 5322 13348
rect 5721 13345 5733 13348
rect 5767 13376 5779 13379
rect 8846 13376 8852 13388
rect 5767 13348 8852 13376
rect 5767 13345 5779 13348
rect 5721 13339 5779 13345
rect 8846 13336 8852 13348
rect 8904 13336 8910 13388
rect 4663 13280 5212 13308
rect 7469 13311 7527 13317
rect 4663 13277 4675 13280
rect 4617 13271 4675 13277
rect 7469 13277 7481 13311
rect 7515 13308 7527 13311
rect 7650 13308 7656 13320
rect 7515 13280 7656 13308
rect 7515 13277 7527 13280
rect 7469 13271 7527 13277
rect 7650 13268 7656 13280
rect 7708 13268 7714 13320
rect 8202 13308 8208 13320
rect 8163 13280 8208 13308
rect 8202 13268 8208 13280
rect 8260 13268 8266 13320
rect 9140 13317 9168 13484
rect 13262 13472 13268 13484
rect 13320 13472 13326 13524
rect 13354 13472 13360 13524
rect 13412 13512 13418 13524
rect 14277 13515 14335 13521
rect 14277 13512 14289 13515
rect 13412 13484 14289 13512
rect 13412 13472 13418 13484
rect 14277 13481 14289 13484
rect 14323 13481 14335 13515
rect 14277 13475 14335 13481
rect 9493 13379 9551 13385
rect 9493 13376 9505 13379
rect 9232 13348 9505 13376
rect 8481 13311 8539 13317
rect 8481 13277 8493 13311
rect 8527 13308 8539 13311
rect 8757 13311 8815 13317
rect 8757 13308 8769 13311
rect 8527 13280 8769 13308
rect 8527 13277 8539 13280
rect 8481 13271 8539 13277
rect 8757 13277 8769 13280
rect 8803 13277 8815 13311
rect 8757 13271 8815 13277
rect 9125 13311 9183 13317
rect 9125 13277 9137 13311
rect 9171 13277 9183 13311
rect 9125 13271 9183 13277
rect 4264 13240 4476 13244
rect 9232 13240 9260 13348
rect 9493 13345 9505 13348
rect 9539 13376 9551 13379
rect 12069 13379 12127 13385
rect 12069 13376 12081 13379
rect 9539 13348 12081 13376
rect 9539 13345 9551 13348
rect 9493 13339 9551 13345
rect 12069 13345 12081 13348
rect 12115 13376 12127 13379
rect 12986 13376 12992 13388
rect 12115 13348 12992 13376
rect 12115 13345 12127 13348
rect 12069 13339 12127 13345
rect 12986 13336 12992 13348
rect 13044 13336 13050 13388
rect 9401 13311 9459 13317
rect 9401 13277 9413 13311
rect 9447 13308 9459 13311
rect 9861 13311 9919 13317
rect 9861 13308 9873 13311
rect 9447 13280 9873 13308
rect 9447 13277 9459 13280
rect 9401 13271 9459 13277
rect 9861 13277 9873 13280
rect 9907 13277 9919 13311
rect 9861 13271 9919 13277
rect 11330 13268 11336 13320
rect 11388 13308 11394 13320
rect 11793 13311 11851 13317
rect 11793 13308 11805 13311
rect 11388 13280 11805 13308
rect 11388 13268 11394 13280
rect 11793 13277 11805 13280
rect 11839 13277 11851 13311
rect 12434 13308 12440 13320
rect 12395 13280 12440 13308
rect 11793 13271 11851 13277
rect 12434 13268 12440 13280
rect 12492 13268 12498 13320
rect 14093 13311 14151 13317
rect 14093 13277 14105 13311
rect 14139 13308 14151 13311
rect 14182 13308 14188 13320
rect 14139 13280 14188 13308
rect 14139 13277 14151 13280
rect 14093 13271 14151 13277
rect 14182 13268 14188 13280
rect 14240 13268 14246 13320
rect 3068 13216 9260 13240
rect 3068 13212 4292 13216
rect 4448 13212 9260 13216
rect 10870 13200 10876 13252
rect 10928 13240 10934 13252
rect 11609 13243 11667 13249
rect 11609 13240 11621 13243
rect 10928 13212 11621 13240
rect 10928 13200 10934 13212
rect 11609 13209 11621 13212
rect 11655 13209 11667 13243
rect 11609 13203 11667 13209
rect 12912 13184 12940 13226
rect 2498 13132 2504 13184
rect 2556 13172 2562 13184
rect 2685 13175 2743 13181
rect 2685 13172 2697 13175
rect 2556 13144 2697 13172
rect 2556 13132 2562 13144
rect 2685 13141 2697 13144
rect 2731 13141 2743 13175
rect 2685 13135 2743 13141
rect 2866 13132 2872 13184
rect 2924 13172 2930 13184
rect 3789 13175 3847 13181
rect 3789 13172 3801 13175
rect 2924 13144 3801 13172
rect 2924 13132 2930 13144
rect 3789 13141 3801 13144
rect 3835 13141 3847 13175
rect 3789 13135 3847 13141
rect 4154 13132 4160 13184
rect 4212 13172 4218 13184
rect 4249 13175 4307 13181
rect 4249 13172 4261 13175
rect 4212 13144 4261 13172
rect 4212 13132 4218 13144
rect 4249 13141 4261 13144
rect 4295 13141 4307 13175
rect 4706 13172 4712 13184
rect 4667 13144 4712 13172
rect 4249 13135 4307 13141
rect 4706 13132 4712 13144
rect 4764 13132 4770 13184
rect 5442 13132 5448 13184
rect 5500 13172 5506 13184
rect 5537 13175 5595 13181
rect 5537 13172 5549 13175
rect 5500 13144 5549 13172
rect 5500 13132 5506 13144
rect 5537 13141 5549 13144
rect 5583 13141 5595 13175
rect 5537 13135 5595 13141
rect 5629 13175 5687 13181
rect 5629 13141 5641 13175
rect 5675 13172 5687 13175
rect 5902 13172 5908 13184
rect 5675 13144 5908 13172
rect 5675 13141 5687 13144
rect 5629 13135 5687 13141
rect 5902 13132 5908 13144
rect 5960 13132 5966 13184
rect 7929 13175 7987 13181
rect 7929 13141 7941 13175
rect 7975 13172 7987 13175
rect 8294 13172 8300 13184
rect 7975 13144 8300 13172
rect 7975 13141 7987 13144
rect 7929 13135 7987 13141
rect 8294 13132 8300 13144
rect 8352 13132 8358 13184
rect 8662 13172 8668 13184
rect 8623 13144 8668 13172
rect 8662 13132 8668 13144
rect 8720 13132 8726 13184
rect 8757 13175 8815 13181
rect 8757 13141 8769 13175
rect 8803 13172 8815 13175
rect 10778 13172 10784 13184
rect 8803 13144 10784 13172
rect 8803 13141 8815 13144
rect 8757 13135 8815 13141
rect 10778 13132 10784 13144
rect 10836 13132 10842 13184
rect 11287 13175 11345 13181
rect 11287 13141 11299 13175
rect 11333 13172 11345 13175
rect 11422 13172 11428 13184
rect 11333 13144 11428 13172
rect 11333 13141 11345 13144
rect 11287 13135 11345 13141
rect 11422 13132 11428 13144
rect 11480 13132 11486 13184
rect 11977 13175 12035 13181
rect 11977 13141 11989 13175
rect 12023 13172 12035 13175
rect 12710 13172 12716 13184
rect 12023 13144 12716 13172
rect 12023 13141 12035 13144
rect 11977 13135 12035 13141
rect 12710 13132 12716 13144
rect 12768 13132 12774 13184
rect 12894 13132 12900 13184
rect 12952 13132 12958 13184
rect 13863 13175 13921 13181
rect 13863 13141 13875 13175
rect 13909 13172 13921 13175
rect 14090 13172 14096 13184
rect 13909 13144 14096 13172
rect 13909 13141 13921 13144
rect 13863 13135 13921 13141
rect 14090 13132 14096 13144
rect 14148 13132 14154 13184
rect 1104 13082 14812 13104
rect 1104 13030 5547 13082
rect 5599 13030 5611 13082
rect 5663 13030 5675 13082
rect 5727 13030 5739 13082
rect 5791 13030 5803 13082
rect 5855 13030 10144 13082
rect 10196 13030 10208 13082
rect 10260 13030 10272 13082
rect 10324 13030 10336 13082
rect 10388 13030 10400 13082
rect 10452 13030 14812 13082
rect 1104 13008 14812 13030
rect 2958 12928 2964 12980
rect 3016 12968 3022 12980
rect 4706 12968 4712 12980
rect 3016 12940 4712 12968
rect 3016 12928 3022 12940
rect 3252 12886 3280 12940
rect 4706 12928 4712 12940
rect 4764 12928 4770 12980
rect 5442 12968 5448 12980
rect 5403 12940 5448 12968
rect 5442 12928 5448 12940
rect 5500 12928 5506 12980
rect 5813 12971 5871 12977
rect 5813 12937 5825 12971
rect 5859 12968 5871 12971
rect 6365 12971 6423 12977
rect 6365 12968 6377 12971
rect 5859 12940 6377 12968
rect 5859 12937 5871 12940
rect 5813 12931 5871 12937
rect 6365 12937 6377 12940
rect 6411 12937 6423 12971
rect 6365 12931 6423 12937
rect 12434 12928 12440 12980
rect 12492 12968 12498 12980
rect 13311 12971 13369 12977
rect 13311 12968 13323 12971
rect 12492 12940 13323 12968
rect 12492 12928 12498 12940
rect 13311 12937 13323 12940
rect 13357 12937 13369 12971
rect 14182 12968 14188 12980
rect 14143 12940 14188 12968
rect 13311 12931 13369 12937
rect 14182 12928 14188 12940
rect 14240 12928 14246 12980
rect 5077 12903 5135 12909
rect 5077 12869 5089 12903
rect 5123 12900 5135 12903
rect 5123 12872 6040 12900
rect 5123 12869 5135 12872
rect 5077 12863 5135 12869
rect 2498 12832 2504 12844
rect 2459 12804 2504 12832
rect 2498 12792 2504 12804
rect 2556 12792 2562 12844
rect 2866 12832 2872 12844
rect 2827 12804 2872 12832
rect 2866 12792 2872 12804
rect 2924 12792 2930 12844
rect 4614 12832 4620 12844
rect 4575 12804 4620 12832
rect 4614 12792 4620 12804
rect 4672 12792 4678 12844
rect 4801 12835 4859 12841
rect 4801 12801 4813 12835
rect 4847 12801 4859 12835
rect 4801 12795 4859 12801
rect 5353 12835 5411 12841
rect 5353 12801 5365 12835
rect 5399 12801 5411 12835
rect 5353 12795 5411 12801
rect 4338 12705 4344 12708
rect 4295 12699 4344 12705
rect 4295 12696 4307 12699
rect 4251 12668 4307 12696
rect 4295 12665 4307 12668
rect 4341 12665 4344 12699
rect 4295 12659 4344 12665
rect 4338 12656 4344 12659
rect 4396 12696 4402 12708
rect 4816 12696 4844 12795
rect 4396 12668 4844 12696
rect 4396 12656 4402 12668
rect 4816 12628 4844 12668
rect 4890 12656 4896 12708
rect 4948 12696 4954 12708
rect 5368 12696 5396 12795
rect 6012 12776 6040 12872
rect 7024 12872 8524 12900
rect 6733 12835 6791 12841
rect 6733 12801 6745 12835
rect 6779 12801 6791 12835
rect 6733 12795 6791 12801
rect 5902 12764 5908 12776
rect 5863 12736 5908 12764
rect 5902 12724 5908 12736
rect 5960 12724 5966 12776
rect 5994 12724 6000 12776
rect 6052 12764 6058 12776
rect 6641 12767 6699 12773
rect 6052 12736 6145 12764
rect 6052 12724 6058 12736
rect 6641 12733 6653 12767
rect 6687 12733 6699 12767
rect 6641 12727 6699 12733
rect 6656 12696 6684 12727
rect 4948 12668 6684 12696
rect 4948 12656 4954 12668
rect 5074 12628 5080 12640
rect 4816 12600 5080 12628
rect 5074 12588 5080 12600
rect 5132 12628 5138 12640
rect 6748 12628 6776 12795
rect 6914 12792 6920 12844
rect 6972 12832 6978 12844
rect 7024 12841 7052 12872
rect 7282 12841 7288 12844
rect 7009 12835 7067 12841
rect 7009 12832 7021 12835
rect 6972 12804 7021 12832
rect 6972 12792 6978 12804
rect 7009 12801 7021 12804
rect 7055 12801 7067 12835
rect 7276 12832 7288 12841
rect 7243 12804 7288 12832
rect 7009 12795 7067 12801
rect 7276 12795 7288 12804
rect 7282 12792 7288 12795
rect 7340 12792 7346 12844
rect 8496 12773 8524 12872
rect 8662 12860 8668 12912
rect 8720 12900 8726 12912
rect 8757 12903 8815 12909
rect 8757 12900 8769 12903
rect 8720 12872 8769 12900
rect 8720 12860 8726 12872
rect 8757 12869 8769 12872
rect 8803 12869 8815 12903
rect 8757 12863 8815 12869
rect 9306 12860 9312 12912
rect 9364 12860 9370 12912
rect 10689 12903 10747 12909
rect 10689 12869 10701 12903
rect 10735 12900 10747 12903
rect 11330 12900 11336 12912
rect 10735 12872 11336 12900
rect 10735 12869 10747 12872
rect 10689 12863 10747 12869
rect 11330 12860 11336 12872
rect 11388 12860 11394 12912
rect 12894 12860 12900 12912
rect 12952 12860 12958 12912
rect 11146 12832 11152 12844
rect 11107 12804 11152 12832
rect 11146 12792 11152 12804
rect 11204 12792 11210 12844
rect 11517 12835 11575 12841
rect 11517 12801 11529 12835
rect 11563 12832 11575 12835
rect 13814 12832 13820 12844
rect 11563 12804 12020 12832
rect 13775 12804 13820 12832
rect 11563 12801 11575 12804
rect 11517 12795 11575 12801
rect 8481 12767 8539 12773
rect 8481 12733 8493 12767
rect 8527 12733 8539 12767
rect 8481 12727 8539 12733
rect 8386 12628 8392 12640
rect 5132 12600 6776 12628
rect 8347 12600 8392 12628
rect 5132 12588 5138 12600
rect 8386 12588 8392 12600
rect 8444 12588 8450 12640
rect 8496 12628 8524 12727
rect 8846 12724 8852 12776
rect 8904 12764 8910 12776
rect 10505 12767 10563 12773
rect 10505 12764 10517 12767
rect 8904 12736 10517 12764
rect 8904 12724 8910 12736
rect 10505 12733 10517 12736
rect 10551 12733 10563 12767
rect 10505 12727 10563 12733
rect 10520 12696 10548 12727
rect 11422 12724 11428 12776
rect 11480 12764 11486 12776
rect 11885 12767 11943 12773
rect 11885 12764 11897 12767
rect 11480 12736 11897 12764
rect 11480 12724 11486 12736
rect 11885 12733 11897 12736
rect 11931 12733 11943 12767
rect 11992 12764 12020 12804
rect 13814 12792 13820 12804
rect 13872 12792 13878 12844
rect 14090 12832 14096 12844
rect 14051 12804 14096 12832
rect 14090 12792 14096 12804
rect 14148 12792 14154 12844
rect 14274 12832 14280 12844
rect 14235 12804 14280 12832
rect 14274 12792 14280 12804
rect 14332 12792 14338 12844
rect 12986 12764 12992 12776
rect 11992 12736 12992 12764
rect 11885 12727 11943 12733
rect 12986 12724 12992 12736
rect 13044 12724 13050 12776
rect 13630 12724 13636 12776
rect 13688 12764 13694 12776
rect 13725 12767 13783 12773
rect 13725 12764 13737 12767
rect 13688 12736 13737 12764
rect 13688 12724 13694 12736
rect 13725 12733 13737 12736
rect 13771 12733 13783 12767
rect 13725 12727 13783 12733
rect 11514 12696 11520 12708
rect 10520 12668 11520 12696
rect 11514 12656 11520 12668
rect 11572 12656 11578 12708
rect 13446 12696 13452 12708
rect 13407 12668 13452 12696
rect 13446 12656 13452 12668
rect 13504 12656 13510 12708
rect 9490 12628 9496 12640
rect 8496 12600 9496 12628
rect 9490 12588 9496 12600
rect 9548 12588 9554 12640
rect 10873 12631 10931 12637
rect 10873 12597 10885 12631
rect 10919 12628 10931 12631
rect 10962 12628 10968 12640
rect 10919 12600 10968 12628
rect 10919 12597 10931 12600
rect 10873 12591 10931 12597
rect 10962 12588 10968 12600
rect 11020 12588 11026 12640
rect 11241 12631 11299 12637
rect 11241 12597 11253 12631
rect 11287 12628 11299 12631
rect 11330 12628 11336 12640
rect 11287 12600 11336 12628
rect 11287 12597 11299 12600
rect 11241 12591 11299 12597
rect 11330 12588 11336 12600
rect 11388 12588 11394 12640
rect 1104 12538 14812 12560
rect 1104 12486 3248 12538
rect 3300 12486 3312 12538
rect 3364 12486 3376 12538
rect 3428 12486 3440 12538
rect 3492 12486 3504 12538
rect 3556 12486 7846 12538
rect 7898 12486 7910 12538
rect 7962 12486 7974 12538
rect 8026 12486 8038 12538
rect 8090 12486 8102 12538
rect 8154 12486 12443 12538
rect 12495 12486 12507 12538
rect 12559 12486 12571 12538
rect 12623 12486 12635 12538
rect 12687 12486 12699 12538
rect 12751 12486 14812 12538
rect 1104 12464 14812 12486
rect 7558 12424 7564 12436
rect 7519 12396 7564 12424
rect 7558 12384 7564 12396
rect 7616 12384 7622 12436
rect 7650 12384 7656 12436
rect 7708 12424 7714 12436
rect 8021 12427 8079 12433
rect 8021 12424 8033 12427
rect 7708 12396 8033 12424
rect 7708 12384 7714 12396
rect 8021 12393 8033 12396
rect 8067 12393 8079 12427
rect 8021 12387 8079 12393
rect 4065 12359 4123 12365
rect 4065 12325 4077 12359
rect 4111 12356 4123 12359
rect 6086 12356 6092 12368
rect 4111 12328 6092 12356
rect 4111 12325 4123 12328
rect 4065 12319 4123 12325
rect 6086 12316 6092 12328
rect 6144 12316 6150 12368
rect 8036 12356 8064 12387
rect 8202 12384 8208 12436
rect 8260 12424 8266 12436
rect 8297 12427 8355 12433
rect 8297 12424 8309 12427
rect 8260 12396 8309 12424
rect 8260 12384 8266 12396
rect 8297 12393 8309 12396
rect 8343 12393 8355 12427
rect 8297 12387 8355 12393
rect 11146 12384 11152 12436
rect 11204 12424 11210 12436
rect 11609 12427 11667 12433
rect 11609 12424 11621 12427
rect 11204 12396 11621 12424
rect 11204 12384 11210 12396
rect 11609 12393 11621 12396
rect 11655 12393 11667 12427
rect 11609 12387 11667 12393
rect 11790 12384 11796 12436
rect 11848 12424 11854 12436
rect 13630 12424 13636 12436
rect 11848 12396 13636 12424
rect 11848 12384 11854 12396
rect 13630 12384 13636 12396
rect 13688 12384 13694 12436
rect 14274 12424 14280 12436
rect 14235 12396 14280 12424
rect 14274 12384 14280 12396
rect 14332 12384 14338 12436
rect 8938 12356 8944 12368
rect 8036 12328 8944 12356
rect 8938 12316 8944 12328
rect 8996 12316 9002 12368
rect 2774 12288 2780 12300
rect 1872 12260 2780 12288
rect 1765 12223 1823 12229
rect 1765 12189 1777 12223
rect 1811 12220 1823 12223
rect 1872 12220 1900 12260
rect 2774 12248 2780 12260
rect 2832 12248 2838 12300
rect 3513 12291 3571 12297
rect 3513 12257 3525 12291
rect 3559 12288 3571 12291
rect 4798 12288 4804 12300
rect 3559 12260 4384 12288
rect 4759 12260 4804 12288
rect 3559 12257 3571 12260
rect 3513 12251 3571 12257
rect 3970 12220 3976 12232
rect 1811 12192 1900 12220
rect 3931 12192 3976 12220
rect 1811 12189 1823 12192
rect 1765 12183 1823 12189
rect 1872 12164 1900 12192
rect 3970 12180 3976 12192
rect 4028 12180 4034 12232
rect 4062 12180 4068 12232
rect 4120 12220 4126 12232
rect 4356 12229 4384 12260
rect 4798 12248 4804 12260
rect 4856 12248 4862 12300
rect 5077 12291 5135 12297
rect 5077 12257 5089 12291
rect 5123 12288 5135 12291
rect 5350 12288 5356 12300
rect 5123 12260 5356 12288
rect 5123 12257 5135 12260
rect 5077 12251 5135 12257
rect 5350 12248 5356 12260
rect 5408 12248 5414 12300
rect 5721 12291 5779 12297
rect 5721 12257 5733 12291
rect 5767 12257 5779 12291
rect 5721 12251 5779 12257
rect 4249 12223 4307 12229
rect 4249 12220 4261 12223
rect 4120 12192 4261 12220
rect 4120 12180 4126 12192
rect 4249 12189 4261 12192
rect 4295 12189 4307 12223
rect 4249 12183 4307 12189
rect 4341 12223 4399 12229
rect 4341 12189 4353 12223
rect 4387 12220 4399 12223
rect 4614 12220 4620 12232
rect 4387 12192 4620 12220
rect 4387 12189 4399 12192
rect 4341 12183 4399 12189
rect 4614 12180 4620 12192
rect 4672 12220 4678 12232
rect 4709 12223 4767 12229
rect 4709 12220 4721 12223
rect 4672 12192 4721 12220
rect 4672 12180 4678 12192
rect 4709 12189 4721 12192
rect 4755 12189 4767 12223
rect 4709 12183 4767 12189
rect 4982 12180 4988 12232
rect 5040 12220 5046 12232
rect 5258 12220 5264 12232
rect 5040 12192 5264 12220
rect 5040 12180 5046 12192
rect 5258 12180 5264 12192
rect 5316 12220 5322 12232
rect 5736 12220 5764 12251
rect 8386 12248 8392 12300
rect 8444 12288 8450 12300
rect 10137 12291 10195 12297
rect 8444 12260 8616 12288
rect 8444 12248 8450 12260
rect 5316 12192 5764 12220
rect 5316 12180 5322 12192
rect 5902 12180 5908 12232
rect 5960 12180 5966 12232
rect 6181 12223 6239 12229
rect 6181 12189 6193 12223
rect 6227 12220 6239 12223
rect 6914 12220 6920 12232
rect 6227 12192 6920 12220
rect 6227 12189 6239 12192
rect 6181 12183 6239 12189
rect 6914 12180 6920 12192
rect 6972 12180 6978 12232
rect 7558 12180 7564 12232
rect 7616 12220 7622 12232
rect 7745 12223 7803 12229
rect 7745 12220 7757 12223
rect 7616 12192 7757 12220
rect 7616 12180 7622 12192
rect 7745 12189 7757 12192
rect 7791 12189 7803 12223
rect 8294 12220 8300 12232
rect 8255 12192 8300 12220
rect 7745 12183 7803 12189
rect 8294 12180 8300 12192
rect 8352 12180 8358 12232
rect 8588 12229 8616 12260
rect 10137 12257 10149 12291
rect 10183 12288 10195 12291
rect 10870 12288 10876 12300
rect 10183 12260 10876 12288
rect 10183 12257 10195 12260
rect 10137 12251 10195 12257
rect 10870 12248 10876 12260
rect 10928 12248 10934 12300
rect 12342 12248 12348 12300
rect 12400 12288 12406 12300
rect 13909 12291 13967 12297
rect 13909 12288 13921 12291
rect 12400 12260 13921 12288
rect 12400 12248 12406 12260
rect 13909 12257 13921 12260
rect 13955 12257 13967 12291
rect 13909 12251 13967 12257
rect 8573 12223 8631 12229
rect 8573 12189 8585 12223
rect 8619 12189 8631 12223
rect 8573 12183 8631 12189
rect 9490 12180 9496 12232
rect 9548 12220 9554 12232
rect 9861 12223 9919 12229
rect 9861 12220 9873 12223
rect 9548 12192 9873 12220
rect 9548 12180 9554 12192
rect 9861 12189 9873 12192
rect 9907 12189 9919 12223
rect 9861 12183 9919 12189
rect 14185 12223 14243 12229
rect 14185 12189 14197 12223
rect 14231 12220 14243 12223
rect 14461 12223 14519 12229
rect 14461 12220 14473 12223
rect 14231 12192 14473 12220
rect 14231 12189 14243 12192
rect 14185 12183 14243 12189
rect 14461 12189 14473 12192
rect 14507 12220 14519 12223
rect 14921 12223 14979 12229
rect 14921 12220 14933 12223
rect 14507 12192 14933 12220
rect 14507 12189 14519 12192
rect 14461 12183 14519 12189
rect 14921 12189 14933 12192
rect 14967 12189 14979 12223
rect 14921 12183 14979 12189
rect 1854 12112 1860 12164
rect 1912 12112 1918 12164
rect 2038 12152 2044 12164
rect 1999 12124 2044 12152
rect 2038 12112 2044 12124
rect 2096 12112 2102 12164
rect 3789 12155 3847 12161
rect 2976 12096 3004 12138
rect 3789 12121 3801 12155
rect 3835 12121 3847 12155
rect 4890 12152 4896 12164
rect 3789 12115 3847 12121
rect 4126 12124 4896 12152
rect 2958 12044 2964 12096
rect 3016 12044 3022 12096
rect 3602 12044 3608 12096
rect 3660 12084 3666 12096
rect 3804 12084 3832 12115
rect 4126 12084 4154 12124
rect 4890 12112 4896 12124
rect 4948 12112 4954 12164
rect 5920 12152 5948 12180
rect 6454 12161 6460 12164
rect 6448 12152 6460 12161
rect 5920 12124 6460 12152
rect 6448 12115 6460 12124
rect 6454 12112 6460 12115
rect 6512 12112 6518 12164
rect 8389 12155 8447 12161
rect 8389 12152 8401 12155
rect 8220 12124 8401 12152
rect 3660 12056 4154 12084
rect 3660 12044 3666 12056
rect 4430 12044 4436 12096
rect 4488 12084 4494 12096
rect 5169 12087 5227 12093
rect 5169 12084 5181 12087
rect 4488 12056 5181 12084
rect 4488 12044 4494 12056
rect 5169 12053 5181 12056
rect 5215 12053 5227 12087
rect 5169 12047 5227 12053
rect 5442 12044 5448 12096
rect 5500 12084 5506 12096
rect 5537 12087 5595 12093
rect 5537 12084 5549 12087
rect 5500 12056 5549 12084
rect 5500 12044 5506 12056
rect 5537 12053 5549 12056
rect 5583 12053 5595 12087
rect 5537 12047 5595 12053
rect 5629 12087 5687 12093
rect 5629 12053 5641 12087
rect 5675 12084 5687 12087
rect 5902 12084 5908 12096
rect 5675 12056 5908 12084
rect 5675 12053 5687 12056
rect 5629 12047 5687 12053
rect 5902 12044 5908 12056
rect 5960 12044 5966 12096
rect 8220 12093 8248 12124
rect 8389 12121 8401 12124
rect 8435 12121 8447 12155
rect 11885 12155 11943 12161
rect 8389 12115 8447 12121
rect 8205 12087 8263 12093
rect 8205 12053 8217 12087
rect 8251 12053 8263 12087
rect 8205 12047 8263 12053
rect 8757 12087 8815 12093
rect 8757 12053 8769 12087
rect 8803 12084 8815 12087
rect 9306 12084 9312 12096
rect 8803 12056 9312 12084
rect 8803 12053 8815 12056
rect 8757 12047 8815 12053
rect 9306 12044 9312 12056
rect 9364 12084 9370 12096
rect 9677 12087 9735 12093
rect 9677 12084 9689 12087
rect 9364 12056 9689 12084
rect 9364 12044 9370 12056
rect 9677 12053 9689 12056
rect 9723 12084 9735 12087
rect 10612 12084 10640 12138
rect 11885 12121 11897 12155
rect 11931 12152 11943 12155
rect 12158 12152 12164 12164
rect 11931 12124 12164 12152
rect 11931 12121 11943 12124
rect 11885 12115 11943 12121
rect 12158 12112 12164 12124
rect 12216 12112 12222 12164
rect 13633 12155 13691 12161
rect 10962 12084 10968 12096
rect 9723 12056 10968 12084
rect 9723 12053 9735 12056
rect 9677 12047 9735 12053
rect 10962 12044 10968 12056
rect 11020 12084 11026 12096
rect 11606 12084 11612 12096
rect 11020 12056 11612 12084
rect 11020 12044 11026 12056
rect 11606 12044 11612 12056
rect 11664 12084 11670 12096
rect 11701 12087 11759 12093
rect 11701 12084 11713 12087
rect 11664 12056 11713 12084
rect 11664 12044 11670 12056
rect 11701 12053 11713 12056
rect 11747 12084 11759 12087
rect 12250 12084 12256 12096
rect 11747 12056 12256 12084
rect 11747 12053 11759 12056
rect 11701 12047 11759 12053
rect 12250 12044 12256 12056
rect 12308 12084 12314 12096
rect 12452 12084 12480 12138
rect 13633 12121 13645 12155
rect 13679 12152 13691 12155
rect 14274 12152 14280 12164
rect 13679 12124 14280 12152
rect 13679 12121 13691 12124
rect 13633 12115 13691 12121
rect 14274 12112 14280 12124
rect 14332 12112 14338 12164
rect 12894 12084 12900 12096
rect 12308 12056 12900 12084
rect 12308 12044 12314 12056
rect 12894 12044 12900 12056
rect 12952 12044 12958 12096
rect 1104 11994 14812 12016
rect 1104 11942 5547 11994
rect 5599 11942 5611 11994
rect 5663 11942 5675 11994
rect 5727 11942 5739 11994
rect 5791 11942 5803 11994
rect 5855 11942 10144 11994
rect 10196 11942 10208 11994
rect 10260 11942 10272 11994
rect 10324 11942 10336 11994
rect 10388 11942 10400 11994
rect 10452 11942 14812 11994
rect 1104 11920 14812 11942
rect 2038 11840 2044 11892
rect 2096 11880 2102 11892
rect 3237 11883 3295 11889
rect 3237 11880 3249 11883
rect 2096 11852 3249 11880
rect 2096 11840 2102 11852
rect 3237 11849 3249 11852
rect 3283 11849 3295 11883
rect 3789 11883 3847 11889
rect 3789 11880 3801 11883
rect 3237 11843 3295 11849
rect 3436 11852 3801 11880
rect 3237 11679 3295 11685
rect 3237 11645 3249 11679
rect 3283 11676 3295 11679
rect 3436 11676 3464 11852
rect 3789 11849 3801 11852
rect 3835 11849 3847 11883
rect 3789 11843 3847 11849
rect 4798 11840 4804 11892
rect 4856 11880 4862 11892
rect 4985 11883 5043 11889
rect 4985 11880 4997 11883
rect 4856 11852 4997 11880
rect 4856 11840 4862 11852
rect 4985 11849 4997 11852
rect 5031 11849 5043 11883
rect 5442 11880 5448 11892
rect 5403 11852 5448 11880
rect 4985 11843 5043 11849
rect 5442 11840 5448 11852
rect 5500 11840 5506 11892
rect 8297 11883 8355 11889
rect 8297 11849 8309 11883
rect 8343 11880 8355 11883
rect 8478 11880 8484 11892
rect 8343 11852 8484 11880
rect 8343 11849 8355 11852
rect 8297 11843 8355 11849
rect 8478 11840 8484 11852
rect 8536 11840 8542 11892
rect 8754 11840 8760 11892
rect 8812 11880 8818 11892
rect 10137 11883 10195 11889
rect 8812 11852 9536 11880
rect 8812 11840 8818 11852
rect 4062 11812 4068 11824
rect 3528 11784 4068 11812
rect 3528 11753 3556 11784
rect 4062 11772 4068 11784
rect 4120 11772 4126 11824
rect 4540 11784 4936 11812
rect 3513 11747 3571 11753
rect 3513 11713 3525 11747
rect 3559 11713 3571 11747
rect 3513 11707 3571 11713
rect 3789 11747 3847 11753
rect 3789 11713 3801 11747
rect 3835 11713 3847 11747
rect 3789 11707 3847 11713
rect 3973 11747 4031 11753
rect 3973 11713 3985 11747
rect 4019 11744 4031 11747
rect 4430 11744 4436 11756
rect 4019 11716 4436 11744
rect 4019 11713 4031 11716
rect 3973 11707 4031 11713
rect 3283 11648 3464 11676
rect 3283 11645 3295 11648
rect 3237 11639 3295 11645
rect 3421 11611 3479 11617
rect 3421 11577 3433 11611
rect 3467 11608 3479 11611
rect 3804 11608 3832 11707
rect 4430 11704 4436 11716
rect 4488 11704 4494 11756
rect 4540 11753 4568 11784
rect 4908 11756 4936 11784
rect 5350 11772 5356 11824
rect 5408 11812 5414 11824
rect 5813 11815 5871 11821
rect 5813 11812 5825 11815
rect 5408 11784 5825 11812
rect 5408 11772 5414 11784
rect 5813 11781 5825 11784
rect 5859 11781 5871 11815
rect 6914 11812 6920 11824
rect 5813 11775 5871 11781
rect 6380 11784 6920 11812
rect 4525 11747 4583 11753
rect 4525 11713 4537 11747
rect 4571 11713 4583 11747
rect 4525 11707 4583 11713
rect 4617 11747 4675 11753
rect 4617 11713 4629 11747
rect 4663 11713 4675 11747
rect 4617 11707 4675 11713
rect 4246 11636 4252 11688
rect 4304 11676 4310 11688
rect 4632 11676 4660 11707
rect 4706 11704 4712 11756
rect 4764 11744 4770 11756
rect 4801 11747 4859 11753
rect 4801 11744 4813 11747
rect 4764 11716 4813 11744
rect 4764 11704 4770 11716
rect 4801 11713 4813 11716
rect 4847 11713 4859 11747
rect 4801 11707 4859 11713
rect 4890 11704 4896 11756
rect 4948 11744 4954 11756
rect 4948 11716 4993 11744
rect 4948 11704 4954 11716
rect 5074 11704 5080 11756
rect 5132 11744 5138 11756
rect 6380 11753 6408 11784
rect 6914 11772 6920 11784
rect 6972 11772 6978 11824
rect 9401 11815 9459 11821
rect 9401 11812 9413 11815
rect 8588 11784 9413 11812
rect 6365 11747 6423 11753
rect 5132 11716 5177 11744
rect 5132 11704 5138 11716
rect 6365 11713 6377 11747
rect 6411 11713 6423 11747
rect 6621 11747 6679 11753
rect 6621 11744 6633 11747
rect 6365 11707 6423 11713
rect 6472 11716 6633 11744
rect 4304 11648 4660 11676
rect 4304 11636 4310 11648
rect 5350 11636 5356 11688
rect 5408 11676 5414 11688
rect 5902 11676 5908 11688
rect 5408 11648 5908 11676
rect 5408 11636 5414 11648
rect 5902 11636 5908 11648
rect 5960 11636 5966 11688
rect 5994 11636 6000 11688
rect 6052 11676 6058 11688
rect 6472 11676 6500 11716
rect 6621 11713 6633 11716
rect 6667 11744 6679 11747
rect 8021 11747 8079 11753
rect 8021 11744 8033 11747
rect 6667 11716 8033 11744
rect 6667 11713 6679 11716
rect 6621 11707 6679 11713
rect 8021 11713 8033 11716
rect 8067 11744 8079 11747
rect 8478 11744 8484 11756
rect 8067 11716 8484 11744
rect 8067 11713 8079 11716
rect 8021 11707 8079 11713
rect 8478 11704 8484 11716
rect 8536 11704 8542 11756
rect 8588 11753 8616 11784
rect 9401 11781 9413 11784
rect 9447 11781 9459 11815
rect 9401 11775 9459 11781
rect 8573 11747 8631 11753
rect 8573 11713 8585 11747
rect 8619 11713 8631 11747
rect 8573 11707 8631 11713
rect 8938 11704 8944 11756
rect 8996 11704 9002 11756
rect 9030 11704 9036 11756
rect 9088 11744 9094 11756
rect 9088 11716 9133 11744
rect 9088 11704 9094 11716
rect 9214 11704 9220 11756
rect 9272 11744 9278 11756
rect 9508 11753 9536 11852
rect 10137 11849 10149 11883
rect 10183 11880 10195 11883
rect 10321 11883 10379 11889
rect 10321 11880 10333 11883
rect 10183 11852 10333 11880
rect 10183 11849 10195 11852
rect 10137 11843 10195 11849
rect 10321 11849 10333 11852
rect 10367 11849 10379 11883
rect 10321 11843 10379 11849
rect 10870 11840 10876 11892
rect 10928 11880 10934 11892
rect 10965 11883 11023 11889
rect 10965 11880 10977 11883
rect 10928 11852 10977 11880
rect 10928 11840 10934 11852
rect 10965 11849 10977 11852
rect 11011 11849 11023 11883
rect 10965 11843 11023 11849
rect 11054 11840 11060 11892
rect 11112 11880 11118 11892
rect 11333 11883 11391 11889
rect 11333 11880 11345 11883
rect 11112 11852 11345 11880
rect 11112 11840 11118 11852
rect 11333 11849 11345 11852
rect 11379 11880 11391 11883
rect 14274 11880 14280 11892
rect 11379 11852 14136 11880
rect 14235 11852 14280 11880
rect 11379 11849 11391 11852
rect 11333 11843 11391 11849
rect 10229 11815 10287 11821
rect 10229 11781 10241 11815
rect 10275 11812 10287 11815
rect 11146 11812 11152 11824
rect 10275 11784 11152 11812
rect 10275 11781 10287 11784
rect 10229 11775 10287 11781
rect 11146 11772 11152 11784
rect 11204 11772 11210 11824
rect 11606 11812 11612 11824
rect 11567 11784 11612 11812
rect 11606 11772 11612 11784
rect 11664 11772 11670 11824
rect 12802 11812 12808 11824
rect 12763 11784 12808 11812
rect 12802 11772 12808 11784
rect 12860 11772 12866 11824
rect 13354 11772 13360 11824
rect 13412 11772 13418 11824
rect 14108 11812 14136 11852
rect 14274 11840 14280 11852
rect 14332 11840 14338 11892
rect 15289 11815 15347 11821
rect 15289 11812 15301 11815
rect 14108 11784 15301 11812
rect 15289 11781 15301 11784
rect 15335 11781 15347 11815
rect 15289 11775 15347 11781
rect 9309 11747 9367 11753
rect 9309 11744 9321 11747
rect 9272 11716 9321 11744
rect 9272 11704 9278 11716
rect 9309 11713 9321 11716
rect 9355 11713 9367 11747
rect 9309 11707 9367 11713
rect 9493 11747 9551 11753
rect 9493 11713 9505 11747
rect 9539 11713 9551 11747
rect 9493 11707 9551 11713
rect 9585 11747 9643 11753
rect 9585 11713 9597 11747
rect 9631 11713 9643 11747
rect 9950 11744 9956 11756
rect 9911 11716 9956 11744
rect 9585 11707 9643 11713
rect 7834 11676 7840 11688
rect 6052 11648 6097 11676
rect 6380 11648 6500 11676
rect 7760 11648 7840 11676
rect 6052 11636 6058 11648
rect 4614 11608 4620 11620
rect 3467 11580 4620 11608
rect 3467 11577 3479 11580
rect 3421 11571 3479 11577
rect 4614 11568 4620 11580
rect 4672 11568 4678 11620
rect 5920 11608 5948 11636
rect 6380 11608 6408 11648
rect 7760 11617 7788 11648
rect 7834 11636 7840 11648
rect 7892 11636 7898 11688
rect 8297 11679 8355 11685
rect 8297 11645 8309 11679
rect 8343 11676 8355 11679
rect 8757 11679 8815 11685
rect 8343 11648 8708 11676
rect 8343 11645 8355 11648
rect 8297 11639 8355 11645
rect 5920 11580 6408 11608
rect 7745 11611 7803 11617
rect 7745 11577 7757 11611
rect 7791 11577 7803 11611
rect 7745 11571 7803 11577
rect 8205 11611 8263 11617
rect 8205 11577 8217 11611
rect 8251 11608 8263 11611
rect 8481 11611 8539 11617
rect 8481 11608 8493 11611
rect 8251 11580 8493 11608
rect 8251 11577 8263 11580
rect 8205 11571 8263 11577
rect 8481 11577 8493 11580
rect 8527 11577 8539 11611
rect 8680 11608 8708 11648
rect 8757 11645 8769 11679
rect 8803 11676 8815 11679
rect 8956 11676 8984 11704
rect 8803 11648 8984 11676
rect 8803 11645 8815 11648
rect 8757 11639 8815 11645
rect 9398 11636 9404 11688
rect 9456 11676 9462 11688
rect 9600 11676 9628 11707
rect 9950 11704 9956 11716
rect 10008 11704 10014 11756
rect 10042 11704 10048 11756
rect 10100 11744 10106 11756
rect 10870 11744 10876 11756
rect 10100 11716 10876 11744
rect 10100 11704 10106 11716
rect 10870 11704 10876 11716
rect 10928 11704 10934 11756
rect 11057 11747 11115 11753
rect 11057 11713 11069 11747
rect 11103 11713 11115 11747
rect 11238 11744 11244 11756
rect 11199 11716 11244 11744
rect 11057 11707 11115 11713
rect 10686 11676 10692 11688
rect 9456 11648 9628 11676
rect 10647 11648 10692 11676
rect 9456 11636 9462 11648
rect 10686 11636 10692 11648
rect 10744 11636 10750 11688
rect 10778 11636 10784 11688
rect 10836 11676 10842 11688
rect 11072 11676 11100 11707
rect 11238 11704 11244 11716
rect 11296 11704 11302 11756
rect 11330 11704 11336 11756
rect 11388 11744 11394 11756
rect 11388 11716 11433 11744
rect 11388 11704 11394 11716
rect 11514 11704 11520 11756
rect 11572 11744 11578 11756
rect 12069 11747 12127 11753
rect 12069 11744 12081 11747
rect 11572 11716 12081 11744
rect 11572 11704 11578 11716
rect 12069 11713 12081 11716
rect 12115 11713 12127 11747
rect 12069 11707 12127 11713
rect 11790 11676 11796 11688
rect 10836 11648 10881 11676
rect 11072 11648 11796 11676
rect 10836 11636 10842 11648
rect 11790 11636 11796 11648
rect 11848 11636 11854 11688
rect 12158 11676 12164 11688
rect 12119 11648 12164 11676
rect 12158 11636 12164 11648
rect 12216 11636 12222 11688
rect 12253 11679 12311 11685
rect 12253 11645 12265 11679
rect 12299 11645 12311 11679
rect 12253 11639 12311 11645
rect 9214 11608 9220 11620
rect 8680 11580 9220 11608
rect 8481 11571 8539 11577
rect 9214 11568 9220 11580
rect 9272 11568 9278 11620
rect 2958 11500 2964 11552
rect 3016 11540 3022 11552
rect 3605 11543 3663 11549
rect 3605 11540 3617 11543
rect 3016 11512 3617 11540
rect 3016 11500 3022 11512
rect 3605 11509 3617 11512
rect 3651 11540 3663 11543
rect 4062 11540 4068 11552
rect 3651 11512 4068 11540
rect 3651 11509 3663 11512
rect 3605 11503 3663 11509
rect 4062 11500 4068 11512
rect 4120 11500 4126 11552
rect 4338 11500 4344 11552
rect 4396 11540 4402 11552
rect 4433 11543 4491 11549
rect 4433 11540 4445 11543
rect 4396 11512 4445 11540
rect 4396 11500 4402 11512
rect 4433 11509 4445 11512
rect 4479 11509 4491 11543
rect 4433 11503 4491 11509
rect 4522 11500 4528 11552
rect 4580 11540 4586 11552
rect 4709 11543 4767 11549
rect 4709 11540 4721 11543
rect 4580 11512 4721 11540
rect 4580 11500 4586 11512
rect 4709 11509 4721 11512
rect 4755 11509 4767 11543
rect 4709 11503 4767 11509
rect 8754 11500 8760 11552
rect 8812 11540 8818 11552
rect 8849 11543 8907 11549
rect 8849 11540 8861 11543
rect 8812 11512 8861 11540
rect 8812 11500 8818 11512
rect 8849 11509 8861 11512
rect 8895 11509 8907 11543
rect 9674 11540 9680 11552
rect 9635 11512 9680 11540
rect 8849 11503 8907 11509
rect 9674 11500 9680 11512
rect 9732 11500 9738 11552
rect 11606 11500 11612 11552
rect 11664 11540 11670 11552
rect 11701 11543 11759 11549
rect 11701 11540 11713 11543
rect 11664 11512 11713 11540
rect 11664 11500 11670 11512
rect 11701 11509 11713 11512
rect 11747 11509 11759 11543
rect 12268 11540 12296 11639
rect 12342 11636 12348 11688
rect 12400 11676 12406 11688
rect 12529 11679 12587 11685
rect 12529 11676 12541 11679
rect 12400 11648 12541 11676
rect 12400 11636 12406 11648
rect 12529 11645 12541 11648
rect 12575 11645 12587 11679
rect 12529 11639 12587 11645
rect 12894 11540 12900 11552
rect 12268 11512 12900 11540
rect 11701 11503 11759 11509
rect 12894 11500 12900 11512
rect 12952 11500 12958 11552
rect 1104 11450 14812 11472
rect 1104 11398 3248 11450
rect 3300 11398 3312 11450
rect 3364 11398 3376 11450
rect 3428 11398 3440 11450
rect 3492 11398 3504 11450
rect 3556 11398 7846 11450
rect 7898 11398 7910 11450
rect 7962 11398 7974 11450
rect 8026 11398 8038 11450
rect 8090 11398 8102 11450
rect 8154 11398 12443 11450
rect 12495 11398 12507 11450
rect 12559 11398 12571 11450
rect 12623 11398 12635 11450
rect 12687 11398 12699 11450
rect 12751 11398 14812 11450
rect 1104 11376 14812 11398
rect 3602 11336 3608 11348
rect 3563 11308 3608 11336
rect 3602 11296 3608 11308
rect 3660 11296 3666 11348
rect 3973 11339 4031 11345
rect 3973 11305 3985 11339
rect 4019 11336 4031 11339
rect 4387 11339 4445 11345
rect 4387 11336 4399 11339
rect 4019 11308 4399 11336
rect 4019 11305 4031 11308
rect 3973 11299 4031 11305
rect 4387 11305 4399 11308
rect 4433 11336 4445 11339
rect 4614 11336 4620 11348
rect 4433 11308 4620 11336
rect 4433 11305 4445 11308
rect 4387 11299 4445 11305
rect 4614 11296 4620 11308
rect 4672 11296 4678 11348
rect 6454 11296 6460 11348
rect 6512 11336 6518 11348
rect 8711 11339 8769 11345
rect 6512 11308 8432 11336
rect 6512 11296 6518 11308
rect 3881 11271 3939 11277
rect 3881 11268 3893 11271
rect 3252 11240 3893 11268
rect 2133 11203 2191 11209
rect 2133 11169 2145 11203
rect 2179 11200 2191 11203
rect 3252 11200 3280 11240
rect 3881 11237 3893 11240
rect 3927 11237 3939 11271
rect 3881 11231 3939 11237
rect 4062 11228 4068 11280
rect 4120 11268 4126 11280
rect 5997 11271 6055 11277
rect 5997 11268 6009 11271
rect 4120 11240 6009 11268
rect 4120 11228 4126 11240
rect 5997 11237 6009 11240
rect 6043 11268 6055 11271
rect 6178 11268 6184 11280
rect 6043 11240 6184 11268
rect 6043 11237 6055 11240
rect 5997 11231 6055 11237
rect 6178 11228 6184 11240
rect 6236 11228 6242 11280
rect 6365 11271 6423 11277
rect 6365 11237 6377 11271
rect 6411 11268 6423 11271
rect 6822 11268 6828 11280
rect 6411 11240 6828 11268
rect 6411 11237 6423 11240
rect 6365 11231 6423 11237
rect 6822 11228 6828 11240
rect 6880 11228 6886 11280
rect 2179 11172 3280 11200
rect 3789 11203 3847 11209
rect 2179 11169 2191 11172
rect 2133 11163 2191 11169
rect 3789 11169 3801 11203
rect 3835 11200 3847 11203
rect 4522 11200 4528 11212
rect 3835 11172 4528 11200
rect 3835 11169 3847 11172
rect 3789 11163 3847 11169
rect 4522 11160 4528 11172
rect 4580 11160 4586 11212
rect 5258 11160 5264 11212
rect 5316 11200 5322 11212
rect 5721 11203 5779 11209
rect 5721 11200 5733 11203
rect 5316 11172 5733 11200
rect 5316 11160 5322 11172
rect 5721 11169 5733 11172
rect 5767 11200 5779 11203
rect 5810 11200 5816 11212
rect 5767 11172 5816 11200
rect 5767 11169 5779 11172
rect 5721 11163 5779 11169
rect 5810 11160 5816 11172
rect 5868 11160 5874 11212
rect 6914 11200 6920 11212
rect 6875 11172 6920 11200
rect 6914 11160 6920 11172
rect 6972 11160 6978 11212
rect 7285 11203 7343 11209
rect 7285 11169 7297 11203
rect 7331 11200 7343 11203
rect 8294 11200 8300 11212
rect 7331 11172 8300 11200
rect 7331 11169 7343 11172
rect 7285 11163 7343 11169
rect 8294 11160 8300 11172
rect 8352 11160 8358 11212
rect 8404 11200 8432 11308
rect 8711 11305 8723 11339
rect 8757 11336 8769 11339
rect 8846 11336 8852 11348
rect 8757 11308 8852 11336
rect 8757 11305 8769 11308
rect 8711 11299 8769 11305
rect 8846 11296 8852 11308
rect 8904 11336 8910 11348
rect 9398 11336 9404 11348
rect 8904 11308 9404 11336
rect 8904 11296 8910 11308
rect 9398 11296 9404 11308
rect 9456 11296 9462 11348
rect 9493 11339 9551 11345
rect 9493 11305 9505 11339
rect 9539 11336 9551 11339
rect 9674 11336 9680 11348
rect 9539 11308 9680 11336
rect 9539 11305 9551 11308
rect 9493 11299 9551 11305
rect 8570 11228 8576 11280
rect 8628 11268 8634 11280
rect 9306 11268 9312 11280
rect 8628 11240 9312 11268
rect 8628 11228 8634 11240
rect 9306 11228 9312 11240
rect 9364 11228 9370 11280
rect 8662 11200 8668 11212
rect 8404 11172 8668 11200
rect 8662 11160 8668 11172
rect 8720 11200 8726 11212
rect 8938 11200 8944 11212
rect 8720 11172 8944 11200
rect 8720 11160 8726 11172
rect 8938 11160 8944 11172
rect 8996 11160 9002 11212
rect 9508 11200 9536 11299
rect 9674 11296 9680 11308
rect 9732 11296 9738 11348
rect 10686 11296 10692 11348
rect 10744 11336 10750 11348
rect 11149 11339 11207 11345
rect 11149 11336 11161 11339
rect 10744 11308 11161 11336
rect 10744 11296 10750 11308
rect 11149 11305 11161 11308
rect 11195 11305 11207 11339
rect 11149 11299 11207 11305
rect 11238 11296 11244 11348
rect 11296 11336 11302 11348
rect 14185 11339 14243 11345
rect 14185 11336 14197 11339
rect 11296 11308 14197 11336
rect 11296 11296 11302 11308
rect 14185 11305 14197 11308
rect 14231 11305 14243 11339
rect 14185 11299 14243 11305
rect 10962 11268 10968 11280
rect 9140 11172 9536 11200
rect 9784 11240 10968 11268
rect 1854 11132 1860 11144
rect 1815 11104 1860 11132
rect 1854 11092 1860 11104
rect 1912 11092 1918 11144
rect 4065 11135 4123 11141
rect 4065 11101 4077 11135
rect 4111 11101 4123 11135
rect 4065 11095 4123 11101
rect 4157 11135 4215 11141
rect 4157 11101 4169 11135
rect 4203 11132 4215 11135
rect 4246 11132 4252 11144
rect 4203 11104 4252 11132
rect 4203 11101 4215 11104
rect 4157 11095 4215 11101
rect 4080 11064 4108 11095
rect 4246 11092 4252 11104
rect 4304 11092 4310 11144
rect 5902 11092 5908 11144
rect 5960 11132 5966 11144
rect 6181 11135 6239 11141
rect 6181 11132 6193 11135
rect 5960 11104 6193 11132
rect 5960 11092 5966 11104
rect 6181 11101 6193 11104
rect 6227 11101 6239 11135
rect 6181 11095 6239 11101
rect 6825 11135 6883 11141
rect 6825 11101 6837 11135
rect 6871 11132 6883 11135
rect 6932 11132 6960 11160
rect 9140 11141 9168 11172
rect 9784 11141 9812 11240
rect 10962 11228 10968 11240
rect 11020 11228 11026 11280
rect 11057 11271 11115 11277
rect 11057 11237 11069 11271
rect 11103 11268 11115 11271
rect 11514 11268 11520 11280
rect 11103 11240 11520 11268
rect 11103 11237 11115 11240
rect 11057 11231 11115 11237
rect 11514 11228 11520 11240
rect 11572 11228 11578 11280
rect 9858 11160 9864 11212
rect 9916 11200 9922 11212
rect 10597 11203 10655 11209
rect 10597 11200 10609 11203
rect 9916 11172 10609 11200
rect 9916 11160 9922 11172
rect 10597 11169 10609 11172
rect 10643 11169 10655 11203
rect 11698 11200 11704 11212
rect 11659 11172 11704 11200
rect 10597 11163 10655 11169
rect 11698 11160 11704 11172
rect 11756 11160 11762 11212
rect 12437 11203 12495 11209
rect 12437 11169 12449 11203
rect 12483 11200 12495 11203
rect 15381 11203 15439 11209
rect 15381 11200 15393 11203
rect 12483 11172 15393 11200
rect 12483 11169 12495 11172
rect 12437 11163 12495 11169
rect 15381 11169 15393 11172
rect 15427 11169 15439 11203
rect 15381 11163 15439 11169
rect 6871 11104 6960 11132
rect 9129 11135 9187 11141
rect 6871 11101 6883 11104
rect 6825 11095 6883 11101
rect 9129 11101 9141 11135
rect 9175 11101 9187 11135
rect 9309 11135 9367 11141
rect 9129 11095 9187 11101
rect 9217 11113 9275 11119
rect 9217 11079 9229 11113
rect 9263 11079 9275 11113
rect 9309 11101 9321 11135
rect 9355 11132 9367 11135
rect 9769 11135 9827 11141
rect 9769 11132 9781 11135
rect 9355 11104 9781 11132
rect 9355 11101 9367 11104
rect 9309 11095 9367 11101
rect 9769 11101 9781 11104
rect 9815 11101 9827 11135
rect 9769 11095 9827 11101
rect 9950 11092 9956 11144
rect 10008 11132 10014 11144
rect 10413 11135 10471 11141
rect 10413 11132 10425 11135
rect 10008 11104 10425 11132
rect 10008 11092 10014 11104
rect 10413 11101 10425 11104
rect 10459 11132 10471 11135
rect 10689 11135 10747 11141
rect 10459 11104 10640 11132
rect 10459 11101 10471 11104
rect 10413 11095 10471 11101
rect 9217 11076 9275 11079
rect 10612 11076 10640 11104
rect 10689 11101 10701 11135
rect 10735 11132 10747 11135
rect 11146 11132 11152 11144
rect 10735 11104 11152 11132
rect 10735 11101 10747 11104
rect 10689 11095 10747 11101
rect 11146 11092 11152 11104
rect 11204 11092 11210 11144
rect 11517 11135 11575 11141
rect 11517 11101 11529 11135
rect 11563 11132 11575 11135
rect 11606 11132 11612 11144
rect 11563 11104 11612 11132
rect 11563 11101 11575 11104
rect 11517 11095 11575 11101
rect 11606 11092 11612 11104
rect 11664 11092 11670 11144
rect 12066 11132 12072 11144
rect 12027 11104 12072 11132
rect 12066 11092 12072 11104
rect 12124 11132 12130 11144
rect 12342 11132 12348 11144
rect 12124 11104 12348 11132
rect 12124 11092 12130 11104
rect 12342 11092 12348 11104
rect 12400 11092 12406 11144
rect 13814 11092 13820 11144
rect 13872 11132 13878 11144
rect 14093 11135 14151 11141
rect 14093 11132 14105 11135
rect 13872 11104 14105 11132
rect 13872 11092 13878 11104
rect 14093 11101 14105 11104
rect 14139 11101 14151 11135
rect 14093 11095 14151 11101
rect 4338 11064 4344 11076
rect 2976 11008 3004 11050
rect 4080 11036 4344 11064
rect 4338 11024 4344 11036
rect 4396 11064 4402 11076
rect 5445 11067 5503 11073
rect 5445 11064 5457 11067
rect 4396 11036 5457 11064
rect 4396 11024 4402 11036
rect 5445 11033 5457 11036
rect 5491 11033 5503 11067
rect 5445 11027 5503 11033
rect 5534 11024 5540 11076
rect 5592 11064 5598 11076
rect 6270 11064 6276 11076
rect 5592 11036 5637 11064
rect 6231 11036 6276 11064
rect 5592 11024 5598 11036
rect 6270 11024 6276 11036
rect 6328 11024 6334 11076
rect 6457 11067 6515 11073
rect 6457 11033 6469 11067
rect 6503 11064 6515 11067
rect 6638 11064 6644 11076
rect 6503 11036 6644 11064
rect 6503 11033 6515 11036
rect 6457 11027 6515 11033
rect 6638 11024 6644 11036
rect 6696 11024 6702 11076
rect 7650 11024 7656 11076
rect 7708 11024 7714 11076
rect 9214 11024 9220 11076
rect 9272 11024 9278 11076
rect 10134 11064 10140 11076
rect 10095 11036 10140 11064
rect 10134 11024 10140 11036
rect 10192 11024 10198 11076
rect 10226 11024 10232 11076
rect 10284 11064 10290 11076
rect 10321 11067 10379 11073
rect 10321 11064 10333 11067
rect 10284 11036 10333 11064
rect 10284 11024 10290 11036
rect 10321 11033 10333 11036
rect 10367 11033 10379 11067
rect 10321 11027 10379 11033
rect 10594 11024 10600 11076
rect 10652 11024 10658 11076
rect 13354 11024 13360 11076
rect 13412 11024 13418 11076
rect 2958 10956 2964 11008
rect 3016 10956 3022 11008
rect 5074 10996 5080 11008
rect 5035 10968 5080 10996
rect 5074 10956 5080 10968
rect 5132 10956 5138 11008
rect 6546 10956 6552 11008
rect 6604 10996 6610 11008
rect 6733 10999 6791 11005
rect 6733 10996 6745 10999
rect 6604 10968 6745 10996
rect 6604 10956 6610 10968
rect 6733 10965 6745 10968
rect 6779 10965 6791 10999
rect 7668 10996 7696 11024
rect 8570 10996 8576 11008
rect 7668 10968 8576 10996
rect 6733 10959 6791 10965
rect 8570 10956 8576 10968
rect 8628 10956 8634 11008
rect 8938 10996 8944 11008
rect 8899 10968 8944 10996
rect 8938 10956 8944 10968
rect 8996 10956 9002 11008
rect 9677 10999 9735 11005
rect 9677 10965 9689 10999
rect 9723 10996 9735 10999
rect 9766 10996 9772 11008
rect 9723 10968 9772 10996
rect 9723 10965 9735 10968
rect 9677 10959 9735 10965
rect 9766 10956 9772 10968
rect 9824 10956 9830 11008
rect 10413 10999 10471 11005
rect 10413 10965 10425 10999
rect 10459 10996 10471 10999
rect 10502 10996 10508 11008
rect 10459 10968 10508 10996
rect 10459 10965 10471 10968
rect 10413 10959 10471 10965
rect 10502 10956 10508 10968
rect 10560 10956 10566 11008
rect 11054 10956 11060 11008
rect 11112 10996 11118 11008
rect 11609 10999 11667 11005
rect 11609 10996 11621 10999
rect 11112 10968 11621 10996
rect 11112 10956 11118 10968
rect 11609 10965 11621 10968
rect 11655 10996 11667 10999
rect 12158 10996 12164 11008
rect 11655 10968 12164 10996
rect 11655 10965 11667 10968
rect 11609 10959 11667 10965
rect 12158 10956 12164 10968
rect 12216 10956 12222 11008
rect 13863 10999 13921 11005
rect 13863 10965 13875 10999
rect 13909 10996 13921 10999
rect 14090 10996 14096 11008
rect 13909 10968 14096 10996
rect 13909 10965 13921 10968
rect 13863 10959 13921 10965
rect 14090 10956 14096 10968
rect 14148 10956 14154 11008
rect 14461 10999 14519 11005
rect 14461 10965 14473 10999
rect 14507 10996 14519 10999
rect 15013 10999 15071 11005
rect 15013 10996 15025 10999
rect 14507 10968 15025 10996
rect 14507 10965 14519 10968
rect 14461 10959 14519 10965
rect 15013 10965 15025 10968
rect 15059 10965 15071 10999
rect 15013 10959 15071 10965
rect 1104 10906 14812 10928
rect 1104 10854 5547 10906
rect 5599 10854 5611 10906
rect 5663 10854 5675 10906
rect 5727 10854 5739 10906
rect 5791 10854 5803 10906
rect 5855 10854 10144 10906
rect 10196 10854 10208 10906
rect 10260 10854 10272 10906
rect 10324 10854 10336 10906
rect 10388 10854 10400 10906
rect 10452 10854 14812 10906
rect 1104 10832 14812 10854
rect 15010 10820 15016 10872
rect 15068 10860 15074 10872
rect 15197 10863 15255 10869
rect 15197 10860 15209 10863
rect 15068 10832 15209 10860
rect 15068 10820 15074 10832
rect 15197 10829 15209 10832
rect 15243 10829 15255 10863
rect 15197 10823 15255 10829
rect 4246 10792 4252 10804
rect 4207 10764 4252 10792
rect 4246 10752 4252 10764
rect 4304 10752 4310 10804
rect 4341 10795 4399 10801
rect 4341 10761 4353 10795
rect 4387 10792 4399 10795
rect 4614 10792 4620 10804
rect 4387 10764 4620 10792
rect 4387 10761 4399 10764
rect 4341 10755 4399 10761
rect 4614 10752 4620 10764
rect 4672 10752 4678 10804
rect 4709 10795 4767 10801
rect 4709 10761 4721 10795
rect 4755 10792 4767 10795
rect 5074 10792 5080 10804
rect 4755 10764 5080 10792
rect 4755 10761 4767 10764
rect 4709 10755 4767 10761
rect 5074 10752 5080 10764
rect 5132 10752 5138 10804
rect 5442 10792 5448 10804
rect 5184 10764 5448 10792
rect 3329 10727 3387 10733
rect 3329 10693 3341 10727
rect 3375 10724 3387 10727
rect 3878 10724 3884 10736
rect 3375 10696 3884 10724
rect 3375 10693 3387 10696
rect 3329 10687 3387 10693
rect 3878 10684 3884 10696
rect 3936 10684 3942 10736
rect 4522 10724 4528 10736
rect 4080 10696 4528 10724
rect 1673 10659 1731 10665
rect 1673 10625 1685 10659
rect 1719 10656 1731 10659
rect 1854 10656 1860 10668
rect 1719 10628 1860 10656
rect 1719 10625 1731 10628
rect 1673 10619 1731 10625
rect 1854 10616 1860 10628
rect 1912 10656 1918 10668
rect 3510 10656 3516 10668
rect 1912 10628 2774 10656
rect 3471 10628 3516 10656
rect 1912 10616 1918 10628
rect 2746 10520 2774 10628
rect 3510 10616 3516 10628
rect 3568 10616 3574 10668
rect 3694 10656 3700 10668
rect 3655 10628 3700 10656
rect 3694 10616 3700 10628
rect 3752 10616 3758 10668
rect 3786 10616 3792 10668
rect 3844 10656 3850 10668
rect 4080 10665 4108 10696
rect 4522 10684 4528 10696
rect 4580 10684 4586 10736
rect 4801 10727 4859 10733
rect 4801 10693 4813 10727
rect 4847 10724 4859 10727
rect 4982 10724 4988 10736
rect 4847 10696 4988 10724
rect 4847 10693 4859 10696
rect 4801 10687 4859 10693
rect 4982 10684 4988 10696
rect 5040 10724 5046 10736
rect 5184 10724 5212 10764
rect 5442 10752 5448 10764
rect 5500 10752 5506 10804
rect 5629 10795 5687 10801
rect 5629 10761 5641 10795
rect 5675 10792 5687 10795
rect 5902 10792 5908 10804
rect 5675 10764 5908 10792
rect 5675 10761 5687 10764
rect 5629 10755 5687 10761
rect 5902 10752 5908 10764
rect 5960 10752 5966 10804
rect 5997 10795 6055 10801
rect 5997 10761 6009 10795
rect 6043 10792 6055 10795
rect 6270 10792 6276 10804
rect 6043 10764 6276 10792
rect 6043 10761 6055 10764
rect 5997 10755 6055 10761
rect 6270 10752 6276 10764
rect 6328 10752 6334 10804
rect 7650 10792 7656 10804
rect 6380 10764 7656 10792
rect 5040 10696 5212 10724
rect 5040 10684 5046 10696
rect 5258 10684 5264 10736
rect 5316 10724 5322 10736
rect 5353 10727 5411 10733
rect 5353 10724 5365 10727
rect 5316 10696 5365 10724
rect 5316 10684 5322 10696
rect 5353 10693 5365 10696
rect 5399 10693 5411 10727
rect 5353 10687 5411 10693
rect 5460 10696 5948 10724
rect 3973 10659 4031 10665
rect 3844 10628 3889 10656
rect 3844 10616 3850 10628
rect 3973 10625 3985 10659
rect 4019 10625 4031 10659
rect 3973 10619 4031 10625
rect 4065 10659 4123 10665
rect 4065 10625 4077 10659
rect 4111 10625 4123 10659
rect 4065 10619 4123 10625
rect 4249 10659 4307 10665
rect 4249 10625 4261 10659
rect 4295 10656 4307 10659
rect 5166 10656 5172 10668
rect 4295 10628 5172 10656
rect 4295 10625 4307 10628
rect 4249 10619 4307 10625
rect 3988 10588 4016 10619
rect 5166 10616 5172 10628
rect 5224 10656 5230 10668
rect 5460 10656 5488 10696
rect 5224 10628 5488 10656
rect 5537 10659 5595 10665
rect 5224 10616 5230 10628
rect 5537 10625 5549 10659
rect 5583 10625 5595 10659
rect 5537 10619 5595 10625
rect 3896 10560 4016 10588
rect 3142 10520 3148 10532
rect 2746 10492 3148 10520
rect 3142 10480 3148 10492
rect 3200 10480 3206 10532
rect 3896 10520 3924 10560
rect 4890 10548 4896 10600
rect 4948 10588 4954 10600
rect 4948 10560 5120 10588
rect 4948 10548 4954 10560
rect 3528 10492 3924 10520
rect 3973 10523 4031 10529
rect 1394 10412 1400 10464
rect 1452 10452 1458 10464
rect 1581 10455 1639 10461
rect 1581 10452 1593 10455
rect 1452 10424 1593 10452
rect 1452 10412 1458 10424
rect 1581 10421 1593 10424
rect 1627 10421 1639 10455
rect 1581 10415 1639 10421
rect 3050 10412 3056 10464
rect 3108 10452 3114 10464
rect 3528 10452 3556 10492
rect 3973 10489 3985 10523
rect 4019 10520 4031 10523
rect 4982 10520 4988 10532
rect 4019 10492 4988 10520
rect 4019 10489 4031 10492
rect 3973 10483 4031 10489
rect 4982 10480 4988 10492
rect 5040 10480 5046 10532
rect 3108 10424 3556 10452
rect 3605 10455 3663 10461
rect 3108 10412 3114 10424
rect 3605 10421 3617 10455
rect 3651 10452 3663 10455
rect 3878 10452 3884 10464
rect 3651 10424 3884 10452
rect 3651 10421 3663 10424
rect 3605 10415 3663 10421
rect 3878 10412 3884 10424
rect 3936 10412 3942 10464
rect 4430 10412 4436 10464
rect 4488 10452 4494 10464
rect 5092 10452 5120 10560
rect 5552 10520 5580 10619
rect 5626 10616 5632 10668
rect 5684 10656 5690 10668
rect 5810 10665 5816 10668
rect 5767 10659 5816 10665
rect 5684 10628 5729 10656
rect 5684 10616 5690 10628
rect 5767 10625 5779 10659
rect 5813 10625 5816 10659
rect 5767 10619 5816 10625
rect 5810 10616 5816 10619
rect 5868 10616 5874 10668
rect 5920 10665 5948 10696
rect 6178 10684 6184 10736
rect 6236 10724 6242 10736
rect 6380 10733 6408 10764
rect 6365 10727 6423 10733
rect 6365 10724 6377 10727
rect 6236 10696 6377 10724
rect 6236 10684 6242 10696
rect 6365 10693 6377 10696
rect 6411 10693 6423 10727
rect 7300 10710 7328 10764
rect 7650 10752 7656 10764
rect 7708 10752 7714 10804
rect 8294 10752 8300 10804
rect 8352 10792 8358 10804
rect 8941 10795 8999 10801
rect 8941 10792 8953 10795
rect 8352 10764 8953 10792
rect 8352 10752 8358 10764
rect 8941 10761 8953 10764
rect 8987 10761 8999 10795
rect 9766 10792 9772 10804
rect 8941 10755 8999 10761
rect 9232 10764 9772 10792
rect 6365 10687 6423 10693
rect 8386 10684 8392 10736
rect 8444 10724 8450 10736
rect 9232 10733 9260 10764
rect 9766 10752 9772 10764
rect 9824 10752 9830 10804
rect 10686 10752 10692 10804
rect 10744 10792 10750 10804
rect 11287 10795 11345 10801
rect 11287 10792 11299 10795
rect 10744 10764 11299 10792
rect 10744 10752 10750 10764
rect 11287 10761 11299 10764
rect 11333 10792 11345 10795
rect 13814 10792 13820 10804
rect 11333 10764 13820 10792
rect 11333 10761 11345 10764
rect 11287 10755 11345 10761
rect 13814 10752 13820 10764
rect 13872 10752 13878 10804
rect 9217 10727 9275 10733
rect 8444 10696 9076 10724
rect 8444 10684 8450 10696
rect 5905 10659 5963 10665
rect 5905 10625 5917 10659
rect 5951 10625 5963 10659
rect 6546 10656 6552 10668
rect 6507 10628 6552 10656
rect 5905 10619 5963 10625
rect 6546 10616 6552 10628
rect 6604 10616 6610 10668
rect 6914 10656 6920 10668
rect 6875 10628 6920 10656
rect 6914 10616 6920 10628
rect 6972 10616 6978 10668
rect 8570 10656 8576 10668
rect 8531 10628 8576 10656
rect 8570 10616 8576 10628
rect 8628 10616 8634 10668
rect 8938 10656 8944 10668
rect 8899 10628 8944 10656
rect 8938 10616 8944 10628
rect 8996 10616 9002 10668
rect 9048 10665 9076 10696
rect 9217 10693 9229 10727
rect 9263 10693 9275 10727
rect 9217 10687 9275 10693
rect 9324 10696 9628 10724
rect 9033 10659 9091 10665
rect 9033 10625 9045 10659
rect 9079 10656 9091 10659
rect 9324 10656 9352 10696
rect 9490 10656 9496 10668
rect 9079 10628 9352 10656
rect 9451 10628 9496 10656
rect 9079 10625 9091 10628
rect 9033 10619 9091 10625
rect 9490 10616 9496 10628
rect 9548 10616 9554 10668
rect 9600 10656 9628 10696
rect 10226 10684 10232 10736
rect 10284 10684 10290 10736
rect 12345 10727 12403 10733
rect 12345 10724 12357 10727
rect 11808 10696 12357 10724
rect 9950 10656 9956 10668
rect 9600 10628 9956 10656
rect 9950 10616 9956 10628
rect 10008 10616 10014 10668
rect 5736 10560 6224 10588
rect 5736 10520 5764 10560
rect 5552 10492 5764 10520
rect 6196 10464 6224 10560
rect 8662 10548 8668 10600
rect 8720 10548 8726 10600
rect 8757 10591 8815 10597
rect 8757 10557 8769 10591
rect 8803 10588 8815 10591
rect 9508 10588 9536 10616
rect 8803 10560 9536 10588
rect 9861 10591 9919 10597
rect 8803 10557 8815 10560
rect 8757 10551 8815 10557
rect 9861 10557 9873 10591
rect 9907 10588 9919 10591
rect 10962 10588 10968 10600
rect 9907 10560 10968 10588
rect 9907 10557 9919 10560
rect 9861 10551 9919 10557
rect 10962 10548 10968 10560
rect 11020 10548 11026 10600
rect 11808 10588 11836 10696
rect 12345 10693 12357 10696
rect 12391 10693 12403 10727
rect 12345 10687 12403 10693
rect 13354 10684 13360 10736
rect 13412 10684 13418 10736
rect 11885 10659 11943 10665
rect 11885 10625 11897 10659
rect 11931 10656 11943 10659
rect 12158 10656 12164 10668
rect 11931 10628 12164 10656
rect 11931 10625 11943 10628
rect 11885 10619 11943 10625
rect 12158 10616 12164 10628
rect 12216 10616 12222 10668
rect 12250 10616 12256 10668
rect 12308 10656 12314 10668
rect 13372 10656 13400 10684
rect 14090 10656 14096 10668
rect 12308 10628 13400 10656
rect 14051 10628 14096 10656
rect 12308 10616 12314 10628
rect 14090 10616 14096 10628
rect 14148 10616 14154 10668
rect 11977 10591 12035 10597
rect 11977 10588 11989 10591
rect 11256 10560 11989 10588
rect 8680 10520 8708 10548
rect 8680 10492 9536 10520
rect 5442 10452 5448 10464
rect 4488 10424 5448 10452
rect 4488 10412 4494 10424
rect 5442 10412 5448 10424
rect 5500 10412 5506 10464
rect 6178 10452 6184 10464
rect 6139 10424 6184 10452
rect 6178 10412 6184 10424
rect 6236 10412 6242 10464
rect 8343 10455 8401 10461
rect 8343 10421 8355 10455
rect 8389 10452 8401 10455
rect 8662 10452 8668 10464
rect 8389 10424 8668 10452
rect 8389 10421 8401 10424
rect 8343 10415 8401 10421
rect 8662 10412 8668 10424
rect 8720 10412 8726 10464
rect 9306 10452 9312 10464
rect 9267 10424 9312 10452
rect 9306 10412 9312 10424
rect 9364 10412 9370 10464
rect 9508 10452 9536 10492
rect 11256 10464 11284 10560
rect 11977 10557 11989 10560
rect 12023 10557 12035 10591
rect 11977 10551 12035 10557
rect 12069 10591 12127 10597
rect 12069 10557 12081 10591
rect 12115 10557 12127 10591
rect 12069 10551 12127 10557
rect 14461 10591 14519 10597
rect 14461 10557 14473 10591
rect 14507 10588 14519 10591
rect 14921 10591 14979 10597
rect 14921 10588 14933 10591
rect 14507 10560 14933 10588
rect 14507 10557 14519 10560
rect 14461 10551 14519 10557
rect 14921 10557 14933 10560
rect 14967 10557 14979 10591
rect 14921 10551 14979 10557
rect 11698 10480 11704 10532
rect 11756 10520 11762 10532
rect 12084 10520 12112 10551
rect 11756 10492 12112 10520
rect 11756 10480 11762 10492
rect 11238 10452 11244 10464
rect 9508 10424 11244 10452
rect 11238 10412 11244 10424
rect 11296 10412 11302 10464
rect 11514 10452 11520 10464
rect 11475 10424 11520 10452
rect 11514 10412 11520 10424
rect 11572 10412 11578 10464
rect 1104 10362 14812 10384
rect 1104 10310 3248 10362
rect 3300 10310 3312 10362
rect 3364 10310 3376 10362
rect 3428 10310 3440 10362
rect 3492 10310 3504 10362
rect 3556 10310 7846 10362
rect 7898 10310 7910 10362
rect 7962 10310 7974 10362
rect 8026 10310 8038 10362
rect 8090 10310 8102 10362
rect 8154 10310 12443 10362
rect 12495 10310 12507 10362
rect 12559 10310 12571 10362
rect 12623 10310 12635 10362
rect 12687 10310 12699 10362
rect 12751 10310 14812 10362
rect 1104 10288 14812 10310
rect 3145 10251 3203 10257
rect 3145 10217 3157 10251
rect 3191 10217 3203 10251
rect 3145 10211 3203 10217
rect 3329 10251 3387 10257
rect 3329 10217 3341 10251
rect 3375 10248 3387 10251
rect 3694 10248 3700 10260
rect 3375 10220 3700 10248
rect 3375 10217 3387 10220
rect 3329 10211 3387 10217
rect 3160 10180 3188 10211
rect 3694 10208 3700 10220
rect 3752 10208 3758 10260
rect 3970 10208 3976 10260
rect 4028 10248 4034 10260
rect 7009 10251 7067 10257
rect 7009 10248 7021 10251
rect 4028 10220 7021 10248
rect 4028 10208 4034 10220
rect 7009 10217 7021 10220
rect 7055 10248 7067 10251
rect 8570 10248 8576 10260
rect 7055 10220 8576 10248
rect 7055 10217 7067 10220
rect 7009 10211 7067 10217
rect 8570 10208 8576 10220
rect 8628 10208 8634 10260
rect 9306 10208 9312 10260
rect 9364 10248 9370 10260
rect 10226 10248 10232 10260
rect 9364 10220 10232 10248
rect 9364 10208 9370 10220
rect 10226 10208 10232 10220
rect 10284 10208 10290 10260
rect 10962 10248 10968 10260
rect 10923 10220 10968 10248
rect 10962 10208 10968 10220
rect 11020 10208 11026 10260
rect 12158 10248 12164 10260
rect 12119 10220 12164 10248
rect 12158 10208 12164 10220
rect 12216 10208 12222 10260
rect 12986 10248 12992 10260
rect 12947 10220 12992 10248
rect 12986 10208 12992 10220
rect 13044 10208 13050 10260
rect 13354 10208 13360 10260
rect 13412 10248 13418 10260
rect 13817 10251 13875 10257
rect 13817 10248 13829 10251
rect 13412 10220 13829 10248
rect 13412 10208 13418 10220
rect 13817 10217 13829 10220
rect 13863 10217 13875 10251
rect 13817 10211 13875 10217
rect 3160 10152 3372 10180
rect 1397 10115 1455 10121
rect 1397 10081 1409 10115
rect 1443 10112 1455 10115
rect 3142 10112 3148 10124
rect 1443 10084 3148 10112
rect 1443 10081 1455 10084
rect 1397 10075 1455 10081
rect 3142 10072 3148 10084
rect 3200 10072 3206 10124
rect 3237 10047 3295 10053
rect 3237 10013 3249 10047
rect 3283 10038 3295 10047
rect 3344 10044 3372 10152
rect 4154 10140 4160 10192
rect 4212 10180 4218 10192
rect 4709 10183 4767 10189
rect 4709 10180 4721 10183
rect 4212 10152 4721 10180
rect 4212 10140 4218 10152
rect 4709 10149 4721 10152
rect 4755 10149 4767 10183
rect 5166 10180 5172 10192
rect 5127 10152 5172 10180
rect 4709 10143 4767 10149
rect 4724 10112 4752 10143
rect 5166 10140 5172 10152
rect 5224 10140 5230 10192
rect 5261 10183 5319 10189
rect 5261 10149 5273 10183
rect 5307 10180 5319 10183
rect 5350 10180 5356 10192
rect 5307 10152 5356 10180
rect 5307 10149 5319 10152
rect 5261 10143 5319 10149
rect 5350 10140 5356 10152
rect 5408 10140 5414 10192
rect 5626 10140 5632 10192
rect 5684 10180 5690 10192
rect 5902 10180 5908 10192
rect 5684 10152 5908 10180
rect 5684 10140 5690 10152
rect 5902 10140 5908 10152
rect 5960 10180 5966 10192
rect 7561 10183 7619 10189
rect 7561 10180 7573 10183
rect 5960 10152 7573 10180
rect 5960 10140 5966 10152
rect 7561 10149 7573 10152
rect 7607 10149 7619 10183
rect 7561 10143 7619 10149
rect 9493 10183 9551 10189
rect 9493 10149 9505 10183
rect 9539 10180 9551 10183
rect 9950 10180 9956 10192
rect 9539 10152 9956 10180
rect 9539 10149 9551 10152
rect 9493 10143 9551 10149
rect 9950 10140 9956 10152
rect 10008 10140 10014 10192
rect 11057 10183 11115 10189
rect 11057 10180 11069 10183
rect 10060 10152 11069 10180
rect 4724 10084 5764 10112
rect 3786 10044 3792 10056
rect 3344 10038 3792 10044
rect 3283 10016 3792 10038
rect 3283 10013 3372 10016
rect 3237 10010 3372 10013
rect 3237 10007 3295 10010
rect 3786 10004 3792 10016
rect 3844 10004 3850 10056
rect 3878 10004 3884 10056
rect 3936 10044 3942 10056
rect 4157 10047 4215 10053
rect 4157 10044 4169 10047
rect 3936 10016 4169 10044
rect 3936 10004 3942 10016
rect 4157 10013 4169 10016
rect 4203 10013 4215 10047
rect 4338 10044 4344 10056
rect 4299 10016 4344 10044
rect 4157 10007 4215 10013
rect 1673 9979 1731 9985
rect 1673 9945 1685 9979
rect 1719 9945 1731 9979
rect 2958 9976 2964 9988
rect 2898 9948 2964 9976
rect 1673 9939 1731 9945
rect 1688 9908 1716 9939
rect 2958 9936 2964 9948
rect 3016 9936 3022 9988
rect 4172 9976 4200 10007
rect 4338 10004 4344 10016
rect 4396 10004 4402 10056
rect 4433 10047 4491 10053
rect 4433 10013 4445 10047
rect 4479 10046 4491 10047
rect 4522 10046 4528 10056
rect 4479 10018 4528 10046
rect 4479 10013 4491 10018
rect 4433 10007 4491 10013
rect 4522 10004 4528 10018
rect 4580 10004 4586 10056
rect 4614 10004 4620 10056
rect 4672 10044 4678 10056
rect 4982 10044 4988 10056
rect 4672 10016 4717 10044
rect 4943 10016 4988 10044
rect 4672 10004 4678 10016
rect 4982 10004 4988 10016
rect 5040 10004 5046 10056
rect 5074 10004 5080 10056
rect 5132 10044 5138 10056
rect 5350 10044 5356 10056
rect 5132 10016 5177 10044
rect 5311 10016 5356 10044
rect 5132 10004 5138 10016
rect 5350 10004 5356 10016
rect 5408 10004 5414 10056
rect 5442 10004 5448 10056
rect 5500 10044 5506 10056
rect 5736 10053 5764 10084
rect 6178 10072 6184 10124
rect 6236 10112 6242 10124
rect 8573 10115 8631 10121
rect 8573 10112 8585 10115
rect 6236 10084 8585 10112
rect 6236 10072 6242 10084
rect 8573 10081 8585 10084
rect 8619 10081 8631 10115
rect 8573 10075 8631 10081
rect 9033 10115 9091 10121
rect 9033 10081 9045 10115
rect 9079 10081 9091 10115
rect 9033 10075 9091 10081
rect 5721 10047 5779 10053
rect 5500 10016 5545 10044
rect 5500 10004 5506 10016
rect 5721 10013 5733 10047
rect 5767 10013 5779 10047
rect 5721 10007 5779 10013
rect 7561 10047 7619 10053
rect 7561 10013 7573 10047
rect 7607 10013 7619 10047
rect 7742 10044 7748 10056
rect 7703 10016 7748 10044
rect 7561 10007 7619 10013
rect 7576 9976 7604 10007
rect 7742 10004 7748 10016
rect 7800 10004 7806 10056
rect 8021 10047 8079 10053
rect 8021 10013 8033 10047
rect 8067 10044 8079 10047
rect 8478 10044 8484 10056
rect 8067 10016 8484 10044
rect 8067 10013 8079 10016
rect 8021 10007 8079 10013
rect 8478 10004 8484 10016
rect 8536 10004 8542 10056
rect 8662 10044 8668 10056
rect 8623 10016 8668 10044
rect 8662 10004 8668 10016
rect 8720 10044 8726 10056
rect 9048 10044 9076 10075
rect 9766 10072 9772 10124
rect 9824 10112 9830 10124
rect 10060 10112 10088 10152
rect 11057 10149 11069 10152
rect 11103 10149 11115 10183
rect 11057 10143 11115 10149
rect 9824 10084 10088 10112
rect 10321 10115 10379 10121
rect 9824 10072 9830 10084
rect 10321 10081 10333 10115
rect 10367 10112 10379 10115
rect 10502 10112 10508 10124
rect 10367 10084 10508 10112
rect 10367 10081 10379 10084
rect 10321 10075 10379 10081
rect 10502 10072 10508 10084
rect 10560 10072 10566 10124
rect 10689 10115 10747 10121
rect 10689 10081 10701 10115
rect 10735 10112 10747 10115
rect 11514 10112 11520 10124
rect 10735 10084 11520 10112
rect 10735 10081 10747 10084
rect 10689 10075 10747 10081
rect 11514 10072 11520 10084
rect 11572 10072 11578 10124
rect 11698 10072 11704 10124
rect 11756 10112 11762 10124
rect 11885 10115 11943 10121
rect 11885 10112 11897 10115
rect 11756 10084 11897 10112
rect 11756 10072 11762 10084
rect 11885 10081 11897 10084
rect 11931 10081 11943 10115
rect 12621 10115 12679 10121
rect 12621 10112 12633 10115
rect 11885 10075 11943 10081
rect 12406 10084 12633 10112
rect 8720 10016 9076 10044
rect 9125 10047 9183 10053
rect 8720 10004 8726 10016
rect 9125 10013 9137 10047
rect 9171 10013 9183 10047
rect 9125 10007 9183 10013
rect 9953 10047 10011 10053
rect 9953 10013 9965 10047
rect 9999 10013 10011 10047
rect 9953 10007 10011 10013
rect 10045 10047 10103 10053
rect 10045 10013 10057 10047
rect 10091 10044 10103 10047
rect 10410 10044 10416 10056
rect 10091 10016 10416 10044
rect 10091 10013 10103 10016
rect 10045 10007 10103 10013
rect 3252 9948 4108 9976
rect 4172 9948 7604 9976
rect 3252 9908 3280 9948
rect 3510 9908 3516 9920
rect 1688 9880 3280 9908
rect 3471 9880 3516 9908
rect 3510 9868 3516 9880
rect 3568 9868 3574 9920
rect 3694 9868 3700 9920
rect 3752 9908 3758 9920
rect 4080 9917 4108 9948
rect 8846 9936 8852 9988
rect 8904 9976 8910 9988
rect 9140 9976 9168 10007
rect 8904 9948 9168 9976
rect 9968 9976 9996 10007
rect 10410 10004 10416 10016
rect 10468 10044 10474 10056
rect 10778 10044 10784 10056
rect 10468 10016 10784 10044
rect 10468 10004 10474 10016
rect 10778 10004 10784 10016
rect 10836 10004 10842 10056
rect 11054 10044 11060 10056
rect 11015 10016 11060 10044
rect 11054 10004 11060 10016
rect 11112 10004 11118 10056
rect 11238 10044 11244 10056
rect 11199 10016 11244 10044
rect 11238 10004 11244 10016
rect 11296 10044 11302 10056
rect 12406 10044 12434 10084
rect 12621 10081 12633 10084
rect 12667 10081 12679 10115
rect 12621 10075 12679 10081
rect 12805 10115 12863 10121
rect 12805 10081 12817 10115
rect 12851 10112 12863 10115
rect 12894 10112 12900 10124
rect 12851 10084 12900 10112
rect 12851 10081 12863 10084
rect 12805 10075 12863 10081
rect 12894 10072 12900 10084
rect 12952 10072 12958 10124
rect 13633 10115 13691 10121
rect 13633 10081 13645 10115
rect 13679 10112 13691 10115
rect 15105 10115 15163 10121
rect 15105 10112 15117 10115
rect 13679 10084 15117 10112
rect 13679 10081 13691 10084
rect 13633 10075 13691 10081
rect 15105 10081 15117 10084
rect 15151 10081 15163 10115
rect 15105 10075 15163 10081
rect 11296 10016 12434 10044
rect 12529 10047 12587 10053
rect 11296 10004 11302 10016
rect 12529 10013 12541 10047
rect 12575 10044 12587 10047
rect 13446 10044 13452 10056
rect 12575 10016 13452 10044
rect 12575 10013 12587 10016
rect 12529 10007 12587 10013
rect 13446 10004 13452 10016
rect 13504 10004 13510 10056
rect 13357 9979 13415 9985
rect 9968 9948 11376 9976
rect 8904 9936 8910 9948
rect 3881 9911 3939 9917
rect 3881 9908 3893 9911
rect 3752 9880 3893 9908
rect 3752 9868 3758 9880
rect 3881 9877 3893 9880
rect 3927 9877 3939 9911
rect 3881 9871 3939 9877
rect 4065 9911 4123 9917
rect 4065 9877 4077 9911
rect 4111 9877 4123 9911
rect 4065 9871 4123 9877
rect 4246 9868 4252 9920
rect 4304 9908 4310 9920
rect 4525 9911 4583 9917
rect 4525 9908 4537 9911
rect 4304 9880 4537 9908
rect 4304 9868 4310 9880
rect 4525 9877 4537 9880
rect 4571 9877 4583 9911
rect 4525 9871 4583 9877
rect 4798 9868 4804 9920
rect 4856 9908 4862 9920
rect 5537 9911 5595 9917
rect 5537 9908 5549 9911
rect 4856 9880 5549 9908
rect 4856 9868 4862 9880
rect 5537 9877 5549 9880
rect 5583 9908 5595 9911
rect 6362 9908 6368 9920
rect 5583 9880 6368 9908
rect 5583 9877 5595 9880
rect 5537 9871 5595 9877
rect 6362 9868 6368 9880
rect 6420 9868 6426 9920
rect 7926 9908 7932 9920
rect 7887 9880 7932 9908
rect 7926 9868 7932 9880
rect 7984 9868 7990 9920
rect 9585 9911 9643 9917
rect 9585 9877 9597 9911
rect 9631 9908 9643 9911
rect 9858 9908 9864 9920
rect 9631 9880 9864 9908
rect 9631 9877 9643 9880
rect 9585 9871 9643 9877
rect 9858 9868 9864 9880
rect 9916 9868 9922 9920
rect 10042 9868 10048 9920
rect 10100 9908 10106 9920
rect 11348 9917 11376 9948
rect 13357 9945 13369 9979
rect 13403 9976 13415 9979
rect 13722 9976 13728 9988
rect 13403 9948 13728 9976
rect 13403 9945 13415 9948
rect 13357 9939 13415 9945
rect 13722 9936 13728 9948
rect 13780 9936 13786 9988
rect 13998 9936 14004 9988
rect 14056 9976 14062 9988
rect 14369 9979 14427 9985
rect 14369 9976 14381 9979
rect 14056 9948 14381 9976
rect 14056 9936 14062 9948
rect 14369 9945 14381 9948
rect 14415 9945 14427 9979
rect 14369 9939 14427 9945
rect 10229 9911 10287 9917
rect 10229 9908 10241 9911
rect 10100 9880 10241 9908
rect 10100 9868 10106 9880
rect 10229 9877 10241 9880
rect 10275 9877 10287 9911
rect 10229 9871 10287 9877
rect 11333 9911 11391 9917
rect 11333 9877 11345 9911
rect 11379 9877 11391 9911
rect 11698 9908 11704 9920
rect 11659 9880 11704 9908
rect 11333 9871 11391 9877
rect 11698 9868 11704 9880
rect 11756 9868 11762 9920
rect 11793 9911 11851 9917
rect 11793 9877 11805 9911
rect 11839 9908 11851 9911
rect 12158 9908 12164 9920
rect 11839 9880 12164 9908
rect 11839 9877 11851 9880
rect 11793 9871 11851 9877
rect 12158 9868 12164 9880
rect 12216 9868 12222 9920
rect 13449 9911 13507 9917
rect 13449 9877 13461 9911
rect 13495 9908 13507 9911
rect 13630 9908 13636 9920
rect 13495 9880 13636 9908
rect 13495 9877 13507 9880
rect 13449 9871 13507 9877
rect 13630 9868 13636 9880
rect 13688 9868 13694 9920
rect 14274 9908 14280 9920
rect 14235 9880 14280 9908
rect 14274 9868 14280 9880
rect 14332 9868 14338 9920
rect 1104 9818 14812 9840
rect 1104 9766 5547 9818
rect 5599 9766 5611 9818
rect 5663 9766 5675 9818
rect 5727 9766 5739 9818
rect 5791 9766 5803 9818
rect 5855 9766 10144 9818
rect 10196 9766 10208 9818
rect 10260 9766 10272 9818
rect 10324 9766 10336 9818
rect 10388 9766 10400 9818
rect 10452 9766 14812 9818
rect 1104 9744 14812 9766
rect 3878 9704 3884 9716
rect 2792 9676 3884 9704
rect 2792 9622 2820 9676
rect 3878 9664 3884 9676
rect 3936 9664 3942 9716
rect 4338 9664 4344 9716
rect 4396 9704 4402 9716
rect 4522 9704 4528 9716
rect 4396 9676 4528 9704
rect 4396 9664 4402 9676
rect 4522 9664 4528 9676
rect 4580 9704 4586 9716
rect 4985 9707 5043 9713
rect 4985 9704 4997 9707
rect 4580 9676 4997 9704
rect 4580 9664 4586 9676
rect 4985 9673 4997 9676
rect 5031 9673 5043 9707
rect 4985 9667 5043 9673
rect 5350 9664 5356 9716
rect 5408 9704 5414 9716
rect 6454 9704 6460 9716
rect 5408 9676 6460 9704
rect 5408 9664 5414 9676
rect 6454 9664 6460 9676
rect 6512 9704 6518 9716
rect 7190 9704 7196 9716
rect 6512 9676 6960 9704
rect 7151 9676 7196 9704
rect 6512 9664 6518 9676
rect 3620 9608 4752 9636
rect 1394 9568 1400 9580
rect 1355 9540 1400 9568
rect 1394 9528 1400 9540
rect 1452 9528 1458 9580
rect 1765 9503 1823 9509
rect 1765 9469 1777 9503
rect 1811 9500 1823 9503
rect 2774 9500 2780 9512
rect 1811 9472 2780 9500
rect 1811 9469 1823 9472
rect 1765 9463 1823 9469
rect 2774 9460 2780 9472
rect 2832 9460 2838 9512
rect 2866 9392 2872 9444
rect 2924 9432 2930 9444
rect 3620 9441 3648 9608
rect 4246 9568 4252 9580
rect 4207 9540 4252 9568
rect 4246 9528 4252 9540
rect 4304 9528 4310 9580
rect 4430 9568 4436 9580
rect 4391 9540 4436 9568
rect 4430 9528 4436 9540
rect 4488 9528 4494 9580
rect 4614 9568 4620 9580
rect 4527 9540 4620 9568
rect 4614 9528 4620 9540
rect 4672 9528 4678 9580
rect 4724 9577 4752 9608
rect 5442 9596 5448 9648
rect 5500 9636 5506 9648
rect 5813 9639 5871 9645
rect 5813 9636 5825 9639
rect 5500 9608 5825 9636
rect 5500 9596 5506 9608
rect 5813 9605 5825 9608
rect 5859 9605 5871 9639
rect 6932 9636 6960 9676
rect 7190 9664 7196 9676
rect 7248 9664 7254 9716
rect 9858 9664 9864 9716
rect 9916 9704 9922 9716
rect 11517 9707 11575 9713
rect 11517 9704 11529 9707
rect 9916 9676 11529 9704
rect 9916 9664 9922 9676
rect 11517 9673 11529 9676
rect 11563 9673 11575 9707
rect 11517 9667 11575 9673
rect 11698 9664 11704 9716
rect 11756 9704 11762 9716
rect 11885 9707 11943 9713
rect 11885 9704 11897 9707
rect 11756 9676 11897 9704
rect 11756 9664 11762 9676
rect 11885 9673 11897 9676
rect 11931 9673 11943 9707
rect 11885 9667 11943 9673
rect 6932 9608 7052 9636
rect 5813 9599 5871 9605
rect 4709 9571 4767 9577
rect 4709 9537 4721 9571
rect 4755 9537 4767 9571
rect 4709 9531 4767 9537
rect 3881 9503 3939 9509
rect 3881 9469 3893 9503
rect 3927 9500 3939 9503
rect 3970 9500 3976 9512
rect 3927 9472 3976 9500
rect 3927 9469 3939 9472
rect 3881 9463 3939 9469
rect 3970 9460 3976 9472
rect 4028 9500 4034 9512
rect 4632 9500 4660 9528
rect 4028 9472 4660 9500
rect 4028 9460 4034 9472
rect 3421 9435 3479 9441
rect 3421 9432 3433 9435
rect 2924 9404 3433 9432
rect 2924 9392 2930 9404
rect 3421 9401 3433 9404
rect 3467 9401 3479 9435
rect 3421 9395 3479 9401
rect 3605 9435 3663 9441
rect 3605 9401 3617 9435
rect 3651 9401 3663 9435
rect 4724 9432 4752 9531
rect 4798 9528 4804 9580
rect 4856 9568 4862 9580
rect 5721 9571 5779 9577
rect 4856 9540 4901 9568
rect 4856 9528 4862 9540
rect 5721 9537 5733 9571
rect 5767 9537 5779 9571
rect 6362 9568 6368 9580
rect 6323 9540 6368 9568
rect 5721 9531 5779 9537
rect 4982 9432 4988 9444
rect 4724 9404 4988 9432
rect 3605 9395 3663 9401
rect 4982 9392 4988 9404
rect 5040 9432 5046 9444
rect 5353 9435 5411 9441
rect 5353 9432 5365 9435
rect 5040 9404 5365 9432
rect 5040 9392 5046 9404
rect 5353 9401 5365 9404
rect 5399 9401 5411 9435
rect 5736 9432 5764 9531
rect 6362 9528 6368 9540
rect 6420 9528 6426 9580
rect 6641 9571 6699 9577
rect 6641 9537 6653 9571
rect 6687 9568 6699 9571
rect 6822 9568 6828 9580
rect 6687 9540 6828 9568
rect 6687 9537 6699 9540
rect 6641 9531 6699 9537
rect 6822 9528 6828 9540
rect 6880 9528 6886 9580
rect 6917 9571 6975 9577
rect 6917 9537 6929 9571
rect 6963 9537 6975 9571
rect 7024 9568 7052 9608
rect 7098 9596 7104 9648
rect 7156 9636 7162 9648
rect 7742 9636 7748 9648
rect 7156 9608 7748 9636
rect 7156 9596 7162 9608
rect 7742 9596 7748 9608
rect 7800 9636 7806 9648
rect 8205 9639 8263 9645
rect 8205 9636 8217 9639
rect 7800 9608 8217 9636
rect 7800 9596 7806 9608
rect 8205 9605 8217 9608
rect 8251 9636 8263 9639
rect 10321 9639 10379 9645
rect 10321 9636 10333 9639
rect 8251 9608 10333 9636
rect 8251 9605 8263 9608
rect 8205 9599 8263 9605
rect 10321 9605 10333 9608
rect 10367 9605 10379 9639
rect 10321 9599 10379 9605
rect 10965 9639 11023 9645
rect 10965 9605 10977 9639
rect 11011 9636 11023 9639
rect 14274 9636 14280 9648
rect 11011 9608 14280 9636
rect 11011 9605 11023 9608
rect 10965 9599 11023 9605
rect 14274 9596 14280 9608
rect 14332 9596 14338 9648
rect 7561 9571 7619 9577
rect 7561 9568 7573 9571
rect 7024 9540 7573 9568
rect 6917 9531 6975 9537
rect 7561 9537 7573 9540
rect 7607 9568 7619 9571
rect 7607 9540 8064 9568
rect 7607 9537 7619 9540
rect 7561 9531 7619 9537
rect 5902 9500 5908 9512
rect 5863 9472 5908 9500
rect 5902 9460 5908 9472
rect 5960 9460 5966 9512
rect 6380 9500 6408 9528
rect 6932 9500 6960 9531
rect 7650 9500 7656 9512
rect 6380 9472 6960 9500
rect 7611 9472 7656 9500
rect 7650 9460 7656 9472
rect 7708 9460 7714 9512
rect 7742 9460 7748 9512
rect 7800 9500 7806 9512
rect 7837 9503 7895 9509
rect 7837 9500 7849 9503
rect 7800 9472 7849 9500
rect 7800 9460 7806 9472
rect 7837 9469 7849 9472
rect 7883 9500 7895 9503
rect 7926 9500 7932 9512
rect 7883 9472 7932 9500
rect 7883 9469 7895 9472
rect 7837 9463 7895 9469
rect 7926 9460 7932 9472
rect 7984 9460 7990 9512
rect 8036 9500 8064 9540
rect 8110 9528 8116 9580
rect 8168 9568 8174 9580
rect 8481 9571 8539 9577
rect 8168 9540 8213 9568
rect 8168 9528 8174 9540
rect 8481 9537 8493 9571
rect 8527 9568 8539 9571
rect 8570 9568 8576 9580
rect 8527 9540 8576 9568
rect 8527 9537 8539 9540
rect 8481 9531 8539 9537
rect 8570 9528 8576 9540
rect 8628 9528 8634 9580
rect 8849 9571 8907 9577
rect 8849 9537 8861 9571
rect 8895 9568 8907 9571
rect 8938 9568 8944 9580
rect 8895 9540 8944 9568
rect 8895 9537 8907 9540
rect 8849 9531 8907 9537
rect 8938 9528 8944 9540
rect 8996 9528 9002 9580
rect 9033 9571 9091 9577
rect 9033 9537 9045 9571
rect 9079 9568 9091 9571
rect 9342 9571 9400 9577
rect 9079 9540 9260 9568
rect 9079 9537 9091 9540
rect 9033 9531 9091 9537
rect 8297 9503 8355 9509
rect 8297 9500 8309 9503
rect 8036 9472 8309 9500
rect 8297 9469 8309 9472
rect 8343 9469 8355 9503
rect 8297 9463 8355 9469
rect 8662 9460 8668 9512
rect 8720 9500 8726 9512
rect 9125 9503 9183 9509
rect 9125 9500 9137 9503
rect 8720 9472 9137 9500
rect 8720 9460 8726 9472
rect 9125 9469 9137 9472
rect 9171 9469 9183 9503
rect 9232 9500 9260 9540
rect 9342 9537 9354 9571
rect 9388 9568 9400 9571
rect 9582 9568 9588 9580
rect 9388 9540 9588 9568
rect 9388 9537 9400 9540
rect 9342 9531 9400 9537
rect 9582 9528 9588 9540
rect 9640 9528 9646 9580
rect 9950 9568 9956 9580
rect 9911 9540 9956 9568
rect 9950 9528 9956 9540
rect 10008 9528 10014 9580
rect 10137 9571 10195 9577
rect 10137 9537 10149 9571
rect 10183 9568 10195 9571
rect 10505 9571 10563 9577
rect 10505 9568 10517 9571
rect 10183 9540 10517 9568
rect 10183 9537 10195 9540
rect 10137 9531 10195 9537
rect 10505 9537 10517 9540
rect 10551 9568 10563 9571
rect 10594 9568 10600 9580
rect 10551 9540 10600 9568
rect 10551 9537 10563 9540
rect 10505 9531 10563 9537
rect 10594 9528 10600 9540
rect 10652 9568 10658 9580
rect 11517 9571 11575 9577
rect 11517 9568 11529 9571
rect 10652 9540 11529 9568
rect 10652 9528 10658 9540
rect 11517 9537 11529 9540
rect 11563 9537 11575 9571
rect 11517 9531 11575 9537
rect 11606 9528 11612 9580
rect 11664 9568 11670 9580
rect 11793 9571 11851 9577
rect 11664 9540 11709 9568
rect 11664 9528 11670 9540
rect 11793 9537 11805 9571
rect 11839 9568 11851 9571
rect 11882 9568 11888 9580
rect 11839 9540 11888 9568
rect 11839 9537 11851 9540
rect 11793 9531 11851 9537
rect 11882 9528 11888 9540
rect 11940 9528 11946 9580
rect 12250 9568 12256 9580
rect 12211 9540 12256 9568
rect 12250 9528 12256 9540
rect 12308 9528 12314 9580
rect 12713 9571 12771 9577
rect 12713 9537 12725 9571
rect 12759 9568 12771 9571
rect 12802 9568 12808 9580
rect 12759 9540 12808 9568
rect 12759 9537 12771 9540
rect 12713 9531 12771 9537
rect 12802 9528 12808 9540
rect 12860 9568 12866 9580
rect 15013 9571 15071 9577
rect 15013 9568 15025 9571
rect 12860 9540 15025 9568
rect 12860 9528 12866 9540
rect 15013 9537 15025 9540
rect 15059 9537 15071 9571
rect 15013 9531 15071 9537
rect 10226 9500 10232 9512
rect 9232 9472 10232 9500
rect 9125 9463 9183 9469
rect 10226 9460 10232 9472
rect 10284 9460 10290 9512
rect 10781 9503 10839 9509
rect 10781 9469 10793 9503
rect 10827 9469 10839 9503
rect 10781 9463 10839 9469
rect 10873 9503 10931 9509
rect 10873 9469 10885 9503
rect 10919 9500 10931 9503
rect 11422 9500 11428 9512
rect 10919 9472 11428 9500
rect 10919 9469 10931 9472
rect 10873 9463 10931 9469
rect 6457 9435 6515 9441
rect 6457 9432 6469 9435
rect 5736 9404 6469 9432
rect 5353 9395 5411 9401
rect 6457 9401 6469 9404
rect 6503 9401 6515 9435
rect 6457 9395 6515 9401
rect 3050 9324 3056 9376
rect 3108 9364 3114 9376
rect 3191 9367 3249 9373
rect 3191 9364 3203 9367
rect 3108 9336 3203 9364
rect 3108 9324 3114 9336
rect 3191 9333 3203 9336
rect 3237 9333 3249 9367
rect 3191 9327 3249 9333
rect 3973 9367 4031 9373
rect 3973 9333 3985 9367
rect 4019 9364 4031 9367
rect 4062 9364 4068 9376
rect 4019 9336 4068 9364
rect 4019 9333 4031 9336
rect 3973 9327 4031 9333
rect 4062 9324 4068 9336
rect 4120 9324 4126 9376
rect 4246 9364 4252 9376
rect 4207 9336 4252 9364
rect 4246 9324 4252 9336
rect 4304 9324 4310 9376
rect 6472 9364 6500 9395
rect 6914 9392 6920 9444
rect 6972 9432 6978 9444
rect 7101 9435 7159 9441
rect 7101 9432 7113 9435
rect 6972 9404 7113 9432
rect 6972 9392 6978 9404
rect 7101 9401 7113 9404
rect 7147 9432 7159 9435
rect 8386 9432 8392 9444
rect 7147 9404 8392 9432
rect 7147 9401 7159 9404
rect 7101 9395 7159 9401
rect 8386 9392 8392 9404
rect 8444 9392 8450 9444
rect 9033 9435 9091 9441
rect 9033 9401 9045 9435
rect 9079 9432 9091 9435
rect 9674 9432 9680 9444
rect 9079 9404 9680 9432
rect 9079 9401 9091 9404
rect 9033 9395 9091 9401
rect 9674 9392 9680 9404
rect 9732 9392 9738 9444
rect 9861 9435 9919 9441
rect 9861 9401 9873 9435
rect 9907 9432 9919 9435
rect 10686 9432 10692 9444
rect 9907 9404 10692 9432
rect 9907 9401 9919 9404
rect 9861 9395 9919 9401
rect 10686 9392 10692 9404
rect 10744 9392 10750 9444
rect 10502 9364 10508 9376
rect 6472 9336 10508 9364
rect 10502 9324 10508 9336
rect 10560 9324 10566 9376
rect 10796 9364 10824 9463
rect 11422 9460 11428 9472
rect 11480 9460 11486 9512
rect 12158 9460 12164 9512
rect 12216 9500 12222 9512
rect 12345 9503 12403 9509
rect 12345 9500 12357 9503
rect 12216 9472 12357 9500
rect 12216 9460 12222 9472
rect 12345 9469 12357 9472
rect 12391 9469 12403 9503
rect 12345 9463 12403 9469
rect 12529 9503 12587 9509
rect 12529 9469 12541 9503
rect 12575 9500 12587 9503
rect 12894 9500 12900 9512
rect 12575 9472 12900 9500
rect 12575 9469 12587 9472
rect 12529 9463 12587 9469
rect 12894 9460 12900 9472
rect 12952 9460 12958 9512
rect 11333 9435 11391 9441
rect 11333 9401 11345 9435
rect 11379 9432 11391 9435
rect 13722 9432 13728 9444
rect 11379 9404 13728 9432
rect 11379 9401 11391 9404
rect 11333 9395 11391 9401
rect 13722 9392 13728 9404
rect 13780 9392 13786 9444
rect 12342 9364 12348 9376
rect 10796 9336 12348 9364
rect 12342 9324 12348 9336
rect 12400 9324 12406 9376
rect 13998 9364 14004 9376
rect 13959 9336 14004 9364
rect 13998 9324 14004 9336
rect 14056 9324 14062 9376
rect 1104 9274 14812 9296
rect 1104 9222 3248 9274
rect 3300 9222 3312 9274
rect 3364 9222 3376 9274
rect 3428 9222 3440 9274
rect 3492 9222 3504 9274
rect 3556 9222 7846 9274
rect 7898 9222 7910 9274
rect 7962 9222 7974 9274
rect 8026 9222 8038 9274
rect 8090 9222 8102 9274
rect 8154 9222 12443 9274
rect 12495 9222 12507 9274
rect 12559 9222 12571 9274
rect 12623 9222 12635 9274
rect 12687 9222 12699 9274
rect 12751 9222 14812 9274
rect 1104 9200 14812 9222
rect 2774 9120 2780 9172
rect 2832 9160 2838 9172
rect 3237 9163 3295 9169
rect 2832 9132 2877 9160
rect 2832 9120 2838 9132
rect 3237 9129 3249 9163
rect 3283 9160 3295 9163
rect 3602 9160 3608 9172
rect 3283 9132 3608 9160
rect 3283 9129 3295 9132
rect 3237 9123 3295 9129
rect 2866 9052 2872 9104
rect 2924 9092 2930 9104
rect 3252 9092 3280 9123
rect 3602 9120 3608 9132
rect 3660 9120 3666 9172
rect 7650 9120 7656 9172
rect 7708 9160 7714 9172
rect 8113 9163 8171 9169
rect 8113 9160 8125 9163
rect 7708 9132 8125 9160
rect 7708 9120 7714 9132
rect 8113 9129 8125 9132
rect 8159 9129 8171 9163
rect 8662 9160 8668 9172
rect 8623 9132 8668 9160
rect 8113 9123 8171 9129
rect 8662 9120 8668 9132
rect 8720 9120 8726 9172
rect 9125 9163 9183 9169
rect 9125 9129 9137 9163
rect 9171 9160 9183 9163
rect 9582 9160 9588 9172
rect 9171 9132 9588 9160
rect 9171 9129 9183 9132
rect 9125 9123 9183 9129
rect 9582 9120 9588 9132
rect 9640 9120 9646 9172
rect 10042 9120 10048 9172
rect 10100 9120 10106 9172
rect 10226 9120 10232 9172
rect 10284 9160 10290 9172
rect 11701 9163 11759 9169
rect 11701 9160 11713 9163
rect 10284 9132 11713 9160
rect 10284 9120 10290 9132
rect 11701 9129 11713 9132
rect 11747 9160 11759 9163
rect 11882 9160 11888 9172
rect 11747 9132 11888 9160
rect 11747 9129 11759 9132
rect 11701 9123 11759 9129
rect 11882 9120 11888 9132
rect 11940 9120 11946 9172
rect 12894 9120 12900 9172
rect 12952 9160 12958 9172
rect 14185 9163 14243 9169
rect 14185 9160 14197 9163
rect 12952 9132 14197 9160
rect 12952 9120 12958 9132
rect 14185 9129 14197 9132
rect 14231 9129 14243 9163
rect 14185 9123 14243 9129
rect 2924 9064 2969 9092
rect 3068 9064 3280 9092
rect 3513 9095 3571 9101
rect 2924 9052 2930 9064
rect 2685 8997 2743 9003
rect 2685 8963 2697 8997
rect 2731 8963 2743 8997
rect 2685 8957 2743 8963
rect 2961 8959 3019 8965
rect 2700 8888 2728 8957
rect 2961 8925 2973 8959
rect 3007 8956 3019 8959
rect 3068 8956 3096 9064
rect 3513 9061 3525 9095
rect 3559 9092 3571 9095
rect 3878 9092 3884 9104
rect 3559 9064 3884 9092
rect 3559 9061 3571 9064
rect 3513 9055 3571 9061
rect 3878 9052 3884 9064
rect 3936 9052 3942 9104
rect 6822 9052 6828 9104
rect 6880 9092 6886 9104
rect 8294 9092 8300 9104
rect 6880 9064 8300 9092
rect 6880 9052 6886 9064
rect 3142 8984 3148 9036
rect 3200 9024 3206 9036
rect 7116 9033 7144 9064
rect 8294 9052 8300 9064
rect 8352 9052 8358 9104
rect 8570 9052 8576 9104
rect 8628 9052 8634 9104
rect 6365 9027 6423 9033
rect 3200 8996 4660 9024
rect 3200 8984 3206 8996
rect 4632 8968 4660 8996
rect 6365 8993 6377 9027
rect 6411 9024 6423 9027
rect 6917 9027 6975 9033
rect 6917 9024 6929 9027
rect 6411 8996 6929 9024
rect 6411 8993 6423 8996
rect 6365 8987 6423 8993
rect 6917 8993 6929 8996
rect 6963 8993 6975 9027
rect 6917 8987 6975 8993
rect 7101 9027 7159 9033
rect 7101 8993 7113 9027
rect 7147 8993 7159 9027
rect 7101 8987 7159 8993
rect 3007 8928 3096 8956
rect 3007 8925 3019 8928
rect 2961 8919 3019 8925
rect 3234 8916 3240 8968
rect 3292 8956 3298 8968
rect 3329 8959 3387 8965
rect 3329 8956 3341 8959
rect 3292 8928 3341 8956
rect 3292 8916 3298 8928
rect 3329 8925 3341 8928
rect 3375 8925 3387 8959
rect 3970 8956 3976 8968
rect 3931 8928 3976 8956
rect 3329 8919 3387 8925
rect 3970 8916 3976 8928
rect 4028 8916 4034 8968
rect 4062 8916 4068 8968
rect 4120 8956 4126 8968
rect 4614 8956 4620 8968
rect 4120 8928 4165 8956
rect 4575 8928 4620 8956
rect 4120 8916 4126 8928
rect 4614 8916 4620 8928
rect 4672 8916 4678 8968
rect 6932 8956 6960 8987
rect 7742 8984 7748 9036
rect 7800 9024 7806 9036
rect 7837 9027 7895 9033
rect 7837 9024 7849 9027
rect 7800 8996 7849 9024
rect 7800 8984 7806 8996
rect 7837 8993 7849 8996
rect 7883 8993 7895 9027
rect 8588 9024 8616 9052
rect 7837 8987 7895 8993
rect 8036 8996 8616 9024
rect 7374 8956 7380 8968
rect 6932 8928 7380 8956
rect 7374 8916 7380 8928
rect 7432 8916 7438 8968
rect 7653 8959 7711 8965
rect 7653 8925 7665 8959
rect 7699 8956 7711 8959
rect 8036 8956 8064 8996
rect 9490 8984 9496 9036
rect 9548 9024 9554 9036
rect 9585 9027 9643 9033
rect 9585 9024 9597 9027
rect 9548 8996 9597 9024
rect 9548 8984 9554 8996
rect 9585 8993 9597 8996
rect 9631 8993 9643 9027
rect 9766 9024 9772 9036
rect 9727 8996 9772 9024
rect 9585 8987 9643 8993
rect 8202 8956 8208 8968
rect 7699 8928 8064 8956
rect 8163 8928 8208 8956
rect 7699 8925 7711 8928
rect 7653 8919 7711 8925
rect 8202 8916 8208 8928
rect 8260 8916 8266 8968
rect 8294 8916 8300 8968
rect 8352 8956 8358 8968
rect 8573 8959 8631 8965
rect 8573 8956 8585 8959
rect 8352 8928 8585 8956
rect 8352 8916 8358 8928
rect 8573 8925 8585 8928
rect 8619 8925 8631 8959
rect 9600 8956 9628 8987
rect 9766 8984 9772 8996
rect 9824 8984 9830 9036
rect 10060 9024 10088 9120
rect 10229 9027 10287 9033
rect 10229 9024 10241 9027
rect 10060 8996 10241 9024
rect 10229 8993 10241 8996
rect 10275 8993 10287 9027
rect 10229 8987 10287 8993
rect 10686 8984 10692 9036
rect 10744 9024 10750 9036
rect 12066 9024 12072 9036
rect 10744 8996 12072 9024
rect 10744 8984 10750 8996
rect 12066 8984 12072 8996
rect 12124 9024 12130 9036
rect 13909 9027 13967 9033
rect 13909 9024 13921 9027
rect 12124 8996 13921 9024
rect 12124 8984 12130 8996
rect 13909 8993 13921 8996
rect 13955 9024 13967 9027
rect 14921 9027 14979 9033
rect 14921 9024 14933 9027
rect 13955 8996 14933 9024
rect 13955 8993 13967 8996
rect 13909 8987 13967 8993
rect 14921 8993 14933 8996
rect 14967 8993 14979 9027
rect 14921 8987 14979 8993
rect 15010 8984 15016 9036
rect 15068 9024 15074 9036
rect 15068 8996 15113 9024
rect 15068 8984 15074 8996
rect 9953 8959 10011 8965
rect 9953 8956 9965 8959
rect 9600 8928 9965 8956
rect 8573 8919 8631 8925
rect 9953 8925 9965 8928
rect 9999 8925 10011 8959
rect 14093 8959 14151 8965
rect 11362 8928 12480 8956
rect 9953 8919 10011 8925
rect 3694 8888 3700 8900
rect 2700 8860 3700 8888
rect 3694 8848 3700 8860
rect 3752 8888 3758 8900
rect 4246 8888 4252 8900
rect 3752 8860 4252 8888
rect 3752 8848 3758 8860
rect 4246 8848 4252 8860
rect 4304 8848 4310 8900
rect 4433 8891 4491 8897
rect 4433 8857 4445 8891
rect 4479 8888 4491 8891
rect 4522 8888 4528 8900
rect 4479 8860 4528 8888
rect 4479 8857 4491 8860
rect 4433 8851 4491 8857
rect 4522 8848 4528 8860
rect 4580 8848 4586 8900
rect 4890 8888 4896 8900
rect 4851 8860 4896 8888
rect 4890 8848 4896 8860
rect 4948 8848 4954 8900
rect 5350 8848 5356 8900
rect 5408 8848 5414 8900
rect 6825 8891 6883 8897
rect 6825 8857 6837 8891
rect 6871 8888 6883 8891
rect 8588 8888 8616 8919
rect 11885 8891 11943 8897
rect 6871 8860 7328 8888
rect 8588 8860 10088 8888
rect 6871 8857 6883 8860
rect 6825 8851 6883 8857
rect 3789 8823 3847 8829
rect 3789 8789 3801 8823
rect 3835 8820 3847 8823
rect 4338 8820 4344 8832
rect 3835 8792 4344 8820
rect 3835 8789 3847 8792
rect 3789 8783 3847 8789
rect 4338 8780 4344 8792
rect 4396 8780 4402 8832
rect 6454 8780 6460 8832
rect 6512 8820 6518 8832
rect 7300 8829 7328 8860
rect 7285 8823 7343 8829
rect 6512 8792 6557 8820
rect 6512 8780 6518 8792
rect 7285 8789 7297 8823
rect 7331 8789 7343 8823
rect 7285 8783 7343 8789
rect 7742 8780 7748 8832
rect 7800 8820 7806 8832
rect 8938 8820 8944 8832
rect 7800 8792 7845 8820
rect 8899 8792 8944 8820
rect 7800 8780 7806 8792
rect 8938 8780 8944 8792
rect 8996 8780 9002 8832
rect 9493 8823 9551 8829
rect 9493 8789 9505 8823
rect 9539 8820 9551 8823
rect 9950 8820 9956 8832
rect 9539 8792 9956 8820
rect 9539 8789 9551 8792
rect 9493 8783 9551 8789
rect 9950 8780 9956 8792
rect 10008 8780 10014 8832
rect 10060 8820 10088 8860
rect 11885 8857 11897 8891
rect 11931 8888 11943 8891
rect 12158 8888 12164 8900
rect 11931 8860 12164 8888
rect 11931 8857 11943 8860
rect 11885 8851 11943 8857
rect 11900 8820 11928 8851
rect 12158 8848 12164 8860
rect 12216 8848 12222 8900
rect 10060 8792 11928 8820
rect 12452 8820 12480 8928
rect 14093 8925 14105 8959
rect 14139 8956 14151 8959
rect 15289 8959 15347 8965
rect 15289 8956 15301 8959
rect 14139 8928 15301 8956
rect 14139 8925 14151 8928
rect 14093 8919 14151 8925
rect 15289 8925 15301 8928
rect 15335 8925 15347 8959
rect 15289 8919 15347 8925
rect 13354 8888 13360 8900
rect 13202 8874 13360 8888
rect 13188 8860 13360 8874
rect 12618 8820 12624 8832
rect 12452 8792 12624 8820
rect 12618 8780 12624 8792
rect 12676 8820 12682 8832
rect 13188 8820 13216 8860
rect 13354 8848 13360 8860
rect 13412 8848 13418 8900
rect 13538 8848 13544 8900
rect 13596 8888 13602 8900
rect 13633 8891 13691 8897
rect 13633 8888 13645 8891
rect 13596 8860 13645 8888
rect 13596 8848 13602 8860
rect 13633 8857 13645 8860
rect 13679 8857 13691 8891
rect 13633 8851 13691 8857
rect 14369 8823 14427 8829
rect 14369 8820 14381 8823
rect 12676 8792 14381 8820
rect 12676 8780 12682 8792
rect 14369 8789 14381 8792
rect 14415 8789 14427 8823
rect 14369 8783 14427 8789
rect 1104 8730 14812 8752
rect 1104 8678 5547 8730
rect 5599 8678 5611 8730
rect 5663 8678 5675 8730
rect 5727 8678 5739 8730
rect 5791 8678 5803 8730
rect 5855 8678 10144 8730
rect 10196 8678 10208 8730
rect 10260 8678 10272 8730
rect 10324 8678 10336 8730
rect 10388 8678 10400 8730
rect 10452 8678 14812 8730
rect 1104 8656 14812 8678
rect 2869 8619 2927 8625
rect 2869 8585 2881 8619
rect 2915 8616 2927 8619
rect 3970 8616 3976 8628
rect 2915 8588 3976 8616
rect 2915 8585 2927 8588
rect 2869 8579 2927 8585
rect 3970 8576 3976 8588
rect 4028 8576 4034 8628
rect 4062 8576 4068 8628
rect 4120 8616 4126 8628
rect 4801 8619 4859 8625
rect 4801 8616 4813 8619
rect 4120 8588 4813 8616
rect 4120 8576 4126 8588
rect 4801 8585 4813 8588
rect 4847 8585 4859 8619
rect 4801 8579 4859 8585
rect 4890 8576 4896 8628
rect 4948 8616 4954 8628
rect 5077 8619 5135 8625
rect 5077 8616 5089 8619
rect 4948 8588 5089 8616
rect 4948 8576 4954 8588
rect 5077 8585 5089 8588
rect 5123 8585 5135 8619
rect 5077 8579 5135 8585
rect 6733 8619 6791 8625
rect 6733 8585 6745 8619
rect 6779 8616 6791 8619
rect 7190 8616 7196 8628
rect 6779 8588 7196 8616
rect 6779 8585 6791 8588
rect 6733 8579 6791 8585
rect 7190 8576 7196 8588
rect 7248 8576 7254 8628
rect 7742 8616 7748 8628
rect 7703 8588 7748 8616
rect 7742 8576 7748 8588
rect 7800 8576 7806 8628
rect 9490 8616 9496 8628
rect 8864 8588 9496 8616
rect 3878 8508 3884 8560
rect 3936 8508 3942 8560
rect 4338 8548 4344 8560
rect 4299 8520 4344 8548
rect 4338 8508 4344 8520
rect 4396 8508 4402 8560
rect 6454 8548 6460 8560
rect 5276 8520 6460 8548
rect 4893 8483 4951 8489
rect 4893 8449 4905 8483
rect 4939 8480 4951 8483
rect 4982 8480 4988 8492
rect 4939 8452 4988 8480
rect 4939 8449 4951 8452
rect 4893 8443 4951 8449
rect 4982 8440 4988 8452
rect 5040 8440 5046 8492
rect 5276 8489 5304 8520
rect 6454 8508 6460 8520
rect 6512 8508 6518 8560
rect 6822 8508 6828 8560
rect 6880 8508 6886 8560
rect 8573 8551 8631 8557
rect 8573 8517 8585 8551
rect 8619 8548 8631 8551
rect 8662 8548 8668 8560
rect 8619 8520 8668 8548
rect 8619 8517 8631 8520
rect 8573 8511 8631 8517
rect 8662 8508 8668 8520
rect 8720 8508 8726 8560
rect 5261 8483 5319 8489
rect 5261 8449 5273 8483
rect 5307 8449 5319 8483
rect 5261 8443 5319 8449
rect 6089 8483 6147 8489
rect 6089 8449 6101 8483
rect 6135 8480 6147 8483
rect 6840 8480 6868 8508
rect 7374 8480 7380 8492
rect 6135 8452 6408 8480
rect 6840 8452 6960 8480
rect 7335 8452 7380 8480
rect 6135 8449 6147 8452
rect 6089 8443 6147 8449
rect 4614 8412 4620 8424
rect 4527 8384 4620 8412
rect 4614 8372 4620 8384
rect 4672 8412 4678 8424
rect 5442 8412 5448 8424
rect 4672 8384 5448 8412
rect 4672 8372 4678 8384
rect 5442 8372 5448 8384
rect 5500 8372 5506 8424
rect 6380 8353 6408 8452
rect 6932 8421 6960 8452
rect 7374 8440 7380 8452
rect 7432 8440 7438 8492
rect 7742 8440 7748 8492
rect 7800 8480 7806 8492
rect 8021 8483 8079 8489
rect 8021 8480 8033 8483
rect 7800 8452 8033 8480
rect 7800 8440 7806 8452
rect 8021 8449 8033 8452
rect 8067 8449 8079 8483
rect 8478 8480 8484 8492
rect 8439 8452 8484 8480
rect 8021 8443 8079 8449
rect 8478 8440 8484 8452
rect 8536 8440 8542 8492
rect 8754 8480 8760 8492
rect 8715 8452 8760 8480
rect 8754 8440 8760 8452
rect 8812 8440 8818 8492
rect 8864 8489 8892 8588
rect 9490 8576 9496 8588
rect 9548 8576 9554 8628
rect 13998 8616 14004 8628
rect 11164 8588 14004 8616
rect 11164 8557 11192 8588
rect 13998 8576 14004 8588
rect 14056 8576 14062 8628
rect 11149 8551 11207 8557
rect 10258 8520 11100 8548
rect 8849 8483 8907 8489
rect 8849 8449 8861 8483
rect 8895 8449 8907 8483
rect 10965 8483 11023 8489
rect 8849 8443 8907 8449
rect 9048 8452 9352 8480
rect 6825 8415 6883 8421
rect 6825 8381 6837 8415
rect 6871 8381 6883 8415
rect 6825 8375 6883 8381
rect 6917 8415 6975 8421
rect 6917 8381 6929 8415
rect 6963 8381 6975 8415
rect 6917 8375 6975 8381
rect 7285 8415 7343 8421
rect 7285 8381 7297 8415
rect 7331 8381 7343 8415
rect 7285 8375 7343 8381
rect 6365 8347 6423 8353
rect 6365 8313 6377 8347
rect 6411 8313 6423 8347
rect 6840 8344 6868 8375
rect 7300 8344 7328 8375
rect 7466 8372 7472 8424
rect 7524 8412 7530 8424
rect 7929 8415 7987 8421
rect 7929 8412 7941 8415
rect 7524 8384 7941 8412
rect 7524 8372 7530 8384
rect 7929 8381 7941 8384
rect 7975 8381 7987 8415
rect 9048 8412 9076 8452
rect 9214 8412 9220 8424
rect 7929 8375 7987 8381
rect 8680 8384 9076 8412
rect 9175 8384 9220 8412
rect 8202 8344 8208 8356
rect 6840 8316 8208 8344
rect 6365 8307 6423 8313
rect 8202 8304 8208 8316
rect 8260 8304 8266 8356
rect 8680 8353 8708 8384
rect 9214 8372 9220 8384
rect 9272 8372 9278 8424
rect 9324 8412 9352 8452
rect 10965 8449 10977 8483
rect 11011 8449 11023 8483
rect 11072 8480 11100 8520
rect 11149 8517 11161 8551
rect 11195 8517 11207 8551
rect 11149 8511 11207 8517
rect 11333 8551 11391 8557
rect 11333 8517 11345 8551
rect 11379 8548 11391 8551
rect 12069 8551 12127 8557
rect 12069 8548 12081 8551
rect 11379 8520 12081 8548
rect 11379 8517 11391 8520
rect 11333 8511 11391 8517
rect 12069 8517 12081 8520
rect 12115 8517 12127 8551
rect 12069 8511 12127 8517
rect 12250 8508 12256 8560
rect 12308 8548 12314 8560
rect 12345 8551 12403 8557
rect 12345 8548 12357 8551
rect 12308 8520 12357 8548
rect 12308 8508 12314 8520
rect 12345 8517 12357 8520
rect 12391 8517 12403 8551
rect 12345 8511 12403 8517
rect 13446 8508 13452 8560
rect 13504 8508 13510 8560
rect 11072 8452 11744 8480
rect 10965 8443 11023 8449
rect 9674 8412 9680 8424
rect 9324 8384 9680 8412
rect 9674 8372 9680 8384
rect 9732 8372 9738 8424
rect 10980 8412 11008 8443
rect 11716 8412 11744 8452
rect 11790 8440 11796 8492
rect 11848 8480 11854 8492
rect 11885 8483 11943 8489
rect 11885 8480 11897 8483
rect 11848 8452 11897 8480
rect 11848 8440 11854 8452
rect 11885 8449 11897 8452
rect 11931 8449 11943 8483
rect 11885 8443 11943 8449
rect 11974 8440 11980 8492
rect 12032 8480 12038 8492
rect 12437 8483 12495 8489
rect 12437 8480 12449 8483
rect 12032 8452 12449 8480
rect 12032 8440 12038 8452
rect 12437 8449 12449 8452
rect 12483 8449 12495 8483
rect 12437 8443 12495 8449
rect 14461 8483 14519 8489
rect 14461 8449 14473 8483
rect 14507 8480 14519 8483
rect 14921 8483 14979 8489
rect 14921 8480 14933 8483
rect 14507 8452 14933 8480
rect 14507 8449 14519 8452
rect 14461 8443 14519 8449
rect 14921 8449 14933 8452
rect 14967 8449 14979 8483
rect 14921 8443 14979 8449
rect 12161 8415 12219 8421
rect 12161 8412 12173 8415
rect 10980 8384 11652 8412
rect 11716 8384 12173 8412
rect 11624 8353 11652 8384
rect 12161 8381 12173 8384
rect 12207 8412 12219 8415
rect 12713 8415 12771 8421
rect 12207 8384 12434 8412
rect 12207 8381 12219 8384
rect 12161 8375 12219 8381
rect 8665 8347 8723 8353
rect 8665 8313 8677 8347
rect 8711 8313 8723 8347
rect 8665 8307 8723 8313
rect 11609 8347 11667 8353
rect 11609 8313 11621 8347
rect 11655 8313 11667 8347
rect 12406 8344 12434 8384
rect 12713 8381 12725 8415
rect 12759 8412 12771 8415
rect 13538 8412 13544 8424
rect 12759 8384 13544 8412
rect 12759 8381 12771 8384
rect 12713 8375 12771 8381
rect 13538 8372 13544 8384
rect 13596 8372 13602 8424
rect 14182 8412 14188 8424
rect 14143 8384 14188 8412
rect 14182 8372 14188 8384
rect 14240 8372 14246 8424
rect 12618 8344 12624 8356
rect 12406 8316 12624 8344
rect 11609 8307 11667 8313
rect 12618 8304 12624 8316
rect 12676 8304 12682 8356
rect 5350 8276 5356 8288
rect 5311 8248 5356 8276
rect 5350 8236 5356 8248
rect 5408 8276 5414 8288
rect 5721 8279 5779 8285
rect 5721 8276 5733 8279
rect 5408 8248 5733 8276
rect 5408 8236 5414 8248
rect 5721 8245 5733 8248
rect 5767 8245 5779 8279
rect 5721 8239 5779 8245
rect 5810 8236 5816 8288
rect 5868 8276 5874 8288
rect 5905 8279 5963 8285
rect 5905 8276 5917 8279
rect 5868 8248 5917 8276
rect 5868 8236 5874 8248
rect 5905 8245 5917 8248
rect 5951 8245 5963 8279
rect 5905 8239 5963 8245
rect 8389 8279 8447 8285
rect 8389 8245 8401 8279
rect 8435 8276 8447 8279
rect 9122 8276 9128 8288
rect 8435 8248 9128 8276
rect 8435 8245 8447 8248
rect 8389 8239 8447 8245
rect 9122 8236 9128 8248
rect 9180 8236 9186 8288
rect 9950 8236 9956 8288
rect 10008 8276 10014 8288
rect 10643 8279 10701 8285
rect 10643 8276 10655 8279
rect 10008 8248 10655 8276
rect 10008 8236 10014 8248
rect 10643 8245 10655 8248
rect 10689 8245 10701 8279
rect 10643 8239 10701 8245
rect 10778 8236 10784 8288
rect 10836 8276 10842 8288
rect 10836 8248 10881 8276
rect 10836 8236 10842 8248
rect 1104 8186 14812 8208
rect 1104 8134 3248 8186
rect 3300 8134 3312 8186
rect 3364 8134 3376 8186
rect 3428 8134 3440 8186
rect 3492 8134 3504 8186
rect 3556 8134 7846 8186
rect 7898 8134 7910 8186
rect 7962 8134 7974 8186
rect 8026 8134 8038 8186
rect 8090 8134 8102 8186
rect 8154 8134 12443 8186
rect 12495 8134 12507 8186
rect 12559 8134 12571 8186
rect 12623 8134 12635 8186
rect 12687 8134 12699 8186
rect 12751 8134 14812 8186
rect 1104 8112 14812 8134
rect 9214 8032 9220 8084
rect 9272 8072 9278 8084
rect 9585 8075 9643 8081
rect 9585 8072 9597 8075
rect 9272 8044 9597 8072
rect 9272 8032 9278 8044
rect 9585 8041 9597 8044
rect 9631 8041 9643 8075
rect 9585 8035 9643 8041
rect 14182 8032 14188 8084
rect 14240 8072 14246 8084
rect 14277 8075 14335 8081
rect 14277 8072 14289 8075
rect 14240 8044 14289 8072
rect 14240 8032 14246 8044
rect 14277 8041 14289 8044
rect 14323 8041 14335 8075
rect 14277 8035 14335 8041
rect 11698 8004 11704 8016
rect 11659 7976 11704 8004
rect 11698 7964 11704 7976
rect 11756 7964 11762 8016
rect 13909 8007 13967 8013
rect 13909 7973 13921 8007
rect 13955 8004 13967 8007
rect 15105 8007 15163 8013
rect 15105 8004 15117 8007
rect 13955 7976 15117 8004
rect 13955 7973 13967 7976
rect 13909 7967 13967 7973
rect 15105 7973 15117 7976
rect 15151 7973 15163 8007
rect 15105 7967 15163 7973
rect 2498 7936 2504 7948
rect 2459 7908 2504 7936
rect 2498 7896 2504 7908
rect 2556 7896 2562 7948
rect 5442 7936 5448 7948
rect 5403 7908 5448 7936
rect 5442 7896 5448 7908
rect 5500 7896 5506 7948
rect 5810 7936 5816 7948
rect 5771 7908 5816 7936
rect 5810 7896 5816 7908
rect 5868 7896 5874 7948
rect 7098 7896 7104 7948
rect 7156 7936 7162 7948
rect 7239 7939 7297 7945
rect 7239 7936 7251 7939
rect 7156 7908 7251 7936
rect 7156 7896 7162 7908
rect 7239 7905 7251 7908
rect 7285 7936 7297 7939
rect 7285 7908 8248 7936
rect 7285 7905 7297 7908
rect 7239 7899 7297 7905
rect 8220 7880 8248 7908
rect 8754 7896 8760 7948
rect 8812 7936 8818 7948
rect 9861 7939 9919 7945
rect 9861 7936 9873 7939
rect 8812 7908 9873 7936
rect 8812 7896 8818 7908
rect 1670 7828 1676 7880
rect 1728 7868 1734 7880
rect 2225 7871 2283 7877
rect 2225 7868 2237 7871
rect 1728 7840 2237 7868
rect 1728 7828 1734 7840
rect 2225 7837 2237 7840
rect 2271 7837 2283 7871
rect 2682 7868 2688 7880
rect 2643 7840 2688 7868
rect 2225 7831 2283 7837
rect 2682 7828 2688 7840
rect 2740 7828 2746 7880
rect 2777 7871 2835 7877
rect 2777 7837 2789 7871
rect 2823 7868 2835 7871
rect 2958 7868 2964 7880
rect 2823 7840 2964 7868
rect 2823 7837 2835 7840
rect 2777 7831 2835 7837
rect 2958 7828 2964 7840
rect 3016 7828 3022 7880
rect 7374 7868 7380 7880
rect 7335 7840 7380 7868
rect 7374 7828 7380 7840
rect 7432 7828 7438 7880
rect 7742 7868 7748 7880
rect 7703 7840 7748 7868
rect 7742 7828 7748 7840
rect 7800 7828 7806 7880
rect 8202 7868 8208 7880
rect 8163 7840 8208 7868
rect 8202 7828 8208 7840
rect 8260 7828 8266 7880
rect 8662 7828 8668 7880
rect 8720 7868 8726 7880
rect 9232 7877 9260 7908
rect 9861 7905 9873 7908
rect 9907 7905 9919 7939
rect 9861 7899 9919 7905
rect 12434 7896 12440 7948
rect 12492 7936 12498 7948
rect 12492 7908 12537 7936
rect 12492 7896 12498 7908
rect 8941 7871 8999 7877
rect 8941 7868 8953 7871
rect 8720 7840 8953 7868
rect 8720 7828 8726 7840
rect 8941 7837 8953 7840
rect 8987 7837 8999 7871
rect 8941 7831 8999 7837
rect 9217 7871 9275 7877
rect 9217 7837 9229 7871
rect 9263 7837 9275 7871
rect 9217 7831 9275 7837
rect 9401 7871 9459 7877
rect 9401 7837 9413 7871
rect 9447 7868 9459 7871
rect 9493 7871 9551 7877
rect 9493 7868 9505 7871
rect 9447 7840 9505 7868
rect 9447 7837 9459 7840
rect 9401 7831 9459 7837
rect 9493 7837 9505 7840
rect 9539 7837 9551 7871
rect 9674 7868 9680 7880
rect 9635 7840 9680 7868
rect 9493 7831 9551 7837
rect 9674 7828 9680 7840
rect 9732 7828 9738 7880
rect 9950 7868 9956 7880
rect 9911 7840 9956 7868
rect 9950 7828 9956 7840
rect 10008 7828 10014 7880
rect 10321 7871 10379 7877
rect 10321 7837 10333 7871
rect 10367 7868 10379 7871
rect 12158 7868 12164 7880
rect 10367 7840 12164 7868
rect 10367 7837 10379 7840
rect 10321 7831 10379 7837
rect 12158 7828 12164 7840
rect 12216 7828 12222 7880
rect 14461 7871 14519 7877
rect 14461 7837 14473 7871
rect 14507 7868 14519 7871
rect 15013 7871 15071 7877
rect 15013 7868 15025 7871
rect 14507 7840 15025 7868
rect 14507 7837 14519 7840
rect 14461 7831 14519 7837
rect 15013 7837 15025 7840
rect 15059 7837 15071 7871
rect 15013 7831 15071 7837
rect 6730 7760 6736 7812
rect 6788 7760 6794 7812
rect 7929 7803 7987 7809
rect 7929 7769 7941 7803
rect 7975 7800 7987 7803
rect 8478 7800 8484 7812
rect 7975 7772 8484 7800
rect 7975 7769 7987 7772
rect 7929 7763 7987 7769
rect 8478 7760 8484 7772
rect 8536 7800 8542 7812
rect 9033 7803 9091 7809
rect 9033 7800 9045 7803
rect 8536 7772 9045 7800
rect 8536 7760 8542 7772
rect 9033 7769 9045 7772
rect 9079 7769 9091 7803
rect 9033 7763 9091 7769
rect 10588 7803 10646 7809
rect 10588 7769 10600 7803
rect 10634 7800 10646 7803
rect 10778 7800 10784 7812
rect 10634 7772 10784 7800
rect 10634 7769 10646 7772
rect 10588 7763 10646 7769
rect 10778 7760 10784 7772
rect 10836 7760 10842 7812
rect 1946 7692 1952 7744
rect 2004 7732 2010 7744
rect 2133 7735 2191 7741
rect 2133 7732 2145 7735
rect 2004 7704 2145 7732
rect 2004 7692 2010 7704
rect 2133 7701 2145 7704
rect 2179 7701 2191 7735
rect 2133 7695 2191 7701
rect 2314 7692 2320 7744
rect 2372 7732 2378 7744
rect 2501 7735 2559 7741
rect 2501 7732 2513 7735
rect 2372 7704 2513 7732
rect 2372 7692 2378 7704
rect 2501 7701 2513 7704
rect 2547 7701 2559 7735
rect 3326 7732 3332 7744
rect 3239 7704 3332 7732
rect 2501 7695 2559 7701
rect 3326 7692 3332 7704
rect 3384 7732 3390 7744
rect 3878 7732 3884 7744
rect 3384 7704 3884 7732
rect 3384 7692 3390 7704
rect 3878 7692 3884 7704
rect 3936 7732 3942 7744
rect 3973 7735 4031 7741
rect 3973 7732 3985 7735
rect 3936 7704 3985 7732
rect 3936 7692 3942 7704
rect 3973 7701 3985 7704
rect 4019 7732 4031 7735
rect 5350 7732 5356 7744
rect 4019 7704 5356 7732
rect 4019 7701 4031 7704
rect 3973 7695 4031 7701
rect 5350 7692 5356 7704
rect 5408 7732 5414 7744
rect 6748 7732 6776 7760
rect 5408 7704 6776 7732
rect 5408 7692 5414 7704
rect 8570 7692 8576 7744
rect 8628 7732 8634 7744
rect 8665 7735 8723 7741
rect 8665 7732 8677 7735
rect 8628 7704 8677 7732
rect 8628 7692 8634 7704
rect 8665 7701 8677 7704
rect 8711 7732 8723 7735
rect 8938 7732 8944 7744
rect 8711 7704 8944 7732
rect 8711 7701 8723 7704
rect 8665 7695 8723 7701
rect 8938 7692 8944 7704
rect 8996 7732 9002 7744
rect 10137 7735 10195 7741
rect 10137 7732 10149 7735
rect 8996 7704 10149 7732
rect 8996 7692 9002 7704
rect 10137 7701 10149 7704
rect 10183 7701 10195 7735
rect 10137 7695 10195 7701
rect 11885 7735 11943 7741
rect 11885 7701 11897 7735
rect 11931 7732 11943 7735
rect 11977 7735 12035 7741
rect 11977 7732 11989 7735
rect 11931 7704 11989 7732
rect 11931 7701 11943 7704
rect 11885 7695 11943 7701
rect 11977 7701 11989 7704
rect 12023 7732 12035 7735
rect 12342 7732 12348 7744
rect 12023 7704 12348 7732
rect 12023 7701 12035 7704
rect 11977 7695 12035 7701
rect 12342 7692 12348 7704
rect 12400 7692 12406 7744
rect 13446 7692 13452 7744
rect 13504 7732 13510 7744
rect 13648 7732 13676 7786
rect 14090 7732 14096 7744
rect 13504 7704 14096 7732
rect 13504 7692 13510 7704
rect 14090 7692 14096 7704
rect 14148 7692 14154 7744
rect 1104 7642 14812 7664
rect 1104 7590 5547 7642
rect 5599 7590 5611 7642
rect 5663 7590 5675 7642
rect 5727 7590 5739 7642
rect 5791 7590 5803 7642
rect 5855 7590 10144 7642
rect 10196 7590 10208 7642
rect 10260 7590 10272 7642
rect 10324 7590 10336 7642
rect 10388 7590 10400 7642
rect 10452 7590 14812 7642
rect 1104 7568 14812 7590
rect 7101 7531 7159 7537
rect 7101 7497 7113 7531
rect 7147 7528 7159 7531
rect 7466 7528 7472 7540
rect 7147 7500 7472 7528
rect 7147 7497 7159 7500
rect 7101 7491 7159 7497
rect 7466 7488 7472 7500
rect 7524 7488 7530 7540
rect 7653 7531 7711 7537
rect 7653 7497 7665 7531
rect 7699 7528 7711 7531
rect 7742 7528 7748 7540
rect 7699 7500 7748 7528
rect 7699 7497 7711 7500
rect 7653 7491 7711 7497
rect 7742 7488 7748 7500
rect 7800 7488 7806 7540
rect 11422 7488 11428 7540
rect 11480 7528 11486 7540
rect 11517 7531 11575 7537
rect 11517 7528 11529 7531
rect 11480 7500 11529 7528
rect 11480 7488 11486 7500
rect 11517 7497 11529 7500
rect 11563 7497 11575 7531
rect 11517 7491 11575 7497
rect 12158 7488 12164 7540
rect 12216 7528 12222 7540
rect 12216 7500 13216 7528
rect 12216 7488 12222 7500
rect 3326 7420 3332 7472
rect 3384 7420 3390 7472
rect 6825 7463 6883 7469
rect 6825 7429 6837 7463
rect 6871 7460 6883 7463
rect 7374 7460 7380 7472
rect 6871 7432 7380 7460
rect 6871 7429 6883 7432
rect 6825 7423 6883 7429
rect 7374 7420 7380 7432
rect 7432 7420 7438 7472
rect 8570 7420 8576 7472
rect 8628 7420 8634 7472
rect 9122 7460 9128 7472
rect 9083 7432 9128 7460
rect 9122 7420 9128 7432
rect 9180 7420 9186 7472
rect 10502 7460 10508 7472
rect 9600 7432 10508 7460
rect 9600 7404 9628 7432
rect 10502 7420 10508 7432
rect 10560 7420 10566 7472
rect 12342 7420 12348 7472
rect 12400 7420 12406 7472
rect 13188 7460 13216 7500
rect 13262 7488 13268 7540
rect 13320 7528 13326 7540
rect 13357 7531 13415 7537
rect 13357 7528 13369 7531
rect 13320 7500 13369 7528
rect 13320 7488 13326 7500
rect 13357 7497 13369 7500
rect 13403 7497 13415 7531
rect 13722 7528 13728 7540
rect 13683 7500 13728 7528
rect 13357 7491 13415 7497
rect 13722 7488 13728 7500
rect 13780 7488 13786 7540
rect 13817 7531 13875 7537
rect 13817 7497 13829 7531
rect 13863 7528 13875 7531
rect 14921 7531 14979 7537
rect 14921 7528 14933 7531
rect 13863 7500 14933 7528
rect 13863 7497 13875 7500
rect 13817 7491 13875 7497
rect 14921 7497 14933 7500
rect 14967 7497 14979 7531
rect 14921 7491 14979 7497
rect 13188 7432 13308 7460
rect 1946 7392 1952 7404
rect 1907 7364 1952 7392
rect 1946 7352 1952 7364
rect 2004 7352 2010 7404
rect 2314 7392 2320 7404
rect 2275 7364 2320 7392
rect 2314 7352 2320 7364
rect 2372 7352 2378 7404
rect 3743 7395 3801 7401
rect 3743 7361 3755 7395
rect 3789 7392 3801 7395
rect 4154 7392 4160 7404
rect 3789 7364 4160 7392
rect 3789 7361 3801 7364
rect 3743 7355 3801 7361
rect 4154 7352 4160 7364
rect 4212 7352 4218 7404
rect 4614 7392 4620 7404
rect 4575 7364 4620 7392
rect 4614 7352 4620 7364
rect 4672 7352 4678 7404
rect 4801 7395 4859 7401
rect 4801 7361 4813 7395
rect 4847 7361 4859 7395
rect 7098 7392 7104 7404
rect 7059 7364 7104 7392
rect 4801 7355 4859 7361
rect 4065 7327 4123 7333
rect 4065 7293 4077 7327
rect 4111 7293 4123 7327
rect 4172 7324 4200 7352
rect 4816 7324 4844 7355
rect 7098 7352 7104 7364
rect 7156 7352 7162 7404
rect 7190 7352 7196 7404
rect 7248 7392 7254 7404
rect 9401 7395 9459 7401
rect 7248 7364 7293 7392
rect 7248 7352 7254 7364
rect 9401 7361 9413 7395
rect 9447 7392 9459 7395
rect 9490 7392 9496 7404
rect 9447 7364 9496 7392
rect 9447 7361 9459 7364
rect 9401 7355 9459 7361
rect 9490 7352 9496 7364
rect 9548 7352 9554 7404
rect 9582 7352 9588 7404
rect 9640 7392 9646 7404
rect 10134 7392 10140 7404
rect 9640 7364 9733 7392
rect 10095 7364 10140 7392
rect 9640 7352 9646 7364
rect 10134 7352 10140 7364
rect 10192 7352 10198 7404
rect 11333 7395 11391 7401
rect 11333 7361 11345 7395
rect 11379 7392 11391 7395
rect 11698 7392 11704 7404
rect 11379 7364 11704 7392
rect 11379 7361 11391 7364
rect 11333 7355 11391 7361
rect 11698 7352 11704 7364
rect 11756 7352 11762 7404
rect 13280 7401 13308 7432
rect 13265 7395 13323 7401
rect 13265 7361 13277 7395
rect 13311 7392 13323 7395
rect 13354 7392 13360 7404
rect 13311 7364 13360 7392
rect 13311 7361 13323 7364
rect 13265 7355 13323 7361
rect 13354 7352 13360 7364
rect 13412 7352 13418 7404
rect 14461 7395 14519 7401
rect 14461 7361 14473 7395
rect 14507 7392 14519 7395
rect 15197 7395 15255 7401
rect 15197 7392 15209 7395
rect 14507 7364 15209 7392
rect 14507 7361 14519 7364
rect 14461 7355 14519 7361
rect 15197 7361 15209 7364
rect 15243 7361 15255 7395
rect 15197 7355 15255 7361
rect 4172 7296 4844 7324
rect 4065 7287 4123 7293
rect 4080 7256 4108 7287
rect 6822 7284 6828 7336
rect 6880 7324 6886 7336
rect 7009 7327 7067 7333
rect 7009 7324 7021 7327
rect 6880 7296 7021 7324
rect 6880 7284 6886 7296
rect 7009 7293 7021 7296
rect 7055 7293 7067 7327
rect 7009 7287 7067 7293
rect 7469 7327 7527 7333
rect 7469 7293 7481 7327
rect 7515 7324 7527 7327
rect 7742 7324 7748 7336
rect 7515 7296 7748 7324
rect 7515 7293 7527 7296
rect 7469 7287 7527 7293
rect 7742 7284 7748 7296
rect 7800 7284 7806 7336
rect 10045 7327 10103 7333
rect 10045 7293 10057 7327
rect 10091 7324 10103 7327
rect 10689 7327 10747 7333
rect 10091 7296 10640 7324
rect 10091 7293 10103 7296
rect 10045 7287 10103 7293
rect 4706 7256 4712 7268
rect 4080 7228 4712 7256
rect 4706 7216 4712 7228
rect 4764 7216 4770 7268
rect 10134 7256 10140 7268
rect 9876 7228 10140 7256
rect 4430 7188 4436 7200
rect 4391 7160 4436 7188
rect 4430 7148 4436 7160
rect 4488 7148 4494 7200
rect 4522 7148 4528 7200
rect 4580 7188 4586 7200
rect 4617 7191 4675 7197
rect 4617 7188 4629 7191
rect 4580 7160 4629 7188
rect 4580 7148 4586 7160
rect 4617 7157 4629 7160
rect 4663 7157 4675 7191
rect 6730 7188 6736 7200
rect 6691 7160 6736 7188
rect 4617 7151 4675 7157
rect 6730 7148 6736 7160
rect 6788 7148 6794 7200
rect 7282 7188 7288 7200
rect 7243 7160 7288 7188
rect 7282 7148 7288 7160
rect 7340 7148 7346 7200
rect 7374 7148 7380 7200
rect 7432 7188 7438 7200
rect 9876 7197 9904 7228
rect 10134 7216 10140 7228
rect 10192 7216 10198 7268
rect 10612 7256 10640 7296
rect 10689 7293 10701 7327
rect 10735 7324 10747 7327
rect 12989 7327 13047 7333
rect 12989 7324 13001 7327
rect 10735 7296 13001 7324
rect 10735 7293 10747 7296
rect 10689 7287 10747 7293
rect 12989 7293 13001 7296
rect 13035 7293 13047 7327
rect 12989 7287 13047 7293
rect 14001 7327 14059 7333
rect 14001 7293 14013 7327
rect 14047 7324 14059 7327
rect 15105 7327 15163 7333
rect 15105 7324 15117 7327
rect 14047 7296 15117 7324
rect 14047 7293 14059 7296
rect 14001 7287 14059 7293
rect 15105 7293 15117 7296
rect 15151 7293 15163 7327
rect 15105 7287 15163 7293
rect 11606 7256 11612 7268
rect 10612 7228 11612 7256
rect 11606 7216 11612 7228
rect 11664 7216 11670 7268
rect 14277 7259 14335 7265
rect 14277 7225 14289 7259
rect 14323 7256 14335 7259
rect 15381 7259 15439 7265
rect 15381 7256 15393 7259
rect 14323 7228 15393 7256
rect 14323 7225 14335 7228
rect 14277 7219 14335 7225
rect 15381 7225 15393 7228
rect 15427 7225 15439 7259
rect 15381 7219 15439 7225
rect 9861 7191 9919 7197
rect 7432 7160 7477 7188
rect 7432 7148 7438 7160
rect 9861 7157 9873 7191
rect 9907 7157 9919 7191
rect 9861 7151 9919 7157
rect 10413 7191 10471 7197
rect 10413 7157 10425 7191
rect 10459 7188 10471 7191
rect 10502 7188 10508 7200
rect 10459 7160 10508 7188
rect 10459 7157 10471 7160
rect 10413 7151 10471 7157
rect 10502 7148 10508 7160
rect 10560 7148 10566 7200
rect 10597 7191 10655 7197
rect 10597 7157 10609 7191
rect 10643 7188 10655 7191
rect 11422 7188 11428 7200
rect 10643 7160 11428 7188
rect 10643 7157 10655 7160
rect 10597 7151 10655 7157
rect 11422 7148 11428 7160
rect 11480 7148 11486 7200
rect 1104 7098 14812 7120
rect 1104 7046 3248 7098
rect 3300 7046 3312 7098
rect 3364 7046 3376 7098
rect 3428 7046 3440 7098
rect 3492 7046 3504 7098
rect 3556 7046 7846 7098
rect 7898 7046 7910 7098
rect 7962 7046 7974 7098
rect 8026 7046 8038 7098
rect 8090 7046 8102 7098
rect 8154 7046 12443 7098
rect 12495 7046 12507 7098
rect 12559 7046 12571 7098
rect 12623 7046 12635 7098
rect 12687 7046 12699 7098
rect 12751 7046 14812 7098
rect 1104 7024 14812 7046
rect 2133 6987 2191 6993
rect 2133 6953 2145 6987
rect 2179 6984 2191 6987
rect 2498 6984 2504 6996
rect 2179 6956 2504 6984
rect 2179 6953 2191 6956
rect 2133 6947 2191 6953
rect 2498 6944 2504 6956
rect 2556 6944 2562 6996
rect 3694 6944 3700 6996
rect 3752 6984 3758 6996
rect 3752 6956 4844 6984
rect 3752 6944 3758 6956
rect 4154 6876 4160 6928
rect 4212 6916 4218 6928
rect 4212 6888 4660 6916
rect 4212 6876 4218 6888
rect 2317 6851 2375 6857
rect 2317 6817 2329 6851
rect 2363 6848 2375 6851
rect 3050 6848 3056 6860
rect 2363 6820 3056 6848
rect 2363 6817 2375 6820
rect 2317 6811 2375 6817
rect 3050 6808 3056 6820
rect 3108 6808 3114 6860
rect 3329 6851 3387 6857
rect 3329 6817 3341 6851
rect 3375 6817 3387 6851
rect 3602 6848 3608 6860
rect 3563 6820 3608 6848
rect 3329 6811 3387 6817
rect 2038 6780 2044 6792
rect 1999 6752 2044 6780
rect 2038 6740 2044 6752
rect 2096 6740 2102 6792
rect 2225 6783 2283 6789
rect 2225 6749 2237 6783
rect 2271 6780 2283 6783
rect 2501 6783 2559 6789
rect 2501 6780 2513 6783
rect 2271 6752 2513 6780
rect 2271 6749 2283 6752
rect 2225 6743 2283 6749
rect 2501 6749 2513 6752
rect 2547 6749 2559 6783
rect 2501 6743 2559 6749
rect 2593 6783 2651 6789
rect 2593 6749 2605 6783
rect 2639 6780 2651 6783
rect 2961 6783 3019 6789
rect 2639 6752 2912 6780
rect 2639 6749 2651 6752
rect 2593 6743 2651 6749
rect 2516 6712 2544 6743
rect 2682 6712 2688 6724
rect 2516 6684 2688 6712
rect 2682 6672 2688 6684
rect 2740 6672 2746 6724
rect 2314 6644 2320 6656
rect 2275 6616 2320 6644
rect 2314 6604 2320 6616
rect 2372 6604 2378 6656
rect 2884 6653 2912 6752
rect 2961 6749 2973 6783
rect 3007 6780 3019 6783
rect 3237 6783 3295 6789
rect 3237 6780 3249 6783
rect 3007 6752 3249 6780
rect 3007 6749 3019 6752
rect 2961 6743 3019 6749
rect 3237 6749 3249 6752
rect 3283 6749 3295 6783
rect 3344 6780 3372 6811
rect 3602 6808 3608 6820
rect 3660 6808 3666 6860
rect 4522 6848 4528 6860
rect 3712 6820 4528 6848
rect 3712 6780 3740 6820
rect 4522 6808 4528 6820
rect 4580 6808 4586 6860
rect 4632 6848 4660 6888
rect 4816 6848 4844 6956
rect 7374 6944 7380 6996
rect 7432 6984 7438 6996
rect 8113 6987 8171 6993
rect 8113 6984 8125 6987
rect 7432 6956 8125 6984
rect 7432 6944 7438 6956
rect 8113 6953 8125 6956
rect 8159 6953 8171 6987
rect 9582 6984 9588 6996
rect 8113 6947 8171 6953
rect 9048 6956 9588 6984
rect 7190 6876 7196 6928
rect 7248 6916 7254 6928
rect 7469 6919 7527 6925
rect 7469 6916 7481 6919
rect 7248 6888 7481 6916
rect 7248 6876 7254 6888
rect 7469 6885 7481 6888
rect 7515 6885 7527 6919
rect 7469 6879 7527 6885
rect 8846 6876 8852 6928
rect 8904 6916 8910 6928
rect 9048 6916 9076 6956
rect 9582 6944 9588 6956
rect 9640 6944 9646 6996
rect 10134 6944 10140 6996
rect 10192 6984 10198 6996
rect 10597 6987 10655 6993
rect 10597 6984 10609 6987
rect 10192 6956 10609 6984
rect 10192 6944 10198 6956
rect 10597 6953 10609 6956
rect 10643 6953 10655 6987
rect 10597 6947 10655 6953
rect 11146 6944 11152 6996
rect 11204 6984 11210 6996
rect 11204 6956 14504 6984
rect 11204 6944 11210 6956
rect 14476 6928 14504 6956
rect 8904 6888 9076 6916
rect 11057 6919 11115 6925
rect 8904 6876 8910 6888
rect 11057 6885 11069 6919
rect 11103 6885 11115 6919
rect 11057 6879 11115 6885
rect 4890 6848 4896 6860
rect 4632 6820 4752 6848
rect 4816 6820 4896 6848
rect 3344 6752 3740 6780
rect 3789 6783 3847 6789
rect 3237 6743 3295 6749
rect 3789 6749 3801 6783
rect 3835 6749 3847 6783
rect 3789 6743 3847 6749
rect 3142 6672 3148 6724
rect 3200 6712 3206 6724
rect 3252 6712 3280 6743
rect 3804 6712 3832 6743
rect 3878 6740 3884 6792
rect 3936 6740 3942 6792
rect 4154 6780 4160 6792
rect 4115 6752 4160 6780
rect 4154 6740 4160 6752
rect 4212 6740 4218 6792
rect 4614 6780 4620 6792
rect 4264 6752 4620 6780
rect 3200 6684 3832 6712
rect 3896 6712 3924 6740
rect 4264 6712 4292 6752
rect 4614 6740 4620 6752
rect 4672 6740 4678 6792
rect 4724 6789 4752 6820
rect 4890 6808 4896 6820
rect 4948 6848 4954 6860
rect 5629 6851 5687 6857
rect 5629 6848 5641 6851
rect 4948 6820 5641 6848
rect 4948 6808 4954 6820
rect 5629 6817 5641 6820
rect 5675 6848 5687 6851
rect 5902 6848 5908 6860
rect 5675 6820 5908 6848
rect 5675 6817 5687 6820
rect 5629 6811 5687 6817
rect 5902 6808 5908 6820
rect 5960 6808 5966 6860
rect 8205 6851 8263 6857
rect 7024 6820 7972 6848
rect 4709 6783 4767 6789
rect 4709 6749 4721 6783
rect 4755 6749 4767 6783
rect 4709 6743 4767 6749
rect 5534 6740 5540 6792
rect 5592 6780 5598 6792
rect 5997 6783 6055 6789
rect 5997 6780 6009 6783
rect 5592 6752 6009 6780
rect 5592 6740 5598 6752
rect 5997 6749 6009 6752
rect 6043 6749 6055 6783
rect 5997 6743 6055 6749
rect 6638 6740 6644 6792
rect 6696 6780 6702 6792
rect 7024 6780 7052 6820
rect 7944 6789 7972 6820
rect 8205 6817 8217 6851
rect 8251 6848 8263 6851
rect 11072 6848 11100 6879
rect 14458 6876 14464 6928
rect 14516 6876 14522 6928
rect 11514 6848 11520 6860
rect 8251 6820 9352 6848
rect 11072 6820 11520 6848
rect 8251 6817 8263 6820
rect 8205 6811 8263 6817
rect 7469 6783 7527 6789
rect 7469 6780 7481 6783
rect 6696 6752 7052 6780
rect 7392 6752 7481 6780
rect 6696 6740 6702 6752
rect 3896 6684 4292 6712
rect 3200 6672 3206 6684
rect 4522 6672 4528 6724
rect 4580 6712 4586 6724
rect 5445 6715 5503 6721
rect 5445 6712 5457 6715
rect 4580 6684 5457 6712
rect 4580 6672 4586 6684
rect 5445 6681 5457 6684
rect 5491 6681 5503 6715
rect 5445 6675 5503 6681
rect 6264 6715 6322 6721
rect 6264 6681 6276 6715
rect 6310 6712 6322 6715
rect 6546 6712 6552 6724
rect 6310 6684 6552 6712
rect 6310 6681 6322 6684
rect 6264 6675 6322 6681
rect 6546 6672 6552 6684
rect 6604 6672 6610 6724
rect 2869 6647 2927 6653
rect 2869 6613 2881 6647
rect 2915 6644 2927 6647
rect 3234 6644 3240 6656
rect 2915 6616 3240 6644
rect 2915 6613 2927 6616
rect 2869 6607 2927 6613
rect 3234 6604 3240 6616
rect 3292 6604 3298 6656
rect 3694 6604 3700 6656
rect 3752 6644 3758 6656
rect 3881 6647 3939 6653
rect 3881 6644 3893 6647
rect 3752 6616 3893 6644
rect 3752 6604 3758 6616
rect 3881 6613 3893 6616
rect 3927 6613 3939 6647
rect 3881 6607 3939 6613
rect 3970 6604 3976 6656
rect 4028 6644 4034 6656
rect 4801 6647 4859 6653
rect 4801 6644 4813 6647
rect 4028 6616 4813 6644
rect 4028 6604 4034 6616
rect 4801 6613 4813 6616
rect 4847 6613 4859 6647
rect 5074 6644 5080 6656
rect 5035 6616 5080 6644
rect 4801 6607 4859 6613
rect 5074 6604 5080 6616
rect 5132 6604 5138 6656
rect 5166 6604 5172 6656
rect 5224 6644 5230 6656
rect 5537 6647 5595 6653
rect 5537 6644 5549 6647
rect 5224 6616 5549 6644
rect 5224 6604 5230 6616
rect 5537 6613 5549 6616
rect 5583 6644 5595 6647
rect 6454 6644 6460 6656
rect 5583 6616 6460 6644
rect 5583 6613 5595 6616
rect 5537 6607 5595 6613
rect 6454 6604 6460 6616
rect 6512 6604 6518 6656
rect 6822 6604 6828 6656
rect 6880 6644 6886 6656
rect 7392 6653 7420 6752
rect 7469 6749 7481 6752
rect 7515 6749 7527 6783
rect 7469 6743 7527 6749
rect 7653 6783 7711 6789
rect 7653 6749 7665 6783
rect 7699 6749 7711 6783
rect 7653 6743 7711 6749
rect 7929 6783 7987 6789
rect 7929 6749 7941 6783
rect 7975 6749 7987 6783
rect 7929 6743 7987 6749
rect 8389 6783 8447 6789
rect 8389 6749 8401 6783
rect 8435 6780 8447 6783
rect 8570 6780 8576 6792
rect 8435 6752 8576 6780
rect 8435 6749 8447 6752
rect 8389 6743 8447 6749
rect 7668 6712 7696 6743
rect 8570 6740 8576 6752
rect 8628 6780 8634 6792
rect 9030 6780 9036 6792
rect 8628 6752 9036 6780
rect 8628 6740 8634 6752
rect 9030 6740 9036 6752
rect 9088 6740 9094 6792
rect 9214 6780 9220 6792
rect 9175 6752 9220 6780
rect 9214 6740 9220 6752
rect 9272 6740 9278 6792
rect 9324 6780 9352 6820
rect 11514 6808 11520 6820
rect 11572 6808 11578 6860
rect 13630 6808 13636 6860
rect 13688 6848 13694 6860
rect 13909 6851 13967 6857
rect 13909 6848 13921 6851
rect 13688 6820 13921 6848
rect 13688 6808 13694 6820
rect 13909 6817 13921 6820
rect 13955 6817 13967 6851
rect 13909 6811 13967 6817
rect 11422 6780 11428 6792
rect 9324 6752 11284 6780
rect 11383 6752 11428 6780
rect 8662 6712 8668 6724
rect 7668 6684 8668 6712
rect 7377 6647 7435 6653
rect 7377 6644 7389 6647
rect 6880 6616 7389 6644
rect 6880 6604 6886 6616
rect 7377 6613 7389 6616
rect 7423 6613 7435 6647
rect 7377 6607 7435 6613
rect 7466 6604 7472 6656
rect 7524 6644 7530 6656
rect 7668 6644 7696 6684
rect 8662 6672 8668 6684
rect 8720 6672 8726 6724
rect 8757 6715 8815 6721
rect 8757 6681 8769 6715
rect 8803 6712 8815 6715
rect 9484 6715 9542 6721
rect 8803 6684 9444 6712
rect 8803 6681 8815 6684
rect 8757 6675 8815 6681
rect 7524 6616 7696 6644
rect 7745 6647 7803 6653
rect 7524 6604 7530 6616
rect 7745 6613 7757 6647
rect 7791 6644 7803 6647
rect 7834 6644 7840 6656
rect 7791 6616 7840 6644
rect 7791 6613 7803 6616
rect 7745 6607 7803 6613
rect 7834 6604 7840 6616
rect 7892 6604 7898 6656
rect 8478 6644 8484 6656
rect 8439 6616 8484 6644
rect 8478 6604 8484 6616
rect 8536 6604 8542 6656
rect 9033 6647 9091 6653
rect 9033 6613 9045 6647
rect 9079 6644 9091 6647
rect 9122 6644 9128 6656
rect 9079 6616 9128 6644
rect 9079 6613 9091 6616
rect 9033 6607 9091 6613
rect 9122 6604 9128 6616
rect 9180 6604 9186 6656
rect 9416 6644 9444 6684
rect 9484 6681 9496 6715
rect 9530 6712 9542 6715
rect 9582 6712 9588 6724
rect 9530 6684 9588 6712
rect 9530 6681 9542 6684
rect 9484 6675 9542 6681
rect 9582 6672 9588 6684
rect 9640 6672 9646 6724
rect 11146 6712 11152 6724
rect 10520 6684 11152 6712
rect 10520 6644 10548 6684
rect 11146 6672 11152 6684
rect 11204 6672 11210 6724
rect 9416 6616 10548 6644
rect 10873 6647 10931 6653
rect 10873 6613 10885 6647
rect 10919 6644 10931 6647
rect 10962 6644 10968 6656
rect 10919 6616 10968 6644
rect 10919 6613 10931 6616
rect 10873 6607 10931 6613
rect 10962 6604 10968 6616
rect 11020 6604 11026 6656
rect 11256 6644 11284 6752
rect 11422 6740 11428 6752
rect 11480 6740 11486 6792
rect 11606 6780 11612 6792
rect 11532 6752 11612 6780
rect 11330 6672 11336 6724
rect 11388 6712 11394 6724
rect 11532 6721 11560 6752
rect 11606 6740 11612 6752
rect 11664 6740 11670 6792
rect 14476 6789 14504 6876
rect 14461 6783 14519 6789
rect 14461 6749 14473 6783
rect 14507 6749 14519 6783
rect 14461 6743 14519 6749
rect 11517 6715 11575 6721
rect 11388 6684 11433 6712
rect 11388 6672 11394 6684
rect 11517 6681 11529 6715
rect 11563 6681 11575 6715
rect 11698 6712 11704 6724
rect 11659 6684 11704 6712
rect 11517 6675 11575 6681
rect 11698 6672 11704 6684
rect 11756 6672 11762 6724
rect 11790 6672 11796 6724
rect 11848 6712 11854 6724
rect 11885 6715 11943 6721
rect 11885 6712 11897 6715
rect 11848 6684 11897 6712
rect 11848 6672 11854 6684
rect 11885 6681 11897 6684
rect 11931 6681 11943 6715
rect 11885 6675 11943 6681
rect 12342 6672 12348 6724
rect 12400 6712 12406 6724
rect 12400 6684 12466 6712
rect 12400 6672 12406 6684
rect 13538 6672 13544 6724
rect 13596 6712 13602 6724
rect 13633 6715 13691 6721
rect 13633 6712 13645 6715
rect 13596 6684 13645 6712
rect 13596 6672 13602 6684
rect 13633 6681 13645 6684
rect 13679 6681 13691 6715
rect 13633 6675 13691 6681
rect 11425 6647 11483 6653
rect 11425 6644 11437 6647
rect 11256 6616 11437 6644
rect 11425 6613 11437 6616
rect 11471 6613 11483 6647
rect 14090 6644 14096 6656
rect 14051 6616 14096 6644
rect 11425 6607 11483 6613
rect 14090 6604 14096 6616
rect 14148 6604 14154 6656
rect 14277 6647 14335 6653
rect 14277 6613 14289 6647
rect 14323 6644 14335 6647
rect 14921 6647 14979 6653
rect 14921 6644 14933 6647
rect 14323 6616 14933 6644
rect 14323 6613 14335 6616
rect 14277 6607 14335 6613
rect 14921 6613 14933 6616
rect 14967 6613 14979 6647
rect 14921 6607 14979 6613
rect 1104 6554 14812 6576
rect 1104 6502 5547 6554
rect 5599 6502 5611 6554
rect 5663 6502 5675 6554
rect 5727 6502 5739 6554
rect 5791 6502 5803 6554
rect 5855 6502 10144 6554
rect 10196 6502 10208 6554
rect 10260 6502 10272 6554
rect 10324 6502 10336 6554
rect 10388 6502 10400 6554
rect 10452 6502 14812 6554
rect 1104 6480 14812 6502
rect 3142 6440 3148 6452
rect 3103 6412 3148 6440
rect 3142 6400 3148 6412
rect 3200 6400 3206 6452
rect 3602 6400 3608 6452
rect 3660 6440 3666 6452
rect 5074 6440 5080 6452
rect 3660 6412 4936 6440
rect 5035 6412 5080 6440
rect 3660 6400 3666 6412
rect 1670 6372 1676 6384
rect 1412 6344 1676 6372
rect 1412 6313 1440 6344
rect 1670 6332 1676 6344
rect 1728 6332 1734 6384
rect 2406 6332 2412 6384
rect 2464 6332 2470 6384
rect 3050 6332 3056 6384
rect 3108 6372 3114 6384
rect 4525 6375 4583 6381
rect 4525 6372 4537 6375
rect 3108 6344 4537 6372
rect 3108 6332 3114 6344
rect 4525 6341 4537 6344
rect 4571 6341 4583 6375
rect 4908 6372 4936 6412
rect 5074 6400 5080 6412
rect 5132 6400 5138 6452
rect 6733 6443 6791 6449
rect 6733 6440 6745 6443
rect 5184 6412 6745 6440
rect 5184 6372 5212 6412
rect 6733 6409 6745 6412
rect 6779 6409 6791 6443
rect 6733 6403 6791 6409
rect 6825 6443 6883 6449
rect 6825 6409 6837 6443
rect 6871 6440 6883 6443
rect 7374 6440 7380 6452
rect 6871 6412 7380 6440
rect 6871 6409 6883 6412
rect 6825 6403 6883 6409
rect 4908 6344 5212 6372
rect 5629 6375 5687 6381
rect 4525 6335 4583 6341
rect 5629 6341 5641 6375
rect 5675 6372 5687 6375
rect 5994 6372 6000 6384
rect 5675 6344 6000 6372
rect 5675 6341 5687 6344
rect 5629 6335 5687 6341
rect 5994 6332 6000 6344
rect 6052 6332 6058 6384
rect 6546 6332 6552 6384
rect 6604 6372 6610 6384
rect 6840 6372 6868 6403
rect 7374 6400 7380 6412
rect 7432 6400 7438 6452
rect 8570 6440 8576 6452
rect 7484 6412 8576 6440
rect 6604 6344 6868 6372
rect 6604 6332 6610 6344
rect 1397 6307 1455 6313
rect 1397 6273 1409 6307
rect 1443 6273 1455 6307
rect 3234 6304 3240 6316
rect 3195 6276 3240 6304
rect 1397 6267 1455 6273
rect 3234 6264 3240 6276
rect 3292 6264 3298 6316
rect 3329 6307 3387 6313
rect 3329 6273 3341 6307
rect 3375 6273 3387 6307
rect 3329 6267 3387 6273
rect 3513 6307 3571 6313
rect 3513 6273 3525 6307
rect 3559 6304 3571 6307
rect 3602 6304 3608 6316
rect 3559 6276 3608 6304
rect 3559 6273 3571 6276
rect 3513 6267 3571 6273
rect 1673 6239 1731 6245
rect 1673 6205 1685 6239
rect 1719 6236 1731 6239
rect 2314 6236 2320 6248
rect 1719 6208 2320 6236
rect 1719 6205 1731 6208
rect 1673 6199 1731 6205
rect 2314 6196 2320 6208
rect 2372 6196 2378 6248
rect 2958 6196 2964 6248
rect 3016 6236 3022 6248
rect 3344 6236 3372 6267
rect 3602 6264 3608 6276
rect 3660 6264 3666 6316
rect 3970 6304 3976 6316
rect 3931 6276 3976 6304
rect 3970 6264 3976 6276
rect 4028 6264 4034 6316
rect 4430 6304 4436 6316
rect 4391 6276 4436 6304
rect 4430 6264 4436 6276
rect 4488 6264 4494 6316
rect 4617 6307 4675 6313
rect 4617 6273 4629 6307
rect 4663 6304 4675 6307
rect 4798 6304 4804 6316
rect 4663 6276 4804 6304
rect 4663 6273 4675 6276
rect 4617 6267 4675 6273
rect 4798 6264 4804 6276
rect 4856 6264 4862 6316
rect 4908 6276 5304 6304
rect 3878 6236 3884 6248
rect 3016 6208 3884 6236
rect 3016 6196 3022 6208
rect 3878 6196 3884 6208
rect 3936 6196 3942 6248
rect 4065 6239 4123 6245
rect 4065 6205 4077 6239
rect 4111 6236 4123 6239
rect 4154 6236 4160 6248
rect 4111 6208 4160 6236
rect 4111 6205 4123 6208
rect 4065 6199 4123 6205
rect 4154 6196 4160 6208
rect 4212 6196 4218 6248
rect 4249 6239 4307 6245
rect 4249 6205 4261 6239
rect 4295 6236 4307 6239
rect 4908 6236 4936 6276
rect 5276 6248 5304 6276
rect 5350 6264 5356 6316
rect 5408 6304 5414 6316
rect 5537 6307 5595 6313
rect 5537 6304 5549 6307
rect 5408 6276 5549 6304
rect 5408 6264 5414 6276
rect 5537 6273 5549 6276
rect 5583 6273 5595 6307
rect 5810 6304 5816 6316
rect 5771 6276 5816 6304
rect 5537 6267 5595 6273
rect 5810 6264 5816 6276
rect 5868 6264 5874 6316
rect 5905 6307 5963 6313
rect 5905 6273 5917 6307
rect 5951 6273 5963 6307
rect 5905 6267 5963 6273
rect 7193 6307 7251 6313
rect 7193 6273 7205 6307
rect 7239 6273 7251 6307
rect 7374 6304 7380 6316
rect 7335 6276 7380 6304
rect 7193 6267 7251 6273
rect 4295 6208 4936 6236
rect 4295 6205 4307 6208
rect 4249 6199 4307 6205
rect 4982 6196 4988 6248
rect 5040 6236 5046 6248
rect 5166 6236 5172 6248
rect 5040 6208 5172 6236
rect 5040 6196 5046 6208
rect 5166 6196 5172 6208
rect 5224 6196 5230 6248
rect 5258 6196 5264 6248
rect 5316 6236 5322 6248
rect 5316 6208 5361 6236
rect 5316 6196 5322 6208
rect 5442 6196 5448 6248
rect 5500 6236 5506 6248
rect 5920 6236 5948 6267
rect 5500 6208 5948 6236
rect 5500 6196 5506 6208
rect 6086 6196 6092 6248
rect 6144 6236 6150 6248
rect 6917 6239 6975 6245
rect 6917 6236 6929 6239
rect 6144 6208 6929 6236
rect 6144 6196 6150 6208
rect 6917 6205 6929 6208
rect 6963 6205 6975 6239
rect 6917 6199 6975 6205
rect 2774 6128 2780 6180
rect 2832 6168 2838 6180
rect 3605 6171 3663 6177
rect 3605 6168 3617 6171
rect 2832 6140 3617 6168
rect 2832 6128 2838 6140
rect 3605 6137 3617 6140
rect 3651 6137 3663 6171
rect 5074 6168 5080 6180
rect 3605 6131 3663 6137
rect 4448 6140 5080 6168
rect 3421 6103 3479 6109
rect 3421 6069 3433 6103
rect 3467 6100 3479 6103
rect 4448 6100 4476 6140
rect 5074 6128 5080 6140
rect 5132 6128 5138 6180
rect 5721 6171 5779 6177
rect 5721 6137 5733 6171
rect 5767 6168 5779 6171
rect 5902 6168 5908 6180
rect 5767 6140 5908 6168
rect 5767 6137 5779 6140
rect 5721 6131 5779 6137
rect 5902 6128 5908 6140
rect 5960 6128 5966 6180
rect 7208 6168 7236 6267
rect 7374 6264 7380 6276
rect 7432 6264 7438 6316
rect 7484 6313 7512 6412
rect 8570 6400 8576 6412
rect 8628 6400 8634 6452
rect 11333 6443 11391 6449
rect 11333 6409 11345 6443
rect 11379 6440 11391 6443
rect 11698 6440 11704 6452
rect 11379 6412 11704 6440
rect 11379 6409 11391 6412
rect 11333 6403 11391 6409
rect 11698 6400 11704 6412
rect 11756 6400 11762 6452
rect 11977 6443 12035 6449
rect 11977 6409 11989 6443
rect 12023 6440 12035 6443
rect 12158 6440 12164 6452
rect 12023 6412 12164 6440
rect 12023 6409 12035 6412
rect 11977 6403 12035 6409
rect 12158 6400 12164 6412
rect 12216 6400 12222 6452
rect 14461 6443 14519 6449
rect 14461 6409 14473 6443
rect 14507 6440 14519 6443
rect 15013 6443 15071 6449
rect 15013 6440 15025 6443
rect 14507 6412 15025 6440
rect 14507 6409 14519 6412
rect 14461 6403 14519 6409
rect 15013 6409 15025 6412
rect 15059 6409 15071 6443
rect 15013 6403 15071 6409
rect 7834 6372 7840 6384
rect 7795 6344 7840 6372
rect 7834 6332 7840 6344
rect 7892 6332 7898 6384
rect 9122 6372 9128 6384
rect 9035 6344 9128 6372
rect 9122 6332 9128 6344
rect 9180 6372 9186 6384
rect 10042 6372 10048 6384
rect 9180 6344 10048 6372
rect 9180 6332 9186 6344
rect 10042 6332 10048 6344
rect 10100 6332 10106 6384
rect 10502 6332 10508 6384
rect 10560 6372 10566 6384
rect 13449 6375 13507 6381
rect 10560 6344 11928 6372
rect 10560 6332 10566 6344
rect 11900 6316 11928 6344
rect 13449 6341 13461 6375
rect 13495 6372 13507 6375
rect 14277 6375 14335 6381
rect 13495 6344 14228 6372
rect 13495 6341 13507 6344
rect 13449 6335 13507 6341
rect 7469 6307 7527 6313
rect 7469 6273 7481 6307
rect 7515 6273 7527 6307
rect 7469 6267 7527 6273
rect 9858 6264 9864 6316
rect 9916 6304 9922 6316
rect 10226 6313 10232 6316
rect 10220 6304 10232 6313
rect 9916 6276 9961 6304
rect 10187 6276 10232 6304
rect 9916 6264 9922 6276
rect 10220 6267 10232 6276
rect 10226 6264 10232 6267
rect 10284 6264 10290 6316
rect 11238 6264 11244 6316
rect 11296 6304 11302 6316
rect 11698 6304 11704 6316
rect 11296 6276 11704 6304
rect 11296 6264 11302 6276
rect 11698 6264 11704 6276
rect 11756 6264 11762 6316
rect 11882 6304 11888 6316
rect 11843 6276 11888 6304
rect 11882 6264 11888 6276
rect 11940 6264 11946 6316
rect 12342 6264 12348 6316
rect 12400 6264 12406 6316
rect 14200 6304 14228 6344
rect 14277 6341 14289 6375
rect 14323 6372 14335 6375
rect 15197 6375 15255 6381
rect 15197 6372 15209 6375
rect 14323 6344 15209 6372
rect 14323 6341 14335 6344
rect 14277 6335 14335 6341
rect 15197 6341 15209 6344
rect 15243 6341 15255 6375
rect 15197 6335 15255 6341
rect 15013 6307 15071 6313
rect 15013 6304 15025 6307
rect 14200 6276 15025 6304
rect 15013 6273 15025 6276
rect 15059 6273 15071 6307
rect 15013 6267 15071 6273
rect 7561 6239 7619 6245
rect 7561 6205 7573 6239
rect 7607 6205 7619 6239
rect 7561 6199 7619 6205
rect 7374 6168 7380 6180
rect 7208 6140 7380 6168
rect 7374 6128 7380 6140
rect 7432 6128 7438 6180
rect 3467 6072 4476 6100
rect 3467 6069 3479 6072
rect 3421 6063 3479 6069
rect 4614 6060 4620 6112
rect 4672 6100 4678 6112
rect 4709 6103 4767 6109
rect 4709 6100 4721 6103
rect 4672 6072 4721 6100
rect 4672 6060 4678 6072
rect 4709 6069 4721 6072
rect 4755 6069 4767 6103
rect 4709 6063 4767 6069
rect 5626 6060 5632 6112
rect 5684 6100 5690 6112
rect 5997 6103 6055 6109
rect 5997 6100 6009 6103
rect 5684 6072 6009 6100
rect 5684 6060 5690 6072
rect 5997 6069 6009 6072
rect 6043 6069 6055 6103
rect 5997 6063 6055 6069
rect 6086 6060 6092 6112
rect 6144 6100 6150 6112
rect 6365 6103 6423 6109
rect 6365 6100 6377 6103
rect 6144 6072 6377 6100
rect 6144 6060 6150 6072
rect 6365 6069 6377 6072
rect 6411 6069 6423 6103
rect 7466 6100 7472 6112
rect 7427 6072 7472 6100
rect 6365 6063 6423 6069
rect 7466 6060 7472 6072
rect 7524 6060 7530 6112
rect 7576 6100 7604 6199
rect 9030 6196 9036 6248
rect 9088 6236 9094 6248
rect 9585 6239 9643 6245
rect 9585 6236 9597 6239
rect 9088 6208 9597 6236
rect 9088 6196 9094 6208
rect 9585 6205 9597 6208
rect 9631 6205 9643 6239
rect 9585 6199 9643 6205
rect 9953 6239 10011 6245
rect 9953 6205 9965 6239
rect 9999 6205 10011 6239
rect 12360 6236 12388 6264
rect 9953 6199 10011 6205
rect 11532 6208 12388 6236
rect 9398 6128 9404 6180
rect 9456 6168 9462 6180
rect 9968 6168 9996 6199
rect 9456 6140 9996 6168
rect 9456 6128 9462 6140
rect 9214 6100 9220 6112
rect 7576 6072 9220 6100
rect 9214 6060 9220 6072
rect 9272 6100 9278 6112
rect 9416 6100 9444 6128
rect 9272 6072 9444 6100
rect 9272 6060 9278 6072
rect 9490 6060 9496 6112
rect 9548 6100 9554 6112
rect 9769 6103 9827 6109
rect 9769 6100 9781 6103
rect 9548 6072 9781 6100
rect 9548 6060 9554 6072
rect 9769 6069 9781 6072
rect 9815 6069 9827 6103
rect 9769 6063 9827 6069
rect 11422 6060 11428 6112
rect 11480 6100 11486 6112
rect 11532 6109 11560 6208
rect 13354 6196 13360 6248
rect 13412 6236 13418 6248
rect 13725 6239 13783 6245
rect 13725 6236 13737 6239
rect 13412 6208 13737 6236
rect 13412 6196 13418 6208
rect 13725 6205 13737 6208
rect 13771 6205 13783 6239
rect 13725 6199 13783 6205
rect 11885 6171 11943 6177
rect 11885 6137 11897 6171
rect 11931 6168 11943 6171
rect 12158 6168 12164 6180
rect 11931 6140 12164 6168
rect 11931 6137 11943 6140
rect 11885 6131 11943 6137
rect 12158 6128 12164 6140
rect 12216 6128 12222 6180
rect 14093 6171 14151 6177
rect 14093 6137 14105 6171
rect 14139 6168 14151 6171
rect 14458 6168 14464 6180
rect 14139 6140 14464 6168
rect 14139 6137 14151 6140
rect 14093 6131 14151 6137
rect 14458 6128 14464 6140
rect 14516 6128 14522 6180
rect 11517 6103 11575 6109
rect 11517 6100 11529 6103
rect 11480 6072 11529 6100
rect 11480 6060 11486 6072
rect 11517 6069 11529 6072
rect 11563 6069 11575 6103
rect 11517 6063 11575 6069
rect 13354 6060 13360 6112
rect 13412 6100 13418 6112
rect 13817 6103 13875 6109
rect 13817 6100 13829 6103
rect 13412 6072 13829 6100
rect 13412 6060 13418 6072
rect 13817 6069 13829 6072
rect 13863 6069 13875 6103
rect 13817 6063 13875 6069
rect 1104 6010 14812 6032
rect 1104 5958 3248 6010
rect 3300 5958 3312 6010
rect 3364 5958 3376 6010
rect 3428 5958 3440 6010
rect 3492 5958 3504 6010
rect 3556 5958 7846 6010
rect 7898 5958 7910 6010
rect 7962 5958 7974 6010
rect 8026 5958 8038 6010
rect 8090 5958 8102 6010
rect 8154 5958 12443 6010
rect 12495 5958 12507 6010
rect 12559 5958 12571 6010
rect 12623 5958 12635 6010
rect 12687 5958 12699 6010
rect 12751 5958 14812 6010
rect 1104 5936 14812 5958
rect 2038 5856 2044 5908
rect 2096 5896 2102 5908
rect 4614 5896 4620 5908
rect 2096 5868 4620 5896
rect 2096 5856 2102 5868
rect 4614 5856 4620 5868
rect 4672 5856 4678 5908
rect 4798 5896 4804 5908
rect 4759 5868 4804 5896
rect 4798 5856 4804 5868
rect 4856 5856 4862 5908
rect 5258 5856 5264 5908
rect 5316 5896 5322 5908
rect 5316 5868 6960 5896
rect 5316 5856 5322 5868
rect 2682 5788 2688 5840
rect 2740 5828 2746 5840
rect 3421 5831 3479 5837
rect 3421 5828 3433 5831
rect 2740 5800 3433 5828
rect 2740 5788 2746 5800
rect 3421 5797 3433 5800
rect 3467 5828 3479 5831
rect 4430 5828 4436 5840
rect 3467 5800 4436 5828
rect 3467 5797 3479 5800
rect 3421 5791 3479 5797
rect 1397 5763 1455 5769
rect 1397 5729 1409 5763
rect 1443 5760 1455 5763
rect 1670 5760 1676 5772
rect 1443 5732 1676 5760
rect 1443 5729 1455 5732
rect 1397 5723 1455 5729
rect 1670 5720 1676 5732
rect 1728 5720 1734 5772
rect 3234 5760 3240 5772
rect 2700 5732 3096 5760
rect 3195 5732 3240 5760
rect 2700 5704 2728 5732
rect 2682 5652 2688 5704
rect 2740 5652 2746 5704
rect 3068 5692 3096 5732
rect 3234 5720 3240 5732
rect 3292 5720 3298 5772
rect 4356 5769 4384 5800
rect 4430 5788 4436 5800
rect 4488 5788 4494 5840
rect 4341 5763 4399 5769
rect 4341 5729 4353 5763
rect 4387 5729 4399 5763
rect 4341 5723 4399 5729
rect 5445 5763 5503 5769
rect 5445 5729 5457 5763
rect 5491 5760 5503 5763
rect 5644 5760 5672 5868
rect 6932 5828 6960 5868
rect 7190 5856 7196 5908
rect 7248 5896 7254 5908
rect 7607 5899 7665 5905
rect 7607 5896 7619 5899
rect 7248 5868 7619 5896
rect 7248 5856 7254 5868
rect 7607 5865 7619 5868
rect 7653 5896 7665 5899
rect 9950 5896 9956 5908
rect 7653 5868 9956 5896
rect 7653 5865 7665 5868
rect 7607 5859 7665 5865
rect 9950 5856 9956 5868
rect 10008 5856 10014 5908
rect 12161 5899 12219 5905
rect 12161 5865 12173 5899
rect 12207 5896 12219 5899
rect 13538 5896 13544 5908
rect 12207 5868 13544 5896
rect 12207 5865 12219 5868
rect 12161 5859 12219 5865
rect 13538 5856 13544 5868
rect 13596 5856 13602 5908
rect 6932 5800 7696 5828
rect 7668 5772 7696 5800
rect 8018 5788 8024 5840
rect 8076 5828 8082 5840
rect 9490 5828 9496 5840
rect 8076 5800 9496 5828
rect 8076 5788 8082 5800
rect 9490 5788 9496 5800
rect 9548 5788 9554 5840
rect 11977 5831 12035 5837
rect 11977 5828 11989 5831
rect 10796 5800 11989 5828
rect 5491 5732 5672 5760
rect 5721 5763 5779 5769
rect 5491 5729 5503 5732
rect 5445 5723 5503 5729
rect 5721 5729 5733 5763
rect 5767 5760 5779 5763
rect 6730 5760 6736 5772
rect 5767 5732 6736 5760
rect 5767 5729 5779 5732
rect 5721 5723 5779 5729
rect 6730 5720 6736 5732
rect 6788 5760 6794 5772
rect 6788 5732 7144 5760
rect 6788 5720 6794 5732
rect 3513 5695 3571 5701
rect 3513 5692 3525 5695
rect 3068 5664 3525 5692
rect 3513 5661 3525 5664
rect 3559 5692 3571 5695
rect 4062 5692 4068 5704
rect 3559 5664 4068 5692
rect 3559 5661 3571 5664
rect 3513 5655 3571 5661
rect 4062 5652 4068 5664
rect 4120 5652 4126 5704
rect 4614 5692 4620 5704
rect 4575 5664 4620 5692
rect 4614 5652 4620 5664
rect 4672 5652 4678 5704
rect 5626 5652 5632 5704
rect 5684 5692 5690 5704
rect 5802 5695 5860 5701
rect 5802 5692 5814 5695
rect 5684 5664 5814 5692
rect 5684 5652 5690 5664
rect 5802 5661 5814 5664
rect 5848 5661 5860 5695
rect 6086 5692 6092 5704
rect 5802 5655 5860 5661
rect 5920 5664 6092 5692
rect 1673 5627 1731 5633
rect 1673 5593 1685 5627
rect 1719 5593 1731 5627
rect 1673 5587 1731 5593
rect 1688 5556 1716 5587
rect 2406 5584 2412 5636
rect 2464 5584 2470 5636
rect 3237 5627 3295 5633
rect 3237 5624 3249 5627
rect 2976 5596 3249 5624
rect 2976 5556 3004 5596
rect 3237 5593 3249 5596
rect 3283 5593 3295 5627
rect 3237 5587 3295 5593
rect 5169 5627 5227 5633
rect 5169 5593 5181 5627
rect 5215 5624 5227 5627
rect 5920 5624 5948 5664
rect 6086 5652 6092 5664
rect 6144 5652 6150 5704
rect 6178 5652 6184 5704
rect 6236 5692 6242 5704
rect 6236 5664 6281 5692
rect 6236 5652 6242 5664
rect 7116 5636 7144 5732
rect 7650 5720 7656 5772
rect 7708 5720 7714 5772
rect 7742 5720 7748 5772
rect 7800 5760 7806 5772
rect 8297 5763 8355 5769
rect 8297 5760 8309 5763
rect 7800 5732 8309 5760
rect 7800 5720 7806 5732
rect 7944 5701 7972 5732
rect 8297 5729 8309 5732
rect 8343 5729 8355 5763
rect 8662 5760 8668 5772
rect 8575 5732 8668 5760
rect 8297 5723 8355 5729
rect 8662 5720 8668 5732
rect 8720 5760 8726 5772
rect 8846 5760 8852 5772
rect 8720 5732 8852 5760
rect 8720 5720 8726 5732
rect 8846 5720 8852 5732
rect 8904 5720 8910 5772
rect 8987 5763 9045 5769
rect 8987 5729 8999 5763
rect 9033 5760 9045 5763
rect 9214 5760 9220 5772
rect 9033 5732 9220 5760
rect 9033 5729 9045 5732
rect 8987 5723 9045 5729
rect 9214 5720 9220 5732
rect 9272 5720 9278 5772
rect 9398 5720 9404 5772
rect 9456 5760 9462 5772
rect 9582 5760 9588 5772
rect 9456 5732 9588 5760
rect 9456 5720 9462 5732
rect 9582 5720 9588 5732
rect 9640 5760 9646 5772
rect 10796 5769 10824 5800
rect 11977 5797 11989 5800
rect 12023 5828 12035 5831
rect 12066 5828 12072 5840
rect 12023 5800 12072 5828
rect 12023 5797 12035 5800
rect 11977 5791 12035 5797
rect 12066 5788 12072 5800
rect 12124 5828 12130 5840
rect 12618 5828 12624 5840
rect 12124 5800 12624 5828
rect 12124 5788 12130 5800
rect 12618 5788 12624 5800
rect 12676 5788 12682 5840
rect 10781 5763 10839 5769
rect 10781 5760 10793 5763
rect 9640 5732 10793 5760
rect 9640 5720 9646 5732
rect 10781 5729 10793 5732
rect 10827 5729 10839 5763
rect 10781 5723 10839 5729
rect 10962 5720 10968 5772
rect 11020 5760 11026 5772
rect 11425 5763 11483 5769
rect 11020 5732 11284 5760
rect 11020 5720 11026 5732
rect 7837 5695 7895 5701
rect 7837 5661 7849 5695
rect 7883 5661 7895 5695
rect 7837 5655 7895 5661
rect 7929 5695 7987 5701
rect 7929 5661 7941 5695
rect 7975 5661 7987 5695
rect 7929 5655 7987 5661
rect 5215 5596 5948 5624
rect 5215 5593 5227 5596
rect 5169 5587 5227 5593
rect 7098 5584 7104 5636
rect 7156 5584 7162 5636
rect 1688 5528 3004 5556
rect 3050 5516 3056 5568
rect 3108 5556 3114 5568
rect 3145 5559 3203 5565
rect 3145 5556 3157 5559
rect 3108 5528 3157 5556
rect 3108 5516 3114 5528
rect 3145 5525 3157 5528
rect 3191 5556 3203 5559
rect 3602 5556 3608 5568
rect 3191 5528 3608 5556
rect 3191 5525 3203 5528
rect 3145 5519 3203 5525
rect 3602 5516 3608 5528
rect 3660 5516 3666 5568
rect 4798 5516 4804 5568
rect 4856 5556 4862 5568
rect 5261 5559 5319 5565
rect 5261 5556 5273 5559
rect 4856 5528 5273 5556
rect 4856 5516 4862 5528
rect 5261 5525 5273 5528
rect 5307 5556 5319 5559
rect 6730 5556 6736 5568
rect 5307 5528 6736 5556
rect 5307 5525 5319 5528
rect 5261 5519 5319 5525
rect 6730 5516 6736 5528
rect 6788 5516 6794 5568
rect 7852 5556 7880 5655
rect 8018 5652 8024 5704
rect 8076 5692 8082 5704
rect 8481 5695 8539 5701
rect 8076 5664 8121 5692
rect 8076 5652 8082 5664
rect 8481 5661 8493 5695
rect 8527 5692 8539 5695
rect 8570 5692 8576 5704
rect 8527 5664 8576 5692
rect 8527 5661 8539 5664
rect 8481 5655 8539 5661
rect 8570 5652 8576 5664
rect 8628 5652 8634 5704
rect 8754 5692 8760 5704
rect 8715 5664 8760 5692
rect 8754 5652 8760 5664
rect 8812 5652 8818 5704
rect 10413 5695 10471 5701
rect 10413 5661 10425 5695
rect 10459 5692 10471 5695
rect 10502 5692 10508 5704
rect 10459 5664 10508 5692
rect 10459 5661 10471 5664
rect 10413 5655 10471 5661
rect 10502 5652 10508 5664
rect 10560 5652 10566 5704
rect 10870 5692 10876 5704
rect 10831 5664 10876 5692
rect 10870 5652 10876 5664
rect 10928 5652 10934 5704
rect 11054 5692 11060 5704
rect 11015 5664 11060 5692
rect 11054 5652 11060 5664
rect 11112 5652 11118 5704
rect 11256 5692 11284 5732
rect 11425 5729 11437 5763
rect 11471 5760 11483 5763
rect 13630 5760 13636 5772
rect 11471 5732 13636 5760
rect 11471 5729 11483 5732
rect 11425 5723 11483 5729
rect 13630 5720 13636 5732
rect 13688 5760 13694 5772
rect 13909 5763 13967 5769
rect 13909 5760 13921 5763
rect 13688 5732 13921 5760
rect 13688 5720 13694 5732
rect 13909 5729 13921 5732
rect 13955 5729 13967 5763
rect 13909 5723 13967 5729
rect 11609 5695 11667 5701
rect 11609 5692 11621 5695
rect 11256 5664 11621 5692
rect 11609 5661 11621 5664
rect 11655 5661 11667 5695
rect 14458 5692 14464 5704
rect 14419 5664 14464 5692
rect 11609 5655 11667 5661
rect 14458 5652 14464 5664
rect 14516 5652 14522 5704
rect 8205 5627 8263 5633
rect 8205 5593 8217 5627
rect 8251 5624 8263 5627
rect 8251 5618 9168 5624
rect 9214 5618 9220 5636
rect 8251 5596 9220 5618
rect 8251 5593 8263 5596
rect 8205 5587 8263 5593
rect 9140 5590 9220 5596
rect 9214 5584 9220 5590
rect 9272 5584 9278 5636
rect 10042 5584 10048 5636
rect 10100 5584 10106 5636
rect 11790 5624 11796 5636
rect 11751 5596 11796 5624
rect 11790 5584 11796 5596
rect 11848 5584 11854 5636
rect 13633 5627 13691 5633
rect 8386 5556 8392 5568
rect 7852 5528 8392 5556
rect 8386 5516 8392 5528
rect 8444 5516 8450 5568
rect 10060 5556 10088 5584
rect 11422 5556 11428 5568
rect 10060 5528 11428 5556
rect 11422 5516 11428 5528
rect 11480 5556 11486 5568
rect 12452 5556 12480 5610
rect 13633 5593 13645 5627
rect 13679 5624 13691 5627
rect 14921 5627 14979 5633
rect 14921 5624 14933 5627
rect 13679 5596 14933 5624
rect 13679 5593 13691 5596
rect 13633 5587 13691 5593
rect 14921 5593 14933 5596
rect 14967 5593 14979 5627
rect 14921 5587 14979 5593
rect 13354 5556 13360 5568
rect 11480 5528 13360 5556
rect 11480 5516 11486 5528
rect 13354 5516 13360 5528
rect 13412 5556 13418 5568
rect 14090 5556 14096 5568
rect 13412 5528 14096 5556
rect 13412 5516 13418 5528
rect 14090 5516 14096 5528
rect 14148 5516 14154 5568
rect 14182 5516 14188 5568
rect 14240 5556 14246 5568
rect 14277 5559 14335 5565
rect 14277 5556 14289 5559
rect 14240 5528 14289 5556
rect 14240 5516 14246 5528
rect 14277 5525 14289 5528
rect 14323 5525 14335 5559
rect 14277 5519 14335 5525
rect 1104 5466 14812 5488
rect 1104 5414 5547 5466
rect 5599 5414 5611 5466
rect 5663 5414 5675 5466
rect 5727 5414 5739 5466
rect 5791 5414 5803 5466
rect 5855 5414 10144 5466
rect 10196 5414 10208 5466
rect 10260 5414 10272 5466
rect 10324 5414 10336 5466
rect 10388 5414 10400 5466
rect 10452 5414 14812 5466
rect 1104 5392 14812 5414
rect 2501 5355 2559 5361
rect 2501 5321 2513 5355
rect 2547 5352 2559 5355
rect 3234 5352 3240 5364
rect 2547 5324 3240 5352
rect 2547 5321 2559 5324
rect 2501 5315 2559 5321
rect 3234 5312 3240 5324
rect 3292 5312 3298 5364
rect 3329 5355 3387 5361
rect 3329 5321 3341 5355
rect 3375 5352 3387 5355
rect 3789 5355 3847 5361
rect 3375 5324 3556 5352
rect 3375 5321 3387 5324
rect 3329 5315 3387 5321
rect 2682 5284 2688 5296
rect 2332 5256 2688 5284
rect 1670 5216 1676 5228
rect 1631 5188 1676 5216
rect 1670 5176 1676 5188
rect 1728 5176 1734 5228
rect 2332 5225 2360 5256
rect 2682 5244 2688 5256
rect 2740 5244 2746 5296
rect 3252 5256 3464 5284
rect 2317 5219 2375 5225
rect 2317 5185 2329 5219
rect 2363 5185 2375 5219
rect 2498 5216 2504 5228
rect 2459 5188 2504 5216
rect 2317 5179 2375 5185
rect 2498 5176 2504 5188
rect 2556 5176 2562 5228
rect 2777 5219 2835 5225
rect 2777 5216 2789 5219
rect 2608 5188 2789 5216
rect 2608 5080 2636 5188
rect 2777 5185 2789 5188
rect 2823 5185 2835 5219
rect 2777 5179 2835 5185
rect 2869 5219 2927 5225
rect 2869 5185 2881 5219
rect 2915 5216 2927 5219
rect 2958 5216 2964 5228
rect 2915 5188 2964 5216
rect 2915 5185 2927 5188
rect 2869 5179 2927 5185
rect 2958 5176 2964 5188
rect 3016 5176 3022 5228
rect 3053 5219 3111 5225
rect 3053 5185 3065 5219
rect 3099 5185 3111 5219
rect 3053 5179 3111 5185
rect 3145 5219 3203 5225
rect 3145 5185 3157 5219
rect 3191 5216 3203 5219
rect 3252 5216 3280 5256
rect 3191 5188 3280 5216
rect 3329 5219 3387 5225
rect 3191 5185 3203 5188
rect 3145 5179 3203 5185
rect 3329 5185 3341 5219
rect 3375 5185 3387 5219
rect 3329 5179 3387 5185
rect 2682 5108 2688 5160
rect 2740 5148 2746 5160
rect 2740 5120 2785 5148
rect 2740 5108 2746 5120
rect 2866 5080 2872 5092
rect 2608 5052 2872 5080
rect 2866 5040 2872 5052
rect 2924 5040 2930 5092
rect 3068 5080 3096 5179
rect 3234 5108 3240 5160
rect 3292 5148 3298 5160
rect 3344 5148 3372 5179
rect 3292 5120 3372 5148
rect 3436 5148 3464 5256
rect 3528 5225 3556 5324
rect 3789 5321 3801 5355
rect 3835 5352 3847 5355
rect 3970 5352 3976 5364
rect 3835 5324 3976 5352
rect 3835 5321 3847 5324
rect 3789 5315 3847 5321
rect 3970 5312 3976 5324
rect 4028 5312 4034 5364
rect 4062 5312 4068 5364
rect 4120 5352 4126 5364
rect 4157 5355 4215 5361
rect 4157 5352 4169 5355
rect 4120 5324 4169 5352
rect 4120 5312 4126 5324
rect 4157 5321 4169 5324
rect 4203 5321 4215 5355
rect 5353 5355 5411 5361
rect 5353 5352 5365 5355
rect 4157 5315 4215 5321
rect 4908 5324 5365 5352
rect 4908 5293 4936 5324
rect 5353 5321 5365 5324
rect 5399 5321 5411 5355
rect 5353 5315 5411 5321
rect 5902 5312 5908 5364
rect 5960 5312 5966 5364
rect 6914 5352 6920 5364
rect 6104 5324 6920 5352
rect 4893 5287 4951 5293
rect 4893 5253 4905 5287
rect 4939 5253 4951 5287
rect 5920 5284 5948 5312
rect 6104 5293 6132 5324
rect 6914 5312 6920 5324
rect 6972 5312 6978 5364
rect 7009 5355 7067 5361
rect 7009 5321 7021 5355
rect 7055 5352 7067 5355
rect 7282 5352 7288 5364
rect 7055 5324 7288 5352
rect 7055 5321 7067 5324
rect 7009 5315 7067 5321
rect 7282 5312 7288 5324
rect 7340 5312 7346 5364
rect 10502 5352 10508 5364
rect 9872 5324 10180 5352
rect 10463 5324 10508 5352
rect 4893 5247 4951 5253
rect 5000 5256 5948 5284
rect 6089 5287 6147 5293
rect 3513 5219 3571 5225
rect 3513 5185 3525 5219
rect 3559 5216 3571 5219
rect 3602 5216 3608 5228
rect 3559 5188 3608 5216
rect 3559 5185 3571 5188
rect 3513 5179 3571 5185
rect 3602 5176 3608 5188
rect 3660 5176 3666 5228
rect 3694 5176 3700 5228
rect 3752 5216 3758 5228
rect 3752 5188 3797 5216
rect 3752 5176 3758 5188
rect 4154 5176 4160 5228
rect 4212 5216 4218 5228
rect 4249 5219 4307 5225
rect 4249 5216 4261 5219
rect 4212 5188 4261 5216
rect 4212 5176 4218 5188
rect 4249 5185 4261 5188
rect 4295 5216 4307 5219
rect 4522 5216 4528 5228
rect 4295 5188 4528 5216
rect 4295 5185 4307 5188
rect 4249 5179 4307 5185
rect 4522 5176 4528 5188
rect 4580 5176 4586 5228
rect 4706 5216 4712 5228
rect 4667 5188 4712 5216
rect 4706 5176 4712 5188
rect 4764 5176 4770 5228
rect 5000 5225 5028 5256
rect 6089 5253 6101 5287
rect 6135 5253 6147 5287
rect 7190 5284 7196 5296
rect 6089 5247 6147 5253
rect 6564 5256 7196 5284
rect 4985 5219 5043 5225
rect 4985 5185 4997 5219
rect 5031 5185 5043 5219
rect 4985 5179 5043 5185
rect 5074 5176 5080 5228
rect 5132 5216 5138 5228
rect 5258 5216 5264 5228
rect 5132 5188 5177 5216
rect 5219 5188 5264 5216
rect 5132 5176 5138 5188
rect 5258 5176 5264 5188
rect 5316 5216 5322 5228
rect 5629 5219 5687 5225
rect 5629 5216 5641 5219
rect 5316 5188 5641 5216
rect 5316 5176 5322 5188
rect 5629 5185 5641 5188
rect 5675 5185 5687 5219
rect 5810 5216 5816 5228
rect 5771 5188 5816 5216
rect 5629 5179 5687 5185
rect 5810 5176 5816 5188
rect 5868 5176 5874 5228
rect 5902 5176 5908 5228
rect 5960 5216 5966 5228
rect 6181 5219 6239 5225
rect 5960 5188 6005 5216
rect 5960 5176 5966 5188
rect 6181 5185 6193 5219
rect 6227 5216 6239 5219
rect 6270 5216 6276 5228
rect 6227 5188 6276 5216
rect 6227 5185 6239 5188
rect 6181 5179 6239 5185
rect 6270 5176 6276 5188
rect 6328 5176 6334 5228
rect 6564 5225 6592 5256
rect 7190 5244 7196 5256
rect 7248 5244 7254 5296
rect 7558 5244 7564 5296
rect 7616 5284 7622 5296
rect 8294 5284 8300 5296
rect 7616 5256 8300 5284
rect 7616 5244 7622 5256
rect 8294 5244 8300 5256
rect 8352 5244 8358 5296
rect 8386 5244 8392 5296
rect 8444 5284 8450 5296
rect 8444 5256 9168 5284
rect 8444 5244 8450 5256
rect 6549 5219 6607 5225
rect 6549 5185 6561 5219
rect 6595 5185 6607 5219
rect 6822 5216 6828 5228
rect 6783 5188 6828 5216
rect 6549 5179 6607 5185
rect 6822 5176 6828 5188
rect 6880 5176 6886 5228
rect 6914 5176 6920 5228
rect 6972 5216 6978 5228
rect 7101 5219 7159 5225
rect 7101 5216 7113 5219
rect 6972 5188 7113 5216
rect 6972 5176 6978 5188
rect 7101 5185 7113 5188
rect 7147 5216 7159 5219
rect 8478 5216 8484 5228
rect 7147 5188 8484 5216
rect 7147 5185 7159 5188
rect 7101 5179 7159 5185
rect 8478 5176 8484 5188
rect 8536 5176 8542 5228
rect 8846 5176 8852 5228
rect 8904 5216 8910 5228
rect 9140 5225 9168 5256
rect 9214 5244 9220 5296
rect 9272 5284 9278 5296
rect 9872 5290 9900 5324
rect 9692 5284 9900 5290
rect 9272 5262 9900 5284
rect 10152 5284 10180 5324
rect 10502 5312 10508 5324
rect 10560 5312 10566 5364
rect 11514 5352 11520 5364
rect 11475 5324 11520 5352
rect 11514 5312 11520 5324
rect 11572 5312 11578 5364
rect 11974 5352 11980 5364
rect 11935 5324 11980 5352
rect 11974 5312 11980 5324
rect 12032 5312 12038 5364
rect 9272 5256 9720 5262
rect 10152 5256 10456 5284
rect 9272 5244 9278 5256
rect 8941 5219 8999 5225
rect 8941 5216 8953 5219
rect 8904 5188 8953 5216
rect 8904 5176 8910 5188
rect 8941 5185 8953 5188
rect 8987 5185 8999 5219
rect 8941 5179 8999 5185
rect 9125 5219 9183 5225
rect 9125 5185 9137 5219
rect 9171 5185 9183 5219
rect 9125 5179 9183 5185
rect 9493 5219 9551 5225
rect 9674 5220 9680 5228
rect 9493 5185 9505 5219
rect 9539 5216 9551 5219
rect 9600 5216 9680 5220
rect 9539 5192 9680 5216
rect 9539 5188 9628 5192
rect 9539 5185 9551 5188
rect 9493 5179 9551 5185
rect 9674 5176 9680 5192
rect 9732 5176 9738 5228
rect 10428 5225 10456 5256
rect 13354 5244 13360 5296
rect 13412 5244 13418 5296
rect 9953 5219 10011 5225
rect 9953 5216 9965 5219
rect 9876 5188 9965 5216
rect 9876 5160 9904 5188
rect 9953 5185 9965 5188
rect 9999 5185 10011 5219
rect 9953 5179 10011 5185
rect 10413 5219 10471 5225
rect 10413 5185 10425 5219
rect 10459 5185 10471 5219
rect 10413 5179 10471 5185
rect 10502 5176 10508 5228
rect 10560 5216 10566 5228
rect 10560 5188 10605 5216
rect 10560 5176 10566 5188
rect 10686 5176 10692 5228
rect 10744 5216 10750 5228
rect 10965 5219 11023 5225
rect 10744 5188 10789 5216
rect 10744 5176 10750 5188
rect 10965 5185 10977 5219
rect 11011 5216 11023 5219
rect 11885 5219 11943 5225
rect 11885 5216 11897 5219
rect 11011 5188 11897 5216
rect 11011 5185 11023 5188
rect 10965 5179 11023 5185
rect 11885 5185 11897 5188
rect 11931 5216 11943 5219
rect 11974 5216 11980 5228
rect 11931 5188 11980 5216
rect 11931 5185 11943 5188
rect 11885 5179 11943 5185
rect 11974 5176 11980 5188
rect 12032 5176 12038 5228
rect 12066 5176 12072 5228
rect 12124 5216 12130 5228
rect 12337 5219 12395 5225
rect 12337 5216 12349 5219
rect 12124 5188 12349 5216
rect 12124 5176 12130 5188
rect 12337 5185 12349 5188
rect 12383 5185 12395 5219
rect 12337 5179 12395 5185
rect 12434 5176 12440 5228
rect 12492 5216 12498 5228
rect 12529 5219 12587 5225
rect 12529 5216 12541 5219
rect 12492 5188 12541 5216
rect 12492 5176 12498 5188
rect 12529 5185 12541 5188
rect 12575 5185 12587 5219
rect 12529 5179 12587 5185
rect 12618 5176 12624 5228
rect 12676 5216 12682 5228
rect 12676 5188 12721 5216
rect 12676 5176 12682 5188
rect 13814 5176 13820 5228
rect 13872 5216 13878 5228
rect 14415 5219 14473 5225
rect 14415 5216 14427 5219
rect 13872 5188 14427 5216
rect 13872 5176 13878 5188
rect 14415 5185 14427 5188
rect 14461 5185 14473 5219
rect 14415 5179 14473 5185
rect 3786 5148 3792 5160
rect 3436 5120 3792 5148
rect 3292 5108 3298 5120
rect 3786 5108 3792 5120
rect 3844 5108 3850 5160
rect 4433 5151 4491 5157
rect 4433 5117 4445 5151
rect 4479 5148 4491 5151
rect 4890 5148 4896 5160
rect 4479 5120 4896 5148
rect 4479 5117 4491 5120
rect 4433 5111 4491 5117
rect 4890 5108 4896 5120
rect 4948 5108 4954 5160
rect 5537 5151 5595 5157
rect 5537 5117 5549 5151
rect 5583 5148 5595 5151
rect 5994 5148 6000 5160
rect 5583 5120 6000 5148
rect 5583 5117 5595 5120
rect 5537 5111 5595 5117
rect 5994 5108 6000 5120
rect 6052 5148 6058 5160
rect 6457 5151 6515 5157
rect 6457 5148 6469 5151
rect 6052 5120 6469 5148
rect 6052 5108 6058 5120
rect 6457 5117 6469 5120
rect 6503 5117 6515 5151
rect 6457 5111 6515 5117
rect 6641 5151 6699 5157
rect 6641 5117 6653 5151
rect 6687 5148 6699 5151
rect 6730 5148 6736 5160
rect 6687 5120 6736 5148
rect 6687 5117 6699 5120
rect 6641 5111 6699 5117
rect 4154 5080 4160 5092
rect 3068 5052 3188 5080
rect 1394 4972 1400 5024
rect 1452 5012 1458 5024
rect 1581 5015 1639 5021
rect 1581 5012 1593 5015
rect 1452 4984 1593 5012
rect 1452 4972 1458 4984
rect 1581 4981 1593 4984
rect 1627 4981 1639 5015
rect 1581 4975 1639 4981
rect 2225 5015 2283 5021
rect 2225 4981 2237 5015
rect 2271 5012 2283 5015
rect 2406 5012 2412 5024
rect 2271 4984 2412 5012
rect 2271 4981 2283 4984
rect 2225 4975 2283 4981
rect 2406 4972 2412 4984
rect 2464 5012 2470 5024
rect 2682 5012 2688 5024
rect 2464 4984 2688 5012
rect 2464 4972 2470 4984
rect 2682 4972 2688 4984
rect 2740 4972 2746 5024
rect 3050 5012 3056 5024
rect 3011 4984 3056 5012
rect 3050 4972 3056 4984
rect 3108 4972 3114 5024
rect 3160 5012 3188 5052
rect 3436 5052 4160 5080
rect 3436 5012 3464 5052
rect 4154 5040 4160 5052
rect 4212 5040 4218 5092
rect 4985 5083 5043 5089
rect 4985 5049 4997 5083
rect 5031 5080 5043 5083
rect 6086 5080 6092 5092
rect 5031 5052 6092 5080
rect 5031 5049 5043 5052
rect 4985 5043 5043 5049
rect 6086 5040 6092 5052
rect 6144 5040 6150 5092
rect 6546 5040 6552 5092
rect 6604 5080 6610 5092
rect 6656 5080 6684 5111
rect 6730 5108 6736 5120
rect 6788 5108 6794 5160
rect 7558 5108 7564 5160
rect 7616 5148 7622 5160
rect 8662 5148 8668 5160
rect 7616 5120 8668 5148
rect 7616 5108 7622 5120
rect 8662 5108 8668 5120
rect 8720 5108 8726 5160
rect 9858 5108 9864 5160
rect 9916 5108 9922 5160
rect 10042 5148 10048 5160
rect 10003 5120 10048 5148
rect 10042 5108 10048 5120
rect 10100 5108 10106 5160
rect 10778 5108 10784 5160
rect 10836 5148 10842 5160
rect 10873 5151 10931 5157
rect 10873 5148 10885 5151
rect 10836 5120 10885 5148
rect 10836 5108 10842 5120
rect 10873 5117 10885 5120
rect 10919 5117 10931 5151
rect 12158 5148 12164 5160
rect 12119 5120 12164 5148
rect 10873 5111 10931 5117
rect 12158 5108 12164 5120
rect 12216 5108 12222 5160
rect 12989 5151 13047 5157
rect 12989 5148 13001 5151
rect 12636 5120 13001 5148
rect 6604 5052 6684 5080
rect 6604 5040 6610 5052
rect 7006 5040 7012 5092
rect 7064 5080 7070 5092
rect 7650 5080 7656 5092
rect 7064 5052 7656 5080
rect 7064 5040 7070 5052
rect 7650 5040 7656 5052
rect 7708 5040 7714 5092
rect 9766 5080 9772 5092
rect 8404 5052 9772 5080
rect 3160 4984 3464 5012
rect 3513 5015 3571 5021
rect 3513 4981 3525 5015
rect 3559 5012 3571 5015
rect 5350 5012 5356 5024
rect 3559 4984 5356 5012
rect 3559 4981 3571 4984
rect 3513 4975 3571 4981
rect 5350 4972 5356 4984
rect 5408 4972 5414 5024
rect 5718 5012 5724 5024
rect 5679 4984 5724 5012
rect 5718 4972 5724 4984
rect 5776 4972 5782 5024
rect 6181 5015 6239 5021
rect 6181 4981 6193 5015
rect 6227 5012 6239 5015
rect 6362 5012 6368 5024
rect 6227 4984 6368 5012
rect 6227 4981 6239 4984
rect 6181 4975 6239 4981
rect 6362 4972 6368 4984
rect 6420 4972 6426 5024
rect 6454 4972 6460 5024
rect 6512 5012 6518 5024
rect 7558 5012 7564 5024
rect 6512 4984 7564 5012
rect 6512 4972 6518 4984
rect 7558 4972 7564 4984
rect 7616 4972 7622 5024
rect 8202 4972 8208 5024
rect 8260 5012 8266 5024
rect 8404 5021 8432 5052
rect 9766 5040 9772 5052
rect 9824 5040 9830 5092
rect 12636 5080 12664 5120
rect 12989 5117 13001 5120
rect 13035 5117 13047 5151
rect 12989 5111 13047 5117
rect 11900 5052 12664 5080
rect 8389 5015 8447 5021
rect 8389 5012 8401 5015
rect 8260 4984 8401 5012
rect 8260 4972 8266 4984
rect 8389 4981 8401 4984
rect 8435 4981 8447 5015
rect 8389 4975 8447 4981
rect 9125 5015 9183 5021
rect 9125 4981 9137 5015
rect 9171 5012 9183 5015
rect 9306 5012 9312 5024
rect 9171 4984 9312 5012
rect 9171 4981 9183 4984
rect 9125 4975 9183 4981
rect 9306 4972 9312 4984
rect 9364 4972 9370 5024
rect 9401 5015 9459 5021
rect 9401 4981 9413 5015
rect 9447 5012 9459 5015
rect 9490 5012 9496 5024
rect 9447 4984 9496 5012
rect 9447 4981 9459 4984
rect 9401 4975 9459 4981
rect 9490 4972 9496 4984
rect 9548 4972 9554 5024
rect 9677 5015 9735 5021
rect 9677 4981 9689 5015
rect 9723 5012 9735 5015
rect 10134 5012 10140 5024
rect 9723 4984 10140 5012
rect 9723 4981 9735 4984
rect 9677 4975 9735 4981
rect 10134 4972 10140 4984
rect 10192 4972 10198 5024
rect 10229 5015 10287 5021
rect 10229 4981 10241 5015
rect 10275 5012 10287 5015
rect 11054 5012 11060 5024
rect 10275 4984 11060 5012
rect 10275 4981 10287 4984
rect 10229 4975 10287 4981
rect 11054 4972 11060 4984
rect 11112 4972 11118 5024
rect 11241 5015 11299 5021
rect 11241 4981 11253 5015
rect 11287 5012 11299 5015
rect 11900 5012 11928 5052
rect 11287 4984 11928 5012
rect 12437 5015 12495 5021
rect 11287 4981 11299 4984
rect 11241 4975 11299 4981
rect 12437 4981 12449 5015
rect 12483 5012 12495 5015
rect 12894 5012 12900 5024
rect 12483 4984 12900 5012
rect 12483 4981 12495 4984
rect 12437 4975 12495 4981
rect 12894 4972 12900 4984
rect 12952 4972 12958 5024
rect 1104 4922 14812 4944
rect 1104 4870 3248 4922
rect 3300 4870 3312 4922
rect 3364 4870 3376 4922
rect 3428 4870 3440 4922
rect 3492 4870 3504 4922
rect 3556 4870 7846 4922
rect 7898 4870 7910 4922
rect 7962 4870 7974 4922
rect 8026 4870 8038 4922
rect 8090 4870 8102 4922
rect 8154 4870 12443 4922
rect 12495 4870 12507 4922
rect 12559 4870 12571 4922
rect 12623 4870 12635 4922
rect 12687 4870 12699 4922
rect 12751 4870 14812 4922
rect 1104 4848 14812 4870
rect 3142 4768 3148 4820
rect 3200 4808 3206 4820
rect 3329 4811 3387 4817
rect 3329 4808 3341 4811
rect 3200 4780 3341 4808
rect 3200 4768 3206 4780
rect 3329 4777 3341 4780
rect 3375 4777 3387 4811
rect 3329 4771 3387 4777
rect 4801 4811 4859 4817
rect 4801 4777 4813 4811
rect 4847 4808 4859 4811
rect 5258 4808 5264 4820
rect 4847 4780 5264 4808
rect 4847 4777 4859 4780
rect 4801 4771 4859 4777
rect 5258 4768 5264 4780
rect 5316 4768 5322 4820
rect 6270 4768 6276 4820
rect 6328 4808 6334 4820
rect 6733 4811 6791 4817
rect 6733 4808 6745 4811
rect 6328 4780 6745 4808
rect 6328 4768 6334 4780
rect 6733 4777 6745 4780
rect 6779 4808 6791 4811
rect 7098 4808 7104 4820
rect 6779 4780 7104 4808
rect 6779 4777 6791 4780
rect 6733 4771 6791 4777
rect 7098 4768 7104 4780
rect 7156 4808 7162 4820
rect 8846 4808 8852 4820
rect 7156 4780 8852 4808
rect 7156 4768 7162 4780
rect 8846 4768 8852 4780
rect 8904 4768 8910 4820
rect 9306 4768 9312 4820
rect 9364 4808 9370 4820
rect 10686 4808 10692 4820
rect 9364 4780 10692 4808
rect 9364 4768 9370 4780
rect 10686 4768 10692 4780
rect 10744 4768 10750 4820
rect 11054 4768 11060 4820
rect 11112 4808 11118 4820
rect 11655 4811 11713 4817
rect 11655 4808 11667 4811
rect 11112 4780 11667 4808
rect 11112 4768 11118 4780
rect 11655 4777 11667 4780
rect 11701 4808 11713 4811
rect 12342 4808 12348 4820
rect 11701 4780 12348 4808
rect 11701 4777 11713 4780
rect 11655 4771 11713 4777
rect 12342 4768 12348 4780
rect 12400 4768 12406 4820
rect 14090 4808 14096 4820
rect 14051 4780 14096 4808
rect 14090 4768 14096 4780
rect 14148 4768 14154 4820
rect 2682 4700 2688 4752
rect 2740 4740 2746 4752
rect 3513 4743 3571 4749
rect 3513 4740 3525 4743
rect 2740 4712 3525 4740
rect 2740 4700 2746 4712
rect 3513 4709 3525 4712
rect 3559 4709 3571 4743
rect 3513 4703 3571 4709
rect 4706 4700 4712 4752
rect 4764 4740 4770 4752
rect 8941 4743 8999 4749
rect 8941 4740 8953 4743
rect 4764 4712 5948 4740
rect 4764 4700 4770 4712
rect 5920 4684 5948 4712
rect 7484 4712 8953 4740
rect 1397 4675 1455 4681
rect 1397 4641 1409 4675
rect 1443 4672 1455 4675
rect 1670 4672 1676 4684
rect 1443 4644 1676 4672
rect 1443 4641 1455 4644
rect 1397 4635 1455 4641
rect 1670 4632 1676 4644
rect 1728 4632 1734 4684
rect 3050 4632 3056 4684
rect 3108 4672 3114 4684
rect 4617 4675 4675 4681
rect 4617 4672 4629 4675
rect 3108 4644 4629 4672
rect 3108 4632 3114 4644
rect 4617 4641 4629 4644
rect 4663 4641 4675 4675
rect 4890 4672 4896 4684
rect 4851 4644 4896 4672
rect 4617 4635 4675 4641
rect 4890 4632 4896 4644
rect 4948 4632 4954 4684
rect 5629 4675 5687 4681
rect 5629 4672 5641 4675
rect 5276 4644 5641 4672
rect 3237 4607 3295 4613
rect 3237 4604 3249 4607
rect 3160 4576 3249 4604
rect 1673 4539 1731 4545
rect 1673 4505 1685 4539
rect 1719 4536 1731 4539
rect 1762 4536 1768 4548
rect 1719 4508 1768 4536
rect 1719 4505 1731 4508
rect 1673 4499 1731 4505
rect 1762 4496 1768 4508
rect 1820 4496 1826 4548
rect 2682 4496 2688 4548
rect 2740 4496 2746 4548
rect 2958 4428 2964 4480
rect 3016 4468 3022 4480
rect 3160 4477 3188 4576
rect 3237 4573 3249 4576
rect 3283 4573 3295 4607
rect 3237 4567 3295 4573
rect 3973 4607 4031 4613
rect 3973 4573 3985 4607
rect 4019 4604 4031 4607
rect 4154 4604 4160 4616
rect 4019 4576 4160 4604
rect 4019 4573 4031 4576
rect 3973 4567 4031 4573
rect 4154 4564 4160 4576
rect 4212 4564 4218 4616
rect 4338 4604 4344 4616
rect 4299 4576 4344 4604
rect 4338 4564 4344 4576
rect 4396 4564 4402 4616
rect 4522 4564 4528 4616
rect 4580 4604 4586 4616
rect 4709 4607 4767 4613
rect 4709 4604 4721 4607
rect 4580 4576 4721 4604
rect 4580 4564 4586 4576
rect 4709 4573 4721 4576
rect 4755 4573 4767 4607
rect 4709 4567 4767 4573
rect 4798 4564 4804 4616
rect 4856 4604 4862 4616
rect 4985 4607 5043 4613
rect 4985 4604 4997 4607
rect 4856 4576 4997 4604
rect 4856 4564 4862 4576
rect 4985 4573 4997 4576
rect 5031 4573 5043 4607
rect 4985 4567 5043 4573
rect 5166 4564 5172 4616
rect 5224 4604 5230 4616
rect 5276 4613 5304 4644
rect 5629 4641 5641 4644
rect 5675 4672 5687 4675
rect 5810 4672 5816 4684
rect 5675 4644 5816 4672
rect 5675 4641 5687 4644
rect 5629 4635 5687 4641
rect 5810 4632 5816 4644
rect 5868 4632 5874 4684
rect 5902 4632 5908 4684
rect 5960 4672 5966 4684
rect 7374 4672 7380 4684
rect 5960 4644 7380 4672
rect 5960 4632 5966 4644
rect 7374 4632 7380 4644
rect 7432 4632 7438 4684
rect 5261 4607 5319 4613
rect 5261 4604 5273 4607
rect 5224 4576 5273 4604
rect 5224 4564 5230 4576
rect 5261 4573 5273 4576
rect 5307 4573 5319 4607
rect 5261 4567 5319 4573
rect 5353 4607 5411 4613
rect 5353 4573 5365 4607
rect 5399 4573 5411 4607
rect 5353 4567 5411 4573
rect 5537 4607 5595 4613
rect 5537 4573 5549 4607
rect 5583 4604 5595 4607
rect 6730 4604 6736 4616
rect 5583 4576 6736 4604
rect 5583 4573 5595 4576
rect 5537 4567 5595 4573
rect 3694 4496 3700 4548
rect 3752 4536 3758 4548
rect 5368 4536 5396 4567
rect 6730 4564 6736 4576
rect 6788 4564 6794 4616
rect 7006 4564 7012 4616
rect 7064 4564 7070 4616
rect 7484 4613 7512 4712
rect 8941 4709 8953 4712
rect 8987 4709 8999 4743
rect 8941 4703 8999 4709
rect 7558 4632 7564 4684
rect 7616 4672 7622 4684
rect 7616 4644 7661 4672
rect 7616 4632 7622 4644
rect 7742 4632 7748 4684
rect 7800 4672 7806 4684
rect 8205 4675 8263 4681
rect 7800 4644 7845 4672
rect 7800 4632 7806 4644
rect 8205 4641 8217 4675
rect 8251 4672 8263 4675
rect 8294 4672 8300 4684
rect 8251 4644 8300 4672
rect 8251 4641 8263 4644
rect 8205 4635 8263 4641
rect 8294 4632 8300 4644
rect 8352 4632 8358 4684
rect 8665 4675 8723 4681
rect 8665 4641 8677 4675
rect 8711 4672 8723 4675
rect 9490 4672 9496 4684
rect 8711 4644 9496 4672
rect 8711 4641 8723 4644
rect 8665 4635 8723 4641
rect 9490 4632 9496 4644
rect 9548 4632 9554 4684
rect 10134 4632 10140 4684
rect 10192 4672 10198 4684
rect 10229 4675 10287 4681
rect 10229 4672 10241 4675
rect 10192 4644 10241 4672
rect 10192 4632 10198 4644
rect 10229 4641 10241 4644
rect 10275 4641 10287 4675
rect 10502 4672 10508 4684
rect 10229 4635 10287 4641
rect 10336 4644 10508 4672
rect 7469 4607 7527 4613
rect 7469 4573 7481 4607
rect 7515 4573 7527 4607
rect 7469 4567 7527 4573
rect 7650 4564 7656 4616
rect 7708 4604 7714 4616
rect 8113 4607 8171 4613
rect 8113 4604 8125 4607
rect 7708 4576 8125 4604
rect 7708 4564 7714 4576
rect 8113 4573 8125 4576
rect 8159 4573 8171 4607
rect 8113 4567 8171 4573
rect 8386 4564 8392 4616
rect 8444 4604 8450 4616
rect 8573 4607 8631 4613
rect 8573 4604 8585 4607
rect 8444 4576 8585 4604
rect 8444 4564 8450 4576
rect 8573 4573 8585 4576
rect 8619 4573 8631 4607
rect 9309 4607 9367 4613
rect 9309 4604 9321 4607
rect 8573 4567 8631 4573
rect 8956 4576 9321 4604
rect 6641 4539 6699 4545
rect 6641 4536 6653 4539
rect 3752 4508 5396 4536
rect 3752 4496 3758 4508
rect 3145 4471 3203 4477
rect 3145 4468 3157 4471
rect 3016 4440 3157 4468
rect 3016 4428 3022 4440
rect 3145 4437 3157 4440
rect 3191 4437 3203 4471
rect 3145 4431 3203 4437
rect 3234 4428 3240 4480
rect 3292 4468 3298 4480
rect 3786 4468 3792 4480
rect 3292 4440 3792 4468
rect 3292 4428 3298 4440
rect 3786 4428 3792 4440
rect 3844 4468 3850 4480
rect 3881 4471 3939 4477
rect 3881 4468 3893 4471
rect 3844 4440 3893 4468
rect 3844 4428 3850 4440
rect 3881 4437 3893 4440
rect 3927 4437 3939 4471
rect 4246 4468 4252 4480
rect 4207 4440 4252 4468
rect 3881 4431 3939 4437
rect 4246 4428 4252 4440
rect 4304 4428 4310 4480
rect 5368 4468 5396 4508
rect 5920 4508 6653 4536
rect 5920 4480 5948 4508
rect 6641 4505 6653 4508
rect 6687 4505 6699 4539
rect 7024 4536 7052 4564
rect 8956 4536 8984 4576
rect 9309 4573 9321 4576
rect 9355 4573 9367 4607
rect 9309 4567 9367 4573
rect 9582 4564 9588 4616
rect 9640 4604 9646 4616
rect 9861 4607 9919 4613
rect 9861 4604 9873 4607
rect 9640 4576 9873 4604
rect 9640 4564 9646 4576
rect 9861 4573 9873 4576
rect 9907 4573 9919 4607
rect 10336 4604 10364 4644
rect 10502 4632 10508 4644
rect 10560 4632 10566 4684
rect 13630 4632 13636 4684
rect 13688 4672 13694 4684
rect 13909 4675 13967 4681
rect 13909 4672 13921 4675
rect 13688 4644 13921 4672
rect 13688 4632 13694 4644
rect 13909 4641 13921 4644
rect 13955 4672 13967 4675
rect 14366 4672 14372 4684
rect 13955 4644 14372 4672
rect 13955 4641 13967 4644
rect 13909 4635 13967 4641
rect 14366 4632 14372 4644
rect 14424 4632 14430 4684
rect 13538 4604 13544 4616
rect 9861 4567 9919 4573
rect 9968 4576 10364 4604
rect 13499 4576 13544 4604
rect 9968 4536 9996 4576
rect 13538 4564 13544 4576
rect 13596 4564 13602 4616
rect 14458 4604 14464 4616
rect 14419 4576 14464 4604
rect 14458 4564 14464 4576
rect 14516 4564 14522 4616
rect 11422 4536 11428 4548
rect 6641 4499 6699 4505
rect 6932 4508 7052 4536
rect 8496 4508 8984 4536
rect 9324 4508 9996 4536
rect 11270 4508 11428 4536
rect 5902 4468 5908 4480
rect 5368 4440 5908 4468
rect 5902 4428 5908 4440
rect 5960 4428 5966 4480
rect 6822 4428 6828 4480
rect 6880 4468 6886 4480
rect 6932 4477 6960 4508
rect 6917 4471 6975 4477
rect 6917 4468 6929 4471
rect 6880 4440 6929 4468
rect 6880 4428 6886 4440
rect 6917 4437 6929 4440
rect 6963 4437 6975 4471
rect 6917 4431 6975 4437
rect 7006 4428 7012 4480
rect 7064 4468 7070 4480
rect 8496 4477 8524 4508
rect 7101 4471 7159 4477
rect 7101 4468 7113 4471
rect 7064 4440 7113 4468
rect 7064 4428 7070 4440
rect 7101 4437 7113 4440
rect 7147 4437 7159 4471
rect 7101 4431 7159 4437
rect 8481 4471 8539 4477
rect 8481 4437 8493 4471
rect 8527 4437 8539 4471
rect 8481 4431 8539 4437
rect 8570 4428 8576 4480
rect 8628 4468 8634 4480
rect 9324 4468 9352 4508
rect 11422 4496 11428 4508
rect 11480 4536 11486 4548
rect 11480 4508 12558 4536
rect 11480 4496 11486 4508
rect 8628 4440 9352 4468
rect 9401 4471 9459 4477
rect 8628 4428 8634 4440
rect 9401 4437 9413 4471
rect 9447 4468 9459 4471
rect 11793 4471 11851 4477
rect 11793 4468 11805 4471
rect 9447 4440 11805 4468
rect 9447 4437 9459 4440
rect 9401 4431 9459 4437
rect 11793 4437 11805 4440
rect 11839 4468 11851 4471
rect 11882 4468 11888 4480
rect 11839 4440 11888 4468
rect 11839 4437 11851 4440
rect 11793 4431 11851 4437
rect 11882 4428 11888 4440
rect 11940 4428 11946 4480
rect 14182 4428 14188 4480
rect 14240 4468 14246 4480
rect 14277 4471 14335 4477
rect 14277 4468 14289 4471
rect 14240 4440 14289 4468
rect 14240 4428 14246 4440
rect 14277 4437 14289 4440
rect 14323 4437 14335 4471
rect 14277 4431 14335 4437
rect 1104 4378 14812 4400
rect 1104 4326 5547 4378
rect 5599 4326 5611 4378
rect 5663 4326 5675 4378
rect 5727 4326 5739 4378
rect 5791 4326 5803 4378
rect 5855 4326 10144 4378
rect 10196 4326 10208 4378
rect 10260 4326 10272 4378
rect 10324 4326 10336 4378
rect 10388 4326 10400 4378
rect 10452 4326 14812 4378
rect 1104 4304 14812 4326
rect 1762 4224 1768 4276
rect 1820 4264 1826 4276
rect 3605 4267 3663 4273
rect 3605 4264 3617 4267
rect 1820 4236 3617 4264
rect 1820 4224 1826 4236
rect 3605 4233 3617 4236
rect 3651 4233 3663 4267
rect 3605 4227 3663 4233
rect 4801 4267 4859 4273
rect 4801 4233 4813 4267
rect 4847 4233 4859 4267
rect 4801 4227 4859 4233
rect 5629 4267 5687 4273
rect 5629 4233 5641 4267
rect 5675 4264 5687 4267
rect 5902 4264 5908 4276
rect 5675 4236 5908 4264
rect 5675 4233 5687 4236
rect 5629 4227 5687 4233
rect 2682 4156 2688 4208
rect 2740 4156 2746 4208
rect 3191 4199 3249 4205
rect 3191 4165 3203 4199
rect 3237 4196 3249 4199
rect 4154 4196 4160 4208
rect 3237 4168 4160 4196
rect 3237 4165 3249 4168
rect 3191 4159 3249 4165
rect 4154 4156 4160 4168
rect 4212 4156 4218 4208
rect 4816 4140 4844 4227
rect 5902 4224 5908 4236
rect 5960 4224 5966 4276
rect 6362 4264 6368 4276
rect 6323 4236 6368 4264
rect 6362 4224 6368 4236
rect 6420 4224 6426 4276
rect 7466 4224 7472 4276
rect 7524 4264 7530 4276
rect 7561 4267 7619 4273
rect 7561 4264 7573 4267
rect 7524 4236 7573 4264
rect 7524 4224 7530 4236
rect 7561 4233 7573 4236
rect 7607 4233 7619 4267
rect 8570 4264 8576 4276
rect 7561 4227 7619 4233
rect 7668 4236 8576 4264
rect 5169 4199 5227 4205
rect 5169 4165 5181 4199
rect 5215 4196 5227 4199
rect 6638 4196 6644 4208
rect 5215 4168 6644 4196
rect 5215 4165 5227 4168
rect 5169 4159 5227 4165
rect 6638 4156 6644 4168
rect 6696 4156 6702 4208
rect 7190 4196 7196 4208
rect 7151 4168 7196 4196
rect 7190 4156 7196 4168
rect 7248 4156 7254 4208
rect 7374 4196 7380 4208
rect 7287 4168 7380 4196
rect 7374 4156 7380 4168
rect 7432 4196 7438 4208
rect 7668 4196 7696 4236
rect 8570 4224 8576 4236
rect 8628 4224 8634 4276
rect 8665 4267 8723 4273
rect 8665 4233 8677 4267
rect 8711 4264 8723 4267
rect 9125 4267 9183 4273
rect 9125 4264 9137 4267
rect 8711 4236 9137 4264
rect 8711 4233 8723 4236
rect 8665 4227 8723 4233
rect 9125 4233 9137 4236
rect 9171 4233 9183 4267
rect 9125 4227 9183 4233
rect 9493 4267 9551 4273
rect 9493 4233 9505 4267
rect 9539 4264 9551 4267
rect 10137 4267 10195 4273
rect 10137 4264 10149 4267
rect 9539 4236 10149 4264
rect 9539 4233 9551 4236
rect 9493 4227 9551 4233
rect 10137 4233 10149 4236
rect 10183 4233 10195 4267
rect 10137 4227 10195 4233
rect 10781 4267 10839 4273
rect 10781 4233 10793 4267
rect 10827 4264 10839 4267
rect 11517 4267 11575 4273
rect 11517 4264 11529 4267
rect 10827 4236 11529 4264
rect 10827 4233 10839 4236
rect 10781 4227 10839 4233
rect 11517 4233 11529 4236
rect 11563 4233 11575 4267
rect 11882 4264 11888 4276
rect 11843 4236 11888 4264
rect 11517 4227 11575 4233
rect 11882 4224 11888 4236
rect 11940 4224 11946 4276
rect 12575 4267 12633 4273
rect 12575 4233 12587 4267
rect 12621 4264 12633 4267
rect 13538 4264 13544 4276
rect 12621 4236 13544 4264
rect 12621 4233 12633 4236
rect 12575 4227 12633 4233
rect 13538 4224 13544 4236
rect 13596 4224 13602 4276
rect 7432 4168 7696 4196
rect 7432 4156 7438 4168
rect 7742 4156 7748 4208
rect 7800 4196 7806 4208
rect 7800 4168 8156 4196
rect 7800 4156 7806 4168
rect 1394 4128 1400 4140
rect 1355 4100 1400 4128
rect 1394 4088 1400 4100
rect 1452 4088 1458 4140
rect 2958 4088 2964 4140
rect 3016 4128 3022 4140
rect 3329 4131 3387 4137
rect 3329 4128 3341 4131
rect 3016 4100 3341 4128
rect 3016 4088 3022 4100
rect 3329 4097 3341 4100
rect 3375 4097 3387 4131
rect 3329 4091 3387 4097
rect 3421 4131 3479 4137
rect 3421 4097 3433 4131
rect 3467 4128 3479 4131
rect 3510 4128 3516 4140
rect 3467 4100 3516 4128
rect 3467 4097 3479 4100
rect 3421 4091 3479 4097
rect 3510 4088 3516 4100
rect 3568 4088 3574 4140
rect 3602 4088 3608 4140
rect 3660 4128 3666 4140
rect 3697 4131 3755 4137
rect 3697 4128 3709 4131
rect 3660 4100 3709 4128
rect 3660 4088 3666 4100
rect 3697 4097 3709 4100
rect 3743 4097 3755 4131
rect 3878 4128 3884 4140
rect 3839 4100 3884 4128
rect 3697 4091 3755 4097
rect 3878 4088 3884 4100
rect 3936 4088 3942 4140
rect 4709 4131 4767 4137
rect 4709 4128 4721 4131
rect 4172 4100 4721 4128
rect 1765 4063 1823 4069
rect 1765 4029 1777 4063
rect 1811 4060 1823 4063
rect 2774 4060 2780 4072
rect 1811 4032 2780 4060
rect 1811 4029 1823 4032
rect 1765 4023 1823 4029
rect 2774 4020 2780 4032
rect 2832 4020 2838 4072
rect 4172 4001 4200 4100
rect 4709 4097 4721 4100
rect 4755 4128 4767 4131
rect 4798 4128 4804 4140
rect 4755 4100 4804 4128
rect 4755 4097 4767 4100
rect 4709 4091 4767 4097
rect 4798 4088 4804 4100
rect 4856 4088 4862 4140
rect 5258 4128 5264 4140
rect 5219 4100 5264 4128
rect 5258 4088 5264 4100
rect 5316 4088 5322 4140
rect 5905 4131 5963 4137
rect 5905 4097 5917 4131
rect 5951 4128 5963 4131
rect 6546 4128 6552 4140
rect 5951 4100 6552 4128
rect 5951 4097 5963 4100
rect 5905 4091 5963 4097
rect 6546 4088 6552 4100
rect 6604 4088 6610 4140
rect 6733 4131 6791 4137
rect 6733 4097 6745 4131
rect 6779 4128 6791 4131
rect 7006 4128 7012 4140
rect 6779 4100 7012 4128
rect 6779 4097 6791 4100
rect 6733 4091 6791 4097
rect 7006 4088 7012 4100
rect 7064 4088 7070 4140
rect 7098 4088 7104 4140
rect 7156 4128 7162 4140
rect 8021 4131 8079 4137
rect 8021 4128 8033 4131
rect 7156 4100 7201 4128
rect 7392 4100 8033 4128
rect 7156 4088 7162 4100
rect 4338 4020 4344 4072
rect 4396 4060 4402 4072
rect 4433 4063 4491 4069
rect 4433 4060 4445 4063
rect 4396 4032 4445 4060
rect 4396 4020 4402 4032
rect 4433 4029 4445 4032
rect 4479 4029 4491 4063
rect 4433 4023 4491 4029
rect 5350 4020 5356 4072
rect 5408 4060 5414 4072
rect 5408 4032 5453 4060
rect 5408 4020 5414 4032
rect 5534 4020 5540 4072
rect 5592 4060 5598 4072
rect 5629 4063 5687 4069
rect 5629 4060 5641 4063
rect 5592 4032 5641 4060
rect 5592 4020 5598 4032
rect 5629 4029 5641 4032
rect 5675 4029 5687 4063
rect 5629 4023 5687 4029
rect 5813 4063 5871 4069
rect 5813 4029 5825 4063
rect 5859 4060 5871 4063
rect 6454 4060 6460 4072
rect 5859 4032 6460 4060
rect 5859 4029 5871 4032
rect 5813 4023 5871 4029
rect 6454 4020 6460 4032
rect 6512 4020 6518 4072
rect 6638 4020 6644 4072
rect 6696 4060 6702 4072
rect 6825 4063 6883 4069
rect 6825 4060 6837 4063
rect 6696 4032 6837 4060
rect 6696 4020 6702 4032
rect 6825 4029 6837 4032
rect 6871 4060 6883 4063
rect 7392 4060 7420 4100
rect 8021 4097 8033 4100
rect 8067 4097 8079 4131
rect 8128 4128 8156 4168
rect 8294 4156 8300 4208
rect 8352 4196 8358 4208
rect 8352 4168 9812 4196
rect 8352 4156 8358 4168
rect 8202 4128 8208 4140
rect 8128 4100 8208 4128
rect 8021 4091 8079 4097
rect 8202 4088 8208 4100
rect 8260 4128 8266 4140
rect 8260 4100 8984 4128
rect 8260 4088 8266 4100
rect 6871 4032 7420 4060
rect 7929 4063 7987 4069
rect 6871 4029 6883 4032
rect 6825 4023 6883 4029
rect 7929 4029 7941 4063
rect 7975 4029 7987 4063
rect 7929 4023 7987 4029
rect 4157 3995 4215 4001
rect 4157 3961 4169 3995
rect 4203 3961 4215 3995
rect 4157 3955 4215 3961
rect 4522 3952 4528 4004
rect 4580 3992 4586 4004
rect 6914 3992 6920 4004
rect 4580 3964 6920 3992
rect 4580 3952 4586 3964
rect 6914 3952 6920 3964
rect 6972 3952 6978 4004
rect 7944 3992 7972 4023
rect 8478 4020 8484 4072
rect 8536 4060 8542 4072
rect 8956 4069 8984 4100
rect 9490 4088 9496 4140
rect 9548 4128 9554 4140
rect 9784 4128 9812 4168
rect 12342 4156 12348 4208
rect 12400 4196 12406 4208
rect 12400 4168 13018 4196
rect 12400 4156 12406 4168
rect 9953 4131 10011 4137
rect 9953 4128 9965 4131
rect 9548 4100 9720 4128
rect 9784 4100 9965 4128
rect 9548 4088 9554 4100
rect 8757 4063 8815 4069
rect 8757 4060 8769 4063
rect 8536 4032 8769 4060
rect 8536 4020 8542 4032
rect 8757 4029 8769 4032
rect 8803 4029 8815 4063
rect 8757 4023 8815 4029
rect 8941 4063 8999 4069
rect 8941 4029 8953 4063
rect 8987 4060 8999 4063
rect 9030 4060 9036 4072
rect 8987 4032 9036 4060
rect 8987 4029 8999 4032
rect 8941 4023 8999 4029
rect 8297 3995 8355 4001
rect 8297 3992 8309 3995
rect 7944 3964 8309 3992
rect 8297 3961 8309 3964
rect 8343 3961 8355 3995
rect 8772 3992 8800 4023
rect 9030 4020 9036 4032
rect 9088 4020 9094 4072
rect 9692 4069 9720 4100
rect 9953 4097 9965 4100
rect 9999 4097 10011 4131
rect 9953 4091 10011 4097
rect 10502 4088 10508 4140
rect 10560 4128 10566 4140
rect 10873 4131 10931 4137
rect 10873 4128 10885 4131
rect 10560 4100 10885 4128
rect 10560 4088 10566 4100
rect 10873 4097 10885 4100
rect 10919 4128 10931 4131
rect 11054 4128 11060 4140
rect 10919 4100 11060 4128
rect 10919 4097 10931 4100
rect 10873 4091 10931 4097
rect 11054 4088 11060 4100
rect 11112 4088 11118 4140
rect 14001 4131 14059 4137
rect 14001 4097 14013 4131
rect 14047 4128 14059 4131
rect 14090 4128 14096 4140
rect 14047 4100 14096 4128
rect 14047 4097 14059 4100
rect 14001 4091 14059 4097
rect 14090 4088 14096 4100
rect 14148 4088 14154 4140
rect 14366 4128 14372 4140
rect 14327 4100 14372 4128
rect 14366 4088 14372 4100
rect 14424 4088 14430 4140
rect 9585 4063 9643 4069
rect 9585 4029 9597 4063
rect 9631 4029 9643 4063
rect 9585 4023 9643 4029
rect 9677 4063 9735 4069
rect 9677 4029 9689 4063
rect 9723 4029 9735 4063
rect 9677 4023 9735 4029
rect 10965 4063 11023 4069
rect 10965 4029 10977 4063
rect 11011 4060 11023 4063
rect 11330 4060 11336 4072
rect 11011 4032 11336 4060
rect 11011 4029 11023 4032
rect 10965 4023 11023 4029
rect 9600 3992 9628 4023
rect 8772 3964 9628 3992
rect 8297 3955 8355 3961
rect 3970 3924 3976 3936
rect 3931 3896 3976 3924
rect 3970 3884 3976 3896
rect 4028 3884 4034 3936
rect 4062 3884 4068 3936
rect 4120 3924 4126 3936
rect 4617 3927 4675 3933
rect 4617 3924 4629 3927
rect 4120 3896 4629 3924
rect 4120 3884 4126 3896
rect 4617 3893 4629 3896
rect 4663 3893 4675 3927
rect 4617 3887 4675 3893
rect 6089 3927 6147 3933
rect 6089 3893 6101 3927
rect 6135 3924 6147 3927
rect 6822 3924 6828 3936
rect 6135 3896 6828 3924
rect 6135 3893 6147 3896
rect 6089 3887 6147 3893
rect 6822 3884 6828 3896
rect 6880 3884 6886 3936
rect 7006 3924 7012 3936
rect 6967 3896 7012 3924
rect 7006 3884 7012 3896
rect 7064 3884 7070 3936
rect 7098 3884 7104 3936
rect 7156 3924 7162 3936
rect 7156 3896 7201 3924
rect 7156 3884 7162 3896
rect 7742 3884 7748 3936
rect 7800 3924 7806 3936
rect 8205 3927 8263 3933
rect 8205 3924 8217 3927
rect 7800 3896 8217 3924
rect 7800 3884 7806 3896
rect 8205 3893 8217 3896
rect 8251 3893 8263 3927
rect 9600 3924 9628 3964
rect 9766 3952 9772 4004
rect 9824 3992 9830 4004
rect 10413 3995 10471 4001
rect 10413 3992 10425 3995
rect 9824 3964 10425 3992
rect 9824 3952 9830 3964
rect 10413 3961 10425 3964
rect 10459 3961 10471 3995
rect 10413 3955 10471 3961
rect 9674 3924 9680 3936
rect 9600 3896 9680 3924
rect 8205 3887 8263 3893
rect 9674 3884 9680 3896
rect 9732 3924 9738 3936
rect 10980 3924 11008 4023
rect 11330 4020 11336 4032
rect 11388 4020 11394 4072
rect 11974 4060 11980 4072
rect 11935 4032 11980 4060
rect 11974 4020 11980 4032
rect 12032 4020 12038 4072
rect 12161 4063 12219 4069
rect 12161 4029 12173 4063
rect 12207 4060 12219 4063
rect 12894 4060 12900 4072
rect 12207 4032 12900 4060
rect 12207 4029 12219 4032
rect 12161 4023 12219 4029
rect 12894 4020 12900 4032
rect 12952 4020 12958 4072
rect 11054 3924 11060 3936
rect 9732 3896 11060 3924
rect 9732 3884 9738 3896
rect 11054 3884 11060 3896
rect 11112 3884 11118 3936
rect 11333 3927 11391 3933
rect 11333 3893 11345 3927
rect 11379 3924 11391 3927
rect 11422 3924 11428 3936
rect 11379 3896 11428 3924
rect 11379 3893 11391 3896
rect 11333 3887 11391 3893
rect 11422 3884 11428 3896
rect 11480 3924 11486 3936
rect 12342 3924 12348 3936
rect 11480 3896 12348 3924
rect 11480 3884 11486 3896
rect 12342 3884 12348 3896
rect 12400 3884 12406 3936
rect 1104 3834 14812 3856
rect 1104 3782 3248 3834
rect 3300 3782 3312 3834
rect 3364 3782 3376 3834
rect 3428 3782 3440 3834
rect 3492 3782 3504 3834
rect 3556 3782 7846 3834
rect 7898 3782 7910 3834
rect 7962 3782 7974 3834
rect 8026 3782 8038 3834
rect 8090 3782 8102 3834
rect 8154 3782 12443 3834
rect 12495 3782 12507 3834
rect 12559 3782 12571 3834
rect 12623 3782 12635 3834
rect 12687 3782 12699 3834
rect 12751 3782 14812 3834
rect 1104 3760 14812 3782
rect 2774 3680 2780 3732
rect 2832 3720 2838 3732
rect 3053 3723 3111 3729
rect 2832 3692 2877 3720
rect 2832 3680 2838 3692
rect 3053 3689 3065 3723
rect 3099 3720 3111 3723
rect 3421 3723 3479 3729
rect 3421 3720 3433 3723
rect 3099 3692 3433 3720
rect 3099 3689 3111 3692
rect 3053 3683 3111 3689
rect 3421 3689 3433 3692
rect 3467 3720 3479 3723
rect 3602 3720 3608 3732
rect 3467 3692 3608 3720
rect 3467 3689 3479 3692
rect 3421 3683 3479 3689
rect 3602 3680 3608 3692
rect 3660 3680 3666 3732
rect 3878 3680 3884 3732
rect 3936 3720 3942 3732
rect 4525 3723 4583 3729
rect 4525 3720 4537 3723
rect 3936 3692 4537 3720
rect 3936 3680 3942 3692
rect 2869 3655 2927 3661
rect 2869 3621 2881 3655
rect 2915 3652 2927 3655
rect 3970 3652 3976 3664
rect 2915 3624 3976 3652
rect 2915 3621 2927 3624
rect 2869 3615 2927 3621
rect 3970 3612 3976 3624
rect 4028 3612 4034 3664
rect 2685 3587 2743 3593
rect 2685 3553 2697 3587
rect 2731 3584 2743 3587
rect 3053 3587 3111 3593
rect 3053 3584 3065 3587
rect 2731 3556 3065 3584
rect 2731 3553 2743 3556
rect 2685 3547 2743 3553
rect 3053 3553 3065 3556
rect 3099 3553 3111 3587
rect 3053 3547 3111 3553
rect 3145 3587 3203 3593
rect 3145 3553 3157 3587
rect 3191 3584 3203 3587
rect 4062 3584 4068 3596
rect 3191 3556 4068 3584
rect 3191 3553 3203 3556
rect 3145 3547 3203 3553
rect 4062 3544 4068 3556
rect 4120 3544 4126 3596
rect 2961 3519 3019 3525
rect 2961 3485 2973 3519
rect 3007 3485 3019 3519
rect 3418 3516 3424 3528
rect 3379 3488 3424 3516
rect 2961 3479 3019 3485
rect 2976 3448 3004 3479
rect 3418 3476 3424 3488
rect 3476 3476 3482 3528
rect 3605 3519 3663 3525
rect 3605 3485 3617 3519
rect 3651 3516 3663 3519
rect 3786 3516 3792 3528
rect 3651 3488 3792 3516
rect 3651 3485 3663 3488
rect 3605 3479 3663 3485
rect 3786 3476 3792 3488
rect 3844 3476 3850 3528
rect 3973 3519 4031 3525
rect 3973 3485 3985 3519
rect 4019 3485 4031 3519
rect 4172 3516 4200 3692
rect 4525 3689 4537 3692
rect 4571 3689 4583 3723
rect 5166 3720 5172 3732
rect 4525 3683 4583 3689
rect 4632 3692 5172 3720
rect 4433 3519 4491 3525
rect 4433 3516 4445 3519
rect 4172 3488 4445 3516
rect 3973 3479 4031 3485
rect 4433 3485 4445 3488
rect 4479 3485 4491 3519
rect 4632 3516 4660 3692
rect 5166 3680 5172 3692
rect 5224 3680 5230 3732
rect 8386 3720 8392 3732
rect 8347 3692 8392 3720
rect 8386 3680 8392 3692
rect 8444 3680 8450 3732
rect 10045 3723 10103 3729
rect 10045 3689 10057 3723
rect 10091 3720 10103 3723
rect 11974 3720 11980 3732
rect 10091 3692 11980 3720
rect 10091 3689 10103 3692
rect 10045 3683 10103 3689
rect 11974 3680 11980 3692
rect 12032 3680 12038 3732
rect 4908 3624 5396 3652
rect 4908 3528 4936 3624
rect 5258 3584 5264 3596
rect 5092 3556 5264 3584
rect 4697 3519 4755 3525
rect 4697 3516 4709 3519
rect 4632 3488 4709 3516
rect 4433 3479 4491 3485
rect 4697 3485 4709 3488
rect 4743 3485 4755 3519
rect 4697 3479 4755 3485
rect 4801 3497 4859 3503
rect 3142 3448 3148 3460
rect 2976 3420 3148 3448
rect 3142 3408 3148 3420
rect 3200 3408 3206 3460
rect 3988 3448 4016 3479
rect 4801 3463 4813 3497
rect 4847 3463 4859 3497
rect 4890 3476 4896 3528
rect 4948 3525 4954 3528
rect 5092 3525 5120 3556
rect 5258 3544 5264 3556
rect 5316 3544 5322 3596
rect 5368 3525 5396 3624
rect 5442 3612 5448 3664
rect 5500 3652 5506 3664
rect 8941 3655 8999 3661
rect 8941 3652 8953 3655
rect 5500 3624 5672 3652
rect 5500 3612 5506 3624
rect 5644 3593 5672 3624
rect 8036 3624 8953 3652
rect 5629 3587 5687 3593
rect 5629 3553 5641 3587
rect 5675 3553 5687 3587
rect 5629 3547 5687 3553
rect 5997 3587 6055 3593
rect 5997 3553 6009 3587
rect 6043 3584 6055 3587
rect 7006 3584 7012 3596
rect 6043 3556 7012 3584
rect 6043 3553 6055 3556
rect 5997 3547 6055 3553
rect 7006 3544 7012 3556
rect 7064 3544 7070 3596
rect 4948 3519 4969 3525
rect 4957 3485 4969 3519
rect 4948 3479 4969 3485
rect 5077 3519 5135 3525
rect 5077 3485 5089 3519
rect 5123 3485 5135 3519
rect 5077 3479 5135 3485
rect 5353 3519 5411 3525
rect 5353 3485 5365 3519
rect 5399 3485 5411 3519
rect 5534 3516 5540 3528
rect 5495 3488 5540 3516
rect 5353 3479 5411 3485
rect 4948 3476 4954 3479
rect 5534 3476 5540 3488
rect 5592 3476 5598 3528
rect 7423 3519 7481 3525
rect 7423 3485 7435 3519
rect 7469 3516 7481 3519
rect 7650 3516 7656 3528
rect 7469 3488 7656 3516
rect 7469 3485 7481 3488
rect 7423 3479 7481 3485
rect 7650 3476 7656 3488
rect 7708 3476 7714 3528
rect 7929 3519 7987 3525
rect 7929 3485 7941 3519
rect 7975 3516 7987 3519
rect 8036 3516 8064 3624
rect 8941 3621 8953 3624
rect 8987 3621 8999 3655
rect 8941 3615 8999 3621
rect 10686 3612 10692 3664
rect 10744 3652 10750 3664
rect 10781 3655 10839 3661
rect 10781 3652 10793 3655
rect 10744 3624 10793 3652
rect 10744 3612 10750 3624
rect 10781 3621 10793 3624
rect 10827 3621 10839 3655
rect 10781 3615 10839 3621
rect 10870 3612 10876 3664
rect 10928 3652 10934 3664
rect 10928 3624 10973 3652
rect 10928 3612 10934 3624
rect 8202 3584 8208 3596
rect 8163 3556 8208 3584
rect 8202 3544 8208 3556
rect 8260 3544 8266 3596
rect 9490 3584 9496 3596
rect 9451 3556 9496 3584
rect 9490 3544 9496 3556
rect 9548 3544 9554 3596
rect 9766 3544 9772 3596
rect 9824 3584 9830 3596
rect 10502 3584 10508 3596
rect 9824 3556 10508 3584
rect 9824 3544 9830 3556
rect 8386 3516 8392 3528
rect 7975 3488 8064 3516
rect 8347 3488 8392 3516
rect 7975 3485 7987 3488
rect 7929 3479 7987 3485
rect 8386 3476 8392 3488
rect 8444 3476 8450 3528
rect 10060 3525 10088 3556
rect 10502 3544 10508 3556
rect 10560 3544 10566 3596
rect 11330 3584 11336 3596
rect 11291 3556 11336 3584
rect 11330 3544 11336 3556
rect 11388 3544 11394 3596
rect 11517 3587 11575 3593
rect 11517 3553 11529 3587
rect 11563 3584 11575 3587
rect 12894 3584 12900 3596
rect 11563 3556 12900 3584
rect 11563 3553 11575 3556
rect 11517 3547 11575 3553
rect 12894 3544 12900 3556
rect 12952 3544 12958 3596
rect 13909 3587 13967 3593
rect 13909 3553 13921 3587
rect 13955 3584 13967 3587
rect 14366 3584 14372 3596
rect 13955 3556 14372 3584
rect 13955 3553 13967 3556
rect 13909 3547 13967 3553
rect 14366 3544 14372 3556
rect 14424 3544 14430 3596
rect 8481 3519 8539 3525
rect 8481 3485 8493 3519
rect 8527 3516 8539 3519
rect 10045 3519 10103 3525
rect 8527 3488 9996 3516
rect 8527 3485 8539 3488
rect 8481 3479 8539 3485
rect 4801 3460 4859 3463
rect 4338 3448 4344 3460
rect 3988 3420 4344 3448
rect 4338 3408 4344 3420
rect 4396 3408 4402 3460
rect 4798 3408 4804 3460
rect 4856 3408 4862 3460
rect 5166 3408 5172 3460
rect 5224 3448 5230 3460
rect 5445 3451 5503 3457
rect 5445 3448 5457 3451
rect 5224 3420 5457 3448
rect 5224 3408 5230 3420
rect 5445 3417 5457 3420
rect 5491 3417 5503 3451
rect 5445 3411 5503 3417
rect 6914 3408 6920 3460
rect 6972 3408 6978 3460
rect 7116 3420 7604 3448
rect 2593 3383 2651 3389
rect 2593 3349 2605 3383
rect 2639 3380 2651 3383
rect 2774 3380 2780 3392
rect 2639 3352 2780 3380
rect 2639 3349 2651 3352
rect 2593 3343 2651 3349
rect 2774 3340 2780 3352
rect 2832 3380 2838 3392
rect 3602 3380 3608 3392
rect 2832 3352 3608 3380
rect 2832 3340 2838 3352
rect 3602 3340 3608 3352
rect 3660 3340 3666 3392
rect 3786 3380 3792 3392
rect 3747 3352 3792 3380
rect 3786 3340 3792 3352
rect 3844 3340 3850 3392
rect 6638 3340 6644 3392
rect 6696 3380 6702 3392
rect 7116 3380 7144 3420
rect 7576 3389 7604 3420
rect 8294 3408 8300 3460
rect 8352 3448 8358 3460
rect 8662 3448 8668 3460
rect 8352 3420 8668 3448
rect 8352 3408 8358 3420
rect 8662 3408 8668 3420
rect 8720 3408 8726 3460
rect 8754 3408 8760 3460
rect 8812 3448 8818 3460
rect 9968 3448 9996 3488
rect 10045 3485 10057 3519
rect 10091 3485 10103 3519
rect 10045 3479 10103 3485
rect 10134 3476 10140 3528
rect 10192 3516 10198 3528
rect 10413 3519 10471 3525
rect 10413 3516 10425 3519
rect 10192 3488 10425 3516
rect 10192 3476 10198 3488
rect 10413 3485 10425 3488
rect 10459 3485 10471 3519
rect 10413 3479 10471 3485
rect 10686 3448 10692 3460
rect 8812 3420 9444 3448
rect 9968 3420 10692 3448
rect 8812 3408 8818 3420
rect 6696 3352 7144 3380
rect 7561 3383 7619 3389
rect 6696 3340 6702 3352
rect 7561 3349 7573 3383
rect 7607 3349 7619 3383
rect 7561 3343 7619 3349
rect 8021 3383 8079 3389
rect 8021 3349 8033 3383
rect 8067 3380 8079 3383
rect 8772 3380 8800 3408
rect 9306 3380 9312 3392
rect 8067 3352 8800 3380
rect 9267 3352 9312 3380
rect 8067 3349 8079 3352
rect 8021 3343 8079 3349
rect 9306 3340 9312 3352
rect 9364 3340 9370 3392
rect 9416 3389 9444 3420
rect 10686 3408 10692 3420
rect 10744 3408 10750 3460
rect 11054 3408 11060 3460
rect 11112 3448 11118 3460
rect 11885 3451 11943 3457
rect 11885 3448 11897 3451
rect 11112 3420 11897 3448
rect 11112 3408 11118 3420
rect 11885 3417 11897 3420
rect 11931 3417 11943 3451
rect 11885 3411 11943 3417
rect 12342 3408 12348 3460
rect 12400 3448 12406 3460
rect 12400 3420 12466 3448
rect 12400 3408 12406 3420
rect 13354 3408 13360 3460
rect 13412 3448 13418 3460
rect 13633 3451 13691 3457
rect 13633 3448 13645 3451
rect 13412 3420 13645 3448
rect 13412 3408 13418 3420
rect 13633 3417 13645 3420
rect 13679 3417 13691 3451
rect 14921 3451 14979 3457
rect 14921 3448 14933 3451
rect 13633 3411 13691 3417
rect 14108 3420 14933 3448
rect 9401 3383 9459 3389
rect 9401 3349 9413 3383
rect 9447 3380 9459 3383
rect 10594 3380 10600 3392
rect 9447 3352 10600 3380
rect 9447 3349 9459 3352
rect 9401 3343 9459 3349
rect 10594 3340 10600 3352
rect 10652 3340 10658 3392
rect 11238 3380 11244 3392
rect 11199 3352 11244 3380
rect 11238 3340 11244 3352
rect 11296 3340 11302 3392
rect 11330 3340 11336 3392
rect 11388 3380 11394 3392
rect 11701 3383 11759 3389
rect 11701 3380 11713 3383
rect 11388 3352 11713 3380
rect 11388 3340 11394 3352
rect 11701 3349 11713 3352
rect 11747 3349 11759 3383
rect 11701 3343 11759 3349
rect 11974 3340 11980 3392
rect 12032 3380 12038 3392
rect 12802 3380 12808 3392
rect 12032 3352 12808 3380
rect 12032 3340 12038 3352
rect 12802 3340 12808 3352
rect 12860 3340 12866 3392
rect 12894 3340 12900 3392
rect 12952 3380 12958 3392
rect 14108 3389 14136 3420
rect 14921 3417 14933 3420
rect 14967 3417 14979 3451
rect 14921 3411 14979 3417
rect 14093 3383 14151 3389
rect 14093 3380 14105 3383
rect 12952 3352 14105 3380
rect 12952 3340 12958 3352
rect 14093 3349 14105 3352
rect 14139 3349 14151 3383
rect 14458 3380 14464 3392
rect 14419 3352 14464 3380
rect 14093 3343 14151 3349
rect 14458 3340 14464 3352
rect 14516 3340 14522 3392
rect 1104 3290 14812 3312
rect 1104 3238 5547 3290
rect 5599 3238 5611 3290
rect 5663 3238 5675 3290
rect 5727 3238 5739 3290
rect 5791 3238 5803 3290
rect 5855 3238 10144 3290
rect 10196 3238 10208 3290
rect 10260 3238 10272 3290
rect 10324 3238 10336 3290
rect 10388 3238 10400 3290
rect 10452 3238 14812 3290
rect 1104 3216 14812 3238
rect 3786 3176 3792 3188
rect 2884 3148 3792 3176
rect 2884 3117 2912 3148
rect 3786 3136 3792 3148
rect 3844 3136 3850 3188
rect 4338 3176 4344 3188
rect 4299 3148 4344 3176
rect 4338 3136 4344 3148
rect 4396 3176 4402 3188
rect 4890 3176 4896 3188
rect 4396 3148 4896 3176
rect 4396 3136 4402 3148
rect 4890 3136 4896 3148
rect 4948 3136 4954 3188
rect 7009 3179 7067 3185
rect 7009 3145 7021 3179
rect 7055 3176 7067 3179
rect 7098 3176 7104 3188
rect 7055 3148 7104 3176
rect 7055 3145 7067 3148
rect 7009 3139 7067 3145
rect 7098 3136 7104 3148
rect 7156 3136 7162 3188
rect 9582 3176 9588 3188
rect 7484 3148 9588 3176
rect 2869 3111 2927 3117
rect 2869 3077 2881 3111
rect 2915 3077 2927 3111
rect 2869 3071 2927 3077
rect 3878 3068 3884 3120
rect 3936 3068 3942 3120
rect 6914 3108 6920 3120
rect 5934 3080 6920 3108
rect 6914 3068 6920 3080
rect 6972 3068 6978 3120
rect 6638 3040 6644 3052
rect 6599 3012 6644 3040
rect 6638 3000 6644 3012
rect 6696 3000 6702 3052
rect 7190 3040 7196 3052
rect 7151 3012 7196 3040
rect 7190 3000 7196 3012
rect 7248 3000 7254 3052
rect 7484 3049 7512 3148
rect 9582 3136 9588 3148
rect 9640 3136 9646 3188
rect 9674 3136 9680 3188
rect 9732 3136 9738 3188
rect 10505 3179 10563 3185
rect 10505 3145 10517 3179
rect 10551 3176 10563 3179
rect 10594 3176 10600 3188
rect 10551 3148 10600 3176
rect 10551 3145 10563 3148
rect 10505 3139 10563 3145
rect 10594 3136 10600 3148
rect 10652 3136 10658 3188
rect 10686 3136 10692 3188
rect 10744 3176 10750 3188
rect 11609 3179 11667 3185
rect 11609 3176 11621 3179
rect 10744 3148 11621 3176
rect 10744 3136 10750 3148
rect 11609 3145 11621 3148
rect 11655 3145 11667 3179
rect 11609 3139 11667 3145
rect 12621 3179 12679 3185
rect 12621 3145 12633 3179
rect 12667 3176 12679 3179
rect 13354 3176 13360 3188
rect 12667 3148 13360 3176
rect 12667 3145 12679 3148
rect 12621 3139 12679 3145
rect 13354 3136 13360 3148
rect 13412 3136 13418 3188
rect 7742 3108 7748 3120
rect 7703 3080 7748 3108
rect 7742 3068 7748 3080
rect 7800 3068 7806 3120
rect 8202 3068 8208 3120
rect 8260 3068 8266 3120
rect 7469 3043 7527 3049
rect 7469 3009 7481 3043
rect 7515 3009 7527 3043
rect 7469 3003 7527 3009
rect 9030 3000 9036 3052
rect 9088 3040 9094 3052
rect 9692 3049 9720 3136
rect 9766 3068 9772 3120
rect 9824 3068 9830 3120
rect 10045 3111 10103 3117
rect 10045 3077 10057 3111
rect 10091 3108 10103 3111
rect 10778 3108 10784 3120
rect 10091 3080 10784 3108
rect 10091 3077 10103 3080
rect 10045 3071 10103 3077
rect 10778 3068 10784 3080
rect 10836 3068 10842 3120
rect 11054 3108 11060 3120
rect 11015 3080 11060 3108
rect 11054 3068 11060 3080
rect 11112 3068 11118 3120
rect 12069 3111 12127 3117
rect 12069 3077 12081 3111
rect 12115 3108 12127 3111
rect 14093 3111 14151 3117
rect 12115 3080 12848 3108
rect 12115 3077 12127 3080
rect 12069 3071 12127 3077
rect 9769 3065 9827 3068
rect 9401 3043 9459 3049
rect 9401 3040 9413 3043
rect 9088 3012 9413 3040
rect 9088 3000 9094 3012
rect 9401 3009 9413 3012
rect 9447 3009 9459 3043
rect 9401 3003 9459 3009
rect 9677 3043 9735 3049
rect 9677 3009 9689 3043
rect 9723 3009 9735 3043
rect 9769 3031 9781 3065
rect 9815 3031 9827 3065
rect 9769 3025 9827 3031
rect 9857 3043 9915 3049
rect 9677 3003 9735 3009
rect 9857 3009 9869 3043
rect 9903 3040 9915 3043
rect 9950 3040 9956 3052
rect 9903 3012 9956 3040
rect 9903 3009 9915 3012
rect 9857 3003 9915 3009
rect 9950 3000 9956 3012
rect 10008 3000 10014 3052
rect 10502 3000 10508 3052
rect 10560 3040 10566 3052
rect 11333 3043 11391 3049
rect 11333 3040 11345 3043
rect 10560 3012 11345 3040
rect 10560 3000 10566 3012
rect 11333 3009 11345 3012
rect 11379 3009 11391 3043
rect 11333 3003 11391 3009
rect 11517 3043 11575 3049
rect 11517 3009 11529 3043
rect 11563 3009 11575 3043
rect 11517 3003 11575 3009
rect 12437 3043 12495 3049
rect 12437 3009 12449 3043
rect 12483 3040 12495 3043
rect 12710 3040 12716 3052
rect 12483 3012 12716 3040
rect 12483 3009 12495 3012
rect 12437 3003 12495 3009
rect 1670 2932 1676 2984
rect 1728 2972 1734 2984
rect 2593 2975 2651 2981
rect 2593 2972 2605 2975
rect 1728 2944 2605 2972
rect 1728 2932 1734 2944
rect 2593 2941 2605 2944
rect 2639 2972 2651 2975
rect 4246 2972 4252 2984
rect 2639 2944 4252 2972
rect 2639 2941 2651 2944
rect 2593 2935 2651 2941
rect 4246 2932 4252 2944
rect 4304 2972 4310 2984
rect 4433 2975 4491 2981
rect 4433 2972 4445 2975
rect 4304 2944 4445 2972
rect 4304 2932 4310 2944
rect 4433 2941 4445 2944
rect 4479 2941 4491 2975
rect 4433 2935 4491 2941
rect 4709 2975 4767 2981
rect 4709 2941 4721 2975
rect 4755 2972 4767 2975
rect 6365 2975 6423 2981
rect 6365 2972 6377 2975
rect 4755 2944 6377 2972
rect 4755 2941 4767 2944
rect 4709 2935 4767 2941
rect 6365 2941 6377 2944
rect 6411 2941 6423 2975
rect 6546 2972 6552 2984
rect 6507 2944 6552 2972
rect 6365 2935 6423 2941
rect 4448 2836 4476 2935
rect 6546 2932 6552 2944
rect 6604 2932 6610 2984
rect 7285 2975 7343 2981
rect 7285 2941 7297 2975
rect 7331 2972 7343 2975
rect 8386 2972 8392 2984
rect 7331 2944 8392 2972
rect 7331 2941 7343 2944
rect 7285 2935 7343 2941
rect 8386 2932 8392 2944
rect 8444 2932 8450 2984
rect 9214 2932 9220 2984
rect 9272 2972 9278 2984
rect 10042 2972 10048 2984
rect 9272 2944 10048 2972
rect 9272 2932 9278 2944
rect 10042 2932 10048 2944
rect 10100 2972 10106 2984
rect 10597 2975 10655 2981
rect 10597 2972 10609 2975
rect 10100 2944 10609 2972
rect 10100 2932 10106 2944
rect 10597 2941 10609 2944
rect 10643 2941 10655 2975
rect 10597 2935 10655 2941
rect 10689 2975 10747 2981
rect 10689 2941 10701 2975
rect 10735 2972 10747 2975
rect 11054 2972 11060 2984
rect 10735 2944 11060 2972
rect 10735 2941 10747 2944
rect 10689 2935 10747 2941
rect 6181 2907 6239 2913
rect 6181 2873 6193 2907
rect 6227 2904 6239 2907
rect 7190 2904 7196 2916
rect 6227 2876 7196 2904
rect 6227 2873 6239 2876
rect 6181 2867 6239 2873
rect 7190 2864 7196 2876
rect 7248 2864 7254 2916
rect 8772 2876 9352 2904
rect 5442 2836 5448 2848
rect 4448 2808 5448 2836
rect 5442 2796 5448 2808
rect 5500 2796 5506 2848
rect 7742 2796 7748 2848
rect 7800 2836 7806 2848
rect 8772 2836 8800 2876
rect 7800 2808 8800 2836
rect 7800 2796 7806 2808
rect 8846 2796 8852 2848
rect 8904 2836 8910 2848
rect 9217 2839 9275 2845
rect 9217 2836 9229 2839
rect 8904 2808 9229 2836
rect 8904 2796 8910 2808
rect 9217 2805 9229 2808
rect 9263 2805 9275 2839
rect 9324 2836 9352 2876
rect 9766 2864 9772 2916
rect 9824 2904 9830 2916
rect 10137 2907 10195 2913
rect 10137 2904 10149 2907
rect 9824 2876 10149 2904
rect 9824 2864 9830 2876
rect 10137 2873 10149 2876
rect 10183 2873 10195 2907
rect 10612 2904 10640 2935
rect 11054 2932 11060 2944
rect 11112 2932 11118 2984
rect 11238 2904 11244 2916
rect 10612 2876 11244 2904
rect 10137 2867 10195 2873
rect 11238 2864 11244 2876
rect 11296 2864 11302 2916
rect 11333 2907 11391 2913
rect 11333 2873 11345 2907
rect 11379 2904 11391 2907
rect 11422 2904 11428 2916
rect 11379 2876 11428 2904
rect 11379 2873 11391 2876
rect 11333 2867 11391 2873
rect 11422 2864 11428 2876
rect 11480 2864 11486 2916
rect 11532 2836 11560 3003
rect 12710 3000 12716 3012
rect 12768 3000 12774 3052
rect 12820 2972 12848 3080
rect 14093 3077 14105 3111
rect 14139 3108 14151 3111
rect 14182 3108 14188 3120
rect 14139 3080 14188 3108
rect 14139 3077 14151 3080
rect 14093 3071 14151 3077
rect 14182 3068 14188 3080
rect 14240 3068 14246 3120
rect 12986 3000 12992 3052
rect 13044 3000 13050 3052
rect 14366 3000 14372 3052
rect 14424 3040 14430 3052
rect 14424 3012 14469 3040
rect 14424 3000 14430 3012
rect 14090 2972 14096 2984
rect 12820 2944 14096 2972
rect 14090 2932 14096 2944
rect 14148 2932 14154 2984
rect 9324 2808 11560 2836
rect 9217 2799 9275 2805
rect 1104 2746 14812 2768
rect 1104 2694 3248 2746
rect 3300 2694 3312 2746
rect 3364 2694 3376 2746
rect 3428 2694 3440 2746
rect 3492 2694 3504 2746
rect 3556 2694 7846 2746
rect 7898 2694 7910 2746
rect 7962 2694 7974 2746
rect 8026 2694 8038 2746
rect 8090 2694 8102 2746
rect 8154 2694 12443 2746
rect 12495 2694 12507 2746
rect 12559 2694 12571 2746
rect 12623 2694 12635 2746
rect 12687 2694 12699 2746
rect 12751 2694 14812 2746
rect 1104 2672 14812 2694
rect 8573 2635 8631 2641
rect 8573 2601 8585 2635
rect 8619 2632 8631 2635
rect 9306 2632 9312 2644
rect 8619 2604 9312 2632
rect 8619 2601 8631 2604
rect 8573 2595 8631 2601
rect 9306 2592 9312 2604
rect 9364 2592 9370 2644
rect 11146 2632 11152 2644
rect 9416 2604 11152 2632
rect 7190 2524 7196 2576
rect 7248 2564 7254 2576
rect 9416 2564 9444 2604
rect 11146 2592 11152 2604
rect 11204 2592 11210 2644
rect 11238 2592 11244 2644
rect 11296 2632 11302 2644
rect 11333 2635 11391 2641
rect 11333 2632 11345 2635
rect 11296 2604 11345 2632
rect 11296 2592 11302 2604
rect 11333 2601 11345 2604
rect 11379 2601 11391 2635
rect 11333 2595 11391 2601
rect 14185 2635 14243 2641
rect 14185 2601 14197 2635
rect 14231 2632 14243 2635
rect 15013 2635 15071 2641
rect 15013 2632 15025 2635
rect 14231 2604 15025 2632
rect 14231 2601 14243 2604
rect 14185 2595 14243 2601
rect 15013 2601 15025 2604
rect 15059 2601 15071 2635
rect 15013 2595 15071 2601
rect 7248 2536 8248 2564
rect 7248 2524 7254 2536
rect 7837 2499 7895 2505
rect 7837 2465 7849 2499
rect 7883 2496 7895 2499
rect 8113 2499 8171 2505
rect 8113 2496 8125 2499
rect 7883 2468 8125 2496
rect 7883 2465 7895 2468
rect 7837 2459 7895 2465
rect 8113 2465 8125 2468
rect 8159 2465 8171 2499
rect 8113 2459 8171 2465
rect 3605 2431 3663 2437
rect 3605 2397 3617 2431
rect 3651 2428 3663 2431
rect 3970 2428 3976 2440
rect 3651 2400 3976 2428
rect 3651 2397 3663 2400
rect 3605 2391 3663 2397
rect 3970 2388 3976 2400
rect 4028 2428 4034 2440
rect 4065 2431 4123 2437
rect 4065 2428 4077 2431
rect 4028 2400 4077 2428
rect 4028 2388 4034 2400
rect 4065 2397 4077 2400
rect 4111 2397 4123 2431
rect 7742 2428 7748 2440
rect 7703 2400 7748 2428
rect 4065 2391 4123 2397
rect 7742 2388 7748 2400
rect 7800 2388 7806 2440
rect 8220 2437 8248 2536
rect 9048 2536 9444 2564
rect 10888 2536 12204 2564
rect 9048 2437 9076 2536
rect 9582 2496 9588 2508
rect 9543 2468 9588 2496
rect 9582 2456 9588 2468
rect 9640 2496 9646 2508
rect 10888 2496 10916 2536
rect 9640 2468 10916 2496
rect 9640 2456 9646 2468
rect 11790 2456 11796 2508
rect 11848 2496 11854 2508
rect 12176 2505 12204 2536
rect 12069 2499 12127 2505
rect 11848 2468 11893 2496
rect 11848 2456 11854 2468
rect 12069 2465 12081 2499
rect 12115 2465 12127 2499
rect 12069 2459 12127 2465
rect 12161 2499 12219 2505
rect 12161 2465 12173 2499
rect 12207 2465 12219 2499
rect 12161 2459 12219 2465
rect 7929 2431 7987 2437
rect 7929 2397 7941 2431
rect 7975 2397 7987 2431
rect 7929 2391 7987 2397
rect 8205 2431 8263 2437
rect 8205 2397 8217 2431
rect 8251 2397 8263 2431
rect 8205 2391 8263 2397
rect 9033 2431 9091 2437
rect 9033 2397 9045 2431
rect 9079 2397 9091 2431
rect 9214 2428 9220 2440
rect 9175 2400 9220 2428
rect 9033 2391 9091 2397
rect 5261 2363 5319 2369
rect 5261 2329 5273 2363
rect 5307 2329 5319 2363
rect 7944 2360 7972 2391
rect 9214 2388 9220 2400
rect 9272 2388 9278 2440
rect 9309 2431 9367 2437
rect 9309 2397 9321 2431
rect 9355 2397 9367 2431
rect 9309 2391 9367 2397
rect 8662 2360 8668 2372
rect 7944 2332 8668 2360
rect 5261 2323 5319 2329
rect 3878 2252 3884 2304
rect 3936 2292 3942 2304
rect 3973 2295 4031 2301
rect 3973 2292 3985 2295
rect 3936 2264 3985 2292
rect 3936 2252 3942 2264
rect 3973 2261 3985 2264
rect 4019 2292 4031 2295
rect 5276 2292 5304 2323
rect 8662 2320 8668 2332
rect 8720 2320 8726 2372
rect 9324 2360 9352 2391
rect 11146 2388 11152 2440
rect 11204 2428 11210 2440
rect 11701 2431 11759 2437
rect 11701 2428 11713 2431
rect 11204 2400 11713 2428
rect 11204 2388 11210 2400
rect 11701 2397 11713 2400
rect 11747 2397 11759 2431
rect 11701 2391 11759 2397
rect 9766 2360 9772 2372
rect 9324 2332 9772 2360
rect 9766 2320 9772 2332
rect 9824 2320 9830 2372
rect 9861 2363 9919 2369
rect 9861 2329 9873 2363
rect 9907 2329 9919 2363
rect 9861 2323 9919 2329
rect 6457 2295 6515 2301
rect 6457 2292 6469 2295
rect 4019 2264 6469 2292
rect 4019 2261 4031 2264
rect 3973 2255 4031 2261
rect 6457 2261 6469 2264
rect 6503 2292 6515 2295
rect 6914 2292 6920 2304
rect 6503 2264 6920 2292
rect 6503 2261 6515 2264
rect 6457 2255 6515 2261
rect 6914 2252 6920 2264
rect 6972 2292 6978 2304
rect 7285 2295 7343 2301
rect 7285 2292 7297 2295
rect 6972 2264 7297 2292
rect 6972 2252 6978 2264
rect 7285 2261 7297 2264
rect 7331 2292 7343 2295
rect 8202 2292 8208 2304
rect 7331 2264 8208 2292
rect 7331 2261 7343 2264
rect 7285 2255 7343 2261
rect 8202 2252 8208 2264
rect 8260 2292 8266 2304
rect 9030 2292 9036 2304
rect 8260 2264 9036 2292
rect 8260 2252 8266 2264
rect 9030 2252 9036 2264
rect 9088 2252 9094 2304
rect 9125 2295 9183 2301
rect 9125 2261 9137 2295
rect 9171 2292 9183 2295
rect 9398 2292 9404 2304
rect 9171 2264 9404 2292
rect 9171 2261 9183 2264
rect 9125 2255 9183 2261
rect 9398 2252 9404 2264
rect 9456 2252 9462 2304
rect 9493 2295 9551 2301
rect 9493 2261 9505 2295
rect 9539 2292 9551 2295
rect 9876 2292 9904 2323
rect 10318 2320 10324 2372
rect 10376 2320 10382 2372
rect 9539 2264 9904 2292
rect 11716 2292 11744 2391
rect 12084 2360 12112 2459
rect 12894 2456 12900 2508
rect 12952 2496 12958 2508
rect 14369 2499 14427 2505
rect 14369 2496 14381 2499
rect 12952 2468 14381 2496
rect 12952 2456 12958 2468
rect 14369 2465 14381 2468
rect 14415 2465 14427 2499
rect 14369 2459 14427 2465
rect 14090 2428 14096 2440
rect 14051 2400 14096 2428
rect 14090 2388 14096 2400
rect 14148 2388 14154 2440
rect 12437 2363 12495 2369
rect 12437 2360 12449 2363
rect 12084 2332 12449 2360
rect 12437 2329 12449 2332
rect 12483 2329 12495 2363
rect 12437 2323 12495 2329
rect 12526 2320 12532 2372
rect 12584 2360 12590 2372
rect 12894 2360 12900 2372
rect 12584 2332 12900 2360
rect 12584 2320 12590 2332
rect 12894 2320 12900 2332
rect 12952 2320 12958 2372
rect 13909 2295 13967 2301
rect 13909 2292 13921 2295
rect 11716 2264 13921 2292
rect 9539 2261 9551 2264
rect 9493 2255 9551 2261
rect 13909 2261 13921 2264
rect 13955 2261 13967 2295
rect 13909 2255 13967 2261
rect 1104 2202 14812 2224
rect 1104 2150 5547 2202
rect 5599 2150 5611 2202
rect 5663 2150 5675 2202
rect 5727 2150 5739 2202
rect 5791 2150 5803 2202
rect 5855 2150 10144 2202
rect 10196 2150 10208 2202
rect 10260 2150 10272 2202
rect 10324 2150 10336 2202
rect 10388 2150 10400 2202
rect 10452 2150 14812 2202
rect 1104 2128 14812 2150
rect 14918 1068 14924 1080
rect 14879 1040 14924 1068
rect 14918 1028 14924 1040
rect 14976 1028 14982 1080
<< via1 >>
rect 14924 15011 14976 15020
rect 14924 14977 14933 15011
rect 14933 14977 14967 15011
rect 14967 14977 14976 15011
rect 14924 14968 14976 14977
rect 3248 13574 3300 13626
rect 3312 13574 3364 13626
rect 3376 13574 3428 13626
rect 3440 13574 3492 13626
rect 3504 13574 3556 13626
rect 7846 13574 7898 13626
rect 7910 13574 7962 13626
rect 7974 13574 8026 13626
rect 8038 13574 8090 13626
rect 8102 13574 8154 13626
rect 12443 13574 12495 13626
rect 12507 13574 12559 13626
rect 12571 13574 12623 13626
rect 12635 13574 12687 13626
rect 12699 13574 12751 13626
rect 2780 13472 2832 13524
rect 7564 13515 7616 13524
rect 7564 13481 7573 13515
rect 7573 13481 7607 13515
rect 7607 13481 7616 13515
rect 7564 13472 7616 13481
rect 8208 13472 8260 13524
rect 2780 13311 2832 13320
rect 2780 13277 2789 13311
rect 2789 13277 2823 13311
rect 2823 13277 2832 13311
rect 2780 13268 2832 13277
rect 3976 13268 4028 13320
rect 4160 13268 4212 13320
rect 4344 13321 4396 13330
rect 4344 13287 4353 13321
rect 4353 13287 4387 13321
rect 4387 13287 4396 13321
rect 4344 13278 4396 13287
rect 4528 13268 4580 13320
rect 8484 13404 8536 13456
rect 5264 13336 5316 13388
rect 8852 13336 8904 13388
rect 7656 13268 7708 13320
rect 8208 13311 8260 13320
rect 8208 13277 8217 13311
rect 8217 13277 8251 13311
rect 8251 13277 8260 13311
rect 8208 13268 8260 13277
rect 13268 13472 13320 13524
rect 13360 13472 13412 13524
rect 12992 13336 13044 13388
rect 11336 13268 11388 13320
rect 12440 13311 12492 13320
rect 12440 13277 12449 13311
rect 12449 13277 12483 13311
rect 12483 13277 12492 13311
rect 12440 13268 12492 13277
rect 14188 13268 14240 13320
rect 10876 13200 10928 13252
rect 2504 13132 2556 13184
rect 2872 13132 2924 13184
rect 4160 13132 4212 13184
rect 4712 13175 4764 13184
rect 4712 13141 4721 13175
rect 4721 13141 4755 13175
rect 4755 13141 4764 13175
rect 4712 13132 4764 13141
rect 5448 13132 5500 13184
rect 5908 13132 5960 13184
rect 8300 13132 8352 13184
rect 8668 13175 8720 13184
rect 8668 13141 8677 13175
rect 8677 13141 8711 13175
rect 8711 13141 8720 13175
rect 8668 13132 8720 13141
rect 10784 13132 10836 13184
rect 11428 13132 11480 13184
rect 12716 13132 12768 13184
rect 12900 13132 12952 13184
rect 14096 13132 14148 13184
rect 5547 13030 5599 13082
rect 5611 13030 5663 13082
rect 5675 13030 5727 13082
rect 5739 13030 5791 13082
rect 5803 13030 5855 13082
rect 10144 13030 10196 13082
rect 10208 13030 10260 13082
rect 10272 13030 10324 13082
rect 10336 13030 10388 13082
rect 10400 13030 10452 13082
rect 2964 12928 3016 12980
rect 4712 12928 4764 12980
rect 5448 12971 5500 12980
rect 5448 12937 5457 12971
rect 5457 12937 5491 12971
rect 5491 12937 5500 12971
rect 5448 12928 5500 12937
rect 12440 12928 12492 12980
rect 14188 12971 14240 12980
rect 14188 12937 14197 12971
rect 14197 12937 14231 12971
rect 14231 12937 14240 12971
rect 14188 12928 14240 12937
rect 2504 12835 2556 12844
rect 2504 12801 2513 12835
rect 2513 12801 2547 12835
rect 2547 12801 2556 12835
rect 2504 12792 2556 12801
rect 2872 12835 2924 12844
rect 2872 12801 2881 12835
rect 2881 12801 2915 12835
rect 2915 12801 2924 12835
rect 2872 12792 2924 12801
rect 4620 12835 4672 12844
rect 4620 12801 4629 12835
rect 4629 12801 4663 12835
rect 4663 12801 4672 12835
rect 4620 12792 4672 12801
rect 4344 12656 4396 12708
rect 4896 12656 4948 12708
rect 5908 12767 5960 12776
rect 5908 12733 5917 12767
rect 5917 12733 5951 12767
rect 5951 12733 5960 12767
rect 5908 12724 5960 12733
rect 6000 12767 6052 12776
rect 6000 12733 6009 12767
rect 6009 12733 6043 12767
rect 6043 12733 6052 12767
rect 6000 12724 6052 12733
rect 5080 12588 5132 12640
rect 6920 12792 6972 12844
rect 7288 12835 7340 12844
rect 7288 12801 7322 12835
rect 7322 12801 7340 12835
rect 7288 12792 7340 12801
rect 8668 12860 8720 12912
rect 9312 12860 9364 12912
rect 11336 12860 11388 12912
rect 12900 12860 12952 12912
rect 11152 12835 11204 12844
rect 11152 12801 11161 12835
rect 11161 12801 11195 12835
rect 11195 12801 11204 12835
rect 11152 12792 11204 12801
rect 13820 12835 13872 12844
rect 8392 12631 8444 12640
rect 8392 12597 8401 12631
rect 8401 12597 8435 12631
rect 8435 12597 8444 12631
rect 8392 12588 8444 12597
rect 8852 12724 8904 12776
rect 11428 12724 11480 12776
rect 13820 12801 13829 12835
rect 13829 12801 13863 12835
rect 13863 12801 13872 12835
rect 13820 12792 13872 12801
rect 14096 12835 14148 12844
rect 14096 12801 14105 12835
rect 14105 12801 14139 12835
rect 14139 12801 14148 12835
rect 14096 12792 14148 12801
rect 14280 12835 14332 12844
rect 14280 12801 14289 12835
rect 14289 12801 14323 12835
rect 14323 12801 14332 12835
rect 14280 12792 14332 12801
rect 12992 12724 13044 12776
rect 13636 12724 13688 12776
rect 11520 12656 11572 12708
rect 13452 12699 13504 12708
rect 13452 12665 13461 12699
rect 13461 12665 13495 12699
rect 13495 12665 13504 12699
rect 13452 12656 13504 12665
rect 9496 12588 9548 12640
rect 10968 12631 11020 12640
rect 10968 12597 10977 12631
rect 10977 12597 11011 12631
rect 11011 12597 11020 12631
rect 10968 12588 11020 12597
rect 11336 12588 11388 12640
rect 3248 12486 3300 12538
rect 3312 12486 3364 12538
rect 3376 12486 3428 12538
rect 3440 12486 3492 12538
rect 3504 12486 3556 12538
rect 7846 12486 7898 12538
rect 7910 12486 7962 12538
rect 7974 12486 8026 12538
rect 8038 12486 8090 12538
rect 8102 12486 8154 12538
rect 12443 12486 12495 12538
rect 12507 12486 12559 12538
rect 12571 12486 12623 12538
rect 12635 12486 12687 12538
rect 12699 12486 12751 12538
rect 7564 12427 7616 12436
rect 7564 12393 7573 12427
rect 7573 12393 7607 12427
rect 7607 12393 7616 12427
rect 7564 12384 7616 12393
rect 7656 12384 7708 12436
rect 6092 12316 6144 12368
rect 8208 12384 8260 12436
rect 11152 12384 11204 12436
rect 11796 12384 11848 12436
rect 13636 12384 13688 12436
rect 14280 12427 14332 12436
rect 14280 12393 14289 12427
rect 14289 12393 14323 12427
rect 14323 12393 14332 12427
rect 14280 12384 14332 12393
rect 8944 12316 8996 12368
rect 2780 12248 2832 12300
rect 4804 12291 4856 12300
rect 3976 12223 4028 12232
rect 3976 12189 3985 12223
rect 3985 12189 4019 12223
rect 4019 12189 4028 12223
rect 3976 12180 4028 12189
rect 4068 12223 4120 12232
rect 4068 12189 4077 12223
rect 4077 12189 4111 12223
rect 4111 12189 4120 12223
rect 4804 12257 4813 12291
rect 4813 12257 4847 12291
rect 4847 12257 4856 12291
rect 4804 12248 4856 12257
rect 5356 12248 5408 12300
rect 4068 12180 4120 12189
rect 4620 12180 4672 12232
rect 4988 12180 5040 12232
rect 5264 12180 5316 12232
rect 8392 12248 8444 12300
rect 5908 12180 5960 12232
rect 6920 12180 6972 12232
rect 7564 12180 7616 12232
rect 8300 12223 8352 12232
rect 8300 12189 8309 12223
rect 8309 12189 8343 12223
rect 8343 12189 8352 12223
rect 8300 12180 8352 12189
rect 10876 12248 10928 12300
rect 12348 12248 12400 12300
rect 9496 12180 9548 12232
rect 1860 12112 1912 12164
rect 2044 12155 2096 12164
rect 2044 12121 2053 12155
rect 2053 12121 2087 12155
rect 2087 12121 2096 12155
rect 2044 12112 2096 12121
rect 2964 12044 3016 12096
rect 3608 12044 3660 12096
rect 4896 12112 4948 12164
rect 6460 12155 6512 12164
rect 6460 12121 6494 12155
rect 6494 12121 6512 12155
rect 6460 12112 6512 12121
rect 4436 12044 4488 12096
rect 5448 12044 5500 12096
rect 5908 12044 5960 12096
rect 9312 12087 9364 12096
rect 9312 12053 9321 12087
rect 9321 12053 9355 12087
rect 9355 12053 9364 12087
rect 9312 12044 9364 12053
rect 12164 12112 12216 12164
rect 10968 12044 11020 12096
rect 11612 12044 11664 12096
rect 12256 12044 12308 12096
rect 14280 12112 14332 12164
rect 12900 12044 12952 12096
rect 5547 11942 5599 11994
rect 5611 11942 5663 11994
rect 5675 11942 5727 11994
rect 5739 11942 5791 11994
rect 5803 11942 5855 11994
rect 10144 11942 10196 11994
rect 10208 11942 10260 11994
rect 10272 11942 10324 11994
rect 10336 11942 10388 11994
rect 10400 11942 10452 11994
rect 2044 11840 2096 11892
rect 4804 11840 4856 11892
rect 5448 11883 5500 11892
rect 5448 11849 5457 11883
rect 5457 11849 5491 11883
rect 5491 11849 5500 11883
rect 5448 11840 5500 11849
rect 8484 11840 8536 11892
rect 8760 11840 8812 11892
rect 4068 11772 4120 11824
rect 4436 11704 4488 11756
rect 5356 11772 5408 11824
rect 4252 11636 4304 11688
rect 4712 11704 4764 11756
rect 4896 11747 4948 11756
rect 4896 11713 4905 11747
rect 4905 11713 4939 11747
rect 4939 11713 4948 11747
rect 4896 11704 4948 11713
rect 5080 11747 5132 11756
rect 5080 11713 5089 11747
rect 5089 11713 5123 11747
rect 5123 11713 5132 11747
rect 6920 11772 6972 11824
rect 5080 11704 5132 11713
rect 5356 11636 5408 11688
rect 5908 11679 5960 11688
rect 5908 11645 5917 11679
rect 5917 11645 5951 11679
rect 5951 11645 5960 11679
rect 5908 11636 5960 11645
rect 6000 11679 6052 11688
rect 6000 11645 6009 11679
rect 6009 11645 6043 11679
rect 6043 11645 6052 11679
rect 8484 11704 8536 11756
rect 8944 11704 8996 11756
rect 9036 11747 9088 11756
rect 9036 11713 9045 11747
rect 9045 11713 9079 11747
rect 9079 11713 9088 11747
rect 9036 11704 9088 11713
rect 9220 11704 9272 11756
rect 10876 11840 10928 11892
rect 11060 11840 11112 11892
rect 14280 11883 14332 11892
rect 11152 11772 11204 11824
rect 11612 11815 11664 11824
rect 11612 11781 11621 11815
rect 11621 11781 11655 11815
rect 11655 11781 11664 11815
rect 11612 11772 11664 11781
rect 12808 11815 12860 11824
rect 12808 11781 12817 11815
rect 12817 11781 12851 11815
rect 12851 11781 12860 11815
rect 12808 11772 12860 11781
rect 13360 11772 13412 11824
rect 14280 11849 14289 11883
rect 14289 11849 14323 11883
rect 14323 11849 14332 11883
rect 14280 11840 14332 11849
rect 9956 11747 10008 11756
rect 7840 11679 7892 11688
rect 6000 11636 6052 11645
rect 4620 11568 4672 11620
rect 7840 11645 7849 11679
rect 7849 11645 7883 11679
rect 7883 11645 7892 11679
rect 7840 11636 7892 11645
rect 9404 11636 9456 11688
rect 9956 11713 9965 11747
rect 9965 11713 9999 11747
rect 9999 11713 10008 11747
rect 9956 11704 10008 11713
rect 10048 11747 10100 11756
rect 10048 11713 10057 11747
rect 10057 11713 10091 11747
rect 10091 11713 10100 11747
rect 10048 11704 10100 11713
rect 10876 11704 10928 11756
rect 11244 11747 11296 11756
rect 10692 11679 10744 11688
rect 10692 11645 10701 11679
rect 10701 11645 10735 11679
rect 10735 11645 10744 11679
rect 10692 11636 10744 11645
rect 10784 11679 10836 11688
rect 10784 11645 10793 11679
rect 10793 11645 10827 11679
rect 10827 11645 10836 11679
rect 11244 11713 11253 11747
rect 11253 11713 11287 11747
rect 11287 11713 11296 11747
rect 11244 11704 11296 11713
rect 11336 11747 11388 11756
rect 11336 11713 11345 11747
rect 11345 11713 11379 11747
rect 11379 11713 11388 11747
rect 11336 11704 11388 11713
rect 11520 11704 11572 11756
rect 10784 11636 10836 11645
rect 11796 11636 11848 11688
rect 12164 11679 12216 11688
rect 12164 11645 12173 11679
rect 12173 11645 12207 11679
rect 12207 11645 12216 11679
rect 12164 11636 12216 11645
rect 9220 11611 9272 11620
rect 9220 11577 9229 11611
rect 9229 11577 9263 11611
rect 9263 11577 9272 11611
rect 9220 11568 9272 11577
rect 2964 11500 3016 11552
rect 4068 11543 4120 11552
rect 4068 11509 4077 11543
rect 4077 11509 4111 11543
rect 4111 11509 4120 11543
rect 4068 11500 4120 11509
rect 4344 11500 4396 11552
rect 4528 11500 4580 11552
rect 8760 11500 8812 11552
rect 9680 11543 9732 11552
rect 9680 11509 9689 11543
rect 9689 11509 9723 11543
rect 9723 11509 9732 11543
rect 9680 11500 9732 11509
rect 11612 11500 11664 11552
rect 12348 11636 12400 11688
rect 12900 11500 12952 11552
rect 3248 11398 3300 11450
rect 3312 11398 3364 11450
rect 3376 11398 3428 11450
rect 3440 11398 3492 11450
rect 3504 11398 3556 11450
rect 7846 11398 7898 11450
rect 7910 11398 7962 11450
rect 7974 11398 8026 11450
rect 8038 11398 8090 11450
rect 8102 11398 8154 11450
rect 12443 11398 12495 11450
rect 12507 11398 12559 11450
rect 12571 11398 12623 11450
rect 12635 11398 12687 11450
rect 12699 11398 12751 11450
rect 3608 11339 3660 11348
rect 3608 11305 3617 11339
rect 3617 11305 3651 11339
rect 3651 11305 3660 11339
rect 3608 11296 3660 11305
rect 4620 11296 4672 11348
rect 6460 11296 6512 11348
rect 4068 11228 4120 11280
rect 6184 11228 6236 11280
rect 6828 11228 6880 11280
rect 4528 11160 4580 11212
rect 5264 11160 5316 11212
rect 5816 11160 5868 11212
rect 6920 11203 6972 11212
rect 6920 11169 6929 11203
rect 6929 11169 6963 11203
rect 6963 11169 6972 11203
rect 6920 11160 6972 11169
rect 8300 11160 8352 11212
rect 8852 11296 8904 11348
rect 9404 11296 9456 11348
rect 8576 11228 8628 11280
rect 9312 11228 9364 11280
rect 8668 11160 8720 11212
rect 8944 11160 8996 11212
rect 9680 11296 9732 11348
rect 10692 11296 10744 11348
rect 11244 11296 11296 11348
rect 1860 11135 1912 11144
rect 1860 11101 1869 11135
rect 1869 11101 1903 11135
rect 1903 11101 1912 11135
rect 1860 11092 1912 11101
rect 4252 11092 4304 11144
rect 5908 11092 5960 11144
rect 10968 11228 11020 11280
rect 11520 11228 11572 11280
rect 9864 11160 9916 11212
rect 11704 11203 11756 11212
rect 11704 11169 11713 11203
rect 11713 11169 11747 11203
rect 11747 11169 11756 11203
rect 11704 11160 11756 11169
rect 9956 11135 10008 11144
rect 9956 11101 9965 11135
rect 9965 11101 9999 11135
rect 9999 11101 10008 11135
rect 9956 11092 10008 11101
rect 11152 11092 11204 11144
rect 11612 11092 11664 11144
rect 12072 11135 12124 11144
rect 12072 11101 12081 11135
rect 12081 11101 12115 11135
rect 12115 11101 12124 11135
rect 12072 11092 12124 11101
rect 12348 11092 12400 11144
rect 13820 11092 13872 11144
rect 4344 11024 4396 11076
rect 5540 11067 5592 11076
rect 5540 11033 5549 11067
rect 5549 11033 5583 11067
rect 5583 11033 5592 11067
rect 6276 11067 6328 11076
rect 5540 11024 5592 11033
rect 6276 11033 6285 11067
rect 6285 11033 6319 11067
rect 6319 11033 6328 11067
rect 6276 11024 6328 11033
rect 6644 11024 6696 11076
rect 7656 11024 7708 11076
rect 9220 11024 9272 11076
rect 10140 11067 10192 11076
rect 10140 11033 10149 11067
rect 10149 11033 10183 11067
rect 10183 11033 10192 11067
rect 10140 11024 10192 11033
rect 10232 11024 10284 11076
rect 10600 11024 10652 11076
rect 13360 11024 13412 11076
rect 2964 10956 3016 11008
rect 5080 10999 5132 11008
rect 5080 10965 5089 10999
rect 5089 10965 5123 10999
rect 5123 10965 5132 10999
rect 5080 10956 5132 10965
rect 6552 10956 6604 11008
rect 8576 10956 8628 11008
rect 8944 10999 8996 11008
rect 8944 10965 8953 10999
rect 8953 10965 8987 10999
rect 8987 10965 8996 10999
rect 8944 10956 8996 10965
rect 9772 10956 9824 11008
rect 10508 10956 10560 11008
rect 11060 10956 11112 11008
rect 12164 10956 12216 11008
rect 14096 10956 14148 11008
rect 5547 10854 5599 10906
rect 5611 10854 5663 10906
rect 5675 10854 5727 10906
rect 5739 10854 5791 10906
rect 5803 10854 5855 10906
rect 10144 10854 10196 10906
rect 10208 10854 10260 10906
rect 10272 10854 10324 10906
rect 10336 10854 10388 10906
rect 10400 10854 10452 10906
rect 15016 10820 15068 10872
rect 4252 10795 4304 10804
rect 4252 10761 4261 10795
rect 4261 10761 4295 10795
rect 4295 10761 4304 10795
rect 4252 10752 4304 10761
rect 4620 10752 4672 10804
rect 5080 10752 5132 10804
rect 3884 10684 3936 10736
rect 1860 10616 1912 10668
rect 3516 10659 3568 10668
rect 3516 10625 3525 10659
rect 3525 10625 3559 10659
rect 3559 10625 3568 10659
rect 3516 10616 3568 10625
rect 3700 10659 3752 10668
rect 3700 10625 3709 10659
rect 3709 10625 3743 10659
rect 3743 10625 3752 10659
rect 3700 10616 3752 10625
rect 3792 10659 3844 10668
rect 3792 10625 3801 10659
rect 3801 10625 3835 10659
rect 3835 10625 3844 10659
rect 4528 10684 4580 10736
rect 4988 10684 5040 10736
rect 5448 10752 5500 10804
rect 5908 10752 5960 10804
rect 6276 10752 6328 10804
rect 5264 10684 5316 10736
rect 3792 10616 3844 10625
rect 5172 10616 5224 10668
rect 3148 10523 3200 10532
rect 3148 10489 3157 10523
rect 3157 10489 3191 10523
rect 3191 10489 3200 10523
rect 3148 10480 3200 10489
rect 4896 10591 4948 10600
rect 4896 10557 4905 10591
rect 4905 10557 4939 10591
rect 4939 10557 4948 10591
rect 4896 10548 4948 10557
rect 1400 10412 1452 10464
rect 3056 10412 3108 10464
rect 4988 10480 5040 10532
rect 3884 10412 3936 10464
rect 4436 10412 4488 10464
rect 5632 10659 5684 10668
rect 5632 10625 5641 10659
rect 5641 10625 5675 10659
rect 5675 10625 5684 10659
rect 5632 10616 5684 10625
rect 5816 10616 5868 10668
rect 6184 10684 6236 10736
rect 7656 10752 7708 10804
rect 8300 10752 8352 10804
rect 8392 10684 8444 10736
rect 9772 10752 9824 10804
rect 10692 10752 10744 10804
rect 13820 10752 13872 10804
rect 6552 10659 6604 10668
rect 6552 10625 6561 10659
rect 6561 10625 6595 10659
rect 6595 10625 6604 10659
rect 6552 10616 6604 10625
rect 6920 10659 6972 10668
rect 6920 10625 6929 10659
rect 6929 10625 6963 10659
rect 6963 10625 6972 10659
rect 6920 10616 6972 10625
rect 8576 10659 8628 10668
rect 8576 10625 8585 10659
rect 8585 10625 8619 10659
rect 8619 10625 8628 10659
rect 8576 10616 8628 10625
rect 8944 10659 8996 10668
rect 8944 10625 8953 10659
rect 8953 10625 8987 10659
rect 8987 10625 8996 10659
rect 8944 10616 8996 10625
rect 9496 10659 9548 10668
rect 9496 10625 9505 10659
rect 9505 10625 9539 10659
rect 9539 10625 9548 10659
rect 9496 10616 9548 10625
rect 10232 10684 10284 10736
rect 9956 10616 10008 10668
rect 8668 10548 8720 10600
rect 10968 10548 11020 10600
rect 13360 10684 13412 10736
rect 12164 10616 12216 10668
rect 12256 10616 12308 10668
rect 14096 10659 14148 10668
rect 14096 10625 14105 10659
rect 14105 10625 14139 10659
rect 14139 10625 14148 10659
rect 14096 10616 14148 10625
rect 5448 10412 5500 10464
rect 6184 10455 6236 10464
rect 6184 10421 6193 10455
rect 6193 10421 6227 10455
rect 6227 10421 6236 10455
rect 6184 10412 6236 10421
rect 8668 10412 8720 10464
rect 9312 10455 9364 10464
rect 9312 10421 9321 10455
rect 9321 10421 9355 10455
rect 9355 10421 9364 10455
rect 9312 10412 9364 10421
rect 11704 10480 11756 10532
rect 11244 10412 11296 10464
rect 11520 10455 11572 10464
rect 11520 10421 11529 10455
rect 11529 10421 11563 10455
rect 11563 10421 11572 10455
rect 11520 10412 11572 10421
rect 3248 10310 3300 10362
rect 3312 10310 3364 10362
rect 3376 10310 3428 10362
rect 3440 10310 3492 10362
rect 3504 10310 3556 10362
rect 7846 10310 7898 10362
rect 7910 10310 7962 10362
rect 7974 10310 8026 10362
rect 8038 10310 8090 10362
rect 8102 10310 8154 10362
rect 12443 10310 12495 10362
rect 12507 10310 12559 10362
rect 12571 10310 12623 10362
rect 12635 10310 12687 10362
rect 12699 10310 12751 10362
rect 3700 10208 3752 10260
rect 3976 10208 4028 10260
rect 8576 10208 8628 10260
rect 9312 10208 9364 10260
rect 10232 10208 10284 10260
rect 10968 10251 11020 10260
rect 10968 10217 10977 10251
rect 10977 10217 11011 10251
rect 11011 10217 11020 10251
rect 10968 10208 11020 10217
rect 12164 10251 12216 10260
rect 12164 10217 12173 10251
rect 12173 10217 12207 10251
rect 12207 10217 12216 10251
rect 12164 10208 12216 10217
rect 12992 10251 13044 10260
rect 12992 10217 13001 10251
rect 13001 10217 13035 10251
rect 13035 10217 13044 10251
rect 12992 10208 13044 10217
rect 13360 10208 13412 10260
rect 3148 10072 3200 10124
rect 4160 10140 4212 10192
rect 5172 10183 5224 10192
rect 5172 10149 5181 10183
rect 5181 10149 5215 10183
rect 5215 10149 5224 10183
rect 5172 10140 5224 10149
rect 5356 10140 5408 10192
rect 5632 10140 5684 10192
rect 5908 10140 5960 10192
rect 9956 10140 10008 10192
rect 3792 10047 3844 10056
rect 3792 10013 3801 10047
rect 3801 10013 3835 10047
rect 3835 10013 3844 10047
rect 3792 10004 3844 10013
rect 3884 10004 3936 10056
rect 4344 10047 4396 10056
rect 2964 9936 3016 9988
rect 4344 10013 4353 10047
rect 4353 10013 4387 10047
rect 4387 10013 4396 10047
rect 4344 10004 4396 10013
rect 4528 10004 4580 10056
rect 4620 10047 4672 10056
rect 4620 10013 4629 10047
rect 4629 10013 4663 10047
rect 4663 10013 4672 10047
rect 4988 10047 5040 10056
rect 4620 10004 4672 10013
rect 4988 10013 4997 10047
rect 4997 10013 5031 10047
rect 5031 10013 5040 10047
rect 4988 10004 5040 10013
rect 5080 10047 5132 10056
rect 5080 10013 5089 10047
rect 5089 10013 5123 10047
rect 5123 10013 5132 10047
rect 5356 10047 5408 10056
rect 5080 10004 5132 10013
rect 5356 10013 5365 10047
rect 5365 10013 5399 10047
rect 5399 10013 5408 10047
rect 5356 10004 5408 10013
rect 5448 10047 5500 10056
rect 5448 10013 5457 10047
rect 5457 10013 5491 10047
rect 5491 10013 5500 10047
rect 6184 10072 6236 10124
rect 5448 10004 5500 10013
rect 7748 10047 7800 10056
rect 7748 10013 7757 10047
rect 7757 10013 7791 10047
rect 7791 10013 7800 10047
rect 7748 10004 7800 10013
rect 8484 10004 8536 10056
rect 8668 10047 8720 10056
rect 8668 10013 8677 10047
rect 8677 10013 8711 10047
rect 8711 10013 8720 10047
rect 9772 10072 9824 10124
rect 10508 10072 10560 10124
rect 11520 10072 11572 10124
rect 11704 10072 11756 10124
rect 8668 10004 8720 10013
rect 3516 9911 3568 9920
rect 3516 9877 3525 9911
rect 3525 9877 3559 9911
rect 3559 9877 3568 9911
rect 3516 9868 3568 9877
rect 3700 9868 3752 9920
rect 8852 9936 8904 9988
rect 10416 10004 10468 10056
rect 10784 10047 10836 10056
rect 10784 10013 10793 10047
rect 10793 10013 10827 10047
rect 10827 10013 10836 10047
rect 10784 10004 10836 10013
rect 11060 10047 11112 10056
rect 11060 10013 11069 10047
rect 11069 10013 11103 10047
rect 11103 10013 11112 10047
rect 11060 10004 11112 10013
rect 11244 10047 11296 10056
rect 11244 10013 11253 10047
rect 11253 10013 11287 10047
rect 11287 10013 11296 10047
rect 12900 10072 12952 10124
rect 11244 10004 11296 10013
rect 13452 10004 13504 10056
rect 4252 9868 4304 9920
rect 4804 9868 4856 9920
rect 6368 9868 6420 9920
rect 7932 9911 7984 9920
rect 7932 9877 7941 9911
rect 7941 9877 7975 9911
rect 7975 9877 7984 9911
rect 7932 9868 7984 9877
rect 9864 9868 9916 9920
rect 10048 9868 10100 9920
rect 13728 9936 13780 9988
rect 14004 9936 14056 9988
rect 11704 9911 11756 9920
rect 11704 9877 11713 9911
rect 11713 9877 11747 9911
rect 11747 9877 11756 9911
rect 11704 9868 11756 9877
rect 12164 9868 12216 9920
rect 13636 9868 13688 9920
rect 14280 9911 14332 9920
rect 14280 9877 14289 9911
rect 14289 9877 14323 9911
rect 14323 9877 14332 9911
rect 14280 9868 14332 9877
rect 5547 9766 5599 9818
rect 5611 9766 5663 9818
rect 5675 9766 5727 9818
rect 5739 9766 5791 9818
rect 5803 9766 5855 9818
rect 10144 9766 10196 9818
rect 10208 9766 10260 9818
rect 10272 9766 10324 9818
rect 10336 9766 10388 9818
rect 10400 9766 10452 9818
rect 3884 9664 3936 9716
rect 4344 9664 4396 9716
rect 4528 9664 4580 9716
rect 5356 9664 5408 9716
rect 6460 9664 6512 9716
rect 7196 9707 7248 9716
rect 1400 9571 1452 9580
rect 1400 9537 1409 9571
rect 1409 9537 1443 9571
rect 1443 9537 1452 9571
rect 1400 9528 1452 9537
rect 2780 9460 2832 9512
rect 2872 9392 2924 9444
rect 4252 9571 4304 9580
rect 4252 9537 4261 9571
rect 4261 9537 4295 9571
rect 4295 9537 4304 9571
rect 4252 9528 4304 9537
rect 4436 9571 4488 9580
rect 4436 9537 4445 9571
rect 4445 9537 4479 9571
rect 4479 9537 4488 9571
rect 4436 9528 4488 9537
rect 4620 9571 4672 9580
rect 4620 9537 4629 9571
rect 4629 9537 4663 9571
rect 4663 9537 4672 9571
rect 4620 9528 4672 9537
rect 5448 9596 5500 9648
rect 7196 9673 7205 9707
rect 7205 9673 7239 9707
rect 7239 9673 7248 9707
rect 7196 9664 7248 9673
rect 9864 9664 9916 9716
rect 11704 9664 11756 9716
rect 3976 9460 4028 9512
rect 4804 9571 4856 9580
rect 4804 9537 4813 9571
rect 4813 9537 4847 9571
rect 4847 9537 4856 9571
rect 4804 9528 4856 9537
rect 6368 9571 6420 9580
rect 4988 9392 5040 9444
rect 6368 9537 6377 9571
rect 6377 9537 6411 9571
rect 6411 9537 6420 9571
rect 6368 9528 6420 9537
rect 6828 9528 6880 9580
rect 7104 9596 7156 9648
rect 7748 9596 7800 9648
rect 14280 9596 14332 9648
rect 5908 9503 5960 9512
rect 5908 9469 5917 9503
rect 5917 9469 5951 9503
rect 5951 9469 5960 9503
rect 5908 9460 5960 9469
rect 7656 9503 7708 9512
rect 7656 9469 7665 9503
rect 7665 9469 7699 9503
rect 7699 9469 7708 9503
rect 7656 9460 7708 9469
rect 7748 9460 7800 9512
rect 7932 9460 7984 9512
rect 8116 9571 8168 9580
rect 8116 9537 8125 9571
rect 8125 9537 8159 9571
rect 8159 9537 8168 9571
rect 8116 9528 8168 9537
rect 8576 9528 8628 9580
rect 8944 9528 8996 9580
rect 8668 9460 8720 9512
rect 9588 9528 9640 9580
rect 9956 9571 10008 9580
rect 9956 9537 9965 9571
rect 9965 9537 9999 9571
rect 9999 9537 10008 9571
rect 9956 9528 10008 9537
rect 10600 9528 10652 9580
rect 11612 9571 11664 9580
rect 11612 9537 11621 9571
rect 11621 9537 11655 9571
rect 11655 9537 11664 9571
rect 11612 9528 11664 9537
rect 11888 9528 11940 9580
rect 12256 9571 12308 9580
rect 12256 9537 12265 9571
rect 12265 9537 12299 9571
rect 12299 9537 12308 9571
rect 12256 9528 12308 9537
rect 12808 9528 12860 9580
rect 10232 9460 10284 9512
rect 3056 9324 3108 9376
rect 4068 9324 4120 9376
rect 4252 9367 4304 9376
rect 4252 9333 4261 9367
rect 4261 9333 4295 9367
rect 4295 9333 4304 9367
rect 4252 9324 4304 9333
rect 6920 9392 6972 9444
rect 8392 9392 8444 9444
rect 9680 9392 9732 9444
rect 10692 9392 10744 9444
rect 10508 9324 10560 9376
rect 11428 9460 11480 9512
rect 12164 9460 12216 9512
rect 12900 9460 12952 9512
rect 13728 9392 13780 9444
rect 12348 9324 12400 9376
rect 14004 9367 14056 9376
rect 14004 9333 14013 9367
rect 14013 9333 14047 9367
rect 14047 9333 14056 9367
rect 14004 9324 14056 9333
rect 3248 9222 3300 9274
rect 3312 9222 3364 9274
rect 3376 9222 3428 9274
rect 3440 9222 3492 9274
rect 3504 9222 3556 9274
rect 7846 9222 7898 9274
rect 7910 9222 7962 9274
rect 7974 9222 8026 9274
rect 8038 9222 8090 9274
rect 8102 9222 8154 9274
rect 12443 9222 12495 9274
rect 12507 9222 12559 9274
rect 12571 9222 12623 9274
rect 12635 9222 12687 9274
rect 12699 9222 12751 9274
rect 2780 9163 2832 9172
rect 2780 9129 2789 9163
rect 2789 9129 2823 9163
rect 2823 9129 2832 9163
rect 2780 9120 2832 9129
rect 2872 9095 2924 9104
rect 2872 9061 2881 9095
rect 2881 9061 2915 9095
rect 2915 9061 2924 9095
rect 3608 9120 3660 9172
rect 7656 9120 7708 9172
rect 8668 9163 8720 9172
rect 8668 9129 8677 9163
rect 8677 9129 8711 9163
rect 8711 9129 8720 9163
rect 8668 9120 8720 9129
rect 9588 9120 9640 9172
rect 10048 9120 10100 9172
rect 10232 9120 10284 9172
rect 11888 9120 11940 9172
rect 12900 9120 12952 9172
rect 2872 9052 2924 9061
rect 3884 9052 3936 9104
rect 6828 9052 6880 9104
rect 3148 8984 3200 9036
rect 8300 9052 8352 9104
rect 8576 9052 8628 9104
rect 3240 8916 3292 8968
rect 3976 8959 4028 8968
rect 3976 8925 3985 8959
rect 3985 8925 4019 8959
rect 4019 8925 4028 8959
rect 3976 8916 4028 8925
rect 4068 8959 4120 8968
rect 4068 8925 4077 8959
rect 4077 8925 4111 8959
rect 4111 8925 4120 8959
rect 4620 8959 4672 8968
rect 4068 8916 4120 8925
rect 4620 8925 4629 8959
rect 4629 8925 4663 8959
rect 4663 8925 4672 8959
rect 4620 8916 4672 8925
rect 7748 8984 7800 9036
rect 7380 8916 7432 8968
rect 9496 8984 9548 9036
rect 9772 9027 9824 9036
rect 8208 8959 8260 8968
rect 8208 8925 8217 8959
rect 8217 8925 8251 8959
rect 8251 8925 8260 8959
rect 8208 8916 8260 8925
rect 8300 8916 8352 8968
rect 9772 8993 9781 9027
rect 9781 8993 9815 9027
rect 9815 8993 9824 9027
rect 9772 8984 9824 8993
rect 10692 8984 10744 9036
rect 12072 8984 12124 9036
rect 15016 9027 15068 9036
rect 15016 8993 15025 9027
rect 15025 8993 15059 9027
rect 15059 8993 15068 9027
rect 15016 8984 15068 8993
rect 3700 8848 3752 8900
rect 4252 8848 4304 8900
rect 4528 8848 4580 8900
rect 4896 8891 4948 8900
rect 4896 8857 4905 8891
rect 4905 8857 4939 8891
rect 4939 8857 4948 8891
rect 4896 8848 4948 8857
rect 5356 8848 5408 8900
rect 4344 8780 4396 8832
rect 6460 8823 6512 8832
rect 6460 8789 6469 8823
rect 6469 8789 6503 8823
rect 6503 8789 6512 8823
rect 6460 8780 6512 8789
rect 7748 8823 7800 8832
rect 7748 8789 7757 8823
rect 7757 8789 7791 8823
rect 7791 8789 7800 8823
rect 8944 8823 8996 8832
rect 7748 8780 7800 8789
rect 8944 8789 8953 8823
rect 8953 8789 8987 8823
rect 8987 8789 8996 8823
rect 8944 8780 8996 8789
rect 9956 8780 10008 8832
rect 12164 8848 12216 8900
rect 12624 8780 12676 8832
rect 13360 8848 13412 8900
rect 13544 8848 13596 8900
rect 5547 8678 5599 8730
rect 5611 8678 5663 8730
rect 5675 8678 5727 8730
rect 5739 8678 5791 8730
rect 5803 8678 5855 8730
rect 10144 8678 10196 8730
rect 10208 8678 10260 8730
rect 10272 8678 10324 8730
rect 10336 8678 10388 8730
rect 10400 8678 10452 8730
rect 3976 8576 4028 8628
rect 4068 8576 4120 8628
rect 4896 8576 4948 8628
rect 7196 8576 7248 8628
rect 7748 8619 7800 8628
rect 7748 8585 7757 8619
rect 7757 8585 7791 8619
rect 7791 8585 7800 8619
rect 7748 8576 7800 8585
rect 3884 8508 3936 8560
rect 4344 8551 4396 8560
rect 4344 8517 4353 8551
rect 4353 8517 4387 8551
rect 4387 8517 4396 8551
rect 4344 8508 4396 8517
rect 4988 8440 5040 8492
rect 6460 8508 6512 8560
rect 6828 8508 6880 8560
rect 8668 8508 8720 8560
rect 7380 8483 7432 8492
rect 4620 8415 4672 8424
rect 4620 8381 4629 8415
rect 4629 8381 4663 8415
rect 4663 8381 4672 8415
rect 4620 8372 4672 8381
rect 5448 8372 5500 8424
rect 7380 8449 7389 8483
rect 7389 8449 7423 8483
rect 7423 8449 7432 8483
rect 7380 8440 7432 8449
rect 7748 8440 7800 8492
rect 8484 8483 8536 8492
rect 8484 8449 8493 8483
rect 8493 8449 8527 8483
rect 8527 8449 8536 8483
rect 8484 8440 8536 8449
rect 8760 8483 8812 8492
rect 8760 8449 8769 8483
rect 8769 8449 8803 8483
rect 8803 8449 8812 8483
rect 8760 8440 8812 8449
rect 9496 8576 9548 8628
rect 14004 8576 14056 8628
rect 7472 8372 7524 8424
rect 9220 8415 9272 8424
rect 8208 8304 8260 8356
rect 9220 8381 9229 8415
rect 9229 8381 9263 8415
rect 9263 8381 9272 8415
rect 9220 8372 9272 8381
rect 12256 8508 12308 8560
rect 13452 8508 13504 8560
rect 9680 8372 9732 8424
rect 11796 8440 11848 8492
rect 11980 8440 12032 8492
rect 13544 8372 13596 8424
rect 14188 8415 14240 8424
rect 14188 8381 14197 8415
rect 14197 8381 14231 8415
rect 14231 8381 14240 8415
rect 14188 8372 14240 8381
rect 12624 8304 12676 8356
rect 5356 8279 5408 8288
rect 5356 8245 5365 8279
rect 5365 8245 5399 8279
rect 5399 8245 5408 8279
rect 5356 8236 5408 8245
rect 5816 8236 5868 8288
rect 9128 8236 9180 8288
rect 9956 8236 10008 8288
rect 10784 8279 10836 8288
rect 10784 8245 10793 8279
rect 10793 8245 10827 8279
rect 10827 8245 10836 8279
rect 10784 8236 10836 8245
rect 3248 8134 3300 8186
rect 3312 8134 3364 8186
rect 3376 8134 3428 8186
rect 3440 8134 3492 8186
rect 3504 8134 3556 8186
rect 7846 8134 7898 8186
rect 7910 8134 7962 8186
rect 7974 8134 8026 8186
rect 8038 8134 8090 8186
rect 8102 8134 8154 8186
rect 12443 8134 12495 8186
rect 12507 8134 12559 8186
rect 12571 8134 12623 8186
rect 12635 8134 12687 8186
rect 12699 8134 12751 8186
rect 9220 8032 9272 8084
rect 14188 8032 14240 8084
rect 11704 8007 11756 8016
rect 11704 7973 11713 8007
rect 11713 7973 11747 8007
rect 11747 7973 11756 8007
rect 11704 7964 11756 7973
rect 2504 7939 2556 7948
rect 2504 7905 2513 7939
rect 2513 7905 2547 7939
rect 2547 7905 2556 7939
rect 2504 7896 2556 7905
rect 5448 7939 5500 7948
rect 5448 7905 5457 7939
rect 5457 7905 5491 7939
rect 5491 7905 5500 7939
rect 5448 7896 5500 7905
rect 5816 7939 5868 7948
rect 5816 7905 5825 7939
rect 5825 7905 5859 7939
rect 5859 7905 5868 7939
rect 5816 7896 5868 7905
rect 7104 7896 7156 7948
rect 8760 7896 8812 7948
rect 1676 7828 1728 7880
rect 2688 7871 2740 7880
rect 2688 7837 2697 7871
rect 2697 7837 2731 7871
rect 2731 7837 2740 7871
rect 2688 7828 2740 7837
rect 2964 7828 3016 7880
rect 7380 7871 7432 7880
rect 7380 7837 7389 7871
rect 7389 7837 7423 7871
rect 7423 7837 7432 7871
rect 7380 7828 7432 7837
rect 7748 7871 7800 7880
rect 7748 7837 7757 7871
rect 7757 7837 7791 7871
rect 7791 7837 7800 7871
rect 7748 7828 7800 7837
rect 8208 7871 8260 7880
rect 8208 7837 8217 7871
rect 8217 7837 8251 7871
rect 8251 7837 8260 7871
rect 8208 7828 8260 7837
rect 8668 7828 8720 7880
rect 12440 7939 12492 7948
rect 12440 7905 12449 7939
rect 12449 7905 12483 7939
rect 12483 7905 12492 7939
rect 12440 7896 12492 7905
rect 9680 7871 9732 7880
rect 9680 7837 9689 7871
rect 9689 7837 9723 7871
rect 9723 7837 9732 7871
rect 9680 7828 9732 7837
rect 9956 7871 10008 7880
rect 9956 7837 9965 7871
rect 9965 7837 9999 7871
rect 9999 7837 10008 7871
rect 9956 7828 10008 7837
rect 12164 7871 12216 7880
rect 12164 7837 12173 7871
rect 12173 7837 12207 7871
rect 12207 7837 12216 7871
rect 12164 7828 12216 7837
rect 6736 7760 6788 7812
rect 8484 7760 8536 7812
rect 10784 7760 10836 7812
rect 1952 7692 2004 7744
rect 2320 7692 2372 7744
rect 3332 7735 3384 7744
rect 3332 7701 3341 7735
rect 3341 7701 3375 7735
rect 3375 7701 3384 7735
rect 3332 7692 3384 7701
rect 3884 7692 3936 7744
rect 5356 7735 5408 7744
rect 5356 7701 5365 7735
rect 5365 7701 5399 7735
rect 5399 7701 5408 7735
rect 5356 7692 5408 7701
rect 8576 7692 8628 7744
rect 8944 7692 8996 7744
rect 12348 7692 12400 7744
rect 13452 7692 13504 7744
rect 14096 7735 14148 7744
rect 14096 7701 14105 7735
rect 14105 7701 14139 7735
rect 14139 7701 14148 7735
rect 14096 7692 14148 7701
rect 5547 7590 5599 7642
rect 5611 7590 5663 7642
rect 5675 7590 5727 7642
rect 5739 7590 5791 7642
rect 5803 7590 5855 7642
rect 10144 7590 10196 7642
rect 10208 7590 10260 7642
rect 10272 7590 10324 7642
rect 10336 7590 10388 7642
rect 10400 7590 10452 7642
rect 7472 7488 7524 7540
rect 7748 7488 7800 7540
rect 11428 7488 11480 7540
rect 12164 7488 12216 7540
rect 3332 7420 3384 7472
rect 7380 7420 7432 7472
rect 8576 7420 8628 7472
rect 9128 7463 9180 7472
rect 9128 7429 9137 7463
rect 9137 7429 9171 7463
rect 9171 7429 9180 7463
rect 9128 7420 9180 7429
rect 10508 7420 10560 7472
rect 12348 7420 12400 7472
rect 13268 7488 13320 7540
rect 13728 7531 13780 7540
rect 13728 7497 13737 7531
rect 13737 7497 13771 7531
rect 13771 7497 13780 7531
rect 13728 7488 13780 7497
rect 1952 7395 2004 7404
rect 1952 7361 1961 7395
rect 1961 7361 1995 7395
rect 1995 7361 2004 7395
rect 1952 7352 2004 7361
rect 2320 7395 2372 7404
rect 2320 7361 2329 7395
rect 2329 7361 2363 7395
rect 2363 7361 2372 7395
rect 2320 7352 2372 7361
rect 4160 7395 4212 7404
rect 4160 7361 4169 7395
rect 4169 7361 4203 7395
rect 4203 7361 4212 7395
rect 4160 7352 4212 7361
rect 4620 7395 4672 7404
rect 4620 7361 4629 7395
rect 4629 7361 4663 7395
rect 4663 7361 4672 7395
rect 4620 7352 4672 7361
rect 7104 7395 7156 7404
rect 7104 7361 7113 7395
rect 7113 7361 7147 7395
rect 7147 7361 7156 7395
rect 7104 7352 7156 7361
rect 7196 7395 7248 7404
rect 7196 7361 7205 7395
rect 7205 7361 7239 7395
rect 7239 7361 7248 7395
rect 7196 7352 7248 7361
rect 9496 7352 9548 7404
rect 9588 7395 9640 7404
rect 9588 7361 9597 7395
rect 9597 7361 9631 7395
rect 9631 7361 9640 7395
rect 10140 7395 10192 7404
rect 9588 7352 9640 7361
rect 10140 7361 10149 7395
rect 10149 7361 10183 7395
rect 10183 7361 10192 7395
rect 10140 7352 10192 7361
rect 11704 7352 11756 7404
rect 13360 7352 13412 7404
rect 6828 7284 6880 7336
rect 7748 7284 7800 7336
rect 4712 7216 4764 7268
rect 4436 7191 4488 7200
rect 4436 7157 4445 7191
rect 4445 7157 4479 7191
rect 4479 7157 4488 7191
rect 4436 7148 4488 7157
rect 4528 7148 4580 7200
rect 6736 7191 6788 7200
rect 6736 7157 6745 7191
rect 6745 7157 6779 7191
rect 6779 7157 6788 7191
rect 6736 7148 6788 7157
rect 7288 7191 7340 7200
rect 7288 7157 7297 7191
rect 7297 7157 7331 7191
rect 7331 7157 7340 7191
rect 7288 7148 7340 7157
rect 7380 7191 7432 7200
rect 7380 7157 7389 7191
rect 7389 7157 7423 7191
rect 7423 7157 7432 7191
rect 10140 7216 10192 7268
rect 11612 7216 11664 7268
rect 7380 7148 7432 7157
rect 10508 7148 10560 7200
rect 11428 7148 11480 7200
rect 3248 7046 3300 7098
rect 3312 7046 3364 7098
rect 3376 7046 3428 7098
rect 3440 7046 3492 7098
rect 3504 7046 3556 7098
rect 7846 7046 7898 7098
rect 7910 7046 7962 7098
rect 7974 7046 8026 7098
rect 8038 7046 8090 7098
rect 8102 7046 8154 7098
rect 12443 7046 12495 7098
rect 12507 7046 12559 7098
rect 12571 7046 12623 7098
rect 12635 7046 12687 7098
rect 12699 7046 12751 7098
rect 2504 6944 2556 6996
rect 3700 6944 3752 6996
rect 4160 6876 4212 6928
rect 3056 6808 3108 6860
rect 3608 6851 3660 6860
rect 2044 6783 2096 6792
rect 2044 6749 2053 6783
rect 2053 6749 2087 6783
rect 2087 6749 2096 6783
rect 2044 6740 2096 6749
rect 2688 6672 2740 6724
rect 2320 6647 2372 6656
rect 2320 6613 2329 6647
rect 2329 6613 2363 6647
rect 2363 6613 2372 6647
rect 2320 6604 2372 6613
rect 3608 6817 3617 6851
rect 3617 6817 3651 6851
rect 3651 6817 3660 6851
rect 3608 6808 3660 6817
rect 4528 6808 4580 6860
rect 7380 6944 7432 6996
rect 7196 6876 7248 6928
rect 8852 6876 8904 6928
rect 9588 6944 9640 6996
rect 10140 6944 10192 6996
rect 11152 6944 11204 6996
rect 3148 6672 3200 6724
rect 3884 6740 3936 6792
rect 4160 6783 4212 6792
rect 4160 6749 4169 6783
rect 4169 6749 4203 6783
rect 4203 6749 4212 6783
rect 4160 6740 4212 6749
rect 4620 6783 4672 6792
rect 4620 6749 4629 6783
rect 4629 6749 4663 6783
rect 4663 6749 4672 6783
rect 4620 6740 4672 6749
rect 4896 6808 4948 6860
rect 5908 6808 5960 6860
rect 5540 6740 5592 6792
rect 6644 6740 6696 6792
rect 14464 6876 14516 6928
rect 4528 6672 4580 6724
rect 6552 6672 6604 6724
rect 3240 6604 3292 6656
rect 3700 6604 3752 6656
rect 3976 6604 4028 6656
rect 5080 6647 5132 6656
rect 5080 6613 5089 6647
rect 5089 6613 5123 6647
rect 5123 6613 5132 6647
rect 5080 6604 5132 6613
rect 5172 6604 5224 6656
rect 6460 6604 6512 6656
rect 6828 6604 6880 6656
rect 8576 6740 8628 6792
rect 9036 6740 9088 6792
rect 9220 6783 9272 6792
rect 9220 6749 9229 6783
rect 9229 6749 9263 6783
rect 9263 6749 9272 6783
rect 9220 6740 9272 6749
rect 11520 6808 11572 6860
rect 13636 6808 13688 6860
rect 11428 6783 11480 6792
rect 7472 6604 7524 6656
rect 8668 6672 8720 6724
rect 7840 6604 7892 6656
rect 8484 6647 8536 6656
rect 8484 6613 8493 6647
rect 8493 6613 8527 6647
rect 8527 6613 8536 6647
rect 8484 6604 8536 6613
rect 9128 6604 9180 6656
rect 9588 6672 9640 6724
rect 11152 6672 11204 6724
rect 10968 6604 11020 6656
rect 11428 6749 11437 6783
rect 11437 6749 11471 6783
rect 11471 6749 11480 6783
rect 11428 6740 11480 6749
rect 11336 6715 11388 6724
rect 11336 6681 11345 6715
rect 11345 6681 11379 6715
rect 11379 6681 11388 6715
rect 11612 6740 11664 6792
rect 11336 6672 11388 6681
rect 11704 6715 11756 6724
rect 11704 6681 11713 6715
rect 11713 6681 11747 6715
rect 11747 6681 11756 6715
rect 11704 6672 11756 6681
rect 11796 6672 11848 6724
rect 12348 6672 12400 6724
rect 13544 6672 13596 6724
rect 14096 6647 14148 6656
rect 14096 6613 14105 6647
rect 14105 6613 14139 6647
rect 14139 6613 14148 6647
rect 14096 6604 14148 6613
rect 5547 6502 5599 6554
rect 5611 6502 5663 6554
rect 5675 6502 5727 6554
rect 5739 6502 5791 6554
rect 5803 6502 5855 6554
rect 10144 6502 10196 6554
rect 10208 6502 10260 6554
rect 10272 6502 10324 6554
rect 10336 6502 10388 6554
rect 10400 6502 10452 6554
rect 3148 6443 3200 6452
rect 3148 6409 3157 6443
rect 3157 6409 3191 6443
rect 3191 6409 3200 6443
rect 3148 6400 3200 6409
rect 3608 6400 3660 6452
rect 5080 6443 5132 6452
rect 1676 6332 1728 6384
rect 2412 6332 2464 6384
rect 3056 6332 3108 6384
rect 5080 6409 5089 6443
rect 5089 6409 5123 6443
rect 5123 6409 5132 6443
rect 5080 6400 5132 6409
rect 6000 6332 6052 6384
rect 6552 6332 6604 6384
rect 7380 6400 7432 6452
rect 3240 6307 3292 6316
rect 3240 6273 3249 6307
rect 3249 6273 3283 6307
rect 3283 6273 3292 6307
rect 3240 6264 3292 6273
rect 2320 6196 2372 6248
rect 2964 6196 3016 6248
rect 3608 6264 3660 6316
rect 3976 6307 4028 6316
rect 3976 6273 3985 6307
rect 3985 6273 4019 6307
rect 4019 6273 4028 6307
rect 3976 6264 4028 6273
rect 4436 6307 4488 6316
rect 4436 6273 4445 6307
rect 4445 6273 4479 6307
rect 4479 6273 4488 6307
rect 4436 6264 4488 6273
rect 4804 6264 4856 6316
rect 3884 6196 3936 6248
rect 4160 6196 4212 6248
rect 5356 6264 5408 6316
rect 5816 6307 5868 6316
rect 5816 6273 5825 6307
rect 5825 6273 5859 6307
rect 5859 6273 5868 6307
rect 5816 6264 5868 6273
rect 7380 6307 7432 6316
rect 4988 6196 5040 6248
rect 5172 6239 5224 6248
rect 5172 6205 5181 6239
rect 5181 6205 5215 6239
rect 5215 6205 5224 6239
rect 5172 6196 5224 6205
rect 5264 6239 5316 6248
rect 5264 6205 5273 6239
rect 5273 6205 5307 6239
rect 5307 6205 5316 6239
rect 5264 6196 5316 6205
rect 5448 6196 5500 6248
rect 6092 6196 6144 6248
rect 2780 6128 2832 6180
rect 5080 6128 5132 6180
rect 5908 6128 5960 6180
rect 7380 6273 7389 6307
rect 7389 6273 7423 6307
rect 7423 6273 7432 6307
rect 7380 6264 7432 6273
rect 8576 6400 8628 6452
rect 11704 6400 11756 6452
rect 12164 6400 12216 6452
rect 7840 6375 7892 6384
rect 7840 6341 7849 6375
rect 7849 6341 7883 6375
rect 7883 6341 7892 6375
rect 7840 6332 7892 6341
rect 9128 6332 9180 6384
rect 10048 6332 10100 6384
rect 10508 6332 10560 6384
rect 9864 6307 9916 6316
rect 9864 6273 9873 6307
rect 9873 6273 9907 6307
rect 9907 6273 9916 6307
rect 10232 6307 10284 6316
rect 9864 6264 9916 6273
rect 10232 6273 10266 6307
rect 10266 6273 10284 6307
rect 10232 6264 10284 6273
rect 11244 6264 11296 6316
rect 11704 6307 11756 6316
rect 11704 6273 11713 6307
rect 11713 6273 11747 6307
rect 11747 6273 11756 6307
rect 11704 6264 11756 6273
rect 11888 6307 11940 6316
rect 11888 6273 11897 6307
rect 11897 6273 11931 6307
rect 11931 6273 11940 6307
rect 11888 6264 11940 6273
rect 12348 6264 12400 6316
rect 7380 6128 7432 6180
rect 4620 6060 4672 6112
rect 5632 6060 5684 6112
rect 6092 6060 6144 6112
rect 7472 6103 7524 6112
rect 7472 6069 7481 6103
rect 7481 6069 7515 6103
rect 7515 6069 7524 6103
rect 7472 6060 7524 6069
rect 9036 6196 9088 6248
rect 9404 6128 9456 6180
rect 9220 6060 9272 6112
rect 9496 6060 9548 6112
rect 11428 6060 11480 6112
rect 13360 6196 13412 6248
rect 12164 6128 12216 6180
rect 14464 6128 14516 6180
rect 13360 6060 13412 6112
rect 3248 5958 3300 6010
rect 3312 5958 3364 6010
rect 3376 5958 3428 6010
rect 3440 5958 3492 6010
rect 3504 5958 3556 6010
rect 7846 5958 7898 6010
rect 7910 5958 7962 6010
rect 7974 5958 8026 6010
rect 8038 5958 8090 6010
rect 8102 5958 8154 6010
rect 12443 5958 12495 6010
rect 12507 5958 12559 6010
rect 12571 5958 12623 6010
rect 12635 5958 12687 6010
rect 12699 5958 12751 6010
rect 2044 5856 2096 5908
rect 4620 5856 4672 5908
rect 4804 5899 4856 5908
rect 4804 5865 4813 5899
rect 4813 5865 4847 5899
rect 4847 5865 4856 5899
rect 4804 5856 4856 5865
rect 5264 5856 5316 5908
rect 2688 5788 2740 5840
rect 1676 5720 1728 5772
rect 3240 5763 3292 5772
rect 2688 5652 2740 5704
rect 3240 5729 3249 5763
rect 3249 5729 3283 5763
rect 3283 5729 3292 5763
rect 3240 5720 3292 5729
rect 4436 5788 4488 5840
rect 7196 5856 7248 5908
rect 9956 5856 10008 5908
rect 13544 5856 13596 5908
rect 8024 5788 8076 5840
rect 9496 5788 9548 5840
rect 6736 5720 6788 5772
rect 4068 5652 4120 5704
rect 4620 5695 4672 5704
rect 4620 5661 4629 5695
rect 4629 5661 4663 5695
rect 4663 5661 4672 5695
rect 4620 5652 4672 5661
rect 5632 5652 5684 5704
rect 2412 5584 2464 5636
rect 6092 5652 6144 5704
rect 6184 5695 6236 5704
rect 6184 5661 6193 5695
rect 6193 5661 6227 5695
rect 6227 5661 6236 5695
rect 6184 5652 6236 5661
rect 7656 5720 7708 5772
rect 7748 5720 7800 5772
rect 8668 5763 8720 5772
rect 8668 5729 8677 5763
rect 8677 5729 8711 5763
rect 8711 5729 8720 5763
rect 8668 5720 8720 5729
rect 8852 5720 8904 5772
rect 9220 5720 9272 5772
rect 9404 5720 9456 5772
rect 9588 5720 9640 5772
rect 12072 5788 12124 5840
rect 12624 5788 12676 5840
rect 10968 5720 11020 5772
rect 7104 5584 7156 5636
rect 3056 5516 3108 5568
rect 3608 5516 3660 5568
rect 4804 5516 4856 5568
rect 6736 5516 6788 5568
rect 8024 5695 8076 5704
rect 8024 5661 8033 5695
rect 8033 5661 8067 5695
rect 8067 5661 8076 5695
rect 8024 5652 8076 5661
rect 8576 5652 8628 5704
rect 8760 5695 8812 5704
rect 8760 5661 8769 5695
rect 8769 5661 8803 5695
rect 8803 5661 8812 5695
rect 8760 5652 8812 5661
rect 10508 5652 10560 5704
rect 10876 5695 10928 5704
rect 10876 5661 10885 5695
rect 10885 5661 10919 5695
rect 10919 5661 10928 5695
rect 10876 5652 10928 5661
rect 11060 5695 11112 5704
rect 11060 5661 11069 5695
rect 11069 5661 11103 5695
rect 11103 5661 11112 5695
rect 11060 5652 11112 5661
rect 13636 5720 13688 5772
rect 14464 5695 14516 5704
rect 14464 5661 14473 5695
rect 14473 5661 14507 5695
rect 14507 5661 14516 5695
rect 14464 5652 14516 5661
rect 9220 5584 9272 5636
rect 10048 5584 10100 5636
rect 11796 5627 11848 5636
rect 11796 5593 11805 5627
rect 11805 5593 11839 5627
rect 11839 5593 11848 5627
rect 11796 5584 11848 5593
rect 8392 5516 8444 5568
rect 11428 5516 11480 5568
rect 13360 5516 13412 5568
rect 14096 5559 14148 5568
rect 14096 5525 14105 5559
rect 14105 5525 14139 5559
rect 14139 5525 14148 5559
rect 14096 5516 14148 5525
rect 14188 5516 14240 5568
rect 5547 5414 5599 5466
rect 5611 5414 5663 5466
rect 5675 5414 5727 5466
rect 5739 5414 5791 5466
rect 5803 5414 5855 5466
rect 10144 5414 10196 5466
rect 10208 5414 10260 5466
rect 10272 5414 10324 5466
rect 10336 5414 10388 5466
rect 10400 5414 10452 5466
rect 3240 5312 3292 5364
rect 1676 5219 1728 5228
rect 1676 5185 1685 5219
rect 1685 5185 1719 5219
rect 1719 5185 1728 5219
rect 1676 5176 1728 5185
rect 2688 5244 2740 5296
rect 2504 5219 2556 5228
rect 2504 5185 2513 5219
rect 2513 5185 2547 5219
rect 2547 5185 2556 5219
rect 2504 5176 2556 5185
rect 2964 5176 3016 5228
rect 2688 5151 2740 5160
rect 2688 5117 2697 5151
rect 2697 5117 2731 5151
rect 2731 5117 2740 5151
rect 2688 5108 2740 5117
rect 2872 5040 2924 5092
rect 3240 5108 3292 5160
rect 3976 5312 4028 5364
rect 4068 5312 4120 5364
rect 5908 5312 5960 5364
rect 6920 5312 6972 5364
rect 7288 5312 7340 5364
rect 10508 5355 10560 5364
rect 3608 5176 3660 5228
rect 3700 5219 3752 5228
rect 3700 5185 3709 5219
rect 3709 5185 3743 5219
rect 3743 5185 3752 5219
rect 3700 5176 3752 5185
rect 4160 5176 4212 5228
rect 4528 5176 4580 5228
rect 4712 5219 4764 5228
rect 4712 5185 4721 5219
rect 4721 5185 4755 5219
rect 4755 5185 4764 5219
rect 4712 5176 4764 5185
rect 5080 5219 5132 5228
rect 5080 5185 5089 5219
rect 5089 5185 5123 5219
rect 5123 5185 5132 5219
rect 5264 5219 5316 5228
rect 5080 5176 5132 5185
rect 5264 5185 5273 5219
rect 5273 5185 5307 5219
rect 5307 5185 5316 5219
rect 5264 5176 5316 5185
rect 5816 5219 5868 5228
rect 5816 5185 5825 5219
rect 5825 5185 5859 5219
rect 5859 5185 5868 5219
rect 5816 5176 5868 5185
rect 5908 5219 5960 5228
rect 5908 5185 5917 5219
rect 5917 5185 5951 5219
rect 5951 5185 5960 5219
rect 5908 5176 5960 5185
rect 6276 5176 6328 5228
rect 7196 5244 7248 5296
rect 7564 5244 7616 5296
rect 8300 5244 8352 5296
rect 8392 5244 8444 5296
rect 6828 5219 6880 5228
rect 6828 5185 6837 5219
rect 6837 5185 6871 5219
rect 6871 5185 6880 5219
rect 6828 5176 6880 5185
rect 6920 5176 6972 5228
rect 8484 5176 8536 5228
rect 8852 5176 8904 5228
rect 9220 5244 9272 5296
rect 10508 5321 10517 5355
rect 10517 5321 10551 5355
rect 10551 5321 10560 5355
rect 10508 5312 10560 5321
rect 11520 5355 11572 5364
rect 11520 5321 11529 5355
rect 11529 5321 11563 5355
rect 11563 5321 11572 5355
rect 11520 5312 11572 5321
rect 11980 5355 12032 5364
rect 11980 5321 11989 5355
rect 11989 5321 12023 5355
rect 12023 5321 12032 5355
rect 11980 5312 12032 5321
rect 9680 5176 9732 5228
rect 13360 5244 13412 5296
rect 10508 5219 10560 5228
rect 10508 5185 10517 5219
rect 10517 5185 10551 5219
rect 10551 5185 10560 5219
rect 10508 5176 10560 5185
rect 10692 5219 10744 5228
rect 10692 5185 10701 5219
rect 10701 5185 10735 5219
rect 10735 5185 10744 5219
rect 10692 5176 10744 5185
rect 11980 5176 12032 5228
rect 12072 5176 12124 5228
rect 12440 5176 12492 5228
rect 12624 5219 12676 5228
rect 12624 5185 12633 5219
rect 12633 5185 12667 5219
rect 12667 5185 12676 5219
rect 12624 5176 12676 5185
rect 13820 5176 13872 5228
rect 3792 5108 3844 5160
rect 4896 5108 4948 5160
rect 6000 5108 6052 5160
rect 1400 4972 1452 5024
rect 2412 4972 2464 5024
rect 2688 4972 2740 5024
rect 3056 5015 3108 5024
rect 3056 4981 3065 5015
rect 3065 4981 3099 5015
rect 3099 4981 3108 5015
rect 3056 4972 3108 4981
rect 4160 5040 4212 5092
rect 6092 5040 6144 5092
rect 6552 5040 6604 5092
rect 6736 5108 6788 5160
rect 7564 5108 7616 5160
rect 8668 5108 8720 5160
rect 9864 5108 9916 5160
rect 10048 5151 10100 5160
rect 10048 5117 10057 5151
rect 10057 5117 10091 5151
rect 10091 5117 10100 5151
rect 10048 5108 10100 5117
rect 10784 5108 10836 5160
rect 12164 5151 12216 5160
rect 12164 5117 12173 5151
rect 12173 5117 12207 5151
rect 12207 5117 12216 5151
rect 12164 5108 12216 5117
rect 7012 5040 7064 5092
rect 7656 5040 7708 5092
rect 5356 4972 5408 5024
rect 5724 5015 5776 5024
rect 5724 4981 5733 5015
rect 5733 4981 5767 5015
rect 5767 4981 5776 5015
rect 5724 4972 5776 4981
rect 6368 4972 6420 5024
rect 6460 4972 6512 5024
rect 7564 4972 7616 5024
rect 8208 4972 8260 5024
rect 9772 5040 9824 5092
rect 9312 4972 9364 5024
rect 9496 4972 9548 5024
rect 10140 4972 10192 5024
rect 11060 4972 11112 5024
rect 12900 4972 12952 5024
rect 3248 4870 3300 4922
rect 3312 4870 3364 4922
rect 3376 4870 3428 4922
rect 3440 4870 3492 4922
rect 3504 4870 3556 4922
rect 7846 4870 7898 4922
rect 7910 4870 7962 4922
rect 7974 4870 8026 4922
rect 8038 4870 8090 4922
rect 8102 4870 8154 4922
rect 12443 4870 12495 4922
rect 12507 4870 12559 4922
rect 12571 4870 12623 4922
rect 12635 4870 12687 4922
rect 12699 4870 12751 4922
rect 3148 4768 3200 4820
rect 5264 4768 5316 4820
rect 6276 4768 6328 4820
rect 7104 4768 7156 4820
rect 8852 4768 8904 4820
rect 9312 4768 9364 4820
rect 10692 4768 10744 4820
rect 11060 4768 11112 4820
rect 12348 4768 12400 4820
rect 14096 4811 14148 4820
rect 14096 4777 14105 4811
rect 14105 4777 14139 4811
rect 14139 4777 14148 4811
rect 14096 4768 14148 4777
rect 2688 4700 2740 4752
rect 4712 4700 4764 4752
rect 1676 4632 1728 4684
rect 3056 4632 3108 4684
rect 4896 4675 4948 4684
rect 4896 4641 4905 4675
rect 4905 4641 4939 4675
rect 4939 4641 4948 4675
rect 4896 4632 4948 4641
rect 1768 4496 1820 4548
rect 2688 4496 2740 4548
rect 2964 4428 3016 4480
rect 4160 4564 4212 4616
rect 4344 4607 4396 4616
rect 4344 4573 4353 4607
rect 4353 4573 4387 4607
rect 4387 4573 4396 4607
rect 4344 4564 4396 4573
rect 4528 4564 4580 4616
rect 4804 4564 4856 4616
rect 5172 4564 5224 4616
rect 5816 4632 5868 4684
rect 5908 4675 5960 4684
rect 5908 4641 5917 4675
rect 5917 4641 5951 4675
rect 5951 4641 5960 4675
rect 5908 4632 5960 4641
rect 7380 4632 7432 4684
rect 3700 4496 3752 4548
rect 6736 4564 6788 4616
rect 7012 4564 7064 4616
rect 7564 4675 7616 4684
rect 7564 4641 7573 4675
rect 7573 4641 7607 4675
rect 7607 4641 7616 4675
rect 7564 4632 7616 4641
rect 7748 4675 7800 4684
rect 7748 4641 7757 4675
rect 7757 4641 7791 4675
rect 7791 4641 7800 4675
rect 7748 4632 7800 4641
rect 8300 4632 8352 4684
rect 9496 4675 9548 4684
rect 9496 4641 9505 4675
rect 9505 4641 9539 4675
rect 9539 4641 9548 4675
rect 9496 4632 9548 4641
rect 10140 4632 10192 4684
rect 7656 4564 7708 4616
rect 8392 4564 8444 4616
rect 3240 4428 3292 4480
rect 3792 4428 3844 4480
rect 4252 4471 4304 4480
rect 4252 4437 4261 4471
rect 4261 4437 4295 4471
rect 4295 4437 4304 4471
rect 4252 4428 4304 4437
rect 9588 4564 9640 4616
rect 10508 4632 10560 4684
rect 13636 4632 13688 4684
rect 14372 4632 14424 4684
rect 13544 4607 13596 4616
rect 13544 4573 13553 4607
rect 13553 4573 13587 4607
rect 13587 4573 13596 4607
rect 13544 4564 13596 4573
rect 14464 4607 14516 4616
rect 14464 4573 14473 4607
rect 14473 4573 14507 4607
rect 14507 4573 14516 4607
rect 14464 4564 14516 4573
rect 5908 4428 5960 4480
rect 6828 4428 6880 4480
rect 7012 4428 7064 4480
rect 8576 4428 8628 4480
rect 11428 4496 11480 4548
rect 11888 4428 11940 4480
rect 14188 4428 14240 4480
rect 5547 4326 5599 4378
rect 5611 4326 5663 4378
rect 5675 4326 5727 4378
rect 5739 4326 5791 4378
rect 5803 4326 5855 4378
rect 10144 4326 10196 4378
rect 10208 4326 10260 4378
rect 10272 4326 10324 4378
rect 10336 4326 10388 4378
rect 10400 4326 10452 4378
rect 1768 4224 1820 4276
rect 2688 4156 2740 4208
rect 4160 4156 4212 4208
rect 5908 4224 5960 4276
rect 6368 4267 6420 4276
rect 6368 4233 6377 4267
rect 6377 4233 6411 4267
rect 6411 4233 6420 4267
rect 6368 4224 6420 4233
rect 7472 4224 7524 4276
rect 6644 4156 6696 4208
rect 7196 4199 7248 4208
rect 7196 4165 7205 4199
rect 7205 4165 7239 4199
rect 7239 4165 7248 4199
rect 7196 4156 7248 4165
rect 7380 4199 7432 4208
rect 7380 4165 7389 4199
rect 7389 4165 7423 4199
rect 7423 4165 7432 4199
rect 8576 4224 8628 4276
rect 11888 4267 11940 4276
rect 11888 4233 11897 4267
rect 11897 4233 11931 4267
rect 11931 4233 11940 4267
rect 11888 4224 11940 4233
rect 13544 4224 13596 4276
rect 7380 4156 7432 4165
rect 7748 4156 7800 4208
rect 1400 4131 1452 4140
rect 1400 4097 1409 4131
rect 1409 4097 1443 4131
rect 1443 4097 1452 4131
rect 1400 4088 1452 4097
rect 2964 4088 3016 4140
rect 3516 4088 3568 4140
rect 3608 4088 3660 4140
rect 3884 4131 3936 4140
rect 3884 4097 3893 4131
rect 3893 4097 3927 4131
rect 3927 4097 3936 4131
rect 3884 4088 3936 4097
rect 2780 4020 2832 4072
rect 4804 4088 4856 4140
rect 5264 4131 5316 4140
rect 5264 4097 5273 4131
rect 5273 4097 5307 4131
rect 5307 4097 5316 4131
rect 5264 4088 5316 4097
rect 6552 4088 6604 4140
rect 7012 4088 7064 4140
rect 7104 4131 7156 4140
rect 7104 4097 7113 4131
rect 7113 4097 7147 4131
rect 7147 4097 7156 4131
rect 7104 4088 7156 4097
rect 4344 4020 4396 4072
rect 5356 4063 5408 4072
rect 5356 4029 5365 4063
rect 5365 4029 5399 4063
rect 5399 4029 5408 4063
rect 5356 4020 5408 4029
rect 5540 4020 5592 4072
rect 6460 4020 6512 4072
rect 6644 4020 6696 4072
rect 8300 4156 8352 4208
rect 8208 4088 8260 4140
rect 4528 3952 4580 4004
rect 6920 3952 6972 4004
rect 8484 4020 8536 4072
rect 9496 4088 9548 4140
rect 12348 4156 12400 4208
rect 9036 4020 9088 4072
rect 10508 4088 10560 4140
rect 11060 4088 11112 4140
rect 14096 4088 14148 4140
rect 14372 4131 14424 4140
rect 14372 4097 14381 4131
rect 14381 4097 14415 4131
rect 14415 4097 14424 4131
rect 14372 4088 14424 4097
rect 3976 3927 4028 3936
rect 3976 3893 3985 3927
rect 3985 3893 4019 3927
rect 4019 3893 4028 3927
rect 3976 3884 4028 3893
rect 4068 3884 4120 3936
rect 6828 3884 6880 3936
rect 7012 3927 7064 3936
rect 7012 3893 7021 3927
rect 7021 3893 7055 3927
rect 7055 3893 7064 3927
rect 7012 3884 7064 3893
rect 7104 3927 7156 3936
rect 7104 3893 7113 3927
rect 7113 3893 7147 3927
rect 7147 3893 7156 3927
rect 7104 3884 7156 3893
rect 7748 3884 7800 3936
rect 9772 3952 9824 4004
rect 9680 3884 9732 3936
rect 11336 4020 11388 4072
rect 11980 4063 12032 4072
rect 11980 4029 11989 4063
rect 11989 4029 12023 4063
rect 12023 4029 12032 4063
rect 11980 4020 12032 4029
rect 12900 4020 12952 4072
rect 11060 3884 11112 3936
rect 11428 3884 11480 3936
rect 12348 3927 12400 3936
rect 12348 3893 12357 3927
rect 12357 3893 12391 3927
rect 12391 3893 12400 3927
rect 12348 3884 12400 3893
rect 3248 3782 3300 3834
rect 3312 3782 3364 3834
rect 3376 3782 3428 3834
rect 3440 3782 3492 3834
rect 3504 3782 3556 3834
rect 7846 3782 7898 3834
rect 7910 3782 7962 3834
rect 7974 3782 8026 3834
rect 8038 3782 8090 3834
rect 8102 3782 8154 3834
rect 12443 3782 12495 3834
rect 12507 3782 12559 3834
rect 12571 3782 12623 3834
rect 12635 3782 12687 3834
rect 12699 3782 12751 3834
rect 2780 3723 2832 3732
rect 2780 3689 2789 3723
rect 2789 3689 2823 3723
rect 2823 3689 2832 3723
rect 2780 3680 2832 3689
rect 3608 3680 3660 3732
rect 3884 3680 3936 3732
rect 3976 3612 4028 3664
rect 4068 3587 4120 3596
rect 4068 3553 4077 3587
rect 4077 3553 4111 3587
rect 4111 3553 4120 3587
rect 4068 3544 4120 3553
rect 3424 3519 3476 3528
rect 3424 3485 3433 3519
rect 3433 3485 3467 3519
rect 3467 3485 3476 3519
rect 3424 3476 3476 3485
rect 3792 3476 3844 3528
rect 5172 3723 5224 3732
rect 5172 3689 5181 3723
rect 5181 3689 5215 3723
rect 5215 3689 5224 3723
rect 5172 3680 5224 3689
rect 8392 3723 8444 3732
rect 8392 3689 8401 3723
rect 8401 3689 8435 3723
rect 8435 3689 8444 3723
rect 8392 3680 8444 3689
rect 11980 3680 12032 3732
rect 3148 3408 3200 3460
rect 4896 3519 4948 3528
rect 5264 3544 5316 3596
rect 5448 3612 5500 3664
rect 7012 3544 7064 3596
rect 4896 3485 4923 3519
rect 4923 3485 4948 3519
rect 4896 3476 4948 3485
rect 5540 3519 5592 3528
rect 5540 3485 5549 3519
rect 5549 3485 5583 3519
rect 5583 3485 5592 3519
rect 5540 3476 5592 3485
rect 7656 3476 7708 3528
rect 10692 3612 10744 3664
rect 10876 3655 10928 3664
rect 10876 3621 10885 3655
rect 10885 3621 10919 3655
rect 10919 3621 10928 3655
rect 10876 3612 10928 3621
rect 8208 3587 8260 3596
rect 8208 3553 8217 3587
rect 8217 3553 8251 3587
rect 8251 3553 8260 3587
rect 8208 3544 8260 3553
rect 9496 3587 9548 3596
rect 9496 3553 9505 3587
rect 9505 3553 9539 3587
rect 9539 3553 9548 3587
rect 9496 3544 9548 3553
rect 9772 3544 9824 3596
rect 10508 3587 10560 3596
rect 8392 3519 8444 3528
rect 8392 3485 8401 3519
rect 8401 3485 8435 3519
rect 8435 3485 8444 3519
rect 8392 3476 8444 3485
rect 10508 3553 10517 3587
rect 10517 3553 10551 3587
rect 10551 3553 10560 3587
rect 10508 3544 10560 3553
rect 11336 3587 11388 3596
rect 11336 3553 11345 3587
rect 11345 3553 11379 3587
rect 11379 3553 11388 3587
rect 11336 3544 11388 3553
rect 12900 3544 12952 3596
rect 14372 3544 14424 3596
rect 4344 3408 4396 3460
rect 4804 3408 4856 3460
rect 5172 3408 5224 3460
rect 6920 3408 6972 3460
rect 2780 3340 2832 3392
rect 3608 3340 3660 3392
rect 3792 3383 3844 3392
rect 3792 3349 3801 3383
rect 3801 3349 3835 3383
rect 3835 3349 3844 3383
rect 3792 3340 3844 3349
rect 6644 3340 6696 3392
rect 8300 3408 8352 3460
rect 8668 3451 8720 3460
rect 8668 3417 8677 3451
rect 8677 3417 8711 3451
rect 8711 3417 8720 3451
rect 8668 3408 8720 3417
rect 8760 3408 8812 3460
rect 10140 3476 10192 3528
rect 9312 3383 9364 3392
rect 9312 3349 9321 3383
rect 9321 3349 9355 3383
rect 9355 3349 9364 3383
rect 9312 3340 9364 3349
rect 10692 3408 10744 3460
rect 11060 3408 11112 3460
rect 12348 3408 12400 3460
rect 13360 3408 13412 3460
rect 10600 3340 10652 3392
rect 11244 3383 11296 3392
rect 11244 3349 11253 3383
rect 11253 3349 11287 3383
rect 11287 3349 11296 3383
rect 11244 3340 11296 3349
rect 11336 3340 11388 3392
rect 11980 3340 12032 3392
rect 12808 3340 12860 3392
rect 12900 3340 12952 3392
rect 14464 3383 14516 3392
rect 14464 3349 14473 3383
rect 14473 3349 14507 3383
rect 14507 3349 14516 3383
rect 14464 3340 14516 3349
rect 5547 3238 5599 3290
rect 5611 3238 5663 3290
rect 5675 3238 5727 3290
rect 5739 3238 5791 3290
rect 5803 3238 5855 3290
rect 10144 3238 10196 3290
rect 10208 3238 10260 3290
rect 10272 3238 10324 3290
rect 10336 3238 10388 3290
rect 10400 3238 10452 3290
rect 3792 3136 3844 3188
rect 4344 3179 4396 3188
rect 4344 3145 4353 3179
rect 4353 3145 4387 3179
rect 4387 3145 4396 3179
rect 4344 3136 4396 3145
rect 4896 3136 4948 3188
rect 7104 3136 7156 3188
rect 3884 3068 3936 3120
rect 6920 3068 6972 3120
rect 6644 3043 6696 3052
rect 6644 3009 6653 3043
rect 6653 3009 6687 3043
rect 6687 3009 6696 3043
rect 6644 3000 6696 3009
rect 7196 3043 7248 3052
rect 7196 3009 7205 3043
rect 7205 3009 7239 3043
rect 7239 3009 7248 3043
rect 7196 3000 7248 3009
rect 9588 3136 9640 3188
rect 9680 3136 9732 3188
rect 10600 3136 10652 3188
rect 10692 3136 10744 3188
rect 13360 3136 13412 3188
rect 7748 3111 7800 3120
rect 7748 3077 7757 3111
rect 7757 3077 7791 3111
rect 7791 3077 7800 3111
rect 7748 3068 7800 3077
rect 8208 3068 8260 3120
rect 9036 3000 9088 3052
rect 9772 3068 9824 3120
rect 10784 3068 10836 3120
rect 11060 3111 11112 3120
rect 11060 3077 11069 3111
rect 11069 3077 11103 3111
rect 11103 3077 11112 3111
rect 11060 3068 11112 3077
rect 9956 3000 10008 3052
rect 10508 3000 10560 3052
rect 1676 2932 1728 2984
rect 4252 2932 4304 2984
rect 6552 2975 6604 2984
rect 6552 2941 6561 2975
rect 6561 2941 6595 2975
rect 6595 2941 6604 2975
rect 6552 2932 6604 2941
rect 8392 2932 8444 2984
rect 9220 2932 9272 2984
rect 10048 2932 10100 2984
rect 7196 2864 7248 2916
rect 5448 2796 5500 2848
rect 7748 2796 7800 2848
rect 8852 2796 8904 2848
rect 9772 2864 9824 2916
rect 11060 2932 11112 2984
rect 11244 2907 11296 2916
rect 11244 2873 11253 2907
rect 11253 2873 11287 2907
rect 11287 2873 11296 2907
rect 11244 2864 11296 2873
rect 11428 2864 11480 2916
rect 12716 3000 12768 3052
rect 14188 3068 14240 3120
rect 12992 3000 13044 3052
rect 14372 3043 14424 3052
rect 14372 3009 14381 3043
rect 14381 3009 14415 3043
rect 14415 3009 14424 3043
rect 14372 3000 14424 3009
rect 14096 2932 14148 2984
rect 3248 2694 3300 2746
rect 3312 2694 3364 2746
rect 3376 2694 3428 2746
rect 3440 2694 3492 2746
rect 3504 2694 3556 2746
rect 7846 2694 7898 2746
rect 7910 2694 7962 2746
rect 7974 2694 8026 2746
rect 8038 2694 8090 2746
rect 8102 2694 8154 2746
rect 12443 2694 12495 2746
rect 12507 2694 12559 2746
rect 12571 2694 12623 2746
rect 12635 2694 12687 2746
rect 12699 2694 12751 2746
rect 9312 2592 9364 2644
rect 7196 2524 7248 2576
rect 11152 2592 11204 2644
rect 11244 2592 11296 2644
rect 3976 2388 4028 2440
rect 7748 2431 7800 2440
rect 7748 2397 7757 2431
rect 7757 2397 7791 2431
rect 7791 2397 7800 2431
rect 7748 2388 7800 2397
rect 9588 2499 9640 2508
rect 9588 2465 9597 2499
rect 9597 2465 9631 2499
rect 9631 2465 9640 2499
rect 9588 2456 9640 2465
rect 11796 2499 11848 2508
rect 11796 2465 11805 2499
rect 11805 2465 11839 2499
rect 11839 2465 11848 2499
rect 11796 2456 11848 2465
rect 9220 2431 9272 2440
rect 9220 2397 9229 2431
rect 9229 2397 9263 2431
rect 9263 2397 9272 2431
rect 9220 2388 9272 2397
rect 3884 2252 3936 2304
rect 8668 2320 8720 2372
rect 11152 2388 11204 2440
rect 9772 2320 9824 2372
rect 6920 2252 6972 2304
rect 8208 2252 8260 2304
rect 9036 2252 9088 2304
rect 9404 2252 9456 2304
rect 10324 2320 10376 2372
rect 12900 2456 12952 2508
rect 14096 2431 14148 2440
rect 14096 2397 14105 2431
rect 14105 2397 14139 2431
rect 14139 2397 14148 2431
rect 14096 2388 14148 2397
rect 12532 2320 12584 2372
rect 12900 2320 12952 2372
rect 5547 2150 5599 2202
rect 5611 2150 5663 2202
rect 5675 2150 5727 2202
rect 5739 2150 5791 2202
rect 5803 2150 5855 2202
rect 10144 2150 10196 2202
rect 10208 2150 10260 2202
rect 10272 2150 10324 2202
rect 10336 2150 10388 2202
rect 10400 2150 10452 2202
rect 14924 1071 14976 1080
rect 14924 1037 14933 1071
rect 14933 1037 14967 1071
rect 14967 1037 14976 1071
rect 14924 1028 14976 1037
<< metal2 >>
rect 2686 15200 2742 16000
rect 8022 15200 8078 16000
rect 13358 15200 13414 16000
rect 2700 13546 2728 15200
rect 8036 13818 8064 15200
rect 8036 13790 8248 13818
rect 3248 13628 3556 13648
rect 3248 13626 3254 13628
rect 3310 13626 3334 13628
rect 3390 13626 3414 13628
rect 3470 13626 3494 13628
rect 3550 13626 3556 13628
rect 3310 13574 3312 13626
rect 3492 13574 3494 13626
rect 3248 13572 3254 13574
rect 3310 13572 3334 13574
rect 3390 13572 3414 13574
rect 3470 13572 3494 13574
rect 3550 13572 3556 13574
rect 3248 13552 3556 13572
rect 7846 13628 8154 13648
rect 7846 13626 7852 13628
rect 7908 13626 7932 13628
rect 7988 13626 8012 13628
rect 8068 13626 8092 13628
rect 8148 13626 8154 13628
rect 7908 13574 7910 13626
rect 8090 13574 8092 13626
rect 7846 13572 7852 13574
rect 7908 13572 7932 13574
rect 7988 13572 8012 13574
rect 8068 13572 8092 13574
rect 8148 13572 8154 13574
rect 7846 13552 8154 13572
rect 2700 13530 2820 13546
rect 8220 13530 8248 13790
rect 12443 13628 12751 13648
rect 12443 13626 12449 13628
rect 12505 13626 12529 13628
rect 12585 13626 12609 13628
rect 12665 13626 12689 13628
rect 12745 13626 12751 13628
rect 12505 13574 12507 13626
rect 12687 13574 12689 13626
rect 12443 13572 12449 13574
rect 12505 13572 12529 13574
rect 12585 13572 12609 13574
rect 12665 13572 12689 13574
rect 12745 13572 12751 13574
rect 12443 13552 12751 13572
rect 13372 13530 13400 15200
rect 14922 15056 14978 15065
rect 14922 14991 14924 15000
rect 14976 14991 14978 15000
rect 14924 14962 14976 14968
rect 2700 13524 2832 13530
rect 2700 13518 2780 13524
rect 2780 13466 2832 13472
rect 7564 13524 7616 13530
rect 7564 13466 7616 13472
rect 8208 13524 8260 13530
rect 8208 13466 8260 13472
rect 13268 13524 13320 13530
rect 13268 13466 13320 13472
rect 13360 13524 13412 13530
rect 13360 13466 13412 13472
rect 5264 13388 5316 13394
rect 4344 13330 4396 13336
rect 5264 13330 5316 13336
rect 2780 13320 2832 13326
rect 2780 13262 2832 13268
rect 3976 13320 4028 13326
rect 3976 13262 4028 13268
rect 4160 13320 4212 13326
rect 4344 13272 4396 13278
rect 4528 13320 4580 13326
rect 4160 13262 4212 13268
rect 2504 13184 2556 13190
rect 2504 13126 2556 13132
rect 2516 12850 2544 13126
rect 2504 12844 2556 12850
rect 2504 12786 2556 12792
rect 2792 12306 2820 13262
rect 2872 13184 2924 13190
rect 2872 13126 2924 13132
rect 2884 12850 2912 13126
rect 2964 12980 3016 12986
rect 2964 12922 3016 12928
rect 2872 12844 2924 12850
rect 2872 12786 2924 12792
rect 2780 12300 2832 12306
rect 2780 12242 2832 12248
rect 1860 12164 1912 12170
rect 1860 12106 1912 12112
rect 2044 12164 2096 12170
rect 2044 12106 2096 12112
rect 1872 11150 1900 12106
rect 2056 11898 2084 12106
rect 2976 12102 3004 12922
rect 3248 12540 3556 12560
rect 3248 12538 3254 12540
rect 3310 12538 3334 12540
rect 3390 12538 3414 12540
rect 3470 12538 3494 12540
rect 3550 12538 3556 12540
rect 3310 12486 3312 12538
rect 3492 12486 3494 12538
rect 3248 12484 3254 12486
rect 3310 12484 3334 12486
rect 3390 12484 3414 12486
rect 3470 12484 3494 12486
rect 3550 12484 3556 12486
rect 3248 12464 3556 12484
rect 3988 12238 4016 13262
rect 4172 13190 4200 13262
rect 4160 13184 4212 13190
rect 4160 13126 4212 13132
rect 4356 12714 4384 13272
rect 4528 13262 4580 13268
rect 4344 12708 4396 12714
rect 4344 12650 4396 12656
rect 3976 12232 4028 12238
rect 3976 12174 4028 12180
rect 4068 12232 4120 12238
rect 4068 12174 4120 12180
rect 2964 12096 3016 12102
rect 2964 12038 3016 12044
rect 3608 12096 3660 12102
rect 3608 12038 3660 12044
rect 2044 11892 2096 11898
rect 2044 11834 2096 11840
rect 2976 11558 3004 12038
rect 2964 11552 3016 11558
rect 2964 11494 3016 11500
rect 1860 11144 1912 11150
rect 1860 11086 1912 11092
rect 1872 10674 1900 11086
rect 2976 11014 3004 11494
rect 3248 11452 3556 11472
rect 3248 11450 3254 11452
rect 3310 11450 3334 11452
rect 3390 11450 3414 11452
rect 3470 11450 3494 11452
rect 3550 11450 3556 11452
rect 3310 11398 3312 11450
rect 3492 11398 3494 11450
rect 3248 11396 3254 11398
rect 3310 11396 3334 11398
rect 3390 11396 3414 11398
rect 3470 11396 3494 11398
rect 3550 11396 3556 11398
rect 3248 11376 3556 11396
rect 3620 11354 3648 12038
rect 4080 11830 4108 12174
rect 4436 12096 4488 12102
rect 4158 12064 4214 12073
rect 4436 12038 4488 12044
rect 4158 11999 4214 12008
rect 4068 11824 4120 11830
rect 4068 11766 4120 11772
rect 4068 11552 4120 11558
rect 4068 11494 4120 11500
rect 3608 11348 3660 11354
rect 3608 11290 3660 11296
rect 4080 11286 4108 11494
rect 4068 11280 4120 11286
rect 4068 11222 4120 11228
rect 2964 11008 3016 11014
rect 2964 10950 3016 10956
rect 1860 10668 1912 10674
rect 1860 10610 1912 10616
rect 1400 10464 1452 10470
rect 1400 10406 1452 10412
rect 1412 9586 1440 10406
rect 2976 9994 3004 10950
rect 3884 10736 3936 10742
rect 3936 10696 4016 10724
rect 3884 10678 3936 10684
rect 3516 10668 3568 10674
rect 3516 10610 3568 10616
rect 3700 10668 3752 10674
rect 3700 10610 3752 10616
rect 3792 10668 3844 10674
rect 3792 10610 3844 10616
rect 3528 10554 3556 10610
rect 3148 10532 3200 10538
rect 3528 10526 3648 10554
rect 3148 10474 3200 10480
rect 3056 10464 3108 10470
rect 3056 10406 3108 10412
rect 3068 10033 3096 10406
rect 3160 10130 3188 10474
rect 3248 10364 3556 10384
rect 3248 10362 3254 10364
rect 3310 10362 3334 10364
rect 3390 10362 3414 10364
rect 3470 10362 3494 10364
rect 3550 10362 3556 10364
rect 3310 10310 3312 10362
rect 3492 10310 3494 10362
rect 3248 10308 3254 10310
rect 3310 10308 3334 10310
rect 3390 10308 3414 10310
rect 3470 10308 3494 10310
rect 3550 10308 3556 10310
rect 3248 10288 3556 10308
rect 3148 10124 3200 10130
rect 3148 10066 3200 10072
rect 3054 10024 3110 10033
rect 2964 9988 3016 9994
rect 3054 9959 3110 9968
rect 2964 9930 3016 9936
rect 2976 9897 3004 9930
rect 2962 9888 3018 9897
rect 2962 9823 3018 9832
rect 1400 9580 1452 9586
rect 1400 9522 1452 9528
rect 2780 9512 2832 9518
rect 2780 9454 2832 9460
rect 2792 9178 2820 9454
rect 2872 9444 2924 9450
rect 2872 9386 2924 9392
rect 2780 9172 2832 9178
rect 2780 9114 2832 9120
rect 2884 9110 2912 9386
rect 3068 9382 3096 9959
rect 3056 9376 3108 9382
rect 3056 9318 3108 9324
rect 2872 9104 2924 9110
rect 2872 9046 2924 9052
rect 3068 8922 3096 9318
rect 3160 9042 3188 10066
rect 3516 9920 3568 9926
rect 3514 9888 3516 9897
rect 3568 9888 3570 9897
rect 3514 9823 3570 9832
rect 3248 9276 3556 9296
rect 3248 9274 3254 9276
rect 3310 9274 3334 9276
rect 3390 9274 3414 9276
rect 3470 9274 3494 9276
rect 3550 9274 3556 9276
rect 3310 9222 3312 9274
rect 3492 9222 3494 9274
rect 3248 9220 3254 9222
rect 3310 9220 3334 9222
rect 3390 9220 3414 9222
rect 3470 9220 3494 9222
rect 3550 9220 3556 9222
rect 3248 9200 3556 9220
rect 3620 9178 3648 10526
rect 3712 10266 3740 10610
rect 3700 10260 3752 10266
rect 3700 10202 3752 10208
rect 3804 10062 3832 10610
rect 3884 10464 3936 10470
rect 3884 10406 3936 10412
rect 3896 10062 3924 10406
rect 3988 10266 4016 10696
rect 3976 10260 4028 10266
rect 3976 10202 4028 10208
rect 4172 10198 4200 11999
rect 4448 11762 4476 12038
rect 4436 11756 4488 11762
rect 4436 11698 4488 11704
rect 4252 11688 4304 11694
rect 4252 11630 4304 11636
rect 4540 11642 4568 13262
rect 4712 13184 4764 13190
rect 4712 13126 4764 13132
rect 4724 12986 4752 13126
rect 4712 12980 4764 12986
rect 4712 12922 4764 12928
rect 4620 12844 4672 12850
rect 4620 12786 4672 12792
rect 4632 12238 4660 12786
rect 4896 12708 4948 12714
rect 4896 12650 4948 12656
rect 4804 12300 4856 12306
rect 4804 12242 4856 12248
rect 4620 12232 4672 12238
rect 4620 12174 4672 12180
rect 4816 11898 4844 12242
rect 4908 12170 4936 12650
rect 5080 12640 5132 12646
rect 5080 12582 5132 12588
rect 4988 12232 5040 12238
rect 4988 12174 5040 12180
rect 4896 12164 4948 12170
rect 4896 12106 4948 12112
rect 4804 11892 4856 11898
rect 4804 11834 4856 11840
rect 4908 11762 4936 12106
rect 4712 11756 4764 11762
rect 4712 11698 4764 11704
rect 4896 11756 4948 11762
rect 4896 11698 4948 11704
rect 4264 11150 4292 11630
rect 4540 11626 4660 11642
rect 4540 11620 4672 11626
rect 4540 11614 4620 11620
rect 4620 11562 4672 11568
rect 4344 11552 4396 11558
rect 4344 11494 4396 11500
rect 4528 11552 4580 11558
rect 4528 11494 4580 11500
rect 4252 11144 4304 11150
rect 4252 11086 4304 11092
rect 4264 10810 4292 11086
rect 4356 11082 4384 11494
rect 4540 11218 4568 11494
rect 4632 11354 4660 11562
rect 4620 11348 4672 11354
rect 4620 11290 4672 11296
rect 4528 11212 4580 11218
rect 4528 11154 4580 11160
rect 4344 11076 4396 11082
rect 4724 11054 4752 11698
rect 5000 11054 5028 12174
rect 5092 11762 5120 12582
rect 5276 12238 5304 13330
rect 5448 13184 5500 13190
rect 5448 13126 5500 13132
rect 5908 13184 5960 13190
rect 5908 13126 5960 13132
rect 5460 12986 5488 13126
rect 5547 13084 5855 13104
rect 5547 13082 5553 13084
rect 5609 13082 5633 13084
rect 5689 13082 5713 13084
rect 5769 13082 5793 13084
rect 5849 13082 5855 13084
rect 5609 13030 5611 13082
rect 5791 13030 5793 13082
rect 5547 13028 5553 13030
rect 5609 13028 5633 13030
rect 5689 13028 5713 13030
rect 5769 13028 5793 13030
rect 5849 13028 5855 13030
rect 5547 13008 5855 13028
rect 5448 12980 5500 12986
rect 5448 12922 5500 12928
rect 5920 12782 5948 13126
rect 6920 12844 6972 12850
rect 6920 12786 6972 12792
rect 7288 12844 7340 12850
rect 7288 12786 7340 12792
rect 5908 12776 5960 12782
rect 5908 12718 5960 12724
rect 6000 12776 6052 12782
rect 6000 12718 6052 12724
rect 5356 12300 5408 12306
rect 5356 12242 5408 12248
rect 5264 12232 5316 12238
rect 5264 12174 5316 12180
rect 5368 11830 5396 12242
rect 5920 12238 5948 12718
rect 5908 12232 5960 12238
rect 5908 12174 5960 12180
rect 5448 12096 5500 12102
rect 5448 12038 5500 12044
rect 5908 12096 5960 12102
rect 5908 12038 5960 12044
rect 5460 11898 5488 12038
rect 5547 11996 5855 12016
rect 5547 11994 5553 11996
rect 5609 11994 5633 11996
rect 5689 11994 5713 11996
rect 5769 11994 5793 11996
rect 5849 11994 5855 11996
rect 5609 11942 5611 11994
rect 5791 11942 5793 11994
rect 5547 11940 5553 11942
rect 5609 11940 5633 11942
rect 5689 11940 5713 11942
rect 5769 11940 5793 11942
rect 5849 11940 5855 11942
rect 5547 11920 5855 11940
rect 5448 11892 5500 11898
rect 5448 11834 5500 11840
rect 5356 11824 5408 11830
rect 5356 11766 5408 11772
rect 5080 11756 5132 11762
rect 5080 11698 5132 11704
rect 5920 11694 5948 12038
rect 6012 11694 6040 12718
rect 6092 12368 6144 12374
rect 6092 12310 6144 12316
rect 5356 11688 5408 11694
rect 5356 11630 5408 11636
rect 5908 11688 5960 11694
rect 5908 11630 5960 11636
rect 6000 11688 6052 11694
rect 6000 11630 6052 11636
rect 5264 11212 5316 11218
rect 5264 11154 5316 11160
rect 4344 11018 4396 11024
rect 4632 11026 4752 11054
rect 4908 11026 5028 11054
rect 4632 10810 4660 11026
rect 4252 10804 4304 10810
rect 4252 10746 4304 10752
rect 4620 10804 4672 10810
rect 4620 10746 4672 10752
rect 4528 10736 4580 10742
rect 4528 10678 4580 10684
rect 4436 10464 4488 10470
rect 4436 10406 4488 10412
rect 4160 10192 4212 10198
rect 4160 10134 4212 10140
rect 3792 10056 3844 10062
rect 3792 9998 3844 10004
rect 3884 10056 3936 10062
rect 3884 9998 3936 10004
rect 4344 10056 4396 10062
rect 4344 9998 4396 10004
rect 3700 9920 3752 9926
rect 3700 9862 3752 9868
rect 4252 9920 4304 9926
rect 4252 9862 4304 9868
rect 3608 9172 3660 9178
rect 3608 9114 3660 9120
rect 3148 9036 3200 9042
rect 3148 8978 3200 8984
rect 3240 8968 3292 8974
rect 3068 8916 3240 8922
rect 3068 8910 3292 8916
rect 3068 8894 3280 8910
rect 3712 8906 3740 9862
rect 3884 9716 3936 9722
rect 3884 9658 3936 9664
rect 3896 9110 3924 9658
rect 4264 9586 4292 9862
rect 4356 9722 4384 9998
rect 4344 9716 4396 9722
rect 4344 9658 4396 9664
rect 4448 9586 4476 10406
rect 4540 10146 4568 10678
rect 4908 10606 4936 11026
rect 5080 11008 5132 11014
rect 5080 10950 5132 10956
rect 5092 10810 5120 10950
rect 5080 10804 5132 10810
rect 5080 10746 5132 10752
rect 5276 10742 5304 11154
rect 4988 10736 5040 10742
rect 5264 10736 5316 10742
rect 5040 10684 5120 10690
rect 4988 10678 5120 10684
rect 5264 10678 5316 10684
rect 5000 10662 5120 10678
rect 4896 10600 4948 10606
rect 4896 10542 4948 10548
rect 4988 10532 5040 10538
rect 4988 10474 5040 10480
rect 4540 10118 4844 10146
rect 4528 10056 4580 10062
rect 4526 10024 4528 10033
rect 4620 10056 4672 10062
rect 4580 10024 4582 10033
rect 4620 9998 4672 10004
rect 4526 9959 4582 9968
rect 4528 9716 4580 9722
rect 4528 9658 4580 9664
rect 4252 9580 4304 9586
rect 4252 9522 4304 9528
rect 4436 9580 4488 9586
rect 4436 9522 4488 9528
rect 3976 9512 4028 9518
rect 3976 9454 4028 9460
rect 3884 9104 3936 9110
rect 3884 9046 3936 9052
rect 3700 8900 3752 8906
rect 3700 8842 3752 8848
rect 3896 8566 3924 9046
rect 3988 8974 4016 9454
rect 4068 9376 4120 9382
rect 4068 9318 4120 9324
rect 4252 9376 4304 9382
rect 4252 9318 4304 9324
rect 4080 8974 4108 9318
rect 3976 8968 4028 8974
rect 3976 8910 4028 8916
rect 4068 8968 4120 8974
rect 4068 8910 4120 8916
rect 3988 8634 4016 8910
rect 4080 8634 4108 8910
rect 4264 8906 4292 9318
rect 4540 8906 4568 9658
rect 4632 9586 4660 9998
rect 4816 9926 4844 10118
rect 5000 10062 5028 10474
rect 5092 10062 5120 10662
rect 5172 10668 5224 10674
rect 5172 10610 5224 10616
rect 5184 10198 5212 10610
rect 5368 10198 5396 11630
rect 6012 11370 6040 11630
rect 5828 11342 6040 11370
rect 5828 11218 5856 11342
rect 5816 11212 5868 11218
rect 5816 11154 5868 11160
rect 5908 11144 5960 11150
rect 5538 11112 5594 11121
rect 5908 11086 5960 11092
rect 5538 11054 5540 11056
rect 5460 11026 5540 11054
rect 5460 10810 5488 11026
rect 5592 11047 5594 11056
rect 5540 11018 5592 11024
rect 5547 10908 5855 10928
rect 5547 10906 5553 10908
rect 5609 10906 5633 10908
rect 5689 10906 5713 10908
rect 5769 10906 5793 10908
rect 5849 10906 5855 10908
rect 5609 10854 5611 10906
rect 5791 10854 5793 10906
rect 5547 10852 5553 10854
rect 5609 10852 5633 10854
rect 5689 10852 5713 10854
rect 5769 10852 5793 10854
rect 5849 10852 5855 10854
rect 5547 10832 5855 10852
rect 5920 10810 5948 11086
rect 6104 11054 6132 12310
rect 6932 12238 6960 12786
rect 6920 12232 6972 12238
rect 6920 12174 6972 12180
rect 6460 12164 6512 12170
rect 6460 12106 6512 12112
rect 6472 11354 6500 12106
rect 6932 11830 6960 12174
rect 6920 11824 6972 11830
rect 6920 11766 6972 11772
rect 6460 11348 6512 11354
rect 6460 11290 6512 11296
rect 6184 11280 6236 11286
rect 6184 11222 6236 11228
rect 6012 11026 6132 11054
rect 5448 10804 5500 10810
rect 5448 10746 5500 10752
rect 5908 10804 5960 10810
rect 5908 10746 5960 10752
rect 6012 10690 6040 11026
rect 6196 10742 6224 11222
rect 6276 11076 6328 11082
rect 6276 11018 6328 11024
rect 6288 10810 6316 11018
rect 6276 10804 6328 10810
rect 6276 10746 6328 10752
rect 5828 10674 6040 10690
rect 6184 10736 6236 10742
rect 6184 10678 6236 10684
rect 5632 10668 5684 10674
rect 5632 10610 5684 10616
rect 5816 10668 6040 10674
rect 5868 10662 6040 10668
rect 5816 10610 5868 10616
rect 5448 10464 5500 10470
rect 5448 10406 5500 10412
rect 5172 10192 5224 10198
rect 5172 10134 5224 10140
rect 5356 10192 5408 10198
rect 5356 10134 5408 10140
rect 5460 10062 5488 10406
rect 5644 10198 5672 10610
rect 6184 10464 6236 10470
rect 6184 10406 6236 10412
rect 5632 10192 5684 10198
rect 5632 10134 5684 10140
rect 5908 10192 5960 10198
rect 5908 10134 5960 10140
rect 4988 10056 5040 10062
rect 4988 9998 5040 10004
rect 5080 10056 5132 10062
rect 5080 9998 5132 10004
rect 5356 10056 5408 10062
rect 5356 9998 5408 10004
rect 5448 10056 5500 10062
rect 5448 9998 5500 10004
rect 4804 9920 4856 9926
rect 4804 9862 4856 9868
rect 4816 9586 4844 9862
rect 5368 9722 5396 9998
rect 5356 9716 5408 9722
rect 5356 9658 5408 9664
rect 5460 9654 5488 9998
rect 5547 9820 5855 9840
rect 5547 9818 5553 9820
rect 5609 9818 5633 9820
rect 5689 9818 5713 9820
rect 5769 9818 5793 9820
rect 5849 9818 5855 9820
rect 5609 9766 5611 9818
rect 5791 9766 5793 9818
rect 5547 9764 5553 9766
rect 5609 9764 5633 9766
rect 5689 9764 5713 9766
rect 5769 9764 5793 9766
rect 5849 9764 5855 9766
rect 5547 9744 5855 9764
rect 5448 9648 5500 9654
rect 5448 9590 5500 9596
rect 4620 9580 4672 9586
rect 4620 9522 4672 9528
rect 4804 9580 4856 9586
rect 4804 9522 4856 9528
rect 5920 9518 5948 10134
rect 6196 10130 6224 10406
rect 6184 10124 6236 10130
rect 6184 10066 6236 10072
rect 6368 9920 6420 9926
rect 6368 9862 6420 9868
rect 6380 9586 6408 9862
rect 6472 9722 6500 11290
rect 6828 11280 6880 11286
rect 6828 11222 6880 11228
rect 6644 11076 6696 11082
rect 6840 11054 6868 11222
rect 6932 11218 6960 11766
rect 6920 11212 6972 11218
rect 6920 11154 6972 11160
rect 7300 11121 7328 12786
rect 7576 12442 7604 13466
rect 8484 13456 8536 13462
rect 8484 13398 8536 13404
rect 7656 13320 7708 13326
rect 7656 13262 7708 13268
rect 8208 13320 8260 13326
rect 8208 13262 8260 13268
rect 7668 12442 7696 13262
rect 7846 12540 8154 12560
rect 7846 12538 7852 12540
rect 7908 12538 7932 12540
rect 7988 12538 8012 12540
rect 8068 12538 8092 12540
rect 8148 12538 8154 12540
rect 7908 12486 7910 12538
rect 8090 12486 8092 12538
rect 7846 12484 7852 12486
rect 7908 12484 7932 12486
rect 7988 12484 8012 12486
rect 8068 12484 8092 12486
rect 8148 12484 8154 12486
rect 7846 12464 8154 12484
rect 8220 12442 8248 13262
rect 8300 13184 8352 13190
rect 8300 13126 8352 13132
rect 7564 12436 7616 12442
rect 7564 12378 7616 12384
rect 7656 12436 7708 12442
rect 7656 12378 7708 12384
rect 8208 12436 8260 12442
rect 8208 12378 8260 12384
rect 7576 12238 7604 12378
rect 8312 12238 8340 13126
rect 8392 12640 8444 12646
rect 8392 12582 8444 12588
rect 8404 12306 8432 12582
rect 8392 12300 8444 12306
rect 8392 12242 8444 12248
rect 7564 12232 7616 12238
rect 7564 12174 7616 12180
rect 8300 12232 8352 12238
rect 8300 12174 8352 12180
rect 8496 11898 8524 13398
rect 8852 13388 8904 13394
rect 8852 13330 8904 13336
rect 12992 13388 13044 13394
rect 12992 13330 13044 13336
rect 8668 13184 8720 13190
rect 8668 13126 8720 13132
rect 8680 12918 8708 13126
rect 8668 12912 8720 12918
rect 8668 12854 8720 12860
rect 8864 12782 8892 13330
rect 11336 13320 11388 13326
rect 11336 13262 11388 13268
rect 12440 13320 12492 13326
rect 12440 13262 12492 13268
rect 10876 13252 10928 13258
rect 10876 13194 10928 13200
rect 10784 13184 10836 13190
rect 10784 13126 10836 13132
rect 10144 13084 10452 13104
rect 10144 13082 10150 13084
rect 10206 13082 10230 13084
rect 10286 13082 10310 13084
rect 10366 13082 10390 13084
rect 10446 13082 10452 13084
rect 10206 13030 10208 13082
rect 10388 13030 10390 13082
rect 10144 13028 10150 13030
rect 10206 13028 10230 13030
rect 10286 13028 10310 13030
rect 10366 13028 10390 13030
rect 10446 13028 10452 13030
rect 10144 13008 10452 13028
rect 9312 12912 9364 12918
rect 9312 12854 9364 12860
rect 8852 12776 8904 12782
rect 8852 12718 8904 12724
rect 8944 12368 8996 12374
rect 8944 12310 8996 12316
rect 8484 11892 8536 11898
rect 8484 11834 8536 11840
rect 8760 11892 8812 11898
rect 8760 11834 8812 11840
rect 7838 11792 7894 11801
rect 7838 11727 7894 11736
rect 8484 11756 8536 11762
rect 7852 11694 7880 11727
rect 8484 11698 8536 11704
rect 7840 11688 7892 11694
rect 7840 11630 7892 11636
rect 8496 11540 8524 11698
rect 8772 11558 8800 11834
rect 8956 11762 8984 12310
rect 9324 12102 9352 12854
rect 9496 12640 9548 12646
rect 9496 12582 9548 12588
rect 9508 12238 9536 12582
rect 9496 12232 9548 12238
rect 9496 12174 9548 12180
rect 9312 12096 9364 12102
rect 9312 12038 9364 12044
rect 9218 11792 9274 11801
rect 8944 11756 8996 11762
rect 8944 11698 8996 11704
rect 9036 11756 9088 11762
rect 9218 11727 9220 11736
rect 9036 11698 9088 11704
rect 9272 11727 9274 11736
rect 9220 11698 9272 11704
rect 8760 11552 8812 11558
rect 8496 11512 8760 11540
rect 7846 11452 8154 11472
rect 7846 11450 7852 11452
rect 7908 11450 7932 11452
rect 7988 11450 8012 11452
rect 8068 11450 8092 11452
rect 8148 11450 8154 11452
rect 7908 11398 7910 11450
rect 8090 11398 8092 11450
rect 7846 11396 7852 11398
rect 7908 11396 7932 11398
rect 7988 11396 8012 11398
rect 8068 11396 8092 11398
rect 8148 11396 8154 11398
rect 7846 11376 8154 11396
rect 8300 11212 8352 11218
rect 8300 11154 8352 11160
rect 7286 11112 7342 11121
rect 8206 11112 8262 11121
rect 6840 11026 6960 11054
rect 7286 11047 7342 11056
rect 7656 11076 7708 11082
rect 6644 11018 6696 11024
rect 6552 11008 6604 11014
rect 6552 10950 6604 10956
rect 6564 10674 6592 10950
rect 6552 10668 6604 10674
rect 6552 10610 6604 10616
rect 6656 10554 6684 11018
rect 6932 10674 6960 11026
rect 8206 11047 8262 11056
rect 7656 11018 7708 11024
rect 7668 10810 7696 11018
rect 7656 10804 7708 10810
rect 7656 10746 7708 10752
rect 6920 10668 6972 10674
rect 6920 10610 6972 10616
rect 6656 10526 6960 10554
rect 6460 9716 6512 9722
rect 6460 9658 6512 9664
rect 6368 9580 6420 9586
rect 6368 9522 6420 9528
rect 6828 9580 6880 9586
rect 6828 9522 6880 9528
rect 5908 9512 5960 9518
rect 5908 9454 5960 9460
rect 4988 9444 5040 9450
rect 4988 9386 5040 9392
rect 4620 8968 4672 8974
rect 4620 8910 4672 8916
rect 4252 8900 4304 8906
rect 4252 8842 4304 8848
rect 4528 8900 4580 8906
rect 4528 8842 4580 8848
rect 4344 8832 4396 8838
rect 4344 8774 4396 8780
rect 3976 8628 4028 8634
rect 3976 8570 4028 8576
rect 4068 8628 4120 8634
rect 4068 8570 4120 8576
rect 4356 8566 4384 8774
rect 3884 8560 3936 8566
rect 3884 8502 3936 8508
rect 4344 8560 4396 8566
rect 4344 8502 4396 8508
rect 3248 8188 3556 8208
rect 3248 8186 3254 8188
rect 3310 8186 3334 8188
rect 3390 8186 3414 8188
rect 3470 8186 3494 8188
rect 3550 8186 3556 8188
rect 3310 8134 3312 8186
rect 3492 8134 3494 8186
rect 3248 8132 3254 8134
rect 3310 8132 3334 8134
rect 3390 8132 3414 8134
rect 3470 8132 3494 8134
rect 3550 8132 3556 8134
rect 3248 8112 3556 8132
rect 2504 7948 2556 7954
rect 2504 7890 2556 7896
rect 1676 7880 1728 7886
rect 1676 7822 1728 7828
rect 1688 6390 1716 7822
rect 1952 7744 2004 7750
rect 1952 7686 2004 7692
rect 2320 7744 2372 7750
rect 2320 7686 2372 7692
rect 1964 7410 1992 7686
rect 2332 7410 2360 7686
rect 1952 7404 2004 7410
rect 1952 7346 2004 7352
rect 2320 7404 2372 7410
rect 2320 7346 2372 7352
rect 2516 7002 2544 7890
rect 2688 7880 2740 7886
rect 2688 7822 2740 7828
rect 2964 7880 3016 7886
rect 2964 7822 3016 7828
rect 2504 6996 2556 7002
rect 2504 6938 2556 6944
rect 2044 6792 2096 6798
rect 2044 6734 2096 6740
rect 1676 6384 1728 6390
rect 1676 6326 1728 6332
rect 1688 5778 1716 6326
rect 2056 5914 2084 6734
rect 2700 6730 2728 7822
rect 2688 6724 2740 6730
rect 2688 6666 2740 6672
rect 2320 6656 2372 6662
rect 2320 6598 2372 6604
rect 2332 6254 2360 6598
rect 2412 6384 2464 6390
rect 2412 6326 2464 6332
rect 2320 6248 2372 6254
rect 2320 6190 2372 6196
rect 2044 5908 2096 5914
rect 2044 5850 2096 5856
rect 1676 5772 1728 5778
rect 1676 5714 1728 5720
rect 1688 5234 1716 5714
rect 2424 5642 2452 6326
rect 2700 5846 2728 6666
rect 2976 6254 3004 7822
rect 3896 7750 3924 8502
rect 4632 8430 4660 8910
rect 4896 8900 4948 8906
rect 4896 8842 4948 8848
rect 4908 8634 4936 8842
rect 4896 8628 4948 8634
rect 4896 8570 4948 8576
rect 5000 8498 5028 9386
rect 6840 9330 6868 9522
rect 6932 9450 6960 10526
rect 7846 10364 8154 10384
rect 7846 10362 7852 10364
rect 7908 10362 7932 10364
rect 7988 10362 8012 10364
rect 8068 10362 8092 10364
rect 8148 10362 8154 10364
rect 7908 10310 7910 10362
rect 8090 10310 8092 10362
rect 7846 10308 7852 10310
rect 7908 10308 7932 10310
rect 7988 10308 8012 10310
rect 8068 10308 8092 10310
rect 8148 10308 8154 10310
rect 7846 10288 8154 10308
rect 7748 10056 7800 10062
rect 7748 9998 7800 10004
rect 7196 9716 7248 9722
rect 7196 9658 7248 9664
rect 7104 9648 7156 9654
rect 7104 9590 7156 9596
rect 6920 9444 6972 9450
rect 6920 9386 6972 9392
rect 7116 9330 7144 9590
rect 6840 9302 7144 9330
rect 6828 9104 6880 9110
rect 6828 9046 6880 9052
rect 5356 8900 5408 8906
rect 5356 8842 5408 8848
rect 4988 8492 5040 8498
rect 4988 8434 5040 8440
rect 4620 8424 4672 8430
rect 4620 8366 4672 8372
rect 5368 8294 5396 8842
rect 6460 8832 6512 8838
rect 6460 8774 6512 8780
rect 5547 8732 5855 8752
rect 5547 8730 5553 8732
rect 5609 8730 5633 8732
rect 5689 8730 5713 8732
rect 5769 8730 5793 8732
rect 5849 8730 5855 8732
rect 5609 8678 5611 8730
rect 5791 8678 5793 8730
rect 5547 8676 5553 8678
rect 5609 8676 5633 8678
rect 5689 8676 5713 8678
rect 5769 8676 5793 8678
rect 5849 8676 5855 8678
rect 5547 8656 5855 8676
rect 6472 8566 6500 8774
rect 6840 8566 6868 9046
rect 7208 8634 7236 9658
rect 7760 9654 7788 9998
rect 7932 9920 7984 9926
rect 7932 9862 7984 9868
rect 7748 9648 7800 9654
rect 7748 9590 7800 9596
rect 7944 9518 7972 9862
rect 8116 9580 8168 9586
rect 8116 9522 8168 9528
rect 7656 9512 7708 9518
rect 7656 9454 7708 9460
rect 7748 9512 7800 9518
rect 7748 9454 7800 9460
rect 7932 9512 7984 9518
rect 7932 9454 7984 9460
rect 8128 9466 8156 9522
rect 8220 9466 8248 11047
rect 8312 10810 8340 11154
rect 8300 10804 8352 10810
rect 8300 10746 8352 10752
rect 8392 10736 8444 10742
rect 8392 10678 8444 10684
rect 7668 9178 7696 9454
rect 7656 9172 7708 9178
rect 7656 9114 7708 9120
rect 7760 9042 7788 9454
rect 8128 9438 8340 9466
rect 8404 9450 8432 10678
rect 8496 10146 8524 11512
rect 8760 11494 8812 11500
rect 8852 11348 8904 11354
rect 8852 11290 8904 11296
rect 8576 11280 8628 11286
rect 8576 11222 8628 11228
rect 8588 11014 8616 11222
rect 8668 11212 8720 11218
rect 8668 11154 8720 11160
rect 8576 11008 8628 11014
rect 8576 10950 8628 10956
rect 8576 10668 8628 10674
rect 8576 10610 8628 10616
rect 8588 10266 8616 10610
rect 8680 10606 8708 11154
rect 8668 10600 8720 10606
rect 8668 10542 8720 10548
rect 8668 10464 8720 10470
rect 8668 10406 8720 10412
rect 8576 10260 8628 10266
rect 8576 10202 8628 10208
rect 8496 10118 8616 10146
rect 8484 10056 8536 10062
rect 8588 10033 8616 10118
rect 8680 10062 8708 10406
rect 8668 10056 8720 10062
rect 8484 9998 8536 10004
rect 8574 10024 8630 10033
rect 7846 9276 8154 9296
rect 7846 9274 7852 9276
rect 7908 9274 7932 9276
rect 7988 9274 8012 9276
rect 8068 9274 8092 9276
rect 8148 9274 8154 9276
rect 7908 9222 7910 9274
rect 8090 9222 8092 9274
rect 7846 9220 7852 9222
rect 7908 9220 7932 9222
rect 7988 9220 8012 9222
rect 8068 9220 8092 9222
rect 8148 9220 8154 9222
rect 7846 9200 8154 9220
rect 8312 9110 8340 9438
rect 8392 9444 8444 9450
rect 8392 9386 8444 9392
rect 8300 9104 8352 9110
rect 8300 9046 8352 9052
rect 7748 9036 7800 9042
rect 7748 8978 7800 8984
rect 8312 8974 8340 9046
rect 7380 8968 7432 8974
rect 7380 8910 7432 8916
rect 8208 8968 8260 8974
rect 8208 8910 8260 8916
rect 8300 8968 8352 8974
rect 8300 8910 8352 8916
rect 7196 8628 7248 8634
rect 7196 8570 7248 8576
rect 6460 8560 6512 8566
rect 6460 8502 6512 8508
rect 6828 8560 6880 8566
rect 6828 8502 6880 8508
rect 5448 8424 5500 8430
rect 5448 8366 5500 8372
rect 5356 8288 5408 8294
rect 5356 8230 5408 8236
rect 5368 7750 5396 8230
rect 5460 7954 5488 8366
rect 5816 8288 5868 8294
rect 5816 8230 5868 8236
rect 5828 7954 5856 8230
rect 5448 7948 5500 7954
rect 5448 7890 5500 7896
rect 5816 7948 5868 7954
rect 5816 7890 5868 7896
rect 6736 7812 6788 7818
rect 6736 7754 6788 7760
rect 3332 7744 3384 7750
rect 3332 7686 3384 7692
rect 3884 7744 3936 7750
rect 3884 7686 3936 7692
rect 5356 7744 5408 7750
rect 5356 7686 5408 7692
rect 3344 7478 3372 7686
rect 5547 7644 5855 7664
rect 5547 7642 5553 7644
rect 5609 7642 5633 7644
rect 5689 7642 5713 7644
rect 5769 7642 5793 7644
rect 5849 7642 5855 7644
rect 5609 7590 5611 7642
rect 5791 7590 5793 7642
rect 5547 7588 5553 7590
rect 5609 7588 5633 7590
rect 5689 7588 5713 7590
rect 5769 7588 5793 7590
rect 5849 7588 5855 7590
rect 5547 7568 5855 7588
rect 3332 7472 3384 7478
rect 3332 7414 3384 7420
rect 4160 7404 4212 7410
rect 4160 7346 4212 7352
rect 4620 7404 4672 7410
rect 4620 7346 4672 7352
rect 3248 7100 3556 7120
rect 3248 7098 3254 7100
rect 3310 7098 3334 7100
rect 3390 7098 3414 7100
rect 3470 7098 3494 7100
rect 3550 7098 3556 7100
rect 3310 7046 3312 7098
rect 3492 7046 3494 7098
rect 3248 7044 3254 7046
rect 3310 7044 3334 7046
rect 3390 7044 3414 7046
rect 3470 7044 3494 7046
rect 3550 7044 3556 7046
rect 3248 7024 3556 7044
rect 3700 6996 3752 7002
rect 3700 6938 3752 6944
rect 3056 6860 3108 6866
rect 3056 6802 3108 6808
rect 3608 6860 3660 6866
rect 3608 6802 3660 6808
rect 3068 6390 3096 6802
rect 3148 6724 3200 6730
rect 3148 6666 3200 6672
rect 3160 6458 3188 6666
rect 3240 6656 3292 6662
rect 3240 6598 3292 6604
rect 3148 6452 3200 6458
rect 3148 6394 3200 6400
rect 3056 6384 3108 6390
rect 3056 6326 3108 6332
rect 3252 6322 3280 6598
rect 3620 6458 3648 6802
rect 3712 6662 3740 6938
rect 4172 6934 4200 7346
rect 4632 7290 4660 7346
rect 4632 7274 4752 7290
rect 4632 7268 4764 7274
rect 4632 7262 4712 7268
rect 4436 7200 4488 7206
rect 4436 7142 4488 7148
rect 4528 7200 4580 7206
rect 4528 7142 4580 7148
rect 4160 6928 4212 6934
rect 4160 6870 4212 6876
rect 4172 6798 4200 6870
rect 3884 6792 3936 6798
rect 3804 6740 3884 6746
rect 3804 6734 3936 6740
rect 4160 6792 4212 6798
rect 4160 6734 4212 6740
rect 3804 6718 3924 6734
rect 3700 6656 3752 6662
rect 3700 6598 3752 6604
rect 3608 6452 3660 6458
rect 3608 6394 3660 6400
rect 3804 6338 3832 6718
rect 4448 6712 4476 7142
rect 4540 6866 4568 7142
rect 4528 6860 4580 6866
rect 4528 6802 4580 6808
rect 4632 6798 4660 7262
rect 4712 7210 4764 7216
rect 6748 7206 6776 7754
rect 6840 7342 6868 8502
rect 7392 8498 7420 8910
rect 7748 8832 7800 8838
rect 7748 8774 7800 8780
rect 7760 8634 7788 8774
rect 7748 8628 7800 8634
rect 7748 8570 7800 8576
rect 7380 8492 7432 8498
rect 7380 8434 7432 8440
rect 7748 8492 7800 8498
rect 7748 8434 7800 8440
rect 7104 7948 7156 7954
rect 7104 7890 7156 7896
rect 7116 7410 7144 7890
rect 7392 7886 7420 8434
rect 7472 8424 7524 8430
rect 7472 8366 7524 8372
rect 7380 7880 7432 7886
rect 7380 7822 7432 7828
rect 7392 7478 7420 7822
rect 7484 7546 7512 8366
rect 7760 7886 7788 8434
rect 8220 8362 8248 8910
rect 8496 8498 8524 9998
rect 8668 9998 8720 10004
rect 8864 9994 8892 11290
rect 8956 11218 8984 11698
rect 9048 11257 9076 11698
rect 9220 11620 9272 11626
rect 9220 11562 9272 11568
rect 9034 11248 9090 11257
rect 8944 11212 8996 11218
rect 9034 11183 9090 11192
rect 8944 11154 8996 11160
rect 9034 11112 9090 11121
rect 9232 11082 9260 11562
rect 9324 11286 9352 12038
rect 9404 11688 9456 11694
rect 9404 11630 9456 11636
rect 9416 11354 9444 11630
rect 9404 11348 9456 11354
rect 9404 11290 9456 11296
rect 9312 11280 9364 11286
rect 9312 11222 9364 11228
rect 9034 11047 9090 11056
rect 9220 11076 9272 11082
rect 8944 11008 8996 11014
rect 8944 10950 8996 10956
rect 8956 10674 8984 10950
rect 8944 10668 8996 10674
rect 8944 10610 8996 10616
rect 8574 9959 8630 9968
rect 8852 9988 8904 9994
rect 8588 9586 8616 9959
rect 8852 9930 8904 9936
rect 8576 9580 8628 9586
rect 8576 9522 8628 9528
rect 8944 9580 8996 9586
rect 9048 9568 9076 11047
rect 9220 11018 9272 11024
rect 9324 10470 9352 11222
rect 9508 10674 9536 12174
rect 10144 11996 10452 12016
rect 10144 11994 10150 11996
rect 10206 11994 10230 11996
rect 10286 11994 10310 11996
rect 10366 11994 10390 11996
rect 10446 11994 10452 11996
rect 10206 11942 10208 11994
rect 10388 11942 10390 11994
rect 10144 11940 10150 11942
rect 10206 11940 10230 11942
rect 10286 11940 10310 11942
rect 10366 11940 10390 11942
rect 10446 11940 10452 11942
rect 10144 11920 10452 11940
rect 9956 11756 10008 11762
rect 9956 11698 10008 11704
rect 10048 11756 10100 11762
rect 10048 11698 10100 11704
rect 9680 11552 9732 11558
rect 9680 11494 9732 11500
rect 9692 11354 9720 11494
rect 9680 11348 9732 11354
rect 9680 11290 9732 11296
rect 9864 11212 9916 11218
rect 9864 11154 9916 11160
rect 9772 11008 9824 11014
rect 9772 10950 9824 10956
rect 9784 10810 9812 10950
rect 9772 10804 9824 10810
rect 9772 10746 9824 10752
rect 9496 10668 9548 10674
rect 9496 10610 9548 10616
rect 9312 10464 9364 10470
rect 9312 10406 9364 10412
rect 9324 10266 9352 10406
rect 9312 10260 9364 10266
rect 9312 10202 9364 10208
rect 8996 9540 9076 9568
rect 8944 9522 8996 9528
rect 8588 9110 8616 9522
rect 8668 9512 8720 9518
rect 8668 9454 8720 9460
rect 8680 9178 8708 9454
rect 8668 9172 8720 9178
rect 8668 9114 8720 9120
rect 8576 9104 8628 9110
rect 8576 9046 8628 9052
rect 8680 8566 8708 9114
rect 9508 9042 9536 10610
rect 9876 10282 9904 11154
rect 9968 11150 9996 11698
rect 10060 11234 10088 11698
rect 10796 11694 10824 13126
rect 10888 12628 10916 13194
rect 11348 13025 11376 13262
rect 11428 13184 11480 13190
rect 11428 13126 11480 13132
rect 11334 13016 11390 13025
rect 11334 12951 11390 12960
rect 11348 12918 11376 12951
rect 11336 12912 11388 12918
rect 11336 12854 11388 12860
rect 11152 12844 11204 12850
rect 11152 12786 11204 12792
rect 10968 12640 11020 12646
rect 10888 12600 10968 12628
rect 10968 12582 11020 12588
rect 10876 12300 10928 12306
rect 10876 12242 10928 12248
rect 10888 11898 10916 12242
rect 10980 12102 11008 12582
rect 11164 12442 11192 12786
rect 11440 12782 11468 13126
rect 12452 12986 12480 13262
rect 12716 13184 12768 13190
rect 12900 13184 12952 13190
rect 12768 13144 12848 13172
rect 12716 13126 12768 13132
rect 12440 12980 12492 12986
rect 12440 12922 12492 12928
rect 11428 12776 11480 12782
rect 11428 12718 11480 12724
rect 11520 12708 11572 12714
rect 11520 12650 11572 12656
rect 11336 12640 11388 12646
rect 11336 12582 11388 12588
rect 11152 12436 11204 12442
rect 11152 12378 11204 12384
rect 10968 12096 11020 12102
rect 10968 12038 11020 12044
rect 10876 11892 10928 11898
rect 10876 11834 10928 11840
rect 11060 11892 11112 11898
rect 11060 11834 11112 11840
rect 10876 11756 10928 11762
rect 10876 11698 10928 11704
rect 10692 11688 10744 11694
rect 10692 11630 10744 11636
rect 10784 11688 10836 11694
rect 10784 11630 10836 11636
rect 10704 11354 10732 11630
rect 10692 11348 10744 11354
rect 10692 11290 10744 11296
rect 10060 11206 10272 11234
rect 9956 11144 10008 11150
rect 9956 11086 10008 11092
rect 10060 10826 10088 11206
rect 10138 11112 10194 11121
rect 10244 11082 10272 11206
rect 10690 11112 10746 11121
rect 10138 11047 10140 11056
rect 10192 11047 10194 11056
rect 10232 11076 10284 11082
rect 10140 11018 10192 11024
rect 10232 11018 10284 11024
rect 10600 11076 10652 11082
rect 10690 11047 10746 11056
rect 10600 11018 10652 11024
rect 10508 11008 10560 11014
rect 10508 10950 10560 10956
rect 10144 10908 10452 10928
rect 10144 10906 10150 10908
rect 10206 10906 10230 10908
rect 10286 10906 10310 10908
rect 10366 10906 10390 10908
rect 10446 10906 10452 10908
rect 10206 10854 10208 10906
rect 10388 10854 10390 10906
rect 10144 10852 10150 10854
rect 10206 10852 10230 10854
rect 10286 10852 10310 10854
rect 10366 10852 10390 10854
rect 10446 10852 10452 10854
rect 10144 10832 10452 10852
rect 9968 10798 10088 10826
rect 9968 10674 9996 10798
rect 10232 10736 10284 10742
rect 10232 10678 10284 10684
rect 9956 10668 10008 10674
rect 9956 10610 10008 10616
rect 9692 10254 9904 10282
rect 10244 10266 10272 10678
rect 10232 10260 10284 10266
rect 9588 9580 9640 9586
rect 9588 9522 9640 9528
rect 9600 9178 9628 9522
rect 9692 9450 9720 10254
rect 10232 10202 10284 10208
rect 9956 10192 10008 10198
rect 9956 10134 10008 10140
rect 9772 10124 9824 10130
rect 9772 10066 9824 10072
rect 9680 9444 9732 9450
rect 9680 9386 9732 9392
rect 9588 9172 9640 9178
rect 9588 9114 9640 9120
rect 9784 9042 9812 10066
rect 9864 9920 9916 9926
rect 9864 9862 9916 9868
rect 9876 9722 9904 9862
rect 9864 9716 9916 9722
rect 9864 9658 9916 9664
rect 9968 9586 9996 10134
rect 10520 10130 10548 10950
rect 10508 10124 10560 10130
rect 10508 10066 10560 10072
rect 10416 10056 10468 10062
rect 10468 10004 10548 10010
rect 10416 9998 10548 10004
rect 10428 9982 10548 9998
rect 10048 9920 10100 9926
rect 10048 9862 10100 9868
rect 9956 9580 10008 9586
rect 9956 9522 10008 9528
rect 10060 9178 10088 9862
rect 10144 9820 10452 9840
rect 10144 9818 10150 9820
rect 10206 9818 10230 9820
rect 10286 9818 10310 9820
rect 10366 9818 10390 9820
rect 10446 9818 10452 9820
rect 10206 9766 10208 9818
rect 10388 9766 10390 9818
rect 10144 9764 10150 9766
rect 10206 9764 10230 9766
rect 10286 9764 10310 9766
rect 10366 9764 10390 9766
rect 10446 9764 10452 9766
rect 10144 9744 10452 9764
rect 10232 9512 10284 9518
rect 10232 9454 10284 9460
rect 10244 9178 10272 9454
rect 10520 9382 10548 9982
rect 10612 9586 10640 11018
rect 10704 10810 10732 11047
rect 10692 10804 10744 10810
rect 10692 10746 10744 10752
rect 10796 10062 10824 11630
rect 10888 10146 10916 11698
rect 11072 11370 11100 11834
rect 11164 11830 11192 12378
rect 11152 11824 11204 11830
rect 11152 11766 11204 11772
rect 10980 11342 11100 11370
rect 10980 11286 11008 11342
rect 10968 11280 11020 11286
rect 10968 11222 11020 11228
rect 11164 11150 11192 11766
rect 11348 11762 11376 12582
rect 11532 12434 11560 12650
rect 12443 12540 12751 12560
rect 12443 12538 12449 12540
rect 12505 12538 12529 12540
rect 12585 12538 12609 12540
rect 12665 12538 12689 12540
rect 12745 12538 12751 12540
rect 12505 12486 12507 12538
rect 12687 12486 12689 12538
rect 12443 12484 12449 12486
rect 12505 12484 12529 12486
rect 12585 12484 12609 12486
rect 12665 12484 12689 12486
rect 12745 12484 12751 12486
rect 12443 12464 12751 12484
rect 11796 12436 11848 12442
rect 11532 12406 11744 12434
rect 11612 12096 11664 12102
rect 11612 12038 11664 12044
rect 11624 11830 11652 12038
rect 11612 11824 11664 11830
rect 11612 11766 11664 11772
rect 11244 11756 11296 11762
rect 11244 11698 11296 11704
rect 11336 11756 11388 11762
rect 11336 11698 11388 11704
rect 11520 11756 11572 11762
rect 11520 11698 11572 11704
rect 11256 11354 11284 11698
rect 11244 11348 11296 11354
rect 11244 11290 11296 11296
rect 11532 11286 11560 11698
rect 11612 11552 11664 11558
rect 11612 11494 11664 11500
rect 11520 11280 11572 11286
rect 11520 11222 11572 11228
rect 11624 11150 11652 11494
rect 11716 11218 11744 12406
rect 11796 12378 11848 12384
rect 11808 11694 11836 12378
rect 12348 12300 12400 12306
rect 12348 12242 12400 12248
rect 12164 12164 12216 12170
rect 12164 12106 12216 12112
rect 12176 11694 12204 12106
rect 12256 12096 12308 12102
rect 12256 12038 12308 12044
rect 11796 11688 11848 11694
rect 11796 11630 11848 11636
rect 12164 11688 12216 11694
rect 12164 11630 12216 11636
rect 11704 11212 11756 11218
rect 11704 11154 11756 11160
rect 11152 11144 11204 11150
rect 11152 11086 11204 11092
rect 11612 11144 11664 11150
rect 11612 11086 11664 11092
rect 11060 11008 11112 11014
rect 11060 10950 11112 10956
rect 10968 10600 11020 10606
rect 10968 10542 11020 10548
rect 10980 10266 11008 10542
rect 10968 10260 11020 10266
rect 10968 10202 11020 10208
rect 10888 10118 11008 10146
rect 10784 10056 10836 10062
rect 10784 9998 10836 10004
rect 10980 9602 11008 10118
rect 11072 10062 11100 10950
rect 11716 10538 11744 11154
rect 11808 11098 11836 11630
rect 12072 11144 12124 11150
rect 11808 11070 11928 11098
rect 12072 11086 12124 11092
rect 11704 10532 11756 10538
rect 11704 10474 11756 10480
rect 11244 10464 11296 10470
rect 11244 10406 11296 10412
rect 11520 10464 11572 10470
rect 11520 10406 11572 10412
rect 11256 10062 11284 10406
rect 11532 10130 11560 10406
rect 11716 10130 11744 10474
rect 11520 10124 11572 10130
rect 11520 10066 11572 10072
rect 11704 10124 11756 10130
rect 11704 10066 11756 10072
rect 11060 10056 11112 10062
rect 11058 10024 11060 10033
rect 11244 10056 11296 10062
rect 11112 10024 11114 10033
rect 11244 9998 11296 10004
rect 11058 9959 11114 9968
rect 11704 9920 11756 9926
rect 11704 9862 11756 9868
rect 11716 9722 11744 9862
rect 11704 9716 11756 9722
rect 11704 9658 11756 9664
rect 10980 9586 11652 9602
rect 11900 9586 11928 11070
rect 10600 9580 10652 9586
rect 10980 9580 11664 9586
rect 10980 9574 11612 9580
rect 10600 9522 10652 9528
rect 11612 9522 11664 9528
rect 11888 9580 11940 9586
rect 11888 9522 11940 9528
rect 11428 9512 11480 9518
rect 11428 9454 11480 9460
rect 10692 9444 10744 9450
rect 10692 9386 10744 9392
rect 10508 9376 10560 9382
rect 10508 9318 10560 9324
rect 10048 9172 10100 9178
rect 10048 9114 10100 9120
rect 10232 9172 10284 9178
rect 10232 9114 10284 9120
rect 10704 9042 10732 9386
rect 9496 9036 9548 9042
rect 9496 8978 9548 8984
rect 9772 9036 9824 9042
rect 9772 8978 9824 8984
rect 10692 9036 10744 9042
rect 10692 8978 10744 8984
rect 8944 8832 8996 8838
rect 8944 8774 8996 8780
rect 8668 8560 8720 8566
rect 8668 8502 8720 8508
rect 8484 8492 8536 8498
rect 8484 8434 8536 8440
rect 8208 8356 8260 8362
rect 8208 8298 8260 8304
rect 7846 8188 8154 8208
rect 7846 8186 7852 8188
rect 7908 8186 7932 8188
rect 7988 8186 8012 8188
rect 8068 8186 8092 8188
rect 8148 8186 8154 8188
rect 7908 8134 7910 8186
rect 8090 8134 8092 8186
rect 7846 8132 7852 8134
rect 7908 8132 7932 8134
rect 7988 8132 8012 8134
rect 8068 8132 8092 8134
rect 8148 8132 8154 8134
rect 7846 8112 8154 8132
rect 8220 7886 8248 8298
rect 7748 7880 7800 7886
rect 7748 7822 7800 7828
rect 8208 7880 8260 7886
rect 8208 7822 8260 7828
rect 7760 7546 7788 7822
rect 8496 7818 8524 8434
rect 8680 7886 8708 8502
rect 8760 8492 8812 8498
rect 8760 8434 8812 8440
rect 8772 7954 8800 8434
rect 8760 7948 8812 7954
rect 8760 7890 8812 7896
rect 8668 7880 8720 7886
rect 8668 7822 8720 7828
rect 8484 7812 8536 7818
rect 8484 7754 8536 7760
rect 8956 7750 8984 8774
rect 9508 8634 9536 8978
rect 9956 8832 10008 8838
rect 9956 8774 10008 8780
rect 9496 8628 9548 8634
rect 9496 8570 9548 8576
rect 9220 8424 9272 8430
rect 9220 8366 9272 8372
rect 9128 8288 9180 8294
rect 9128 8230 9180 8236
rect 8576 7744 8628 7750
rect 8576 7686 8628 7692
rect 8944 7744 8996 7750
rect 8944 7686 8996 7692
rect 7472 7540 7524 7546
rect 7472 7482 7524 7488
rect 7748 7540 7800 7546
rect 7748 7482 7800 7488
rect 8588 7478 8616 7686
rect 9140 7478 9168 8230
rect 9232 8090 9260 8366
rect 9220 8084 9272 8090
rect 9220 8026 9272 8032
rect 7380 7472 7432 7478
rect 7380 7414 7432 7420
rect 8576 7472 8628 7478
rect 8576 7414 8628 7420
rect 9128 7472 9180 7478
rect 9128 7414 9180 7420
rect 7104 7404 7156 7410
rect 7104 7346 7156 7352
rect 7196 7404 7248 7410
rect 7196 7346 7248 7352
rect 6828 7336 6880 7342
rect 6828 7278 6880 7284
rect 6736 7200 6788 7206
rect 6736 7142 6788 7148
rect 4896 6860 4948 6866
rect 4896 6802 4948 6808
rect 5908 6860 5960 6866
rect 5908 6802 5960 6808
rect 4620 6792 4672 6798
rect 4620 6734 4672 6740
rect 4528 6724 4580 6730
rect 4448 6684 4528 6712
rect 4528 6666 4580 6672
rect 3976 6656 4028 6662
rect 3620 6322 3832 6338
rect 3240 6316 3292 6322
rect 3240 6258 3292 6264
rect 3608 6316 3832 6322
rect 3660 6310 3832 6316
rect 3896 6616 3976 6644
rect 3608 6258 3660 6264
rect 2964 6248 3016 6254
rect 2964 6190 3016 6196
rect 2780 6180 2832 6186
rect 2780 6122 2832 6128
rect 2688 5840 2740 5846
rect 2688 5782 2740 5788
rect 2688 5704 2740 5710
rect 2608 5664 2688 5692
rect 2412 5636 2464 5642
rect 2412 5578 2464 5584
rect 1676 5228 1728 5234
rect 1676 5170 1728 5176
rect 1400 5024 1452 5030
rect 1400 4966 1452 4972
rect 1412 4146 1440 4966
rect 1688 4690 1716 5170
rect 2424 5030 2452 5578
rect 2502 5536 2558 5545
rect 2502 5471 2558 5480
rect 2516 5234 2544 5471
rect 2504 5228 2556 5234
rect 2504 5170 2556 5176
rect 2608 5148 2636 5664
rect 2688 5646 2740 5652
rect 2688 5296 2740 5302
rect 2792 5250 2820 6122
rect 3248 6012 3556 6032
rect 3248 6010 3254 6012
rect 3310 6010 3334 6012
rect 3390 6010 3414 6012
rect 3470 6010 3494 6012
rect 3550 6010 3556 6012
rect 3310 5958 3312 6010
rect 3492 5958 3494 6010
rect 3248 5956 3254 5958
rect 3310 5956 3334 5958
rect 3390 5956 3414 5958
rect 3470 5956 3494 5958
rect 3550 5956 3556 5958
rect 3248 5936 3556 5956
rect 3240 5772 3292 5778
rect 3240 5714 3292 5720
rect 3056 5568 3108 5574
rect 2740 5244 2820 5250
rect 2688 5238 2820 5244
rect 2700 5222 2820 5238
rect 2884 5516 3056 5522
rect 2884 5510 3108 5516
rect 2884 5494 3096 5510
rect 2688 5160 2740 5166
rect 2608 5120 2688 5148
rect 2688 5102 2740 5108
rect 2884 5098 2912 5494
rect 3252 5370 3280 5714
rect 3620 5574 3648 6258
rect 3896 6254 3924 6616
rect 3976 6598 4028 6604
rect 3976 6316 4028 6322
rect 3976 6258 4028 6264
rect 4436 6316 4488 6322
rect 4436 6258 4488 6264
rect 4804 6316 4856 6322
rect 4804 6258 4856 6264
rect 3884 6248 3936 6254
rect 3884 6190 3936 6196
rect 3608 5568 3660 5574
rect 3608 5510 3660 5516
rect 3988 5370 4016 6258
rect 4160 6248 4212 6254
rect 4160 6190 4212 6196
rect 4068 5704 4120 5710
rect 4068 5646 4120 5652
rect 4080 5370 4108 5646
rect 3240 5364 3292 5370
rect 3240 5306 3292 5312
rect 3976 5364 4028 5370
rect 3976 5306 4028 5312
rect 4068 5364 4120 5370
rect 4068 5306 4120 5312
rect 4172 5234 4200 6190
rect 4448 5846 4476 6258
rect 4620 6112 4672 6118
rect 4620 6054 4672 6060
rect 4632 5914 4660 6054
rect 4816 5914 4844 6258
rect 4620 5908 4672 5914
rect 4620 5850 4672 5856
rect 4804 5908 4856 5914
rect 4804 5850 4856 5856
rect 4436 5840 4488 5846
rect 4436 5782 4488 5788
rect 4620 5704 4672 5710
rect 4620 5646 4672 5652
rect 4632 5545 4660 5646
rect 4804 5568 4856 5574
rect 4618 5536 4674 5545
rect 4804 5510 4856 5516
rect 4618 5471 4674 5480
rect 2964 5228 3016 5234
rect 2964 5170 3016 5176
rect 3608 5228 3660 5234
rect 3608 5170 3660 5176
rect 3700 5228 3752 5234
rect 3700 5170 3752 5176
rect 4160 5228 4212 5234
rect 4160 5170 4212 5176
rect 4528 5228 4580 5234
rect 4528 5170 4580 5176
rect 4712 5228 4764 5234
rect 4712 5170 4764 5176
rect 2872 5092 2924 5098
rect 2872 5034 2924 5040
rect 2412 5024 2464 5030
rect 2412 4966 2464 4972
rect 2688 5024 2740 5030
rect 2688 4966 2740 4972
rect 2700 4758 2728 4966
rect 2688 4752 2740 4758
rect 2688 4694 2740 4700
rect 1676 4684 1728 4690
rect 1676 4626 1728 4632
rect 1400 4140 1452 4146
rect 1400 4082 1452 4088
rect 1688 2990 1716 4626
rect 2700 4554 2728 4694
rect 1768 4548 1820 4554
rect 1768 4490 1820 4496
rect 2688 4548 2740 4554
rect 2688 4490 2740 4496
rect 1780 4282 1808 4490
rect 1768 4276 1820 4282
rect 1768 4218 1820 4224
rect 2700 4214 2728 4490
rect 2976 4486 3004 5170
rect 3240 5160 3292 5166
rect 3160 5120 3240 5148
rect 3056 5024 3108 5030
rect 3056 4966 3108 4972
rect 3068 4690 3096 4966
rect 3160 4826 3188 5120
rect 3240 5102 3292 5108
rect 3248 4924 3556 4944
rect 3248 4922 3254 4924
rect 3310 4922 3334 4924
rect 3390 4922 3414 4924
rect 3470 4922 3494 4924
rect 3550 4922 3556 4924
rect 3310 4870 3312 4922
rect 3492 4870 3494 4922
rect 3248 4868 3254 4870
rect 3310 4868 3334 4870
rect 3390 4868 3414 4870
rect 3470 4868 3494 4870
rect 3550 4868 3556 4870
rect 3248 4848 3556 4868
rect 3148 4820 3200 4826
rect 3148 4762 3200 4768
rect 3056 4684 3108 4690
rect 3056 4626 3108 4632
rect 2964 4480 3016 4486
rect 3240 4480 3292 4486
rect 2964 4422 3016 4428
rect 3160 4440 3240 4468
rect 2688 4208 2740 4214
rect 2688 4150 2740 4156
rect 2700 3618 2728 4150
rect 2976 4146 3004 4422
rect 2964 4140 3016 4146
rect 2964 4082 3016 4088
rect 2780 4072 2832 4078
rect 2780 4014 2832 4020
rect 2792 3738 2820 4014
rect 2780 3732 2832 3738
rect 2780 3674 2832 3680
rect 2700 3590 2820 3618
rect 2792 3398 2820 3590
rect 3160 3466 3188 4440
rect 3240 4422 3292 4428
rect 3620 4146 3648 5170
rect 3712 4554 3740 5170
rect 3792 5160 3844 5166
rect 3792 5102 3844 5108
rect 3700 4548 3752 4554
rect 3700 4490 3752 4496
rect 3804 4486 3832 5102
rect 4160 5092 4212 5098
rect 4160 5034 4212 5040
rect 4172 4622 4200 5034
rect 4342 4720 4398 4729
rect 4342 4655 4398 4664
rect 4356 4622 4384 4655
rect 4540 4622 4568 5170
rect 4724 4758 4752 5170
rect 4712 4752 4764 4758
rect 4712 4694 4764 4700
rect 4816 4622 4844 5510
rect 4908 5166 4936 6802
rect 5540 6792 5592 6798
rect 5460 6740 5540 6746
rect 5460 6734 5592 6740
rect 5460 6718 5580 6734
rect 5080 6656 5132 6662
rect 5080 6598 5132 6604
rect 5172 6656 5224 6662
rect 5172 6598 5224 6604
rect 5092 6458 5120 6598
rect 5080 6452 5132 6458
rect 5080 6394 5132 6400
rect 5184 6254 5212 6598
rect 5356 6316 5408 6322
rect 5356 6258 5408 6264
rect 4988 6248 5040 6254
rect 4988 6190 5040 6196
rect 5172 6248 5224 6254
rect 5172 6190 5224 6196
rect 5264 6248 5316 6254
rect 5264 6190 5316 6196
rect 4896 5160 4948 5166
rect 4896 5102 4948 5108
rect 5000 4706 5028 6190
rect 5080 6180 5132 6186
rect 5080 6122 5132 6128
rect 5092 5234 5120 6122
rect 5276 5914 5304 6190
rect 5264 5908 5316 5914
rect 5264 5850 5316 5856
rect 5276 5386 5304 5850
rect 5184 5358 5304 5386
rect 5080 5228 5132 5234
rect 5080 5170 5132 5176
rect 4908 4690 5028 4706
rect 4896 4684 5028 4690
rect 4948 4678 5028 4684
rect 5184 4706 5212 5358
rect 5264 5228 5316 5234
rect 5264 5170 5316 5176
rect 5276 4826 5304 5170
rect 5368 5030 5396 6258
rect 5460 6254 5488 6718
rect 5547 6556 5855 6576
rect 5547 6554 5553 6556
rect 5609 6554 5633 6556
rect 5689 6554 5713 6556
rect 5769 6554 5793 6556
rect 5849 6554 5855 6556
rect 5609 6502 5611 6554
rect 5791 6502 5793 6554
rect 5547 6500 5553 6502
rect 5609 6500 5633 6502
rect 5689 6500 5713 6502
rect 5769 6500 5793 6502
rect 5849 6500 5855 6502
rect 5547 6480 5855 6500
rect 5920 6474 5948 6802
rect 6644 6792 6696 6798
rect 6644 6734 6696 6740
rect 6552 6724 6604 6730
rect 6552 6666 6604 6672
rect 6460 6656 6512 6662
rect 6460 6598 6512 6604
rect 5920 6446 6132 6474
rect 5920 6338 5948 6446
rect 5828 6322 5948 6338
rect 6000 6384 6052 6390
rect 6000 6326 6052 6332
rect 5816 6316 5948 6322
rect 5868 6310 5948 6316
rect 5816 6258 5868 6264
rect 5448 6248 5500 6254
rect 5448 6190 5500 6196
rect 5356 5024 5408 5030
rect 5356 4966 5408 4972
rect 5264 4820 5316 4826
rect 5264 4762 5316 4768
rect 5184 4678 5304 4706
rect 4896 4626 4948 4632
rect 4160 4616 4212 4622
rect 4160 4558 4212 4564
rect 4344 4616 4396 4622
rect 4344 4558 4396 4564
rect 4528 4616 4580 4622
rect 4528 4558 4580 4564
rect 4804 4616 4856 4622
rect 4804 4558 4856 4564
rect 5172 4616 5224 4622
rect 5172 4558 5224 4564
rect 3792 4480 3844 4486
rect 3792 4422 3844 4428
rect 4172 4214 4200 4558
rect 4252 4480 4304 4486
rect 4252 4422 4304 4428
rect 4160 4208 4212 4214
rect 4160 4150 4212 4156
rect 3516 4140 3568 4146
rect 3516 4082 3568 4088
rect 3608 4140 3660 4146
rect 3608 4082 3660 4088
rect 3884 4140 3936 4146
rect 3884 4082 3936 4088
rect 3528 4026 3556 4082
rect 3528 3998 3648 4026
rect 3248 3836 3556 3856
rect 3248 3834 3254 3836
rect 3310 3834 3334 3836
rect 3390 3834 3414 3836
rect 3470 3834 3494 3836
rect 3550 3834 3556 3836
rect 3310 3782 3312 3834
rect 3492 3782 3494 3834
rect 3248 3780 3254 3782
rect 3310 3780 3334 3782
rect 3390 3780 3414 3782
rect 3470 3780 3494 3782
rect 3550 3780 3556 3782
rect 3248 3760 3556 3780
rect 3620 3738 3648 3998
rect 3896 3738 3924 4082
rect 3976 3936 4028 3942
rect 3976 3878 4028 3884
rect 4068 3936 4120 3942
rect 4172 3913 4200 4150
rect 4068 3878 4120 3884
rect 4158 3904 4214 3913
rect 3608 3732 3660 3738
rect 3608 3674 3660 3680
rect 3884 3732 3936 3738
rect 3884 3674 3936 3680
rect 3988 3670 4016 3878
rect 3976 3664 4028 3670
rect 3790 3632 3846 3641
rect 3976 3606 4028 3612
rect 4080 3602 4108 3878
rect 4158 3839 4214 3848
rect 3790 3567 3846 3576
rect 4068 3596 4120 3602
rect 3804 3534 3832 3567
rect 4068 3538 4120 3544
rect 3424 3528 3476 3534
rect 3422 3496 3424 3505
rect 3792 3528 3844 3534
rect 3476 3496 3478 3505
rect 3148 3460 3200 3466
rect 3792 3470 3844 3476
rect 3422 3431 3478 3440
rect 3148 3402 3200 3408
rect 2780 3392 2832 3398
rect 2780 3334 2832 3340
rect 3608 3392 3660 3398
rect 3608 3334 3660 3340
rect 3792 3392 3844 3398
rect 3792 3334 3844 3340
rect 3620 3074 3648 3334
rect 3804 3194 3832 3334
rect 3792 3188 3844 3194
rect 3792 3130 3844 3136
rect 3884 3120 3936 3126
rect 3620 3068 3884 3074
rect 3620 3062 3936 3068
rect 3620 3046 3924 3062
rect 1676 2984 1728 2990
rect 1676 2926 1728 2932
rect 3248 2748 3556 2768
rect 3248 2746 3254 2748
rect 3310 2746 3334 2748
rect 3390 2746 3414 2748
rect 3470 2746 3494 2748
rect 3550 2746 3556 2748
rect 3310 2694 3312 2746
rect 3492 2694 3494 2746
rect 3248 2692 3254 2694
rect 3310 2692 3334 2694
rect 3390 2692 3414 2694
rect 3470 2692 3494 2694
rect 3550 2692 3556 2694
rect 3248 2672 3556 2692
rect 3896 2310 3924 3046
rect 4264 2990 4292 4422
rect 4540 4185 4568 4558
rect 4526 4176 4582 4185
rect 4526 4111 4582 4120
rect 4804 4140 4856 4146
rect 4804 4082 4856 4088
rect 4344 4072 4396 4078
rect 4344 4014 4396 4020
rect 4526 4040 4582 4049
rect 4356 3466 4384 4014
rect 4526 3975 4528 3984
rect 4580 3975 4582 3984
rect 4528 3946 4580 3952
rect 4816 3466 4844 4082
rect 5184 3738 5212 4558
rect 5276 4146 5304 4678
rect 5264 4140 5316 4146
rect 5264 4082 5316 4088
rect 5172 3732 5224 3738
rect 5172 3674 5224 3680
rect 5276 3641 5304 4082
rect 5368 4078 5396 4966
rect 5356 4072 5408 4078
rect 5356 4014 5408 4020
rect 5460 3670 5488 6190
rect 5908 6180 5960 6186
rect 5908 6122 5960 6128
rect 5632 6112 5684 6118
rect 5632 6054 5684 6060
rect 5644 5710 5672 6054
rect 5632 5704 5684 5710
rect 5632 5646 5684 5652
rect 5547 5468 5855 5488
rect 5547 5466 5553 5468
rect 5609 5466 5633 5468
rect 5689 5466 5713 5468
rect 5769 5466 5793 5468
rect 5849 5466 5855 5468
rect 5609 5414 5611 5466
rect 5791 5414 5793 5466
rect 5547 5412 5553 5414
rect 5609 5412 5633 5414
rect 5689 5412 5713 5414
rect 5769 5412 5793 5414
rect 5849 5412 5855 5414
rect 5547 5392 5855 5412
rect 5920 5370 5948 6122
rect 5908 5364 5960 5370
rect 5908 5306 5960 5312
rect 5722 5264 5778 5273
rect 5722 5199 5778 5208
rect 5816 5228 5868 5234
rect 5736 5030 5764 5199
rect 5816 5170 5868 5176
rect 5908 5228 5960 5234
rect 5908 5170 5960 5176
rect 5724 5024 5776 5030
rect 5724 4966 5776 4972
rect 5828 4690 5856 5170
rect 5920 4690 5948 5170
rect 6012 5166 6040 6326
rect 6104 6254 6132 6446
rect 6092 6248 6144 6254
rect 6092 6190 6144 6196
rect 6092 6112 6144 6118
rect 6092 6054 6144 6060
rect 6104 5710 6132 6054
rect 6092 5704 6144 5710
rect 6092 5646 6144 5652
rect 6184 5704 6236 5710
rect 6184 5646 6236 5652
rect 6000 5160 6052 5166
rect 6196 5114 6224 5646
rect 6276 5228 6328 5234
rect 6276 5170 6328 5176
rect 6000 5102 6052 5108
rect 6104 5098 6224 5114
rect 6092 5092 6224 5098
rect 6144 5086 6224 5092
rect 6092 5034 6144 5040
rect 6288 4826 6316 5170
rect 6472 5030 6500 6598
rect 6564 6390 6592 6666
rect 6552 6384 6604 6390
rect 6552 6326 6604 6332
rect 6564 5098 6592 6326
rect 6552 5092 6604 5098
rect 6552 5034 6604 5040
rect 6368 5024 6420 5030
rect 6368 4966 6420 4972
rect 6460 5024 6512 5030
rect 6460 4966 6512 4972
rect 6276 4820 6328 4826
rect 6276 4762 6328 4768
rect 5816 4684 5868 4690
rect 5816 4626 5868 4632
rect 5908 4684 5960 4690
rect 5908 4626 5960 4632
rect 5908 4480 5960 4486
rect 5908 4422 5960 4428
rect 5547 4380 5855 4400
rect 5547 4378 5553 4380
rect 5609 4378 5633 4380
rect 5689 4378 5713 4380
rect 5769 4378 5793 4380
rect 5849 4378 5855 4380
rect 5609 4326 5611 4378
rect 5791 4326 5793 4378
rect 5547 4324 5553 4326
rect 5609 4324 5633 4326
rect 5689 4324 5713 4326
rect 5769 4324 5793 4326
rect 5849 4324 5855 4326
rect 5547 4304 5855 4324
rect 5920 4282 5948 4422
rect 6380 4282 6408 4966
rect 5908 4276 5960 4282
rect 5908 4218 5960 4224
rect 6368 4276 6420 4282
rect 6368 4218 6420 4224
rect 5538 4176 5594 4185
rect 5538 4111 5594 4120
rect 5552 4078 5580 4111
rect 6472 4078 6500 4966
rect 6564 4146 6592 5034
rect 6656 4570 6684 6734
rect 6748 5778 6776 7142
rect 7208 6934 7236 7346
rect 7748 7336 7800 7342
rect 7748 7278 7800 7284
rect 7288 7200 7340 7206
rect 7288 7142 7340 7148
rect 7380 7200 7432 7206
rect 7380 7142 7432 7148
rect 7196 6928 7248 6934
rect 7196 6870 7248 6876
rect 6828 6656 6880 6662
rect 6828 6598 6880 6604
rect 6736 5772 6788 5778
rect 6736 5714 6788 5720
rect 6736 5568 6788 5574
rect 6736 5510 6788 5516
rect 6748 5166 6776 5510
rect 6840 5234 6868 6598
rect 7196 5908 7248 5914
rect 7196 5850 7248 5856
rect 7104 5636 7156 5642
rect 7104 5578 7156 5584
rect 6932 5370 7052 5386
rect 6920 5364 7052 5370
rect 6972 5358 7052 5364
rect 6920 5306 6972 5312
rect 6828 5228 6880 5234
rect 6828 5170 6880 5176
rect 6920 5228 6972 5234
rect 6920 5170 6972 5176
rect 6736 5160 6788 5166
rect 6736 5102 6788 5108
rect 6736 4616 6788 4622
rect 6656 4564 6736 4570
rect 6656 4558 6788 4564
rect 6656 4542 6776 4558
rect 6656 4214 6684 4542
rect 6828 4480 6880 4486
rect 6828 4422 6880 4428
rect 6644 4208 6696 4214
rect 6644 4150 6696 4156
rect 6552 4140 6604 4146
rect 6552 4082 6604 4088
rect 6656 4078 6684 4150
rect 5540 4072 5592 4078
rect 5540 4014 5592 4020
rect 6460 4072 6512 4078
rect 6644 4072 6696 4078
rect 6460 4014 6512 4020
rect 6564 4020 6644 4026
rect 6564 4014 6696 4020
rect 6564 3998 6684 4014
rect 5538 3904 5594 3913
rect 5538 3839 5594 3848
rect 5448 3664 5500 3670
rect 5262 3632 5318 3641
rect 5448 3606 5500 3612
rect 5262 3567 5264 3576
rect 5316 3567 5318 3576
rect 5264 3538 5316 3544
rect 4896 3528 4948 3534
rect 5276 3507 5304 3538
rect 4896 3470 4948 3476
rect 5170 3496 5226 3505
rect 4344 3460 4396 3466
rect 4344 3402 4396 3408
rect 4804 3460 4856 3466
rect 4804 3402 4856 3408
rect 4356 3194 4384 3402
rect 4908 3194 4936 3470
rect 5170 3431 5172 3440
rect 5224 3431 5226 3440
rect 5172 3402 5224 3408
rect 4344 3188 4396 3194
rect 4344 3130 4396 3136
rect 4896 3188 4948 3194
rect 4896 3130 4948 3136
rect 4252 2984 4304 2990
rect 4252 2926 4304 2932
rect 5460 2854 5488 3606
rect 5552 3534 5580 3839
rect 5540 3528 5592 3534
rect 5540 3470 5592 3476
rect 5547 3292 5855 3312
rect 5547 3290 5553 3292
rect 5609 3290 5633 3292
rect 5689 3290 5713 3292
rect 5769 3290 5793 3292
rect 5849 3290 5855 3292
rect 5609 3238 5611 3290
rect 5791 3238 5793 3290
rect 5547 3236 5553 3238
rect 5609 3236 5633 3238
rect 5689 3236 5713 3238
rect 5769 3236 5793 3238
rect 5849 3236 5855 3238
rect 5547 3216 5855 3236
rect 6564 2990 6592 3998
rect 6840 3942 6868 4422
rect 6932 4010 6960 5170
rect 7024 5098 7052 5358
rect 7012 5092 7064 5098
rect 7012 5034 7064 5040
rect 7116 4978 7144 5578
rect 7208 5302 7236 5850
rect 7300 5370 7328 7142
rect 7392 7002 7420 7142
rect 7380 6996 7432 7002
rect 7380 6938 7432 6944
rect 7472 6656 7524 6662
rect 7472 6598 7524 6604
rect 7484 6474 7512 6598
rect 7392 6458 7512 6474
rect 7380 6452 7512 6458
rect 7432 6446 7512 6452
rect 7380 6394 7432 6400
rect 7380 6316 7432 6322
rect 7432 6276 7604 6304
rect 7380 6258 7432 6264
rect 7380 6180 7432 6186
rect 7380 6122 7432 6128
rect 7288 5364 7340 5370
rect 7288 5306 7340 5312
rect 7196 5296 7248 5302
rect 7196 5238 7248 5244
rect 7024 4950 7144 4978
rect 7024 4622 7052 4950
rect 7104 4820 7156 4826
rect 7104 4762 7156 4768
rect 7012 4616 7064 4622
rect 7012 4558 7064 4564
rect 7012 4480 7064 4486
rect 7012 4422 7064 4428
rect 7024 4146 7052 4422
rect 7116 4146 7144 4762
rect 7392 4690 7420 6122
rect 7472 6112 7524 6118
rect 7472 6054 7524 6060
rect 7380 4684 7432 4690
rect 7380 4626 7432 4632
rect 7392 4214 7420 4626
rect 7484 4282 7512 6054
rect 7576 5302 7604 6276
rect 7760 5778 7788 7278
rect 7846 7100 8154 7120
rect 7846 7098 7852 7100
rect 7908 7098 7932 7100
rect 7988 7098 8012 7100
rect 8068 7098 8092 7100
rect 8148 7098 8154 7100
rect 7908 7046 7910 7098
rect 8090 7046 8092 7098
rect 7846 7044 7852 7046
rect 7908 7044 7932 7046
rect 7988 7044 8012 7046
rect 8068 7044 8092 7046
rect 8148 7044 8154 7046
rect 7846 7024 8154 7044
rect 8588 6798 8616 7414
rect 9508 7410 9536 8570
rect 9680 8424 9732 8430
rect 9680 8366 9732 8372
rect 9692 7886 9720 8366
rect 9968 8294 9996 8774
rect 10144 8732 10452 8752
rect 10144 8730 10150 8732
rect 10206 8730 10230 8732
rect 10286 8730 10310 8732
rect 10366 8730 10390 8732
rect 10446 8730 10452 8732
rect 10206 8678 10208 8730
rect 10388 8678 10390 8730
rect 10144 8676 10150 8678
rect 10206 8676 10230 8678
rect 10286 8676 10310 8678
rect 10366 8676 10390 8678
rect 10446 8676 10452 8678
rect 10144 8656 10452 8676
rect 9956 8288 10008 8294
rect 9956 8230 10008 8236
rect 10784 8288 10836 8294
rect 10784 8230 10836 8236
rect 9968 7886 9996 8230
rect 9680 7880 9732 7886
rect 9680 7822 9732 7828
rect 9956 7880 10008 7886
rect 9956 7822 10008 7828
rect 10796 7818 10824 8230
rect 10784 7812 10836 7818
rect 10784 7754 10836 7760
rect 10144 7644 10452 7664
rect 10144 7642 10150 7644
rect 10206 7642 10230 7644
rect 10286 7642 10310 7644
rect 10366 7642 10390 7644
rect 10446 7642 10452 7644
rect 10206 7590 10208 7642
rect 10388 7590 10390 7642
rect 10144 7588 10150 7590
rect 10206 7588 10230 7590
rect 10286 7588 10310 7590
rect 10366 7588 10390 7590
rect 10446 7588 10452 7590
rect 10144 7568 10452 7588
rect 11440 7546 11468 9454
rect 11900 9178 11928 9522
rect 11888 9172 11940 9178
rect 11888 9114 11940 9120
rect 11900 8514 11928 9114
rect 12084 9042 12112 11086
rect 12176 11014 12204 11630
rect 12164 11008 12216 11014
rect 12164 10950 12216 10956
rect 12268 10674 12296 12038
rect 12360 11694 12388 12242
rect 12820 11830 12848 13144
rect 12900 13126 12952 13132
rect 12912 12918 12940 13126
rect 12900 12912 12952 12918
rect 12900 12854 12952 12860
rect 12912 12102 12940 12854
rect 13004 12782 13032 13330
rect 12992 12776 13044 12782
rect 12992 12718 13044 12724
rect 12900 12096 12952 12102
rect 12900 12038 12952 12044
rect 12808 11824 12860 11830
rect 12808 11766 12860 11772
rect 12348 11688 12400 11694
rect 12348 11630 12400 11636
rect 12360 11150 12388 11630
rect 12900 11552 12952 11558
rect 12900 11494 12952 11500
rect 12443 11452 12751 11472
rect 12443 11450 12449 11452
rect 12505 11450 12529 11452
rect 12585 11450 12609 11452
rect 12665 11450 12689 11452
rect 12745 11450 12751 11452
rect 12505 11398 12507 11450
rect 12687 11398 12689 11450
rect 12443 11396 12449 11398
rect 12505 11396 12529 11398
rect 12585 11396 12609 11398
rect 12665 11396 12689 11398
rect 12745 11396 12751 11398
rect 12443 11376 12751 11396
rect 12348 11144 12400 11150
rect 12348 11086 12400 11092
rect 12164 10668 12216 10674
rect 12164 10610 12216 10616
rect 12256 10668 12308 10674
rect 12256 10610 12308 10616
rect 12176 10266 12204 10610
rect 12443 10364 12751 10384
rect 12443 10362 12449 10364
rect 12505 10362 12529 10364
rect 12585 10362 12609 10364
rect 12665 10362 12689 10364
rect 12745 10362 12751 10364
rect 12505 10310 12507 10362
rect 12687 10310 12689 10362
rect 12443 10308 12449 10310
rect 12505 10308 12529 10310
rect 12585 10308 12609 10310
rect 12665 10308 12689 10310
rect 12745 10308 12751 10310
rect 12443 10288 12751 10308
rect 12164 10260 12216 10266
rect 12164 10202 12216 10208
rect 12912 10130 12940 11494
rect 13004 10266 13032 12718
rect 12992 10260 13044 10266
rect 12992 10202 13044 10208
rect 12900 10124 12952 10130
rect 12900 10066 12952 10072
rect 12164 9920 12216 9926
rect 12164 9862 12216 9868
rect 12176 9518 12204 9862
rect 12256 9580 12308 9586
rect 12256 9522 12308 9528
rect 12808 9580 12860 9586
rect 12808 9522 12860 9528
rect 12164 9512 12216 9518
rect 12164 9454 12216 9460
rect 12072 9036 12124 9042
rect 12072 8978 12124 8984
rect 12176 8906 12204 9454
rect 12164 8900 12216 8906
rect 12164 8842 12216 8848
rect 12268 8566 12296 9522
rect 12348 9376 12400 9382
rect 12348 9318 12400 9324
rect 12256 8560 12308 8566
rect 11900 8498 12020 8514
rect 12256 8502 12308 8508
rect 11796 8492 11848 8498
rect 11900 8492 12032 8498
rect 11900 8486 11980 8492
rect 11796 8434 11848 8440
rect 11980 8434 12032 8440
rect 11808 8106 11836 8434
rect 11716 8078 11836 8106
rect 11716 8022 11744 8078
rect 11704 8016 11756 8022
rect 12360 7970 12388 9318
rect 12443 9276 12751 9296
rect 12443 9274 12449 9276
rect 12505 9274 12529 9276
rect 12585 9274 12609 9276
rect 12665 9274 12689 9276
rect 12745 9274 12751 9276
rect 12505 9222 12507 9274
rect 12687 9222 12689 9274
rect 12443 9220 12449 9222
rect 12505 9220 12529 9222
rect 12585 9220 12609 9222
rect 12665 9220 12689 9222
rect 12745 9220 12751 9222
rect 12443 9200 12751 9220
rect 12624 8832 12676 8838
rect 12624 8774 12676 8780
rect 12636 8362 12664 8774
rect 12624 8356 12676 8362
rect 12624 8298 12676 8304
rect 12443 8188 12751 8208
rect 12443 8186 12449 8188
rect 12505 8186 12529 8188
rect 12585 8186 12609 8188
rect 12665 8186 12689 8188
rect 12745 8186 12751 8188
rect 12505 8134 12507 8186
rect 12687 8134 12689 8186
rect 12443 8132 12449 8134
rect 12505 8132 12529 8134
rect 12585 8132 12609 8134
rect 12665 8132 12689 8134
rect 12745 8132 12751 8134
rect 12443 8112 12751 8132
rect 11704 7958 11756 7964
rect 11428 7540 11480 7546
rect 11428 7482 11480 7488
rect 10508 7472 10560 7478
rect 10508 7414 10560 7420
rect 9496 7404 9548 7410
rect 9496 7346 9548 7352
rect 9588 7404 9640 7410
rect 9588 7346 9640 7352
rect 10140 7404 10192 7410
rect 10140 7346 10192 7352
rect 9600 7002 9628 7346
rect 10152 7274 10180 7346
rect 10140 7268 10192 7274
rect 10140 7210 10192 7216
rect 10152 7002 10180 7210
rect 10520 7206 10548 7414
rect 11716 7410 11744 7958
rect 12268 7954 12480 7970
rect 12268 7948 12492 7954
rect 12268 7942 12440 7948
rect 12164 7880 12216 7886
rect 12164 7822 12216 7828
rect 12176 7546 12204 7822
rect 12164 7540 12216 7546
rect 12084 7500 12164 7528
rect 11704 7404 11756 7410
rect 11704 7346 11756 7352
rect 11612 7268 11664 7274
rect 11612 7210 11664 7216
rect 10508 7200 10560 7206
rect 10508 7142 10560 7148
rect 11428 7200 11480 7206
rect 11428 7142 11480 7148
rect 9588 6996 9640 7002
rect 9588 6938 9640 6944
rect 10140 6996 10192 7002
rect 10140 6938 10192 6944
rect 8852 6928 8904 6934
rect 8852 6870 8904 6876
rect 8576 6792 8628 6798
rect 8576 6734 8628 6740
rect 8668 6724 8720 6730
rect 8720 6684 8800 6712
rect 8668 6666 8720 6672
rect 7840 6656 7892 6662
rect 7840 6598 7892 6604
rect 8484 6656 8536 6662
rect 8484 6598 8536 6604
rect 7852 6390 7880 6598
rect 7840 6384 7892 6390
rect 7840 6326 7892 6332
rect 7846 6012 8154 6032
rect 7846 6010 7852 6012
rect 7908 6010 7932 6012
rect 7988 6010 8012 6012
rect 8068 6010 8092 6012
rect 8148 6010 8154 6012
rect 7908 5958 7910 6010
rect 8090 5958 8092 6010
rect 7846 5956 7852 5958
rect 7908 5956 7932 5958
rect 7988 5956 8012 5958
rect 8068 5956 8092 5958
rect 8148 5956 8154 5958
rect 7846 5936 8154 5956
rect 8024 5840 8076 5846
rect 8024 5782 8076 5788
rect 7656 5772 7708 5778
rect 7656 5714 7708 5720
rect 7748 5772 7800 5778
rect 7748 5714 7800 5720
rect 7668 5658 7696 5714
rect 8036 5710 8064 5782
rect 8024 5704 8076 5710
rect 7668 5630 7788 5658
rect 8024 5646 8076 5652
rect 7564 5296 7616 5302
rect 7564 5238 7616 5244
rect 7564 5160 7616 5166
rect 7564 5102 7616 5108
rect 7576 5030 7604 5102
rect 7656 5092 7708 5098
rect 7656 5034 7708 5040
rect 7564 5024 7616 5030
rect 7564 4966 7616 4972
rect 7576 4690 7604 4966
rect 7564 4684 7616 4690
rect 7564 4626 7616 4632
rect 7668 4622 7696 5034
rect 7760 4690 7788 5630
rect 8392 5568 8444 5574
rect 8392 5510 8444 5516
rect 8404 5302 8432 5510
rect 8300 5296 8352 5302
rect 8300 5238 8352 5244
rect 8392 5296 8444 5302
rect 8392 5238 8444 5244
rect 8208 5024 8260 5030
rect 8208 4966 8260 4972
rect 7846 4924 8154 4944
rect 7846 4922 7852 4924
rect 7908 4922 7932 4924
rect 7988 4922 8012 4924
rect 8068 4922 8092 4924
rect 8148 4922 8154 4924
rect 7908 4870 7910 4922
rect 8090 4870 8092 4922
rect 7846 4868 7852 4870
rect 7908 4868 7932 4870
rect 7988 4868 8012 4870
rect 8068 4868 8092 4870
rect 8148 4868 8154 4870
rect 7846 4848 8154 4868
rect 8220 4729 8248 4966
rect 8206 4720 8262 4729
rect 7748 4684 7800 4690
rect 8312 4690 8340 5238
rect 8206 4655 8262 4664
rect 8300 4684 8352 4690
rect 7748 4626 7800 4632
rect 8300 4626 8352 4632
rect 7656 4616 7708 4622
rect 7656 4558 7708 4564
rect 7472 4276 7524 4282
rect 7472 4218 7524 4224
rect 7196 4208 7248 4214
rect 7196 4150 7248 4156
rect 7380 4208 7432 4214
rect 7380 4150 7432 4156
rect 7012 4140 7064 4146
rect 7012 4082 7064 4088
rect 7104 4140 7156 4146
rect 7104 4082 7156 4088
rect 6920 4004 6972 4010
rect 6920 3946 6972 3952
rect 6828 3936 6880 3942
rect 7012 3936 7064 3942
rect 6880 3884 6960 3890
rect 6828 3878 6960 3884
rect 7012 3878 7064 3884
rect 7104 3936 7156 3942
rect 7104 3878 7156 3884
rect 6840 3862 6960 3878
rect 6932 3466 6960 3862
rect 7024 3602 7052 3878
rect 7012 3596 7064 3602
rect 7012 3538 7064 3544
rect 6920 3460 6972 3466
rect 6920 3402 6972 3408
rect 6644 3392 6696 3398
rect 6644 3334 6696 3340
rect 6656 3058 6684 3334
rect 6932 3126 6960 3402
rect 7116 3194 7144 3878
rect 7104 3188 7156 3194
rect 7104 3130 7156 3136
rect 6920 3120 6972 3126
rect 6920 3062 6972 3068
rect 6644 3052 6696 3058
rect 6644 2994 6696 3000
rect 6552 2984 6604 2990
rect 6552 2926 6604 2932
rect 5448 2848 5500 2854
rect 5448 2790 5500 2796
rect 3976 2440 4028 2446
rect 3976 2382 4028 2388
rect 3884 2304 3936 2310
rect 3884 2246 3936 2252
rect 3988 800 4016 2382
rect 6932 2310 6960 3062
rect 7208 3058 7236 4150
rect 7668 3534 7696 4558
rect 7760 4214 7788 4626
rect 8312 4214 8340 4626
rect 8404 4622 8432 5238
rect 8496 5234 8524 6598
rect 8576 6452 8628 6458
rect 8576 6394 8628 6400
rect 8588 5817 8616 6394
rect 8574 5808 8630 5817
rect 8574 5743 8630 5752
rect 8668 5772 8720 5778
rect 8668 5714 8720 5720
rect 8576 5704 8628 5710
rect 8576 5646 8628 5652
rect 8484 5228 8536 5234
rect 8484 5170 8536 5176
rect 8588 5114 8616 5646
rect 8680 5166 8708 5714
rect 8772 5710 8800 6684
rect 8864 5778 8892 6870
rect 9036 6792 9088 6798
rect 9220 6792 9272 6798
rect 9088 6752 9168 6780
rect 9036 6734 9088 6740
rect 9140 6662 9168 6752
rect 9220 6734 9272 6740
rect 9128 6656 9180 6662
rect 9128 6598 9180 6604
rect 9140 6390 9168 6598
rect 9128 6384 9180 6390
rect 9128 6326 9180 6332
rect 9036 6248 9088 6254
rect 9036 6190 9088 6196
rect 8852 5772 8904 5778
rect 8852 5714 8904 5720
rect 8760 5704 8812 5710
rect 8760 5646 8812 5652
rect 8850 5672 8906 5681
rect 8496 5086 8616 5114
rect 8668 5160 8720 5166
rect 8668 5102 8720 5108
rect 8392 4616 8444 4622
rect 8392 4558 8444 4564
rect 7748 4208 7800 4214
rect 7748 4150 7800 4156
rect 8300 4208 8352 4214
rect 8300 4150 8352 4156
rect 8208 4140 8260 4146
rect 8208 4082 8260 4088
rect 7748 3936 7800 3942
rect 7748 3878 7800 3884
rect 7656 3528 7708 3534
rect 7656 3470 7708 3476
rect 7196 3052 7248 3058
rect 7196 2994 7248 3000
rect 7208 2922 7236 2994
rect 7668 2938 7696 3470
rect 7760 3126 7788 3878
rect 7846 3836 8154 3856
rect 7846 3834 7852 3836
rect 7908 3834 7932 3836
rect 7988 3834 8012 3836
rect 8068 3834 8092 3836
rect 8148 3834 8154 3836
rect 7908 3782 7910 3834
rect 8090 3782 8092 3834
rect 7846 3780 7852 3782
rect 7908 3780 7932 3782
rect 7988 3780 8012 3782
rect 8068 3780 8092 3782
rect 8148 3780 8154 3782
rect 7846 3760 8154 3780
rect 8220 3602 8248 4082
rect 8208 3596 8260 3602
rect 8208 3538 8260 3544
rect 8312 3466 8340 4150
rect 8404 3738 8432 4558
rect 8496 4185 8524 5086
rect 8576 4480 8628 4486
rect 8576 4422 8628 4428
rect 8588 4282 8616 4422
rect 8576 4276 8628 4282
rect 8576 4218 8628 4224
rect 8482 4176 8538 4185
rect 8482 4111 8538 4120
rect 8496 4078 8524 4111
rect 8484 4072 8536 4078
rect 8484 4014 8536 4020
rect 8392 3732 8444 3738
rect 8392 3674 8444 3680
rect 8392 3528 8444 3534
rect 8392 3470 8444 3476
rect 8300 3460 8352 3466
rect 8300 3402 8352 3408
rect 7748 3120 7800 3126
rect 7748 3062 7800 3068
rect 8208 3120 8260 3126
rect 8208 3062 8260 3068
rect 7196 2916 7248 2922
rect 7668 2910 7788 2938
rect 7196 2858 7248 2864
rect 7208 2582 7236 2858
rect 7760 2854 7788 2910
rect 7748 2848 7800 2854
rect 7748 2790 7800 2796
rect 7196 2576 7248 2582
rect 7196 2518 7248 2524
rect 7760 2446 7788 2790
rect 7846 2748 8154 2768
rect 7846 2746 7852 2748
rect 7908 2746 7932 2748
rect 7988 2746 8012 2748
rect 8068 2746 8092 2748
rect 8148 2746 8154 2748
rect 7908 2694 7910 2746
rect 8090 2694 8092 2746
rect 7846 2692 7852 2694
rect 7908 2692 7932 2694
rect 7988 2692 8012 2694
rect 8068 2692 8092 2694
rect 8148 2692 8154 2694
rect 7846 2672 8154 2692
rect 7748 2440 7800 2446
rect 7748 2382 7800 2388
rect 8220 2310 8248 3062
rect 8404 2990 8432 3470
rect 8772 3466 8800 5646
rect 8850 5607 8906 5616
rect 8864 5234 8892 5607
rect 8852 5228 8904 5234
rect 8852 5170 8904 5176
rect 8864 4826 8892 5170
rect 8852 4820 8904 4826
rect 8852 4762 8904 4768
rect 9048 4078 9076 6190
rect 9232 6118 9260 6734
rect 9600 6730 9628 6938
rect 9588 6724 9640 6730
rect 9588 6666 9640 6672
rect 10144 6556 10452 6576
rect 10144 6554 10150 6556
rect 10206 6554 10230 6556
rect 10286 6554 10310 6556
rect 10366 6554 10390 6556
rect 10446 6554 10452 6556
rect 10206 6502 10208 6554
rect 10388 6502 10390 6554
rect 10144 6500 10150 6502
rect 10206 6500 10230 6502
rect 10286 6500 10310 6502
rect 10366 6500 10390 6502
rect 10446 6500 10452 6502
rect 10144 6480 10452 6500
rect 10520 6390 10548 7142
rect 11152 6996 11204 7002
rect 11152 6938 11204 6944
rect 11164 6730 11192 6938
rect 11440 6798 11468 7142
rect 11520 6860 11572 6866
rect 11520 6802 11572 6808
rect 11428 6792 11480 6798
rect 11428 6734 11480 6740
rect 11152 6724 11204 6730
rect 11152 6666 11204 6672
rect 11336 6724 11388 6730
rect 11336 6666 11388 6672
rect 10968 6656 11020 6662
rect 10968 6598 11020 6604
rect 10048 6384 10100 6390
rect 10508 6384 10560 6390
rect 10048 6326 10100 6332
rect 10230 6352 10286 6361
rect 9864 6316 9916 6322
rect 9864 6258 9916 6264
rect 9404 6180 9456 6186
rect 9404 6122 9456 6128
rect 9220 6112 9272 6118
rect 9220 6054 9272 6060
rect 9218 5808 9274 5817
rect 9416 5778 9444 6122
rect 9496 6112 9548 6118
rect 9496 6054 9548 6060
rect 9508 5846 9536 6054
rect 9496 5840 9548 5846
rect 9876 5817 9904 6258
rect 9956 5908 10008 5914
rect 9956 5850 10008 5856
rect 9496 5782 9548 5788
rect 9862 5808 9918 5817
rect 9218 5743 9220 5752
rect 9272 5743 9274 5752
rect 9404 5772 9456 5778
rect 9220 5714 9272 5720
rect 9404 5714 9456 5720
rect 9220 5636 9272 5642
rect 9220 5578 9272 5584
rect 9232 5302 9260 5578
rect 9220 5296 9272 5302
rect 9220 5238 9272 5244
rect 9508 5030 9536 5782
rect 9588 5772 9640 5778
rect 9862 5743 9918 5752
rect 9588 5714 9640 5720
rect 9312 5024 9364 5030
rect 9312 4966 9364 4972
rect 9496 5024 9548 5030
rect 9496 4966 9548 4972
rect 9324 4826 9352 4966
rect 9312 4820 9364 4826
rect 9312 4762 9364 4768
rect 9496 4684 9548 4690
rect 9496 4626 9548 4632
rect 9508 4146 9536 4626
rect 9600 4622 9628 5714
rect 9680 5228 9732 5234
rect 9680 5170 9732 5176
rect 9588 4616 9640 4622
rect 9588 4558 9640 4564
rect 9496 4140 9548 4146
rect 9496 4082 9548 4088
rect 9036 4072 9088 4078
rect 9036 4014 9088 4020
rect 9508 3602 9536 4082
rect 9496 3596 9548 3602
rect 9496 3538 9548 3544
rect 8668 3460 8720 3466
rect 8668 3402 8720 3408
rect 8760 3460 8812 3466
rect 8760 3402 8812 3408
rect 8392 2984 8444 2990
rect 8392 2926 8444 2932
rect 8680 2836 8708 3402
rect 9312 3392 9364 3398
rect 9312 3334 9364 3340
rect 9036 3052 9088 3058
rect 9036 2994 9088 3000
rect 8852 2848 8904 2854
rect 8680 2808 8852 2836
rect 8680 2378 8708 2808
rect 8852 2790 8904 2796
rect 9048 2417 9076 2994
rect 9220 2984 9272 2990
rect 9220 2926 9272 2932
rect 9232 2446 9260 2926
rect 9324 2650 9352 3334
rect 9600 3194 9628 4558
rect 9692 4026 9720 5170
rect 9876 5166 9904 5743
rect 9864 5160 9916 5166
rect 9770 5128 9826 5137
rect 9968 5148 9996 5850
rect 10060 5642 10088 6326
rect 10508 6326 10560 6332
rect 10230 6287 10232 6296
rect 10284 6287 10286 6296
rect 10232 6258 10284 6264
rect 10980 5778 11008 6598
rect 11348 6361 11376 6666
rect 11334 6352 11390 6361
rect 11244 6316 11296 6322
rect 11334 6287 11390 6296
rect 11244 6258 11296 6264
rect 10968 5772 11020 5778
rect 10968 5714 11020 5720
rect 10508 5704 10560 5710
rect 10876 5704 10928 5710
rect 10508 5646 10560 5652
rect 10874 5672 10876 5681
rect 11060 5704 11112 5710
rect 10928 5672 10930 5681
rect 10048 5636 10100 5642
rect 10048 5578 10100 5584
rect 10144 5468 10452 5488
rect 10144 5466 10150 5468
rect 10206 5466 10230 5468
rect 10286 5466 10310 5468
rect 10366 5466 10390 5468
rect 10446 5466 10452 5468
rect 10206 5414 10208 5466
rect 10388 5414 10390 5466
rect 10144 5412 10150 5414
rect 10206 5412 10230 5414
rect 10286 5412 10310 5414
rect 10366 5412 10390 5414
rect 10446 5412 10452 5414
rect 10144 5392 10452 5412
rect 10520 5370 10548 5646
rect 11060 5646 11112 5652
rect 10874 5607 10930 5616
rect 10508 5364 10560 5370
rect 10508 5306 10560 5312
rect 10508 5228 10560 5234
rect 10508 5170 10560 5176
rect 10692 5228 10744 5234
rect 10692 5170 10744 5176
rect 10048 5160 10100 5166
rect 9968 5120 10048 5148
rect 9864 5102 9916 5108
rect 10048 5102 10100 5108
rect 9770 5063 9772 5072
rect 9824 5063 9826 5072
rect 9772 5034 9824 5040
rect 10140 5024 10192 5030
rect 10140 4966 10192 4972
rect 10152 4690 10180 4966
rect 10520 4690 10548 5170
rect 10704 4826 10732 5170
rect 10784 5160 10836 5166
rect 10784 5102 10836 5108
rect 10692 4820 10744 4826
rect 10692 4762 10744 4768
rect 10140 4684 10192 4690
rect 10140 4626 10192 4632
rect 10508 4684 10560 4690
rect 10508 4626 10560 4632
rect 10144 4380 10452 4400
rect 10144 4378 10150 4380
rect 10206 4378 10230 4380
rect 10286 4378 10310 4380
rect 10366 4378 10390 4380
rect 10446 4378 10452 4380
rect 10206 4326 10208 4378
rect 10388 4326 10390 4378
rect 10144 4324 10150 4326
rect 10206 4324 10230 4326
rect 10286 4324 10310 4326
rect 10366 4324 10390 4326
rect 10446 4324 10452 4326
rect 10144 4304 10452 4324
rect 10508 4140 10560 4146
rect 10508 4082 10560 4088
rect 9692 4010 9812 4026
rect 9692 4004 9824 4010
rect 9692 3998 9772 4004
rect 9772 3946 9824 3952
rect 9680 3936 9732 3942
rect 9680 3878 9732 3884
rect 9692 3194 9720 3878
rect 10520 3602 10548 4082
rect 10692 3664 10744 3670
rect 10690 3632 10692 3641
rect 10744 3632 10746 3641
rect 9772 3596 9824 3602
rect 9772 3538 9824 3544
rect 10508 3596 10560 3602
rect 10690 3567 10746 3576
rect 10508 3538 10560 3544
rect 9588 3188 9640 3194
rect 9588 3130 9640 3136
rect 9680 3188 9732 3194
rect 9680 3130 9732 3136
rect 9312 2644 9364 2650
rect 9312 2586 9364 2592
rect 9600 2514 9628 3130
rect 9784 3126 9812 3538
rect 10140 3528 10192 3534
rect 10060 3476 10140 3482
rect 10060 3470 10192 3476
rect 10060 3454 10180 3470
rect 9772 3120 9824 3126
rect 9772 3062 9824 3068
rect 9954 3088 10010 3097
rect 9876 3032 9954 3040
rect 9876 3012 9956 3032
rect 9772 2916 9824 2922
rect 9772 2858 9824 2864
rect 9588 2508 9640 2514
rect 9588 2450 9640 2456
rect 9220 2440 9272 2446
rect 9034 2408 9090 2417
rect 8668 2372 8720 2378
rect 9220 2382 9272 2388
rect 9784 2378 9812 2858
rect 9034 2343 9090 2352
rect 9772 2372 9824 2378
rect 8668 2314 8720 2320
rect 9048 2310 9076 2343
rect 9772 2314 9824 2320
rect 6920 2304 6972 2310
rect 6920 2246 6972 2252
rect 8208 2304 8260 2310
rect 8208 2246 8260 2252
rect 9036 2304 9088 2310
rect 9036 2246 9088 2252
rect 9404 2304 9456 2310
rect 9876 2258 9904 3012
rect 10008 3023 10010 3032
rect 9956 2994 10008 3000
rect 10060 2990 10088 3454
rect 10144 3292 10452 3312
rect 10144 3290 10150 3292
rect 10206 3290 10230 3292
rect 10286 3290 10310 3292
rect 10366 3290 10390 3292
rect 10446 3290 10452 3292
rect 10206 3238 10208 3290
rect 10388 3238 10390 3290
rect 10144 3236 10150 3238
rect 10206 3236 10230 3238
rect 10286 3236 10310 3238
rect 10366 3236 10390 3238
rect 10446 3236 10452 3238
rect 10144 3216 10452 3236
rect 10520 3058 10548 3538
rect 10692 3460 10744 3466
rect 10692 3402 10744 3408
rect 10600 3392 10652 3398
rect 10598 3360 10600 3369
rect 10652 3360 10654 3369
rect 10598 3295 10654 3304
rect 10704 3194 10732 3402
rect 10600 3188 10652 3194
rect 10600 3130 10652 3136
rect 10692 3188 10744 3194
rect 10692 3130 10744 3136
rect 10508 3052 10560 3058
rect 10508 2994 10560 3000
rect 10048 2984 10100 2990
rect 10612 2972 10640 3130
rect 10796 3126 10824 5102
rect 11072 5030 11100 5646
rect 11060 5024 11112 5030
rect 11060 4966 11112 4972
rect 11060 4820 11112 4826
rect 11060 4762 11112 4768
rect 11072 4146 11100 4762
rect 11060 4140 11112 4146
rect 11060 4082 11112 4088
rect 11060 3936 11112 3942
rect 11060 3878 11112 3884
rect 10876 3664 10928 3670
rect 10876 3606 10928 3612
rect 10784 3120 10836 3126
rect 10784 3062 10836 3068
rect 10888 2972 10916 3606
rect 11072 3466 11100 3878
rect 11060 3460 11112 3466
rect 11060 3402 11112 3408
rect 11072 3126 11100 3402
rect 11256 3398 11284 6258
rect 11348 4078 11376 6287
rect 11428 6112 11480 6118
rect 11428 6054 11480 6060
rect 11440 5574 11468 6054
rect 11428 5568 11480 5574
rect 11428 5510 11480 5516
rect 11440 4554 11468 5510
rect 11532 5370 11560 6802
rect 11624 6798 11652 7210
rect 11612 6792 11664 6798
rect 11612 6734 11664 6740
rect 11704 6724 11756 6730
rect 11704 6666 11756 6672
rect 11796 6724 11848 6730
rect 11796 6666 11848 6672
rect 11716 6458 11744 6666
rect 11704 6452 11756 6458
rect 11704 6394 11756 6400
rect 11704 6316 11756 6322
rect 11808 6304 11836 6666
rect 11756 6276 11836 6304
rect 11888 6316 11940 6322
rect 11704 6258 11756 6264
rect 11888 6258 11940 6264
rect 11796 5636 11848 5642
rect 11796 5578 11848 5584
rect 11520 5364 11572 5370
rect 11520 5306 11572 5312
rect 11808 5137 11836 5578
rect 11794 5128 11850 5137
rect 11794 5063 11850 5072
rect 11428 4548 11480 4554
rect 11428 4490 11480 4496
rect 11336 4072 11388 4078
rect 11336 4014 11388 4020
rect 11440 3942 11468 4490
rect 11900 4486 11928 6258
rect 12084 5846 12112 7500
rect 12164 7482 12216 7488
rect 12268 6474 12296 7942
rect 12440 7890 12492 7896
rect 12348 7744 12400 7750
rect 12348 7686 12400 7692
rect 12360 7478 12388 7686
rect 12348 7472 12400 7478
rect 12348 7414 12400 7420
rect 12360 6730 12388 7414
rect 12443 7100 12751 7120
rect 12443 7098 12449 7100
rect 12505 7098 12529 7100
rect 12585 7098 12609 7100
rect 12665 7098 12689 7100
rect 12745 7098 12751 7100
rect 12505 7046 12507 7098
rect 12687 7046 12689 7098
rect 12443 7044 12449 7046
rect 12505 7044 12529 7046
rect 12585 7044 12609 7046
rect 12665 7044 12689 7046
rect 12745 7044 12751 7046
rect 12443 7024 12751 7044
rect 12348 6724 12400 6730
rect 12348 6666 12400 6672
rect 12176 6458 12296 6474
rect 12164 6452 12296 6458
rect 12216 6446 12296 6452
rect 12164 6394 12216 6400
rect 12360 6322 12388 6666
rect 12348 6316 12400 6322
rect 12348 6258 12400 6264
rect 12164 6180 12216 6186
rect 12164 6122 12216 6128
rect 12072 5840 12124 5846
rect 12072 5782 12124 5788
rect 11980 5364 12032 5370
rect 12084 5352 12112 5782
rect 12032 5324 12112 5352
rect 11980 5306 12032 5312
rect 11978 5264 12034 5273
rect 11978 5199 11980 5208
rect 12032 5199 12034 5208
rect 12072 5228 12124 5234
rect 11980 5170 12032 5176
rect 12072 5170 12124 5176
rect 11888 4480 11940 4486
rect 11888 4422 11940 4428
rect 11900 4282 11928 4422
rect 11888 4276 11940 4282
rect 11888 4218 11940 4224
rect 11980 4072 12032 4078
rect 11980 4014 12032 4020
rect 11428 3936 11480 3942
rect 11428 3878 11480 3884
rect 11334 3632 11390 3641
rect 11334 3567 11336 3576
rect 11388 3567 11390 3576
rect 11336 3538 11388 3544
rect 11244 3392 11296 3398
rect 11242 3360 11244 3369
rect 11336 3392 11388 3398
rect 11296 3360 11298 3369
rect 11440 3380 11468 3878
rect 11992 3738 12020 4014
rect 11980 3732 12032 3738
rect 11980 3674 12032 3680
rect 11388 3352 11468 3380
rect 11980 3392 12032 3398
rect 11336 3334 11388 3340
rect 11980 3334 12032 3340
rect 11242 3295 11298 3304
rect 11060 3120 11112 3126
rect 11060 3062 11112 3068
rect 11072 2990 11100 3062
rect 10612 2944 10916 2972
rect 11060 2984 11112 2990
rect 10048 2926 10100 2932
rect 11060 2926 11112 2932
rect 11244 2916 11296 2922
rect 11244 2858 11296 2864
rect 11256 2650 11284 2858
rect 11152 2644 11204 2650
rect 11152 2586 11204 2592
rect 11244 2644 11296 2650
rect 11244 2586 11296 2592
rect 11164 2446 11192 2586
rect 11152 2440 11204 2446
rect 10322 2408 10378 2417
rect 11348 2417 11376 3334
rect 11428 2916 11480 2922
rect 11428 2858 11480 2864
rect 11440 2774 11468 2858
rect 11440 2746 11836 2774
rect 11808 2514 11836 2746
rect 11796 2508 11848 2514
rect 11796 2450 11848 2456
rect 11152 2382 11204 2388
rect 11334 2408 11390 2417
rect 10322 2343 10324 2352
rect 10376 2343 10378 2352
rect 11334 2343 11390 2352
rect 10324 2314 10376 2320
rect 9456 2252 9904 2258
rect 9404 2246 9904 2252
rect 9416 2230 9904 2246
rect 5547 2204 5855 2224
rect 5547 2202 5553 2204
rect 5609 2202 5633 2204
rect 5689 2202 5713 2204
rect 5769 2202 5793 2204
rect 5849 2202 5855 2204
rect 5609 2150 5611 2202
rect 5791 2150 5793 2202
rect 5547 2148 5553 2150
rect 5609 2148 5633 2150
rect 5689 2148 5713 2150
rect 5769 2148 5793 2150
rect 5849 2148 5855 2150
rect 5547 2128 5855 2148
rect 10144 2204 10452 2224
rect 10144 2202 10150 2204
rect 10206 2202 10230 2204
rect 10286 2202 10310 2204
rect 10366 2202 10390 2204
rect 10446 2202 10452 2204
rect 10206 2150 10208 2202
rect 10388 2150 10390 2202
rect 10144 2148 10150 2150
rect 10206 2148 10230 2150
rect 10286 2148 10310 2150
rect 10366 2148 10390 2150
rect 10446 2148 10452 2150
rect 10144 2128 10452 2148
rect 11992 800 12020 3334
rect 12084 3097 12112 5170
rect 12176 5166 12204 6122
rect 12443 6012 12751 6032
rect 12443 6010 12449 6012
rect 12505 6010 12529 6012
rect 12585 6010 12609 6012
rect 12665 6010 12689 6012
rect 12745 6010 12751 6012
rect 12505 5958 12507 6010
rect 12687 5958 12689 6010
rect 12443 5956 12449 5958
rect 12505 5956 12529 5958
rect 12585 5956 12609 5958
rect 12665 5956 12689 5958
rect 12745 5956 12751 5958
rect 12443 5936 12751 5956
rect 12624 5840 12676 5846
rect 12624 5782 12676 5788
rect 12636 5234 12664 5782
rect 12440 5228 12492 5234
rect 12360 5188 12440 5216
rect 12164 5160 12216 5166
rect 12164 5102 12216 5108
rect 12360 4826 12388 5188
rect 12440 5170 12492 5176
rect 12624 5228 12676 5234
rect 12624 5170 12676 5176
rect 12443 4924 12751 4944
rect 12443 4922 12449 4924
rect 12505 4922 12529 4924
rect 12585 4922 12609 4924
rect 12665 4922 12689 4924
rect 12745 4922 12751 4924
rect 12505 4870 12507 4922
rect 12687 4870 12689 4922
rect 12443 4868 12449 4870
rect 12505 4868 12529 4870
rect 12585 4868 12609 4870
rect 12665 4868 12689 4870
rect 12745 4868 12751 4870
rect 12443 4848 12751 4868
rect 12348 4820 12400 4826
rect 12348 4762 12400 4768
rect 12348 4208 12400 4214
rect 12348 4150 12400 4156
rect 12360 3942 12388 4150
rect 12348 3936 12400 3942
rect 12348 3878 12400 3884
rect 12360 3466 12388 3878
rect 12443 3836 12751 3856
rect 12443 3834 12449 3836
rect 12505 3834 12529 3836
rect 12585 3834 12609 3836
rect 12665 3834 12689 3836
rect 12745 3834 12751 3836
rect 12505 3782 12507 3834
rect 12687 3782 12689 3834
rect 12443 3780 12449 3782
rect 12505 3780 12529 3782
rect 12585 3780 12609 3782
rect 12665 3780 12689 3782
rect 12745 3780 12751 3782
rect 12443 3760 12751 3780
rect 12348 3460 12400 3466
rect 12348 3402 12400 3408
rect 12070 3088 12126 3097
rect 12070 3023 12126 3032
rect 12360 2360 12388 3402
rect 12820 3398 12848 9522
rect 12912 9518 12940 10066
rect 12900 9512 12952 9518
rect 12900 9454 12952 9460
rect 12912 9178 12940 9454
rect 12900 9172 12952 9178
rect 12900 9114 12952 9120
rect 13280 7546 13308 13466
rect 14188 13320 14240 13326
rect 14188 13262 14240 13268
rect 14096 13184 14148 13190
rect 14096 13126 14148 13132
rect 14108 12850 14136 13126
rect 14200 12986 14228 13262
rect 14188 12980 14240 12986
rect 14188 12922 14240 12928
rect 13820 12844 13872 12850
rect 13820 12786 13872 12792
rect 14096 12844 14148 12850
rect 14096 12786 14148 12792
rect 14280 12844 14332 12850
rect 14280 12786 14332 12792
rect 13636 12776 13688 12782
rect 13636 12718 13688 12724
rect 13452 12708 13504 12714
rect 13452 12650 13504 12656
rect 13360 11824 13412 11830
rect 13360 11766 13412 11772
rect 13372 11082 13400 11766
rect 13360 11076 13412 11082
rect 13360 11018 13412 11024
rect 13372 10742 13400 11018
rect 13360 10736 13412 10742
rect 13360 10678 13412 10684
rect 13372 10266 13400 10678
rect 13360 10260 13412 10266
rect 13360 10202 13412 10208
rect 13372 8906 13400 10202
rect 13464 10062 13492 12650
rect 13648 12442 13676 12718
rect 13636 12436 13688 12442
rect 13636 12378 13688 12384
rect 13832 11150 13860 12786
rect 14292 12442 14320 12786
rect 14280 12436 14332 12442
rect 14280 12378 14332 12384
rect 14280 12164 14332 12170
rect 14280 12106 14332 12112
rect 14292 11898 14320 12106
rect 14280 11892 14332 11898
rect 14280 11834 14332 11840
rect 13820 11144 13872 11150
rect 13820 11086 13872 11092
rect 13832 10810 13860 11086
rect 14096 11008 14148 11014
rect 14096 10950 14148 10956
rect 15014 10976 15070 10985
rect 13820 10804 13872 10810
rect 13820 10746 13872 10752
rect 14108 10674 14136 10950
rect 15014 10911 15070 10920
rect 15028 10878 15056 10911
rect 15016 10872 15068 10878
rect 15016 10814 15068 10820
rect 14096 10668 14148 10674
rect 14096 10610 14148 10616
rect 13452 10056 13504 10062
rect 13452 9998 13504 10004
rect 13728 9988 13780 9994
rect 13728 9930 13780 9936
rect 14004 9988 14056 9994
rect 14004 9930 14056 9936
rect 13636 9920 13688 9926
rect 13636 9862 13688 9868
rect 13360 8900 13412 8906
rect 13360 8842 13412 8848
rect 13544 8900 13596 8906
rect 13544 8842 13596 8848
rect 13372 8548 13400 8842
rect 13452 8560 13504 8566
rect 13372 8520 13452 8548
rect 13452 8502 13504 8508
rect 13464 7750 13492 8502
rect 13556 8430 13584 8842
rect 13544 8424 13596 8430
rect 13544 8366 13596 8372
rect 13452 7744 13504 7750
rect 13452 7686 13504 7692
rect 13268 7540 13320 7546
rect 13268 7482 13320 7488
rect 13360 7404 13412 7410
rect 13360 7346 13412 7352
rect 13372 6254 13400 7346
rect 13648 6866 13676 9862
rect 13740 9450 13768 9930
rect 13728 9444 13780 9450
rect 13728 9386 13780 9392
rect 13740 7546 13768 9386
rect 14016 9382 14044 9930
rect 14280 9920 14332 9926
rect 14280 9862 14332 9868
rect 14292 9654 14320 9862
rect 14280 9648 14332 9654
rect 14280 9590 14332 9596
rect 14004 9376 14056 9382
rect 14004 9318 14056 9324
rect 14016 8634 14044 9318
rect 15014 9072 15070 9081
rect 15014 9007 15016 9016
rect 15068 9007 15070 9016
rect 15016 8978 15068 8984
rect 14004 8628 14056 8634
rect 14004 8570 14056 8576
rect 14188 8424 14240 8430
rect 14188 8366 14240 8372
rect 14200 8090 14228 8366
rect 14188 8084 14240 8090
rect 14188 8026 14240 8032
rect 14096 7744 14148 7750
rect 14096 7686 14148 7692
rect 13728 7540 13780 7546
rect 13728 7482 13780 7488
rect 13636 6860 13688 6866
rect 13636 6802 13688 6808
rect 13544 6724 13596 6730
rect 13544 6666 13596 6672
rect 13360 6248 13412 6254
rect 13360 6190 13412 6196
rect 13360 6112 13412 6118
rect 13360 6054 13412 6060
rect 13372 5574 13400 6054
rect 13556 5914 13584 6666
rect 13544 5908 13596 5914
rect 13544 5850 13596 5856
rect 13648 5778 13676 6802
rect 14108 6662 14136 7686
rect 14462 7032 14518 7041
rect 14462 6967 14518 6976
rect 14476 6934 14504 6967
rect 14464 6928 14516 6934
rect 14464 6870 14516 6876
rect 14096 6656 14148 6662
rect 14096 6598 14148 6604
rect 13636 5772 13688 5778
rect 13636 5714 13688 5720
rect 13360 5568 13412 5574
rect 13360 5510 13412 5516
rect 13372 5302 13400 5510
rect 13360 5296 13412 5302
rect 13360 5238 13412 5244
rect 12900 5024 12952 5030
rect 12900 4966 12952 4972
rect 12912 4078 12940 4966
rect 13648 4690 13676 5714
rect 14108 5574 14136 6598
rect 14464 6180 14516 6186
rect 14464 6122 14516 6128
rect 14476 5710 14504 6122
rect 14464 5704 14516 5710
rect 14464 5646 14516 5652
rect 14096 5568 14148 5574
rect 14096 5510 14148 5516
rect 14188 5568 14240 5574
rect 14188 5510 14240 5516
rect 13818 5264 13874 5273
rect 13818 5199 13820 5208
rect 13872 5199 13874 5208
rect 13820 5170 13872 5176
rect 14108 4826 14136 5510
rect 14096 4820 14148 4826
rect 14096 4762 14148 4768
rect 13636 4684 13688 4690
rect 13636 4626 13688 4632
rect 13544 4616 13596 4622
rect 14200 4570 14228 5510
rect 14476 5001 14504 5646
rect 14462 4992 14518 5001
rect 14462 4927 14518 4936
rect 14372 4684 14424 4690
rect 14372 4626 14424 4632
rect 13544 4558 13596 4564
rect 13556 4282 13584 4558
rect 14108 4542 14228 4570
rect 13544 4276 13596 4282
rect 13544 4218 13596 4224
rect 14108 4146 14136 4542
rect 14188 4480 14240 4486
rect 14188 4422 14240 4428
rect 14096 4140 14148 4146
rect 14096 4082 14148 4088
rect 12900 4072 12952 4078
rect 12900 4014 12952 4020
rect 12912 3602 12940 4014
rect 12900 3596 12952 3602
rect 12900 3538 12952 3544
rect 13360 3460 13412 3466
rect 13360 3402 13412 3408
rect 12808 3392 12860 3398
rect 12808 3334 12860 3340
rect 12900 3392 12952 3398
rect 12900 3334 12952 3340
rect 12912 3210 12940 3334
rect 12728 3182 12940 3210
rect 13372 3194 13400 3402
rect 13360 3188 13412 3194
rect 12728 3058 12756 3182
rect 13360 3130 13412 3136
rect 14200 3126 14228 4422
rect 14384 4146 14412 4626
rect 14464 4616 14516 4622
rect 14464 4558 14516 4564
rect 14372 4140 14424 4146
rect 14372 4082 14424 4088
rect 14384 3602 14412 4082
rect 14372 3596 14424 3602
rect 14372 3538 14424 3544
rect 14188 3120 14240 3126
rect 14188 3062 14240 3068
rect 14384 3058 14412 3538
rect 14476 3398 14504 4558
rect 14464 3392 14516 3398
rect 14464 3334 14516 3340
rect 12716 3052 12768 3058
rect 12992 3052 13044 3058
rect 12716 2994 12768 3000
rect 12912 3012 12992 3040
rect 12443 2748 12751 2768
rect 12443 2746 12449 2748
rect 12505 2746 12529 2748
rect 12585 2746 12609 2748
rect 12665 2746 12689 2748
rect 12745 2746 12751 2748
rect 12505 2694 12507 2746
rect 12687 2694 12689 2746
rect 12443 2692 12449 2694
rect 12505 2692 12529 2694
rect 12585 2692 12609 2694
rect 12665 2692 12689 2694
rect 12745 2692 12751 2694
rect 12443 2672 12751 2692
rect 12912 2514 12940 3012
rect 12992 2994 13044 3000
rect 14372 3052 14424 3058
rect 14372 2994 14424 3000
rect 14096 2984 14148 2990
rect 14476 2961 14504 3334
rect 14096 2926 14148 2932
rect 14462 2952 14518 2961
rect 12900 2508 12952 2514
rect 12900 2450 12952 2456
rect 12912 2378 12940 2450
rect 14108 2446 14136 2926
rect 14462 2887 14518 2896
rect 14096 2440 14148 2446
rect 14096 2382 14148 2388
rect 12532 2372 12584 2378
rect 12360 2332 12532 2360
rect 12532 2314 12584 2320
rect 12900 2372 12952 2378
rect 12900 2314 12952 2320
rect 14924 1080 14976 1086
rect 14922 1048 14924 1057
rect 14976 1048 14978 1057
rect 14922 983 14978 992
rect 3974 0 4030 800
rect 11978 0 12034 800
<< via2 >>
rect 3254 13626 3310 13628
rect 3334 13626 3390 13628
rect 3414 13626 3470 13628
rect 3494 13626 3550 13628
rect 3254 13574 3300 13626
rect 3300 13574 3310 13626
rect 3334 13574 3364 13626
rect 3364 13574 3376 13626
rect 3376 13574 3390 13626
rect 3414 13574 3428 13626
rect 3428 13574 3440 13626
rect 3440 13574 3470 13626
rect 3494 13574 3504 13626
rect 3504 13574 3550 13626
rect 3254 13572 3310 13574
rect 3334 13572 3390 13574
rect 3414 13572 3470 13574
rect 3494 13572 3550 13574
rect 7852 13626 7908 13628
rect 7932 13626 7988 13628
rect 8012 13626 8068 13628
rect 8092 13626 8148 13628
rect 7852 13574 7898 13626
rect 7898 13574 7908 13626
rect 7932 13574 7962 13626
rect 7962 13574 7974 13626
rect 7974 13574 7988 13626
rect 8012 13574 8026 13626
rect 8026 13574 8038 13626
rect 8038 13574 8068 13626
rect 8092 13574 8102 13626
rect 8102 13574 8148 13626
rect 7852 13572 7908 13574
rect 7932 13572 7988 13574
rect 8012 13572 8068 13574
rect 8092 13572 8148 13574
rect 12449 13626 12505 13628
rect 12529 13626 12585 13628
rect 12609 13626 12665 13628
rect 12689 13626 12745 13628
rect 12449 13574 12495 13626
rect 12495 13574 12505 13626
rect 12529 13574 12559 13626
rect 12559 13574 12571 13626
rect 12571 13574 12585 13626
rect 12609 13574 12623 13626
rect 12623 13574 12635 13626
rect 12635 13574 12665 13626
rect 12689 13574 12699 13626
rect 12699 13574 12745 13626
rect 12449 13572 12505 13574
rect 12529 13572 12585 13574
rect 12609 13572 12665 13574
rect 12689 13572 12745 13574
rect 14922 15020 14978 15056
rect 14922 15000 14924 15020
rect 14924 15000 14976 15020
rect 14976 15000 14978 15020
rect 3254 12538 3310 12540
rect 3334 12538 3390 12540
rect 3414 12538 3470 12540
rect 3494 12538 3550 12540
rect 3254 12486 3300 12538
rect 3300 12486 3310 12538
rect 3334 12486 3364 12538
rect 3364 12486 3376 12538
rect 3376 12486 3390 12538
rect 3414 12486 3428 12538
rect 3428 12486 3440 12538
rect 3440 12486 3470 12538
rect 3494 12486 3504 12538
rect 3504 12486 3550 12538
rect 3254 12484 3310 12486
rect 3334 12484 3390 12486
rect 3414 12484 3470 12486
rect 3494 12484 3550 12486
rect 3254 11450 3310 11452
rect 3334 11450 3390 11452
rect 3414 11450 3470 11452
rect 3494 11450 3550 11452
rect 3254 11398 3300 11450
rect 3300 11398 3310 11450
rect 3334 11398 3364 11450
rect 3364 11398 3376 11450
rect 3376 11398 3390 11450
rect 3414 11398 3428 11450
rect 3428 11398 3440 11450
rect 3440 11398 3470 11450
rect 3494 11398 3504 11450
rect 3504 11398 3550 11450
rect 3254 11396 3310 11398
rect 3334 11396 3390 11398
rect 3414 11396 3470 11398
rect 3494 11396 3550 11398
rect 4158 12008 4214 12064
rect 3254 10362 3310 10364
rect 3334 10362 3390 10364
rect 3414 10362 3470 10364
rect 3494 10362 3550 10364
rect 3254 10310 3300 10362
rect 3300 10310 3310 10362
rect 3334 10310 3364 10362
rect 3364 10310 3376 10362
rect 3376 10310 3390 10362
rect 3414 10310 3428 10362
rect 3428 10310 3440 10362
rect 3440 10310 3470 10362
rect 3494 10310 3504 10362
rect 3504 10310 3550 10362
rect 3254 10308 3310 10310
rect 3334 10308 3390 10310
rect 3414 10308 3470 10310
rect 3494 10308 3550 10310
rect 3054 9968 3110 10024
rect 2962 9832 3018 9888
rect 3514 9868 3516 9888
rect 3516 9868 3568 9888
rect 3568 9868 3570 9888
rect 3514 9832 3570 9868
rect 3254 9274 3310 9276
rect 3334 9274 3390 9276
rect 3414 9274 3470 9276
rect 3494 9274 3550 9276
rect 3254 9222 3300 9274
rect 3300 9222 3310 9274
rect 3334 9222 3364 9274
rect 3364 9222 3376 9274
rect 3376 9222 3390 9274
rect 3414 9222 3428 9274
rect 3428 9222 3440 9274
rect 3440 9222 3470 9274
rect 3494 9222 3504 9274
rect 3504 9222 3550 9274
rect 3254 9220 3310 9222
rect 3334 9220 3390 9222
rect 3414 9220 3470 9222
rect 3494 9220 3550 9222
rect 5553 13082 5609 13084
rect 5633 13082 5689 13084
rect 5713 13082 5769 13084
rect 5793 13082 5849 13084
rect 5553 13030 5599 13082
rect 5599 13030 5609 13082
rect 5633 13030 5663 13082
rect 5663 13030 5675 13082
rect 5675 13030 5689 13082
rect 5713 13030 5727 13082
rect 5727 13030 5739 13082
rect 5739 13030 5769 13082
rect 5793 13030 5803 13082
rect 5803 13030 5849 13082
rect 5553 13028 5609 13030
rect 5633 13028 5689 13030
rect 5713 13028 5769 13030
rect 5793 13028 5849 13030
rect 5553 11994 5609 11996
rect 5633 11994 5689 11996
rect 5713 11994 5769 11996
rect 5793 11994 5849 11996
rect 5553 11942 5599 11994
rect 5599 11942 5609 11994
rect 5633 11942 5663 11994
rect 5663 11942 5675 11994
rect 5675 11942 5689 11994
rect 5713 11942 5727 11994
rect 5727 11942 5739 11994
rect 5739 11942 5769 11994
rect 5793 11942 5803 11994
rect 5803 11942 5849 11994
rect 5553 11940 5609 11942
rect 5633 11940 5689 11942
rect 5713 11940 5769 11942
rect 5793 11940 5849 11942
rect 4526 10004 4528 10024
rect 4528 10004 4580 10024
rect 4580 10004 4582 10024
rect 4526 9968 4582 10004
rect 5538 11076 5594 11112
rect 5538 11056 5540 11076
rect 5540 11056 5592 11076
rect 5592 11056 5594 11076
rect 5553 10906 5609 10908
rect 5633 10906 5689 10908
rect 5713 10906 5769 10908
rect 5793 10906 5849 10908
rect 5553 10854 5599 10906
rect 5599 10854 5609 10906
rect 5633 10854 5663 10906
rect 5663 10854 5675 10906
rect 5675 10854 5689 10906
rect 5713 10854 5727 10906
rect 5727 10854 5739 10906
rect 5739 10854 5769 10906
rect 5793 10854 5803 10906
rect 5803 10854 5849 10906
rect 5553 10852 5609 10854
rect 5633 10852 5689 10854
rect 5713 10852 5769 10854
rect 5793 10852 5849 10854
rect 5553 9818 5609 9820
rect 5633 9818 5689 9820
rect 5713 9818 5769 9820
rect 5793 9818 5849 9820
rect 5553 9766 5599 9818
rect 5599 9766 5609 9818
rect 5633 9766 5663 9818
rect 5663 9766 5675 9818
rect 5675 9766 5689 9818
rect 5713 9766 5727 9818
rect 5727 9766 5739 9818
rect 5739 9766 5769 9818
rect 5793 9766 5803 9818
rect 5803 9766 5849 9818
rect 5553 9764 5609 9766
rect 5633 9764 5689 9766
rect 5713 9764 5769 9766
rect 5793 9764 5849 9766
rect 7852 12538 7908 12540
rect 7932 12538 7988 12540
rect 8012 12538 8068 12540
rect 8092 12538 8148 12540
rect 7852 12486 7898 12538
rect 7898 12486 7908 12538
rect 7932 12486 7962 12538
rect 7962 12486 7974 12538
rect 7974 12486 7988 12538
rect 8012 12486 8026 12538
rect 8026 12486 8038 12538
rect 8038 12486 8068 12538
rect 8092 12486 8102 12538
rect 8102 12486 8148 12538
rect 7852 12484 7908 12486
rect 7932 12484 7988 12486
rect 8012 12484 8068 12486
rect 8092 12484 8148 12486
rect 10150 13082 10206 13084
rect 10230 13082 10286 13084
rect 10310 13082 10366 13084
rect 10390 13082 10446 13084
rect 10150 13030 10196 13082
rect 10196 13030 10206 13082
rect 10230 13030 10260 13082
rect 10260 13030 10272 13082
rect 10272 13030 10286 13082
rect 10310 13030 10324 13082
rect 10324 13030 10336 13082
rect 10336 13030 10366 13082
rect 10390 13030 10400 13082
rect 10400 13030 10446 13082
rect 10150 13028 10206 13030
rect 10230 13028 10286 13030
rect 10310 13028 10366 13030
rect 10390 13028 10446 13030
rect 7838 11736 7894 11792
rect 9218 11756 9274 11792
rect 9218 11736 9220 11756
rect 9220 11736 9272 11756
rect 9272 11736 9274 11756
rect 7852 11450 7908 11452
rect 7932 11450 7988 11452
rect 8012 11450 8068 11452
rect 8092 11450 8148 11452
rect 7852 11398 7898 11450
rect 7898 11398 7908 11450
rect 7932 11398 7962 11450
rect 7962 11398 7974 11450
rect 7974 11398 7988 11450
rect 8012 11398 8026 11450
rect 8026 11398 8038 11450
rect 8038 11398 8068 11450
rect 8092 11398 8102 11450
rect 8102 11398 8148 11450
rect 7852 11396 7908 11398
rect 7932 11396 7988 11398
rect 8012 11396 8068 11398
rect 8092 11396 8148 11398
rect 7286 11056 7342 11112
rect 8206 11056 8262 11112
rect 3254 8186 3310 8188
rect 3334 8186 3390 8188
rect 3414 8186 3470 8188
rect 3494 8186 3550 8188
rect 3254 8134 3300 8186
rect 3300 8134 3310 8186
rect 3334 8134 3364 8186
rect 3364 8134 3376 8186
rect 3376 8134 3390 8186
rect 3414 8134 3428 8186
rect 3428 8134 3440 8186
rect 3440 8134 3470 8186
rect 3494 8134 3504 8186
rect 3504 8134 3550 8186
rect 3254 8132 3310 8134
rect 3334 8132 3390 8134
rect 3414 8132 3470 8134
rect 3494 8132 3550 8134
rect 7852 10362 7908 10364
rect 7932 10362 7988 10364
rect 8012 10362 8068 10364
rect 8092 10362 8148 10364
rect 7852 10310 7898 10362
rect 7898 10310 7908 10362
rect 7932 10310 7962 10362
rect 7962 10310 7974 10362
rect 7974 10310 7988 10362
rect 8012 10310 8026 10362
rect 8026 10310 8038 10362
rect 8038 10310 8068 10362
rect 8092 10310 8102 10362
rect 8102 10310 8148 10362
rect 7852 10308 7908 10310
rect 7932 10308 7988 10310
rect 8012 10308 8068 10310
rect 8092 10308 8148 10310
rect 5553 8730 5609 8732
rect 5633 8730 5689 8732
rect 5713 8730 5769 8732
rect 5793 8730 5849 8732
rect 5553 8678 5599 8730
rect 5599 8678 5609 8730
rect 5633 8678 5663 8730
rect 5663 8678 5675 8730
rect 5675 8678 5689 8730
rect 5713 8678 5727 8730
rect 5727 8678 5739 8730
rect 5739 8678 5769 8730
rect 5793 8678 5803 8730
rect 5803 8678 5849 8730
rect 5553 8676 5609 8678
rect 5633 8676 5689 8678
rect 5713 8676 5769 8678
rect 5793 8676 5849 8678
rect 7852 9274 7908 9276
rect 7932 9274 7988 9276
rect 8012 9274 8068 9276
rect 8092 9274 8148 9276
rect 7852 9222 7898 9274
rect 7898 9222 7908 9274
rect 7932 9222 7962 9274
rect 7962 9222 7974 9274
rect 7974 9222 7988 9274
rect 8012 9222 8026 9274
rect 8026 9222 8038 9274
rect 8038 9222 8068 9274
rect 8092 9222 8102 9274
rect 8102 9222 8148 9274
rect 7852 9220 7908 9222
rect 7932 9220 7988 9222
rect 8012 9220 8068 9222
rect 8092 9220 8148 9222
rect 5553 7642 5609 7644
rect 5633 7642 5689 7644
rect 5713 7642 5769 7644
rect 5793 7642 5849 7644
rect 5553 7590 5599 7642
rect 5599 7590 5609 7642
rect 5633 7590 5663 7642
rect 5663 7590 5675 7642
rect 5675 7590 5689 7642
rect 5713 7590 5727 7642
rect 5727 7590 5739 7642
rect 5739 7590 5769 7642
rect 5793 7590 5803 7642
rect 5803 7590 5849 7642
rect 5553 7588 5609 7590
rect 5633 7588 5689 7590
rect 5713 7588 5769 7590
rect 5793 7588 5849 7590
rect 3254 7098 3310 7100
rect 3334 7098 3390 7100
rect 3414 7098 3470 7100
rect 3494 7098 3550 7100
rect 3254 7046 3300 7098
rect 3300 7046 3310 7098
rect 3334 7046 3364 7098
rect 3364 7046 3376 7098
rect 3376 7046 3390 7098
rect 3414 7046 3428 7098
rect 3428 7046 3440 7098
rect 3440 7046 3470 7098
rect 3494 7046 3504 7098
rect 3504 7046 3550 7098
rect 3254 7044 3310 7046
rect 3334 7044 3390 7046
rect 3414 7044 3470 7046
rect 3494 7044 3550 7046
rect 8574 9968 8630 10024
rect 9034 11192 9090 11248
rect 9034 11056 9090 11112
rect 10150 11994 10206 11996
rect 10230 11994 10286 11996
rect 10310 11994 10366 11996
rect 10390 11994 10446 11996
rect 10150 11942 10196 11994
rect 10196 11942 10206 11994
rect 10230 11942 10260 11994
rect 10260 11942 10272 11994
rect 10272 11942 10286 11994
rect 10310 11942 10324 11994
rect 10324 11942 10336 11994
rect 10336 11942 10366 11994
rect 10390 11942 10400 11994
rect 10400 11942 10446 11994
rect 10150 11940 10206 11942
rect 10230 11940 10286 11942
rect 10310 11940 10366 11942
rect 10390 11940 10446 11942
rect 11334 12960 11390 13016
rect 10138 11076 10194 11112
rect 10138 11056 10140 11076
rect 10140 11056 10192 11076
rect 10192 11056 10194 11076
rect 10690 11056 10746 11112
rect 10150 10906 10206 10908
rect 10230 10906 10286 10908
rect 10310 10906 10366 10908
rect 10390 10906 10446 10908
rect 10150 10854 10196 10906
rect 10196 10854 10206 10906
rect 10230 10854 10260 10906
rect 10260 10854 10272 10906
rect 10272 10854 10286 10906
rect 10310 10854 10324 10906
rect 10324 10854 10336 10906
rect 10336 10854 10366 10906
rect 10390 10854 10400 10906
rect 10400 10854 10446 10906
rect 10150 10852 10206 10854
rect 10230 10852 10286 10854
rect 10310 10852 10366 10854
rect 10390 10852 10446 10854
rect 10150 9818 10206 9820
rect 10230 9818 10286 9820
rect 10310 9818 10366 9820
rect 10390 9818 10446 9820
rect 10150 9766 10196 9818
rect 10196 9766 10206 9818
rect 10230 9766 10260 9818
rect 10260 9766 10272 9818
rect 10272 9766 10286 9818
rect 10310 9766 10324 9818
rect 10324 9766 10336 9818
rect 10336 9766 10366 9818
rect 10390 9766 10400 9818
rect 10400 9766 10446 9818
rect 10150 9764 10206 9766
rect 10230 9764 10286 9766
rect 10310 9764 10366 9766
rect 10390 9764 10446 9766
rect 12449 12538 12505 12540
rect 12529 12538 12585 12540
rect 12609 12538 12665 12540
rect 12689 12538 12745 12540
rect 12449 12486 12495 12538
rect 12495 12486 12505 12538
rect 12529 12486 12559 12538
rect 12559 12486 12571 12538
rect 12571 12486 12585 12538
rect 12609 12486 12623 12538
rect 12623 12486 12635 12538
rect 12635 12486 12665 12538
rect 12689 12486 12699 12538
rect 12699 12486 12745 12538
rect 12449 12484 12505 12486
rect 12529 12484 12585 12486
rect 12609 12484 12665 12486
rect 12689 12484 12745 12486
rect 11058 10004 11060 10024
rect 11060 10004 11112 10024
rect 11112 10004 11114 10024
rect 11058 9968 11114 10004
rect 7852 8186 7908 8188
rect 7932 8186 7988 8188
rect 8012 8186 8068 8188
rect 8092 8186 8148 8188
rect 7852 8134 7898 8186
rect 7898 8134 7908 8186
rect 7932 8134 7962 8186
rect 7962 8134 7974 8186
rect 7974 8134 7988 8186
rect 8012 8134 8026 8186
rect 8026 8134 8038 8186
rect 8038 8134 8068 8186
rect 8092 8134 8102 8186
rect 8102 8134 8148 8186
rect 7852 8132 7908 8134
rect 7932 8132 7988 8134
rect 8012 8132 8068 8134
rect 8092 8132 8148 8134
rect 2502 5480 2558 5536
rect 3254 6010 3310 6012
rect 3334 6010 3390 6012
rect 3414 6010 3470 6012
rect 3494 6010 3550 6012
rect 3254 5958 3300 6010
rect 3300 5958 3310 6010
rect 3334 5958 3364 6010
rect 3364 5958 3376 6010
rect 3376 5958 3390 6010
rect 3414 5958 3428 6010
rect 3428 5958 3440 6010
rect 3440 5958 3470 6010
rect 3494 5958 3504 6010
rect 3504 5958 3550 6010
rect 3254 5956 3310 5958
rect 3334 5956 3390 5958
rect 3414 5956 3470 5958
rect 3494 5956 3550 5958
rect 4618 5480 4674 5536
rect 3254 4922 3310 4924
rect 3334 4922 3390 4924
rect 3414 4922 3470 4924
rect 3494 4922 3550 4924
rect 3254 4870 3300 4922
rect 3300 4870 3310 4922
rect 3334 4870 3364 4922
rect 3364 4870 3376 4922
rect 3376 4870 3390 4922
rect 3414 4870 3428 4922
rect 3428 4870 3440 4922
rect 3440 4870 3470 4922
rect 3494 4870 3504 4922
rect 3504 4870 3550 4922
rect 3254 4868 3310 4870
rect 3334 4868 3390 4870
rect 3414 4868 3470 4870
rect 3494 4868 3550 4870
rect 4342 4664 4398 4720
rect 5553 6554 5609 6556
rect 5633 6554 5689 6556
rect 5713 6554 5769 6556
rect 5793 6554 5849 6556
rect 5553 6502 5599 6554
rect 5599 6502 5609 6554
rect 5633 6502 5663 6554
rect 5663 6502 5675 6554
rect 5675 6502 5689 6554
rect 5713 6502 5727 6554
rect 5727 6502 5739 6554
rect 5739 6502 5769 6554
rect 5793 6502 5803 6554
rect 5803 6502 5849 6554
rect 5553 6500 5609 6502
rect 5633 6500 5689 6502
rect 5713 6500 5769 6502
rect 5793 6500 5849 6502
rect 3254 3834 3310 3836
rect 3334 3834 3390 3836
rect 3414 3834 3470 3836
rect 3494 3834 3550 3836
rect 3254 3782 3300 3834
rect 3300 3782 3310 3834
rect 3334 3782 3364 3834
rect 3364 3782 3376 3834
rect 3376 3782 3390 3834
rect 3414 3782 3428 3834
rect 3428 3782 3440 3834
rect 3440 3782 3470 3834
rect 3494 3782 3504 3834
rect 3504 3782 3550 3834
rect 3254 3780 3310 3782
rect 3334 3780 3390 3782
rect 3414 3780 3470 3782
rect 3494 3780 3550 3782
rect 3790 3576 3846 3632
rect 4158 3848 4214 3904
rect 3422 3476 3424 3496
rect 3424 3476 3476 3496
rect 3476 3476 3478 3496
rect 3422 3440 3478 3476
rect 3254 2746 3310 2748
rect 3334 2746 3390 2748
rect 3414 2746 3470 2748
rect 3494 2746 3550 2748
rect 3254 2694 3300 2746
rect 3300 2694 3310 2746
rect 3334 2694 3364 2746
rect 3364 2694 3376 2746
rect 3376 2694 3390 2746
rect 3414 2694 3428 2746
rect 3428 2694 3440 2746
rect 3440 2694 3470 2746
rect 3494 2694 3504 2746
rect 3504 2694 3550 2746
rect 3254 2692 3310 2694
rect 3334 2692 3390 2694
rect 3414 2692 3470 2694
rect 3494 2692 3550 2694
rect 4526 4120 4582 4176
rect 4526 4004 4582 4040
rect 4526 3984 4528 4004
rect 4528 3984 4580 4004
rect 4580 3984 4582 4004
rect 5553 5466 5609 5468
rect 5633 5466 5689 5468
rect 5713 5466 5769 5468
rect 5793 5466 5849 5468
rect 5553 5414 5599 5466
rect 5599 5414 5609 5466
rect 5633 5414 5663 5466
rect 5663 5414 5675 5466
rect 5675 5414 5689 5466
rect 5713 5414 5727 5466
rect 5727 5414 5739 5466
rect 5739 5414 5769 5466
rect 5793 5414 5803 5466
rect 5803 5414 5849 5466
rect 5553 5412 5609 5414
rect 5633 5412 5689 5414
rect 5713 5412 5769 5414
rect 5793 5412 5849 5414
rect 5722 5208 5778 5264
rect 5553 4378 5609 4380
rect 5633 4378 5689 4380
rect 5713 4378 5769 4380
rect 5793 4378 5849 4380
rect 5553 4326 5599 4378
rect 5599 4326 5609 4378
rect 5633 4326 5663 4378
rect 5663 4326 5675 4378
rect 5675 4326 5689 4378
rect 5713 4326 5727 4378
rect 5727 4326 5739 4378
rect 5739 4326 5769 4378
rect 5793 4326 5803 4378
rect 5803 4326 5849 4378
rect 5553 4324 5609 4326
rect 5633 4324 5689 4326
rect 5713 4324 5769 4326
rect 5793 4324 5849 4326
rect 5538 4120 5594 4176
rect 5538 3848 5594 3904
rect 5262 3596 5318 3632
rect 5262 3576 5264 3596
rect 5264 3576 5316 3596
rect 5316 3576 5318 3596
rect 5170 3460 5226 3496
rect 5170 3440 5172 3460
rect 5172 3440 5224 3460
rect 5224 3440 5226 3460
rect 5553 3290 5609 3292
rect 5633 3290 5689 3292
rect 5713 3290 5769 3292
rect 5793 3290 5849 3292
rect 5553 3238 5599 3290
rect 5599 3238 5609 3290
rect 5633 3238 5663 3290
rect 5663 3238 5675 3290
rect 5675 3238 5689 3290
rect 5713 3238 5727 3290
rect 5727 3238 5739 3290
rect 5739 3238 5769 3290
rect 5793 3238 5803 3290
rect 5803 3238 5849 3290
rect 5553 3236 5609 3238
rect 5633 3236 5689 3238
rect 5713 3236 5769 3238
rect 5793 3236 5849 3238
rect 7852 7098 7908 7100
rect 7932 7098 7988 7100
rect 8012 7098 8068 7100
rect 8092 7098 8148 7100
rect 7852 7046 7898 7098
rect 7898 7046 7908 7098
rect 7932 7046 7962 7098
rect 7962 7046 7974 7098
rect 7974 7046 7988 7098
rect 8012 7046 8026 7098
rect 8026 7046 8038 7098
rect 8038 7046 8068 7098
rect 8092 7046 8102 7098
rect 8102 7046 8148 7098
rect 7852 7044 7908 7046
rect 7932 7044 7988 7046
rect 8012 7044 8068 7046
rect 8092 7044 8148 7046
rect 10150 8730 10206 8732
rect 10230 8730 10286 8732
rect 10310 8730 10366 8732
rect 10390 8730 10446 8732
rect 10150 8678 10196 8730
rect 10196 8678 10206 8730
rect 10230 8678 10260 8730
rect 10260 8678 10272 8730
rect 10272 8678 10286 8730
rect 10310 8678 10324 8730
rect 10324 8678 10336 8730
rect 10336 8678 10366 8730
rect 10390 8678 10400 8730
rect 10400 8678 10446 8730
rect 10150 8676 10206 8678
rect 10230 8676 10286 8678
rect 10310 8676 10366 8678
rect 10390 8676 10446 8678
rect 10150 7642 10206 7644
rect 10230 7642 10286 7644
rect 10310 7642 10366 7644
rect 10390 7642 10446 7644
rect 10150 7590 10196 7642
rect 10196 7590 10206 7642
rect 10230 7590 10260 7642
rect 10260 7590 10272 7642
rect 10272 7590 10286 7642
rect 10310 7590 10324 7642
rect 10324 7590 10336 7642
rect 10336 7590 10366 7642
rect 10390 7590 10400 7642
rect 10400 7590 10446 7642
rect 10150 7588 10206 7590
rect 10230 7588 10286 7590
rect 10310 7588 10366 7590
rect 10390 7588 10446 7590
rect 12449 11450 12505 11452
rect 12529 11450 12585 11452
rect 12609 11450 12665 11452
rect 12689 11450 12745 11452
rect 12449 11398 12495 11450
rect 12495 11398 12505 11450
rect 12529 11398 12559 11450
rect 12559 11398 12571 11450
rect 12571 11398 12585 11450
rect 12609 11398 12623 11450
rect 12623 11398 12635 11450
rect 12635 11398 12665 11450
rect 12689 11398 12699 11450
rect 12699 11398 12745 11450
rect 12449 11396 12505 11398
rect 12529 11396 12585 11398
rect 12609 11396 12665 11398
rect 12689 11396 12745 11398
rect 12449 10362 12505 10364
rect 12529 10362 12585 10364
rect 12609 10362 12665 10364
rect 12689 10362 12745 10364
rect 12449 10310 12495 10362
rect 12495 10310 12505 10362
rect 12529 10310 12559 10362
rect 12559 10310 12571 10362
rect 12571 10310 12585 10362
rect 12609 10310 12623 10362
rect 12623 10310 12635 10362
rect 12635 10310 12665 10362
rect 12689 10310 12699 10362
rect 12699 10310 12745 10362
rect 12449 10308 12505 10310
rect 12529 10308 12585 10310
rect 12609 10308 12665 10310
rect 12689 10308 12745 10310
rect 12449 9274 12505 9276
rect 12529 9274 12585 9276
rect 12609 9274 12665 9276
rect 12689 9274 12745 9276
rect 12449 9222 12495 9274
rect 12495 9222 12505 9274
rect 12529 9222 12559 9274
rect 12559 9222 12571 9274
rect 12571 9222 12585 9274
rect 12609 9222 12623 9274
rect 12623 9222 12635 9274
rect 12635 9222 12665 9274
rect 12689 9222 12699 9274
rect 12699 9222 12745 9274
rect 12449 9220 12505 9222
rect 12529 9220 12585 9222
rect 12609 9220 12665 9222
rect 12689 9220 12745 9222
rect 12449 8186 12505 8188
rect 12529 8186 12585 8188
rect 12609 8186 12665 8188
rect 12689 8186 12745 8188
rect 12449 8134 12495 8186
rect 12495 8134 12505 8186
rect 12529 8134 12559 8186
rect 12559 8134 12571 8186
rect 12571 8134 12585 8186
rect 12609 8134 12623 8186
rect 12623 8134 12635 8186
rect 12635 8134 12665 8186
rect 12689 8134 12699 8186
rect 12699 8134 12745 8186
rect 12449 8132 12505 8134
rect 12529 8132 12585 8134
rect 12609 8132 12665 8134
rect 12689 8132 12745 8134
rect 7852 6010 7908 6012
rect 7932 6010 7988 6012
rect 8012 6010 8068 6012
rect 8092 6010 8148 6012
rect 7852 5958 7898 6010
rect 7898 5958 7908 6010
rect 7932 5958 7962 6010
rect 7962 5958 7974 6010
rect 7974 5958 7988 6010
rect 8012 5958 8026 6010
rect 8026 5958 8038 6010
rect 8038 5958 8068 6010
rect 8092 5958 8102 6010
rect 8102 5958 8148 6010
rect 7852 5956 7908 5958
rect 7932 5956 7988 5958
rect 8012 5956 8068 5958
rect 8092 5956 8148 5958
rect 7852 4922 7908 4924
rect 7932 4922 7988 4924
rect 8012 4922 8068 4924
rect 8092 4922 8148 4924
rect 7852 4870 7898 4922
rect 7898 4870 7908 4922
rect 7932 4870 7962 4922
rect 7962 4870 7974 4922
rect 7974 4870 7988 4922
rect 8012 4870 8026 4922
rect 8026 4870 8038 4922
rect 8038 4870 8068 4922
rect 8092 4870 8102 4922
rect 8102 4870 8148 4922
rect 7852 4868 7908 4870
rect 7932 4868 7988 4870
rect 8012 4868 8068 4870
rect 8092 4868 8148 4870
rect 8206 4664 8262 4720
rect 8574 5752 8630 5808
rect 7852 3834 7908 3836
rect 7932 3834 7988 3836
rect 8012 3834 8068 3836
rect 8092 3834 8148 3836
rect 7852 3782 7898 3834
rect 7898 3782 7908 3834
rect 7932 3782 7962 3834
rect 7962 3782 7974 3834
rect 7974 3782 7988 3834
rect 8012 3782 8026 3834
rect 8026 3782 8038 3834
rect 8038 3782 8068 3834
rect 8092 3782 8102 3834
rect 8102 3782 8148 3834
rect 7852 3780 7908 3782
rect 7932 3780 7988 3782
rect 8012 3780 8068 3782
rect 8092 3780 8148 3782
rect 8482 4120 8538 4176
rect 7852 2746 7908 2748
rect 7932 2746 7988 2748
rect 8012 2746 8068 2748
rect 8092 2746 8148 2748
rect 7852 2694 7898 2746
rect 7898 2694 7908 2746
rect 7932 2694 7962 2746
rect 7962 2694 7974 2746
rect 7974 2694 7988 2746
rect 8012 2694 8026 2746
rect 8026 2694 8038 2746
rect 8038 2694 8068 2746
rect 8092 2694 8102 2746
rect 8102 2694 8148 2746
rect 7852 2692 7908 2694
rect 7932 2692 7988 2694
rect 8012 2692 8068 2694
rect 8092 2692 8148 2694
rect 8850 5616 8906 5672
rect 10150 6554 10206 6556
rect 10230 6554 10286 6556
rect 10310 6554 10366 6556
rect 10390 6554 10446 6556
rect 10150 6502 10196 6554
rect 10196 6502 10206 6554
rect 10230 6502 10260 6554
rect 10260 6502 10272 6554
rect 10272 6502 10286 6554
rect 10310 6502 10324 6554
rect 10324 6502 10336 6554
rect 10336 6502 10366 6554
rect 10390 6502 10400 6554
rect 10400 6502 10446 6554
rect 10150 6500 10206 6502
rect 10230 6500 10286 6502
rect 10310 6500 10366 6502
rect 10390 6500 10446 6502
rect 9218 5772 9274 5808
rect 9218 5752 9220 5772
rect 9220 5752 9272 5772
rect 9272 5752 9274 5772
rect 9862 5752 9918 5808
rect 9770 5092 9826 5128
rect 10230 6316 10286 6352
rect 10230 6296 10232 6316
rect 10232 6296 10284 6316
rect 10284 6296 10286 6316
rect 11334 6296 11390 6352
rect 10874 5652 10876 5672
rect 10876 5652 10928 5672
rect 10928 5652 10930 5672
rect 10150 5466 10206 5468
rect 10230 5466 10286 5468
rect 10310 5466 10366 5468
rect 10390 5466 10446 5468
rect 10150 5414 10196 5466
rect 10196 5414 10206 5466
rect 10230 5414 10260 5466
rect 10260 5414 10272 5466
rect 10272 5414 10286 5466
rect 10310 5414 10324 5466
rect 10324 5414 10336 5466
rect 10336 5414 10366 5466
rect 10390 5414 10400 5466
rect 10400 5414 10446 5466
rect 10150 5412 10206 5414
rect 10230 5412 10286 5414
rect 10310 5412 10366 5414
rect 10390 5412 10446 5414
rect 10874 5616 10930 5652
rect 9770 5072 9772 5092
rect 9772 5072 9824 5092
rect 9824 5072 9826 5092
rect 10150 4378 10206 4380
rect 10230 4378 10286 4380
rect 10310 4378 10366 4380
rect 10390 4378 10446 4380
rect 10150 4326 10196 4378
rect 10196 4326 10206 4378
rect 10230 4326 10260 4378
rect 10260 4326 10272 4378
rect 10272 4326 10286 4378
rect 10310 4326 10324 4378
rect 10324 4326 10336 4378
rect 10336 4326 10366 4378
rect 10390 4326 10400 4378
rect 10400 4326 10446 4378
rect 10150 4324 10206 4326
rect 10230 4324 10286 4326
rect 10310 4324 10366 4326
rect 10390 4324 10446 4326
rect 10690 3612 10692 3632
rect 10692 3612 10744 3632
rect 10744 3612 10746 3632
rect 10690 3576 10746 3612
rect 9954 3052 10010 3088
rect 9954 3032 9956 3052
rect 9956 3032 10008 3052
rect 10008 3032 10010 3052
rect 9034 2352 9090 2408
rect 10150 3290 10206 3292
rect 10230 3290 10286 3292
rect 10310 3290 10366 3292
rect 10390 3290 10446 3292
rect 10150 3238 10196 3290
rect 10196 3238 10206 3290
rect 10230 3238 10260 3290
rect 10260 3238 10272 3290
rect 10272 3238 10286 3290
rect 10310 3238 10324 3290
rect 10324 3238 10336 3290
rect 10336 3238 10366 3290
rect 10390 3238 10400 3290
rect 10400 3238 10446 3290
rect 10150 3236 10206 3238
rect 10230 3236 10286 3238
rect 10310 3236 10366 3238
rect 10390 3236 10446 3238
rect 10598 3340 10600 3360
rect 10600 3340 10652 3360
rect 10652 3340 10654 3360
rect 10598 3304 10654 3340
rect 11794 5072 11850 5128
rect 12449 7098 12505 7100
rect 12529 7098 12585 7100
rect 12609 7098 12665 7100
rect 12689 7098 12745 7100
rect 12449 7046 12495 7098
rect 12495 7046 12505 7098
rect 12529 7046 12559 7098
rect 12559 7046 12571 7098
rect 12571 7046 12585 7098
rect 12609 7046 12623 7098
rect 12623 7046 12635 7098
rect 12635 7046 12665 7098
rect 12689 7046 12699 7098
rect 12699 7046 12745 7098
rect 12449 7044 12505 7046
rect 12529 7044 12585 7046
rect 12609 7044 12665 7046
rect 12689 7044 12745 7046
rect 11978 5228 12034 5264
rect 11978 5208 11980 5228
rect 11980 5208 12032 5228
rect 12032 5208 12034 5228
rect 11334 3596 11390 3632
rect 11334 3576 11336 3596
rect 11336 3576 11388 3596
rect 11388 3576 11390 3596
rect 11242 3340 11244 3360
rect 11244 3340 11296 3360
rect 11296 3340 11298 3360
rect 11242 3304 11298 3340
rect 10322 2372 10378 2408
rect 10322 2352 10324 2372
rect 10324 2352 10376 2372
rect 10376 2352 10378 2372
rect 11334 2352 11390 2408
rect 5553 2202 5609 2204
rect 5633 2202 5689 2204
rect 5713 2202 5769 2204
rect 5793 2202 5849 2204
rect 5553 2150 5599 2202
rect 5599 2150 5609 2202
rect 5633 2150 5663 2202
rect 5663 2150 5675 2202
rect 5675 2150 5689 2202
rect 5713 2150 5727 2202
rect 5727 2150 5739 2202
rect 5739 2150 5769 2202
rect 5793 2150 5803 2202
rect 5803 2150 5849 2202
rect 5553 2148 5609 2150
rect 5633 2148 5689 2150
rect 5713 2148 5769 2150
rect 5793 2148 5849 2150
rect 10150 2202 10206 2204
rect 10230 2202 10286 2204
rect 10310 2202 10366 2204
rect 10390 2202 10446 2204
rect 10150 2150 10196 2202
rect 10196 2150 10206 2202
rect 10230 2150 10260 2202
rect 10260 2150 10272 2202
rect 10272 2150 10286 2202
rect 10310 2150 10324 2202
rect 10324 2150 10336 2202
rect 10336 2150 10366 2202
rect 10390 2150 10400 2202
rect 10400 2150 10446 2202
rect 10150 2148 10206 2150
rect 10230 2148 10286 2150
rect 10310 2148 10366 2150
rect 10390 2148 10446 2150
rect 12449 6010 12505 6012
rect 12529 6010 12585 6012
rect 12609 6010 12665 6012
rect 12689 6010 12745 6012
rect 12449 5958 12495 6010
rect 12495 5958 12505 6010
rect 12529 5958 12559 6010
rect 12559 5958 12571 6010
rect 12571 5958 12585 6010
rect 12609 5958 12623 6010
rect 12623 5958 12635 6010
rect 12635 5958 12665 6010
rect 12689 5958 12699 6010
rect 12699 5958 12745 6010
rect 12449 5956 12505 5958
rect 12529 5956 12585 5958
rect 12609 5956 12665 5958
rect 12689 5956 12745 5958
rect 12449 4922 12505 4924
rect 12529 4922 12585 4924
rect 12609 4922 12665 4924
rect 12689 4922 12745 4924
rect 12449 4870 12495 4922
rect 12495 4870 12505 4922
rect 12529 4870 12559 4922
rect 12559 4870 12571 4922
rect 12571 4870 12585 4922
rect 12609 4870 12623 4922
rect 12623 4870 12635 4922
rect 12635 4870 12665 4922
rect 12689 4870 12699 4922
rect 12699 4870 12745 4922
rect 12449 4868 12505 4870
rect 12529 4868 12585 4870
rect 12609 4868 12665 4870
rect 12689 4868 12745 4870
rect 12449 3834 12505 3836
rect 12529 3834 12585 3836
rect 12609 3834 12665 3836
rect 12689 3834 12745 3836
rect 12449 3782 12495 3834
rect 12495 3782 12505 3834
rect 12529 3782 12559 3834
rect 12559 3782 12571 3834
rect 12571 3782 12585 3834
rect 12609 3782 12623 3834
rect 12623 3782 12635 3834
rect 12635 3782 12665 3834
rect 12689 3782 12699 3834
rect 12699 3782 12745 3834
rect 12449 3780 12505 3782
rect 12529 3780 12585 3782
rect 12609 3780 12665 3782
rect 12689 3780 12745 3782
rect 12070 3032 12126 3088
rect 15014 10920 15070 10976
rect 15014 9036 15070 9072
rect 15014 9016 15016 9036
rect 15016 9016 15068 9036
rect 15068 9016 15070 9036
rect 14462 6976 14518 7032
rect 13818 5228 13874 5264
rect 13818 5208 13820 5228
rect 13820 5208 13872 5228
rect 13872 5208 13874 5228
rect 14462 4936 14518 4992
rect 12449 2746 12505 2748
rect 12529 2746 12585 2748
rect 12609 2746 12665 2748
rect 12689 2746 12745 2748
rect 12449 2694 12495 2746
rect 12495 2694 12505 2746
rect 12529 2694 12559 2746
rect 12559 2694 12571 2746
rect 12571 2694 12585 2746
rect 12609 2694 12623 2746
rect 12623 2694 12635 2746
rect 12635 2694 12665 2746
rect 12689 2694 12699 2746
rect 12699 2694 12745 2746
rect 12449 2692 12505 2694
rect 12529 2692 12585 2694
rect 12609 2692 12665 2694
rect 12689 2692 12745 2694
rect 14462 2896 14518 2952
rect 14922 1028 14924 1048
rect 14924 1028 14976 1048
rect 14976 1028 14978 1048
rect 14922 992 14978 1028
<< metal3 >>
rect 14917 15058 14983 15061
rect 15200 15058 16000 15088
rect 14917 15056 16000 15058
rect 14917 15000 14922 15056
rect 14978 15000 16000 15056
rect 14917 14998 16000 15000
rect 14917 14995 14983 14998
rect 15200 14968 16000 14998
rect 3242 13632 3562 13633
rect 3242 13568 3250 13632
rect 3314 13568 3330 13632
rect 3394 13568 3410 13632
rect 3474 13568 3490 13632
rect 3554 13568 3562 13632
rect 3242 13567 3562 13568
rect 7840 13632 8160 13633
rect 7840 13568 7848 13632
rect 7912 13568 7928 13632
rect 7992 13568 8008 13632
rect 8072 13568 8088 13632
rect 8152 13568 8160 13632
rect 7840 13567 8160 13568
rect 12437 13632 12757 13633
rect 12437 13568 12445 13632
rect 12509 13568 12525 13632
rect 12589 13568 12605 13632
rect 12669 13568 12685 13632
rect 12749 13568 12757 13632
rect 12437 13567 12757 13568
rect 5541 13088 5861 13089
rect 5541 13024 5549 13088
rect 5613 13024 5629 13088
rect 5693 13024 5709 13088
rect 5773 13024 5789 13088
rect 5853 13024 5861 13088
rect 5541 13023 5861 13024
rect 10138 13088 10458 13089
rect 10138 13024 10146 13088
rect 10210 13024 10226 13088
rect 10290 13024 10306 13088
rect 10370 13024 10386 13088
rect 10450 13024 10458 13088
rect 10138 13023 10458 13024
rect 11329 13018 11395 13021
rect 15200 13018 16000 13048
rect 11329 13016 16000 13018
rect 11329 12960 11334 13016
rect 11390 12960 16000 13016
rect 11329 12958 16000 12960
rect 11329 12955 11395 12958
rect 15200 12928 16000 12958
rect 3242 12544 3562 12545
rect 3242 12480 3250 12544
rect 3314 12480 3330 12544
rect 3394 12480 3410 12544
rect 3474 12480 3490 12544
rect 3554 12480 3562 12544
rect 3242 12479 3562 12480
rect 7840 12544 8160 12545
rect 7840 12480 7848 12544
rect 7912 12480 7928 12544
rect 7992 12480 8008 12544
rect 8072 12480 8088 12544
rect 8152 12480 8160 12544
rect 7840 12479 8160 12480
rect 12437 12544 12757 12545
rect 12437 12480 12445 12544
rect 12509 12480 12525 12544
rect 12589 12480 12605 12544
rect 12669 12480 12685 12544
rect 12749 12480 12757 12544
rect 12437 12479 12757 12480
rect 0 12066 800 12096
rect 4153 12066 4219 12069
rect 0 12064 4219 12066
rect 0 12008 4158 12064
rect 4214 12008 4219 12064
rect 0 12006 4219 12008
rect 0 11976 800 12006
rect 4153 12003 4219 12006
rect 5541 12000 5861 12001
rect 5541 11936 5549 12000
rect 5613 11936 5629 12000
rect 5693 11936 5709 12000
rect 5773 11936 5789 12000
rect 5853 11936 5861 12000
rect 5541 11935 5861 11936
rect 10138 12000 10458 12001
rect 10138 11936 10146 12000
rect 10210 11936 10226 12000
rect 10290 11936 10306 12000
rect 10370 11936 10386 12000
rect 10450 11936 10458 12000
rect 10138 11935 10458 11936
rect 7833 11794 7899 11797
rect 9213 11794 9279 11797
rect 7833 11792 9279 11794
rect 7833 11736 7838 11792
rect 7894 11736 9218 11792
rect 9274 11736 9279 11792
rect 7833 11734 9279 11736
rect 7833 11731 7899 11734
rect 9213 11731 9279 11734
rect 3242 11456 3562 11457
rect 3242 11392 3250 11456
rect 3314 11392 3330 11456
rect 3394 11392 3410 11456
rect 3474 11392 3490 11456
rect 3554 11392 3562 11456
rect 3242 11391 3562 11392
rect 7840 11456 8160 11457
rect 7840 11392 7848 11456
rect 7912 11392 7928 11456
rect 7992 11392 8008 11456
rect 8072 11392 8088 11456
rect 8152 11392 8160 11456
rect 7840 11391 8160 11392
rect 12437 11456 12757 11457
rect 12437 11392 12445 11456
rect 12509 11392 12525 11456
rect 12589 11392 12605 11456
rect 12669 11392 12685 11456
rect 12749 11392 12757 11456
rect 12437 11391 12757 11392
rect 9029 11250 9095 11253
rect 8894 11248 9095 11250
rect 8894 11192 9034 11248
rect 9090 11192 9095 11248
rect 8894 11190 9095 11192
rect 5533 11114 5599 11117
rect 7281 11114 7347 11117
rect 8201 11114 8267 11117
rect 8894 11114 8954 11190
rect 9029 11187 9095 11190
rect 5533 11112 8954 11114
rect 5533 11056 5538 11112
rect 5594 11056 7286 11112
rect 7342 11056 8206 11112
rect 8262 11056 8954 11112
rect 5533 11054 8954 11056
rect 9029 11114 9095 11117
rect 10133 11114 10199 11117
rect 10685 11114 10751 11117
rect 9029 11112 10751 11114
rect 9029 11056 9034 11112
rect 9090 11056 10138 11112
rect 10194 11056 10690 11112
rect 10746 11056 10751 11112
rect 9029 11054 10751 11056
rect 5533 11051 5599 11054
rect 7281 11051 7347 11054
rect 8201 11051 8267 11054
rect 9029 11051 9095 11054
rect 10133 11051 10199 11054
rect 10685 11051 10751 11054
rect 15009 10978 15075 10981
rect 15200 10978 16000 11008
rect 15009 10976 16000 10978
rect 15009 10920 15014 10976
rect 15070 10920 16000 10976
rect 15009 10918 16000 10920
rect 15009 10915 15075 10918
rect 5541 10912 5861 10913
rect 5541 10848 5549 10912
rect 5613 10848 5629 10912
rect 5693 10848 5709 10912
rect 5773 10848 5789 10912
rect 5853 10848 5861 10912
rect 5541 10847 5861 10848
rect 10138 10912 10458 10913
rect 10138 10848 10146 10912
rect 10210 10848 10226 10912
rect 10290 10848 10306 10912
rect 10370 10848 10386 10912
rect 10450 10848 10458 10912
rect 15200 10888 16000 10918
rect 10138 10847 10458 10848
rect 3242 10368 3562 10369
rect 3242 10304 3250 10368
rect 3314 10304 3330 10368
rect 3394 10304 3410 10368
rect 3474 10304 3490 10368
rect 3554 10304 3562 10368
rect 3242 10303 3562 10304
rect 7840 10368 8160 10369
rect 7840 10304 7848 10368
rect 7912 10304 7928 10368
rect 7992 10304 8008 10368
rect 8072 10304 8088 10368
rect 8152 10304 8160 10368
rect 7840 10303 8160 10304
rect 12437 10368 12757 10369
rect 12437 10304 12445 10368
rect 12509 10304 12525 10368
rect 12589 10304 12605 10368
rect 12669 10304 12685 10368
rect 12749 10304 12757 10368
rect 12437 10303 12757 10304
rect 3049 10026 3115 10029
rect 4521 10026 4587 10029
rect 3049 10024 4587 10026
rect 3049 9968 3054 10024
rect 3110 9968 4526 10024
rect 4582 9968 4587 10024
rect 3049 9966 4587 9968
rect 3049 9963 3115 9966
rect 4521 9963 4587 9966
rect 8569 10026 8635 10029
rect 11053 10026 11119 10029
rect 8569 10024 11119 10026
rect 8569 9968 8574 10024
rect 8630 9968 11058 10024
rect 11114 9968 11119 10024
rect 8569 9966 11119 9968
rect 8569 9963 8635 9966
rect 11053 9963 11119 9966
rect 2957 9890 3023 9893
rect 3509 9890 3575 9893
rect 2957 9888 3575 9890
rect 2957 9832 2962 9888
rect 3018 9832 3514 9888
rect 3570 9832 3575 9888
rect 2957 9830 3575 9832
rect 2957 9827 3023 9830
rect 3509 9827 3575 9830
rect 5541 9824 5861 9825
rect 5541 9760 5549 9824
rect 5613 9760 5629 9824
rect 5693 9760 5709 9824
rect 5773 9760 5789 9824
rect 5853 9760 5861 9824
rect 5541 9759 5861 9760
rect 10138 9824 10458 9825
rect 10138 9760 10146 9824
rect 10210 9760 10226 9824
rect 10290 9760 10306 9824
rect 10370 9760 10386 9824
rect 10450 9760 10458 9824
rect 10138 9759 10458 9760
rect 3242 9280 3562 9281
rect 3242 9216 3250 9280
rect 3314 9216 3330 9280
rect 3394 9216 3410 9280
rect 3474 9216 3490 9280
rect 3554 9216 3562 9280
rect 3242 9215 3562 9216
rect 7840 9280 8160 9281
rect 7840 9216 7848 9280
rect 7912 9216 7928 9280
rect 7992 9216 8008 9280
rect 8072 9216 8088 9280
rect 8152 9216 8160 9280
rect 7840 9215 8160 9216
rect 12437 9280 12757 9281
rect 12437 9216 12445 9280
rect 12509 9216 12525 9280
rect 12589 9216 12605 9280
rect 12669 9216 12685 9280
rect 12749 9216 12757 9280
rect 12437 9215 12757 9216
rect 15009 9074 15075 9077
rect 15200 9074 16000 9104
rect 15009 9072 16000 9074
rect 15009 9016 15014 9072
rect 15070 9016 16000 9072
rect 15009 9014 16000 9016
rect 15009 9011 15075 9014
rect 15200 8984 16000 9014
rect 5541 8736 5861 8737
rect 5541 8672 5549 8736
rect 5613 8672 5629 8736
rect 5693 8672 5709 8736
rect 5773 8672 5789 8736
rect 5853 8672 5861 8736
rect 5541 8671 5861 8672
rect 10138 8736 10458 8737
rect 10138 8672 10146 8736
rect 10210 8672 10226 8736
rect 10290 8672 10306 8736
rect 10370 8672 10386 8736
rect 10450 8672 10458 8736
rect 10138 8671 10458 8672
rect 3242 8192 3562 8193
rect 3242 8128 3250 8192
rect 3314 8128 3330 8192
rect 3394 8128 3410 8192
rect 3474 8128 3490 8192
rect 3554 8128 3562 8192
rect 3242 8127 3562 8128
rect 7840 8192 8160 8193
rect 7840 8128 7848 8192
rect 7912 8128 7928 8192
rect 7992 8128 8008 8192
rect 8072 8128 8088 8192
rect 8152 8128 8160 8192
rect 7840 8127 8160 8128
rect 12437 8192 12757 8193
rect 12437 8128 12445 8192
rect 12509 8128 12525 8192
rect 12589 8128 12605 8192
rect 12669 8128 12685 8192
rect 12749 8128 12757 8192
rect 12437 8127 12757 8128
rect 5541 7648 5861 7649
rect 5541 7584 5549 7648
rect 5613 7584 5629 7648
rect 5693 7584 5709 7648
rect 5773 7584 5789 7648
rect 5853 7584 5861 7648
rect 5541 7583 5861 7584
rect 10138 7648 10458 7649
rect 10138 7584 10146 7648
rect 10210 7584 10226 7648
rect 10290 7584 10306 7648
rect 10370 7584 10386 7648
rect 10450 7584 10458 7648
rect 10138 7583 10458 7584
rect 3242 7104 3562 7105
rect 3242 7040 3250 7104
rect 3314 7040 3330 7104
rect 3394 7040 3410 7104
rect 3474 7040 3490 7104
rect 3554 7040 3562 7104
rect 3242 7039 3562 7040
rect 7840 7104 8160 7105
rect 7840 7040 7848 7104
rect 7912 7040 7928 7104
rect 7992 7040 8008 7104
rect 8072 7040 8088 7104
rect 8152 7040 8160 7104
rect 7840 7039 8160 7040
rect 12437 7104 12757 7105
rect 12437 7040 12445 7104
rect 12509 7040 12525 7104
rect 12589 7040 12605 7104
rect 12669 7040 12685 7104
rect 12749 7040 12757 7104
rect 12437 7039 12757 7040
rect 14457 7034 14523 7037
rect 15200 7034 16000 7064
rect 14457 7032 16000 7034
rect 14457 6976 14462 7032
rect 14518 6976 16000 7032
rect 14457 6974 16000 6976
rect 14457 6971 14523 6974
rect 15200 6944 16000 6974
rect 5541 6560 5861 6561
rect 5541 6496 5549 6560
rect 5613 6496 5629 6560
rect 5693 6496 5709 6560
rect 5773 6496 5789 6560
rect 5853 6496 5861 6560
rect 5541 6495 5861 6496
rect 10138 6560 10458 6561
rect 10138 6496 10146 6560
rect 10210 6496 10226 6560
rect 10290 6496 10306 6560
rect 10370 6496 10386 6560
rect 10450 6496 10458 6560
rect 10138 6495 10458 6496
rect 10225 6354 10291 6357
rect 11329 6354 11395 6357
rect 10225 6352 11395 6354
rect 10225 6296 10230 6352
rect 10286 6296 11334 6352
rect 11390 6296 11395 6352
rect 10225 6294 11395 6296
rect 10225 6291 10291 6294
rect 11329 6291 11395 6294
rect 3242 6016 3562 6017
rect 3242 5952 3250 6016
rect 3314 5952 3330 6016
rect 3394 5952 3410 6016
rect 3474 5952 3490 6016
rect 3554 5952 3562 6016
rect 3242 5951 3562 5952
rect 7840 6016 8160 6017
rect 7840 5952 7848 6016
rect 7912 5952 7928 6016
rect 7992 5952 8008 6016
rect 8072 5952 8088 6016
rect 8152 5952 8160 6016
rect 7840 5951 8160 5952
rect 12437 6016 12757 6017
rect 12437 5952 12445 6016
rect 12509 5952 12525 6016
rect 12589 5952 12605 6016
rect 12669 5952 12685 6016
rect 12749 5952 12757 6016
rect 12437 5951 12757 5952
rect 8569 5810 8635 5813
rect 9213 5810 9279 5813
rect 9857 5810 9923 5813
rect 8569 5808 8770 5810
rect 8569 5752 8574 5808
rect 8630 5752 8770 5808
rect 8569 5750 8770 5752
rect 8569 5747 8635 5750
rect 8710 5674 8770 5750
rect 9213 5808 9923 5810
rect 9213 5752 9218 5808
rect 9274 5752 9862 5808
rect 9918 5752 9923 5808
rect 9213 5750 9923 5752
rect 9213 5747 9279 5750
rect 9857 5747 9923 5750
rect 8845 5674 8911 5677
rect 10869 5674 10935 5677
rect 8710 5672 10935 5674
rect 8710 5616 8850 5672
rect 8906 5616 10874 5672
rect 10930 5616 10935 5672
rect 8710 5614 10935 5616
rect 8845 5611 8911 5614
rect 10869 5611 10935 5614
rect 2497 5538 2563 5541
rect 4613 5538 4679 5541
rect 2497 5536 4722 5538
rect 2497 5480 2502 5536
rect 2558 5480 4618 5536
rect 4674 5480 4722 5536
rect 2497 5478 4722 5480
rect 2497 5475 2563 5478
rect 4613 5475 4722 5478
rect 4662 5266 4722 5475
rect 5541 5472 5861 5473
rect 5541 5408 5549 5472
rect 5613 5408 5629 5472
rect 5693 5408 5709 5472
rect 5773 5408 5789 5472
rect 5853 5408 5861 5472
rect 5541 5407 5861 5408
rect 10138 5472 10458 5473
rect 10138 5408 10146 5472
rect 10210 5408 10226 5472
rect 10290 5408 10306 5472
rect 10370 5408 10386 5472
rect 10450 5408 10458 5472
rect 10138 5407 10458 5408
rect 5717 5266 5783 5269
rect 4662 5264 5783 5266
rect 4662 5208 5722 5264
rect 5778 5208 5783 5264
rect 4662 5206 5783 5208
rect 5717 5203 5783 5206
rect 11973 5266 12039 5269
rect 13813 5266 13879 5269
rect 11973 5264 13879 5266
rect 11973 5208 11978 5264
rect 12034 5208 13818 5264
rect 13874 5208 13879 5264
rect 11973 5206 13879 5208
rect 11973 5203 12039 5206
rect 13813 5203 13879 5206
rect 9765 5130 9831 5133
rect 11789 5130 11855 5133
rect 9765 5128 11855 5130
rect 9765 5072 9770 5128
rect 9826 5072 11794 5128
rect 11850 5072 11855 5128
rect 9765 5070 11855 5072
rect 9765 5067 9831 5070
rect 11789 5067 11855 5070
rect 14457 4994 14523 4997
rect 15200 4994 16000 5024
rect 14457 4992 16000 4994
rect 14457 4936 14462 4992
rect 14518 4936 16000 4992
rect 14457 4934 16000 4936
rect 14457 4931 14523 4934
rect 3242 4928 3562 4929
rect 3242 4864 3250 4928
rect 3314 4864 3330 4928
rect 3394 4864 3410 4928
rect 3474 4864 3490 4928
rect 3554 4864 3562 4928
rect 3242 4863 3562 4864
rect 7840 4928 8160 4929
rect 7840 4864 7848 4928
rect 7912 4864 7928 4928
rect 7992 4864 8008 4928
rect 8072 4864 8088 4928
rect 8152 4864 8160 4928
rect 7840 4863 8160 4864
rect 12437 4928 12757 4929
rect 12437 4864 12445 4928
rect 12509 4864 12525 4928
rect 12589 4864 12605 4928
rect 12669 4864 12685 4928
rect 12749 4864 12757 4928
rect 15200 4904 16000 4934
rect 12437 4863 12757 4864
rect 4337 4722 4403 4725
rect 8201 4722 8267 4725
rect 4337 4720 8267 4722
rect 4337 4664 4342 4720
rect 4398 4664 8206 4720
rect 8262 4664 8267 4720
rect 4337 4662 8267 4664
rect 4337 4659 4403 4662
rect 8201 4659 8267 4662
rect 5541 4384 5861 4385
rect 5541 4320 5549 4384
rect 5613 4320 5629 4384
rect 5693 4320 5709 4384
rect 5773 4320 5789 4384
rect 5853 4320 5861 4384
rect 5541 4319 5861 4320
rect 10138 4384 10458 4385
rect 10138 4320 10146 4384
rect 10210 4320 10226 4384
rect 10290 4320 10306 4384
rect 10370 4320 10386 4384
rect 10450 4320 10458 4384
rect 10138 4319 10458 4320
rect 4521 4178 4587 4181
rect 5533 4178 5599 4181
rect 8477 4178 8543 4181
rect 4521 4176 8543 4178
rect 4521 4120 4526 4176
rect 4582 4120 5538 4176
rect 5594 4120 8482 4176
rect 8538 4120 8543 4176
rect 4521 4118 8543 4120
rect 4521 4115 4587 4118
rect 5533 4115 5599 4118
rect 8477 4115 8543 4118
rect 0 4042 800 4072
rect 4521 4042 4587 4045
rect 0 4040 4587 4042
rect 0 3984 4526 4040
rect 4582 3984 4587 4040
rect 0 3982 4587 3984
rect 0 3952 800 3982
rect 4521 3979 4587 3982
rect 4153 3906 4219 3909
rect 5533 3906 5599 3909
rect 4153 3904 5599 3906
rect 4153 3848 4158 3904
rect 4214 3848 5538 3904
rect 5594 3848 5599 3904
rect 4153 3846 5599 3848
rect 4153 3843 4219 3846
rect 5533 3843 5599 3846
rect 3242 3840 3562 3841
rect 3242 3776 3250 3840
rect 3314 3776 3330 3840
rect 3394 3776 3410 3840
rect 3474 3776 3490 3840
rect 3554 3776 3562 3840
rect 3242 3775 3562 3776
rect 7840 3840 8160 3841
rect 7840 3776 7848 3840
rect 7912 3776 7928 3840
rect 7992 3776 8008 3840
rect 8072 3776 8088 3840
rect 8152 3776 8160 3840
rect 7840 3775 8160 3776
rect 12437 3840 12757 3841
rect 12437 3776 12445 3840
rect 12509 3776 12525 3840
rect 12589 3776 12605 3840
rect 12669 3776 12685 3840
rect 12749 3776 12757 3840
rect 12437 3775 12757 3776
rect 3785 3634 3851 3637
rect 5257 3634 5323 3637
rect 3785 3632 5323 3634
rect 3785 3576 3790 3632
rect 3846 3576 5262 3632
rect 5318 3576 5323 3632
rect 3785 3574 5323 3576
rect 3785 3571 3851 3574
rect 5257 3571 5323 3574
rect 10685 3634 10751 3637
rect 11329 3634 11395 3637
rect 10685 3632 11395 3634
rect 10685 3576 10690 3632
rect 10746 3576 11334 3632
rect 11390 3576 11395 3632
rect 10685 3574 11395 3576
rect 10685 3571 10751 3574
rect 11329 3571 11395 3574
rect 3417 3498 3483 3501
rect 5165 3498 5231 3501
rect 3417 3496 5231 3498
rect 3417 3440 3422 3496
rect 3478 3440 5170 3496
rect 5226 3440 5231 3496
rect 3417 3438 5231 3440
rect 3417 3435 3483 3438
rect 5165 3435 5231 3438
rect 10593 3362 10659 3365
rect 11237 3362 11303 3365
rect 10593 3360 11303 3362
rect 10593 3304 10598 3360
rect 10654 3304 11242 3360
rect 11298 3304 11303 3360
rect 10593 3302 11303 3304
rect 10593 3299 10659 3302
rect 11237 3299 11303 3302
rect 5541 3296 5861 3297
rect 5541 3232 5549 3296
rect 5613 3232 5629 3296
rect 5693 3232 5709 3296
rect 5773 3232 5789 3296
rect 5853 3232 5861 3296
rect 5541 3231 5861 3232
rect 10138 3296 10458 3297
rect 10138 3232 10146 3296
rect 10210 3232 10226 3296
rect 10290 3232 10306 3296
rect 10370 3232 10386 3296
rect 10450 3232 10458 3296
rect 10138 3231 10458 3232
rect 9949 3090 10015 3093
rect 12065 3090 12131 3093
rect 9949 3088 12131 3090
rect 9949 3032 9954 3088
rect 10010 3032 12070 3088
rect 12126 3032 12131 3088
rect 9949 3030 12131 3032
rect 9949 3027 10015 3030
rect 12065 3027 12131 3030
rect 14457 2954 14523 2957
rect 15200 2954 16000 2984
rect 14457 2952 16000 2954
rect 14457 2896 14462 2952
rect 14518 2896 16000 2952
rect 14457 2894 16000 2896
rect 14457 2891 14523 2894
rect 15200 2864 16000 2894
rect 3242 2752 3562 2753
rect 3242 2688 3250 2752
rect 3314 2688 3330 2752
rect 3394 2688 3410 2752
rect 3474 2688 3490 2752
rect 3554 2688 3562 2752
rect 3242 2687 3562 2688
rect 7840 2752 8160 2753
rect 7840 2688 7848 2752
rect 7912 2688 7928 2752
rect 7992 2688 8008 2752
rect 8072 2688 8088 2752
rect 8152 2688 8160 2752
rect 7840 2687 8160 2688
rect 12437 2752 12757 2753
rect 12437 2688 12445 2752
rect 12509 2688 12525 2752
rect 12589 2688 12605 2752
rect 12669 2688 12685 2752
rect 12749 2688 12757 2752
rect 12437 2687 12757 2688
rect 9029 2410 9095 2413
rect 10317 2410 10383 2413
rect 11329 2410 11395 2413
rect 9029 2408 11395 2410
rect 9029 2352 9034 2408
rect 9090 2352 10322 2408
rect 10378 2352 11334 2408
rect 11390 2352 11395 2408
rect 9029 2350 11395 2352
rect 9029 2347 9095 2350
rect 10317 2347 10383 2350
rect 11329 2347 11395 2350
rect 5541 2208 5861 2209
rect 5541 2144 5549 2208
rect 5613 2144 5629 2208
rect 5693 2144 5709 2208
rect 5773 2144 5789 2208
rect 5853 2144 5861 2208
rect 5541 2143 5861 2144
rect 10138 2208 10458 2209
rect 10138 2144 10146 2208
rect 10210 2144 10226 2208
rect 10290 2144 10306 2208
rect 10370 2144 10386 2208
rect 10450 2144 10458 2208
rect 10138 2143 10458 2144
rect 14917 1050 14983 1053
rect 15200 1050 16000 1080
rect 14917 1048 16000 1050
rect 14917 992 14922 1048
rect 14978 992 16000 1048
rect 14917 990 16000 992
rect 14917 987 14983 990
rect 15200 960 16000 990
<< via3 >>
rect 3250 13628 3314 13632
rect 3250 13572 3254 13628
rect 3254 13572 3310 13628
rect 3310 13572 3314 13628
rect 3250 13568 3314 13572
rect 3330 13628 3394 13632
rect 3330 13572 3334 13628
rect 3334 13572 3390 13628
rect 3390 13572 3394 13628
rect 3330 13568 3394 13572
rect 3410 13628 3474 13632
rect 3410 13572 3414 13628
rect 3414 13572 3470 13628
rect 3470 13572 3474 13628
rect 3410 13568 3474 13572
rect 3490 13628 3554 13632
rect 3490 13572 3494 13628
rect 3494 13572 3550 13628
rect 3550 13572 3554 13628
rect 3490 13568 3554 13572
rect 7848 13628 7912 13632
rect 7848 13572 7852 13628
rect 7852 13572 7908 13628
rect 7908 13572 7912 13628
rect 7848 13568 7912 13572
rect 7928 13628 7992 13632
rect 7928 13572 7932 13628
rect 7932 13572 7988 13628
rect 7988 13572 7992 13628
rect 7928 13568 7992 13572
rect 8008 13628 8072 13632
rect 8008 13572 8012 13628
rect 8012 13572 8068 13628
rect 8068 13572 8072 13628
rect 8008 13568 8072 13572
rect 8088 13628 8152 13632
rect 8088 13572 8092 13628
rect 8092 13572 8148 13628
rect 8148 13572 8152 13628
rect 8088 13568 8152 13572
rect 12445 13628 12509 13632
rect 12445 13572 12449 13628
rect 12449 13572 12505 13628
rect 12505 13572 12509 13628
rect 12445 13568 12509 13572
rect 12525 13628 12589 13632
rect 12525 13572 12529 13628
rect 12529 13572 12585 13628
rect 12585 13572 12589 13628
rect 12525 13568 12589 13572
rect 12605 13628 12669 13632
rect 12605 13572 12609 13628
rect 12609 13572 12665 13628
rect 12665 13572 12669 13628
rect 12605 13568 12669 13572
rect 12685 13628 12749 13632
rect 12685 13572 12689 13628
rect 12689 13572 12745 13628
rect 12745 13572 12749 13628
rect 12685 13568 12749 13572
rect 5549 13084 5613 13088
rect 5549 13028 5553 13084
rect 5553 13028 5609 13084
rect 5609 13028 5613 13084
rect 5549 13024 5613 13028
rect 5629 13084 5693 13088
rect 5629 13028 5633 13084
rect 5633 13028 5689 13084
rect 5689 13028 5693 13084
rect 5629 13024 5693 13028
rect 5709 13084 5773 13088
rect 5709 13028 5713 13084
rect 5713 13028 5769 13084
rect 5769 13028 5773 13084
rect 5709 13024 5773 13028
rect 5789 13084 5853 13088
rect 5789 13028 5793 13084
rect 5793 13028 5849 13084
rect 5849 13028 5853 13084
rect 5789 13024 5853 13028
rect 10146 13084 10210 13088
rect 10146 13028 10150 13084
rect 10150 13028 10206 13084
rect 10206 13028 10210 13084
rect 10146 13024 10210 13028
rect 10226 13084 10290 13088
rect 10226 13028 10230 13084
rect 10230 13028 10286 13084
rect 10286 13028 10290 13084
rect 10226 13024 10290 13028
rect 10306 13084 10370 13088
rect 10306 13028 10310 13084
rect 10310 13028 10366 13084
rect 10366 13028 10370 13084
rect 10306 13024 10370 13028
rect 10386 13084 10450 13088
rect 10386 13028 10390 13084
rect 10390 13028 10446 13084
rect 10446 13028 10450 13084
rect 10386 13024 10450 13028
rect 3250 12540 3314 12544
rect 3250 12484 3254 12540
rect 3254 12484 3310 12540
rect 3310 12484 3314 12540
rect 3250 12480 3314 12484
rect 3330 12540 3394 12544
rect 3330 12484 3334 12540
rect 3334 12484 3390 12540
rect 3390 12484 3394 12540
rect 3330 12480 3394 12484
rect 3410 12540 3474 12544
rect 3410 12484 3414 12540
rect 3414 12484 3470 12540
rect 3470 12484 3474 12540
rect 3410 12480 3474 12484
rect 3490 12540 3554 12544
rect 3490 12484 3494 12540
rect 3494 12484 3550 12540
rect 3550 12484 3554 12540
rect 3490 12480 3554 12484
rect 7848 12540 7912 12544
rect 7848 12484 7852 12540
rect 7852 12484 7908 12540
rect 7908 12484 7912 12540
rect 7848 12480 7912 12484
rect 7928 12540 7992 12544
rect 7928 12484 7932 12540
rect 7932 12484 7988 12540
rect 7988 12484 7992 12540
rect 7928 12480 7992 12484
rect 8008 12540 8072 12544
rect 8008 12484 8012 12540
rect 8012 12484 8068 12540
rect 8068 12484 8072 12540
rect 8008 12480 8072 12484
rect 8088 12540 8152 12544
rect 8088 12484 8092 12540
rect 8092 12484 8148 12540
rect 8148 12484 8152 12540
rect 8088 12480 8152 12484
rect 12445 12540 12509 12544
rect 12445 12484 12449 12540
rect 12449 12484 12505 12540
rect 12505 12484 12509 12540
rect 12445 12480 12509 12484
rect 12525 12540 12589 12544
rect 12525 12484 12529 12540
rect 12529 12484 12585 12540
rect 12585 12484 12589 12540
rect 12525 12480 12589 12484
rect 12605 12540 12669 12544
rect 12605 12484 12609 12540
rect 12609 12484 12665 12540
rect 12665 12484 12669 12540
rect 12605 12480 12669 12484
rect 12685 12540 12749 12544
rect 12685 12484 12689 12540
rect 12689 12484 12745 12540
rect 12745 12484 12749 12540
rect 12685 12480 12749 12484
rect 5549 11996 5613 12000
rect 5549 11940 5553 11996
rect 5553 11940 5609 11996
rect 5609 11940 5613 11996
rect 5549 11936 5613 11940
rect 5629 11996 5693 12000
rect 5629 11940 5633 11996
rect 5633 11940 5689 11996
rect 5689 11940 5693 11996
rect 5629 11936 5693 11940
rect 5709 11996 5773 12000
rect 5709 11940 5713 11996
rect 5713 11940 5769 11996
rect 5769 11940 5773 11996
rect 5709 11936 5773 11940
rect 5789 11996 5853 12000
rect 5789 11940 5793 11996
rect 5793 11940 5849 11996
rect 5849 11940 5853 11996
rect 5789 11936 5853 11940
rect 10146 11996 10210 12000
rect 10146 11940 10150 11996
rect 10150 11940 10206 11996
rect 10206 11940 10210 11996
rect 10146 11936 10210 11940
rect 10226 11996 10290 12000
rect 10226 11940 10230 11996
rect 10230 11940 10286 11996
rect 10286 11940 10290 11996
rect 10226 11936 10290 11940
rect 10306 11996 10370 12000
rect 10306 11940 10310 11996
rect 10310 11940 10366 11996
rect 10366 11940 10370 11996
rect 10306 11936 10370 11940
rect 10386 11996 10450 12000
rect 10386 11940 10390 11996
rect 10390 11940 10446 11996
rect 10446 11940 10450 11996
rect 10386 11936 10450 11940
rect 3250 11452 3314 11456
rect 3250 11396 3254 11452
rect 3254 11396 3310 11452
rect 3310 11396 3314 11452
rect 3250 11392 3314 11396
rect 3330 11452 3394 11456
rect 3330 11396 3334 11452
rect 3334 11396 3390 11452
rect 3390 11396 3394 11452
rect 3330 11392 3394 11396
rect 3410 11452 3474 11456
rect 3410 11396 3414 11452
rect 3414 11396 3470 11452
rect 3470 11396 3474 11452
rect 3410 11392 3474 11396
rect 3490 11452 3554 11456
rect 3490 11396 3494 11452
rect 3494 11396 3550 11452
rect 3550 11396 3554 11452
rect 3490 11392 3554 11396
rect 7848 11452 7912 11456
rect 7848 11396 7852 11452
rect 7852 11396 7908 11452
rect 7908 11396 7912 11452
rect 7848 11392 7912 11396
rect 7928 11452 7992 11456
rect 7928 11396 7932 11452
rect 7932 11396 7988 11452
rect 7988 11396 7992 11452
rect 7928 11392 7992 11396
rect 8008 11452 8072 11456
rect 8008 11396 8012 11452
rect 8012 11396 8068 11452
rect 8068 11396 8072 11452
rect 8008 11392 8072 11396
rect 8088 11452 8152 11456
rect 8088 11396 8092 11452
rect 8092 11396 8148 11452
rect 8148 11396 8152 11452
rect 8088 11392 8152 11396
rect 12445 11452 12509 11456
rect 12445 11396 12449 11452
rect 12449 11396 12505 11452
rect 12505 11396 12509 11452
rect 12445 11392 12509 11396
rect 12525 11452 12589 11456
rect 12525 11396 12529 11452
rect 12529 11396 12585 11452
rect 12585 11396 12589 11452
rect 12525 11392 12589 11396
rect 12605 11452 12669 11456
rect 12605 11396 12609 11452
rect 12609 11396 12665 11452
rect 12665 11396 12669 11452
rect 12605 11392 12669 11396
rect 12685 11452 12749 11456
rect 12685 11396 12689 11452
rect 12689 11396 12745 11452
rect 12745 11396 12749 11452
rect 12685 11392 12749 11396
rect 5549 10908 5613 10912
rect 5549 10852 5553 10908
rect 5553 10852 5609 10908
rect 5609 10852 5613 10908
rect 5549 10848 5613 10852
rect 5629 10908 5693 10912
rect 5629 10852 5633 10908
rect 5633 10852 5689 10908
rect 5689 10852 5693 10908
rect 5629 10848 5693 10852
rect 5709 10908 5773 10912
rect 5709 10852 5713 10908
rect 5713 10852 5769 10908
rect 5769 10852 5773 10908
rect 5709 10848 5773 10852
rect 5789 10908 5853 10912
rect 5789 10852 5793 10908
rect 5793 10852 5849 10908
rect 5849 10852 5853 10908
rect 5789 10848 5853 10852
rect 10146 10908 10210 10912
rect 10146 10852 10150 10908
rect 10150 10852 10206 10908
rect 10206 10852 10210 10908
rect 10146 10848 10210 10852
rect 10226 10908 10290 10912
rect 10226 10852 10230 10908
rect 10230 10852 10286 10908
rect 10286 10852 10290 10908
rect 10226 10848 10290 10852
rect 10306 10908 10370 10912
rect 10306 10852 10310 10908
rect 10310 10852 10366 10908
rect 10366 10852 10370 10908
rect 10306 10848 10370 10852
rect 10386 10908 10450 10912
rect 10386 10852 10390 10908
rect 10390 10852 10446 10908
rect 10446 10852 10450 10908
rect 10386 10848 10450 10852
rect 3250 10364 3314 10368
rect 3250 10308 3254 10364
rect 3254 10308 3310 10364
rect 3310 10308 3314 10364
rect 3250 10304 3314 10308
rect 3330 10364 3394 10368
rect 3330 10308 3334 10364
rect 3334 10308 3390 10364
rect 3390 10308 3394 10364
rect 3330 10304 3394 10308
rect 3410 10364 3474 10368
rect 3410 10308 3414 10364
rect 3414 10308 3470 10364
rect 3470 10308 3474 10364
rect 3410 10304 3474 10308
rect 3490 10364 3554 10368
rect 3490 10308 3494 10364
rect 3494 10308 3550 10364
rect 3550 10308 3554 10364
rect 3490 10304 3554 10308
rect 7848 10364 7912 10368
rect 7848 10308 7852 10364
rect 7852 10308 7908 10364
rect 7908 10308 7912 10364
rect 7848 10304 7912 10308
rect 7928 10364 7992 10368
rect 7928 10308 7932 10364
rect 7932 10308 7988 10364
rect 7988 10308 7992 10364
rect 7928 10304 7992 10308
rect 8008 10364 8072 10368
rect 8008 10308 8012 10364
rect 8012 10308 8068 10364
rect 8068 10308 8072 10364
rect 8008 10304 8072 10308
rect 8088 10364 8152 10368
rect 8088 10308 8092 10364
rect 8092 10308 8148 10364
rect 8148 10308 8152 10364
rect 8088 10304 8152 10308
rect 12445 10364 12509 10368
rect 12445 10308 12449 10364
rect 12449 10308 12505 10364
rect 12505 10308 12509 10364
rect 12445 10304 12509 10308
rect 12525 10364 12589 10368
rect 12525 10308 12529 10364
rect 12529 10308 12585 10364
rect 12585 10308 12589 10364
rect 12525 10304 12589 10308
rect 12605 10364 12669 10368
rect 12605 10308 12609 10364
rect 12609 10308 12665 10364
rect 12665 10308 12669 10364
rect 12605 10304 12669 10308
rect 12685 10364 12749 10368
rect 12685 10308 12689 10364
rect 12689 10308 12745 10364
rect 12745 10308 12749 10364
rect 12685 10304 12749 10308
rect 5549 9820 5613 9824
rect 5549 9764 5553 9820
rect 5553 9764 5609 9820
rect 5609 9764 5613 9820
rect 5549 9760 5613 9764
rect 5629 9820 5693 9824
rect 5629 9764 5633 9820
rect 5633 9764 5689 9820
rect 5689 9764 5693 9820
rect 5629 9760 5693 9764
rect 5709 9820 5773 9824
rect 5709 9764 5713 9820
rect 5713 9764 5769 9820
rect 5769 9764 5773 9820
rect 5709 9760 5773 9764
rect 5789 9820 5853 9824
rect 5789 9764 5793 9820
rect 5793 9764 5849 9820
rect 5849 9764 5853 9820
rect 5789 9760 5853 9764
rect 10146 9820 10210 9824
rect 10146 9764 10150 9820
rect 10150 9764 10206 9820
rect 10206 9764 10210 9820
rect 10146 9760 10210 9764
rect 10226 9820 10290 9824
rect 10226 9764 10230 9820
rect 10230 9764 10286 9820
rect 10286 9764 10290 9820
rect 10226 9760 10290 9764
rect 10306 9820 10370 9824
rect 10306 9764 10310 9820
rect 10310 9764 10366 9820
rect 10366 9764 10370 9820
rect 10306 9760 10370 9764
rect 10386 9820 10450 9824
rect 10386 9764 10390 9820
rect 10390 9764 10446 9820
rect 10446 9764 10450 9820
rect 10386 9760 10450 9764
rect 3250 9276 3314 9280
rect 3250 9220 3254 9276
rect 3254 9220 3310 9276
rect 3310 9220 3314 9276
rect 3250 9216 3314 9220
rect 3330 9276 3394 9280
rect 3330 9220 3334 9276
rect 3334 9220 3390 9276
rect 3390 9220 3394 9276
rect 3330 9216 3394 9220
rect 3410 9276 3474 9280
rect 3410 9220 3414 9276
rect 3414 9220 3470 9276
rect 3470 9220 3474 9276
rect 3410 9216 3474 9220
rect 3490 9276 3554 9280
rect 3490 9220 3494 9276
rect 3494 9220 3550 9276
rect 3550 9220 3554 9276
rect 3490 9216 3554 9220
rect 7848 9276 7912 9280
rect 7848 9220 7852 9276
rect 7852 9220 7908 9276
rect 7908 9220 7912 9276
rect 7848 9216 7912 9220
rect 7928 9276 7992 9280
rect 7928 9220 7932 9276
rect 7932 9220 7988 9276
rect 7988 9220 7992 9276
rect 7928 9216 7992 9220
rect 8008 9276 8072 9280
rect 8008 9220 8012 9276
rect 8012 9220 8068 9276
rect 8068 9220 8072 9276
rect 8008 9216 8072 9220
rect 8088 9276 8152 9280
rect 8088 9220 8092 9276
rect 8092 9220 8148 9276
rect 8148 9220 8152 9276
rect 8088 9216 8152 9220
rect 12445 9276 12509 9280
rect 12445 9220 12449 9276
rect 12449 9220 12505 9276
rect 12505 9220 12509 9276
rect 12445 9216 12509 9220
rect 12525 9276 12589 9280
rect 12525 9220 12529 9276
rect 12529 9220 12585 9276
rect 12585 9220 12589 9276
rect 12525 9216 12589 9220
rect 12605 9276 12669 9280
rect 12605 9220 12609 9276
rect 12609 9220 12665 9276
rect 12665 9220 12669 9276
rect 12605 9216 12669 9220
rect 12685 9276 12749 9280
rect 12685 9220 12689 9276
rect 12689 9220 12745 9276
rect 12745 9220 12749 9276
rect 12685 9216 12749 9220
rect 5549 8732 5613 8736
rect 5549 8676 5553 8732
rect 5553 8676 5609 8732
rect 5609 8676 5613 8732
rect 5549 8672 5613 8676
rect 5629 8732 5693 8736
rect 5629 8676 5633 8732
rect 5633 8676 5689 8732
rect 5689 8676 5693 8732
rect 5629 8672 5693 8676
rect 5709 8732 5773 8736
rect 5709 8676 5713 8732
rect 5713 8676 5769 8732
rect 5769 8676 5773 8732
rect 5709 8672 5773 8676
rect 5789 8732 5853 8736
rect 5789 8676 5793 8732
rect 5793 8676 5849 8732
rect 5849 8676 5853 8732
rect 5789 8672 5853 8676
rect 10146 8732 10210 8736
rect 10146 8676 10150 8732
rect 10150 8676 10206 8732
rect 10206 8676 10210 8732
rect 10146 8672 10210 8676
rect 10226 8732 10290 8736
rect 10226 8676 10230 8732
rect 10230 8676 10286 8732
rect 10286 8676 10290 8732
rect 10226 8672 10290 8676
rect 10306 8732 10370 8736
rect 10306 8676 10310 8732
rect 10310 8676 10366 8732
rect 10366 8676 10370 8732
rect 10306 8672 10370 8676
rect 10386 8732 10450 8736
rect 10386 8676 10390 8732
rect 10390 8676 10446 8732
rect 10446 8676 10450 8732
rect 10386 8672 10450 8676
rect 3250 8188 3314 8192
rect 3250 8132 3254 8188
rect 3254 8132 3310 8188
rect 3310 8132 3314 8188
rect 3250 8128 3314 8132
rect 3330 8188 3394 8192
rect 3330 8132 3334 8188
rect 3334 8132 3390 8188
rect 3390 8132 3394 8188
rect 3330 8128 3394 8132
rect 3410 8188 3474 8192
rect 3410 8132 3414 8188
rect 3414 8132 3470 8188
rect 3470 8132 3474 8188
rect 3410 8128 3474 8132
rect 3490 8188 3554 8192
rect 3490 8132 3494 8188
rect 3494 8132 3550 8188
rect 3550 8132 3554 8188
rect 3490 8128 3554 8132
rect 7848 8188 7912 8192
rect 7848 8132 7852 8188
rect 7852 8132 7908 8188
rect 7908 8132 7912 8188
rect 7848 8128 7912 8132
rect 7928 8188 7992 8192
rect 7928 8132 7932 8188
rect 7932 8132 7988 8188
rect 7988 8132 7992 8188
rect 7928 8128 7992 8132
rect 8008 8188 8072 8192
rect 8008 8132 8012 8188
rect 8012 8132 8068 8188
rect 8068 8132 8072 8188
rect 8008 8128 8072 8132
rect 8088 8188 8152 8192
rect 8088 8132 8092 8188
rect 8092 8132 8148 8188
rect 8148 8132 8152 8188
rect 8088 8128 8152 8132
rect 12445 8188 12509 8192
rect 12445 8132 12449 8188
rect 12449 8132 12505 8188
rect 12505 8132 12509 8188
rect 12445 8128 12509 8132
rect 12525 8188 12589 8192
rect 12525 8132 12529 8188
rect 12529 8132 12585 8188
rect 12585 8132 12589 8188
rect 12525 8128 12589 8132
rect 12605 8188 12669 8192
rect 12605 8132 12609 8188
rect 12609 8132 12665 8188
rect 12665 8132 12669 8188
rect 12605 8128 12669 8132
rect 12685 8188 12749 8192
rect 12685 8132 12689 8188
rect 12689 8132 12745 8188
rect 12745 8132 12749 8188
rect 12685 8128 12749 8132
rect 5549 7644 5613 7648
rect 5549 7588 5553 7644
rect 5553 7588 5609 7644
rect 5609 7588 5613 7644
rect 5549 7584 5613 7588
rect 5629 7644 5693 7648
rect 5629 7588 5633 7644
rect 5633 7588 5689 7644
rect 5689 7588 5693 7644
rect 5629 7584 5693 7588
rect 5709 7644 5773 7648
rect 5709 7588 5713 7644
rect 5713 7588 5769 7644
rect 5769 7588 5773 7644
rect 5709 7584 5773 7588
rect 5789 7644 5853 7648
rect 5789 7588 5793 7644
rect 5793 7588 5849 7644
rect 5849 7588 5853 7644
rect 5789 7584 5853 7588
rect 10146 7644 10210 7648
rect 10146 7588 10150 7644
rect 10150 7588 10206 7644
rect 10206 7588 10210 7644
rect 10146 7584 10210 7588
rect 10226 7644 10290 7648
rect 10226 7588 10230 7644
rect 10230 7588 10286 7644
rect 10286 7588 10290 7644
rect 10226 7584 10290 7588
rect 10306 7644 10370 7648
rect 10306 7588 10310 7644
rect 10310 7588 10366 7644
rect 10366 7588 10370 7644
rect 10306 7584 10370 7588
rect 10386 7644 10450 7648
rect 10386 7588 10390 7644
rect 10390 7588 10446 7644
rect 10446 7588 10450 7644
rect 10386 7584 10450 7588
rect 3250 7100 3314 7104
rect 3250 7044 3254 7100
rect 3254 7044 3310 7100
rect 3310 7044 3314 7100
rect 3250 7040 3314 7044
rect 3330 7100 3394 7104
rect 3330 7044 3334 7100
rect 3334 7044 3390 7100
rect 3390 7044 3394 7100
rect 3330 7040 3394 7044
rect 3410 7100 3474 7104
rect 3410 7044 3414 7100
rect 3414 7044 3470 7100
rect 3470 7044 3474 7100
rect 3410 7040 3474 7044
rect 3490 7100 3554 7104
rect 3490 7044 3494 7100
rect 3494 7044 3550 7100
rect 3550 7044 3554 7100
rect 3490 7040 3554 7044
rect 7848 7100 7912 7104
rect 7848 7044 7852 7100
rect 7852 7044 7908 7100
rect 7908 7044 7912 7100
rect 7848 7040 7912 7044
rect 7928 7100 7992 7104
rect 7928 7044 7932 7100
rect 7932 7044 7988 7100
rect 7988 7044 7992 7100
rect 7928 7040 7992 7044
rect 8008 7100 8072 7104
rect 8008 7044 8012 7100
rect 8012 7044 8068 7100
rect 8068 7044 8072 7100
rect 8008 7040 8072 7044
rect 8088 7100 8152 7104
rect 8088 7044 8092 7100
rect 8092 7044 8148 7100
rect 8148 7044 8152 7100
rect 8088 7040 8152 7044
rect 12445 7100 12509 7104
rect 12445 7044 12449 7100
rect 12449 7044 12505 7100
rect 12505 7044 12509 7100
rect 12445 7040 12509 7044
rect 12525 7100 12589 7104
rect 12525 7044 12529 7100
rect 12529 7044 12585 7100
rect 12585 7044 12589 7100
rect 12525 7040 12589 7044
rect 12605 7100 12669 7104
rect 12605 7044 12609 7100
rect 12609 7044 12665 7100
rect 12665 7044 12669 7100
rect 12605 7040 12669 7044
rect 12685 7100 12749 7104
rect 12685 7044 12689 7100
rect 12689 7044 12745 7100
rect 12745 7044 12749 7100
rect 12685 7040 12749 7044
rect 5549 6556 5613 6560
rect 5549 6500 5553 6556
rect 5553 6500 5609 6556
rect 5609 6500 5613 6556
rect 5549 6496 5613 6500
rect 5629 6556 5693 6560
rect 5629 6500 5633 6556
rect 5633 6500 5689 6556
rect 5689 6500 5693 6556
rect 5629 6496 5693 6500
rect 5709 6556 5773 6560
rect 5709 6500 5713 6556
rect 5713 6500 5769 6556
rect 5769 6500 5773 6556
rect 5709 6496 5773 6500
rect 5789 6556 5853 6560
rect 5789 6500 5793 6556
rect 5793 6500 5849 6556
rect 5849 6500 5853 6556
rect 5789 6496 5853 6500
rect 10146 6556 10210 6560
rect 10146 6500 10150 6556
rect 10150 6500 10206 6556
rect 10206 6500 10210 6556
rect 10146 6496 10210 6500
rect 10226 6556 10290 6560
rect 10226 6500 10230 6556
rect 10230 6500 10286 6556
rect 10286 6500 10290 6556
rect 10226 6496 10290 6500
rect 10306 6556 10370 6560
rect 10306 6500 10310 6556
rect 10310 6500 10366 6556
rect 10366 6500 10370 6556
rect 10306 6496 10370 6500
rect 10386 6556 10450 6560
rect 10386 6500 10390 6556
rect 10390 6500 10446 6556
rect 10446 6500 10450 6556
rect 10386 6496 10450 6500
rect 3250 6012 3314 6016
rect 3250 5956 3254 6012
rect 3254 5956 3310 6012
rect 3310 5956 3314 6012
rect 3250 5952 3314 5956
rect 3330 6012 3394 6016
rect 3330 5956 3334 6012
rect 3334 5956 3390 6012
rect 3390 5956 3394 6012
rect 3330 5952 3394 5956
rect 3410 6012 3474 6016
rect 3410 5956 3414 6012
rect 3414 5956 3470 6012
rect 3470 5956 3474 6012
rect 3410 5952 3474 5956
rect 3490 6012 3554 6016
rect 3490 5956 3494 6012
rect 3494 5956 3550 6012
rect 3550 5956 3554 6012
rect 3490 5952 3554 5956
rect 7848 6012 7912 6016
rect 7848 5956 7852 6012
rect 7852 5956 7908 6012
rect 7908 5956 7912 6012
rect 7848 5952 7912 5956
rect 7928 6012 7992 6016
rect 7928 5956 7932 6012
rect 7932 5956 7988 6012
rect 7988 5956 7992 6012
rect 7928 5952 7992 5956
rect 8008 6012 8072 6016
rect 8008 5956 8012 6012
rect 8012 5956 8068 6012
rect 8068 5956 8072 6012
rect 8008 5952 8072 5956
rect 8088 6012 8152 6016
rect 8088 5956 8092 6012
rect 8092 5956 8148 6012
rect 8148 5956 8152 6012
rect 8088 5952 8152 5956
rect 12445 6012 12509 6016
rect 12445 5956 12449 6012
rect 12449 5956 12505 6012
rect 12505 5956 12509 6012
rect 12445 5952 12509 5956
rect 12525 6012 12589 6016
rect 12525 5956 12529 6012
rect 12529 5956 12585 6012
rect 12585 5956 12589 6012
rect 12525 5952 12589 5956
rect 12605 6012 12669 6016
rect 12605 5956 12609 6012
rect 12609 5956 12665 6012
rect 12665 5956 12669 6012
rect 12605 5952 12669 5956
rect 12685 6012 12749 6016
rect 12685 5956 12689 6012
rect 12689 5956 12745 6012
rect 12745 5956 12749 6012
rect 12685 5952 12749 5956
rect 5549 5468 5613 5472
rect 5549 5412 5553 5468
rect 5553 5412 5609 5468
rect 5609 5412 5613 5468
rect 5549 5408 5613 5412
rect 5629 5468 5693 5472
rect 5629 5412 5633 5468
rect 5633 5412 5689 5468
rect 5689 5412 5693 5468
rect 5629 5408 5693 5412
rect 5709 5468 5773 5472
rect 5709 5412 5713 5468
rect 5713 5412 5769 5468
rect 5769 5412 5773 5468
rect 5709 5408 5773 5412
rect 5789 5468 5853 5472
rect 5789 5412 5793 5468
rect 5793 5412 5849 5468
rect 5849 5412 5853 5468
rect 5789 5408 5853 5412
rect 10146 5468 10210 5472
rect 10146 5412 10150 5468
rect 10150 5412 10206 5468
rect 10206 5412 10210 5468
rect 10146 5408 10210 5412
rect 10226 5468 10290 5472
rect 10226 5412 10230 5468
rect 10230 5412 10286 5468
rect 10286 5412 10290 5468
rect 10226 5408 10290 5412
rect 10306 5468 10370 5472
rect 10306 5412 10310 5468
rect 10310 5412 10366 5468
rect 10366 5412 10370 5468
rect 10306 5408 10370 5412
rect 10386 5468 10450 5472
rect 10386 5412 10390 5468
rect 10390 5412 10446 5468
rect 10446 5412 10450 5468
rect 10386 5408 10450 5412
rect 3250 4924 3314 4928
rect 3250 4868 3254 4924
rect 3254 4868 3310 4924
rect 3310 4868 3314 4924
rect 3250 4864 3314 4868
rect 3330 4924 3394 4928
rect 3330 4868 3334 4924
rect 3334 4868 3390 4924
rect 3390 4868 3394 4924
rect 3330 4864 3394 4868
rect 3410 4924 3474 4928
rect 3410 4868 3414 4924
rect 3414 4868 3470 4924
rect 3470 4868 3474 4924
rect 3410 4864 3474 4868
rect 3490 4924 3554 4928
rect 3490 4868 3494 4924
rect 3494 4868 3550 4924
rect 3550 4868 3554 4924
rect 3490 4864 3554 4868
rect 7848 4924 7912 4928
rect 7848 4868 7852 4924
rect 7852 4868 7908 4924
rect 7908 4868 7912 4924
rect 7848 4864 7912 4868
rect 7928 4924 7992 4928
rect 7928 4868 7932 4924
rect 7932 4868 7988 4924
rect 7988 4868 7992 4924
rect 7928 4864 7992 4868
rect 8008 4924 8072 4928
rect 8008 4868 8012 4924
rect 8012 4868 8068 4924
rect 8068 4868 8072 4924
rect 8008 4864 8072 4868
rect 8088 4924 8152 4928
rect 8088 4868 8092 4924
rect 8092 4868 8148 4924
rect 8148 4868 8152 4924
rect 8088 4864 8152 4868
rect 12445 4924 12509 4928
rect 12445 4868 12449 4924
rect 12449 4868 12505 4924
rect 12505 4868 12509 4924
rect 12445 4864 12509 4868
rect 12525 4924 12589 4928
rect 12525 4868 12529 4924
rect 12529 4868 12585 4924
rect 12585 4868 12589 4924
rect 12525 4864 12589 4868
rect 12605 4924 12669 4928
rect 12605 4868 12609 4924
rect 12609 4868 12665 4924
rect 12665 4868 12669 4924
rect 12605 4864 12669 4868
rect 12685 4924 12749 4928
rect 12685 4868 12689 4924
rect 12689 4868 12745 4924
rect 12745 4868 12749 4924
rect 12685 4864 12749 4868
rect 5549 4380 5613 4384
rect 5549 4324 5553 4380
rect 5553 4324 5609 4380
rect 5609 4324 5613 4380
rect 5549 4320 5613 4324
rect 5629 4380 5693 4384
rect 5629 4324 5633 4380
rect 5633 4324 5689 4380
rect 5689 4324 5693 4380
rect 5629 4320 5693 4324
rect 5709 4380 5773 4384
rect 5709 4324 5713 4380
rect 5713 4324 5769 4380
rect 5769 4324 5773 4380
rect 5709 4320 5773 4324
rect 5789 4380 5853 4384
rect 5789 4324 5793 4380
rect 5793 4324 5849 4380
rect 5849 4324 5853 4380
rect 5789 4320 5853 4324
rect 10146 4380 10210 4384
rect 10146 4324 10150 4380
rect 10150 4324 10206 4380
rect 10206 4324 10210 4380
rect 10146 4320 10210 4324
rect 10226 4380 10290 4384
rect 10226 4324 10230 4380
rect 10230 4324 10286 4380
rect 10286 4324 10290 4380
rect 10226 4320 10290 4324
rect 10306 4380 10370 4384
rect 10306 4324 10310 4380
rect 10310 4324 10366 4380
rect 10366 4324 10370 4380
rect 10306 4320 10370 4324
rect 10386 4380 10450 4384
rect 10386 4324 10390 4380
rect 10390 4324 10446 4380
rect 10446 4324 10450 4380
rect 10386 4320 10450 4324
rect 3250 3836 3314 3840
rect 3250 3780 3254 3836
rect 3254 3780 3310 3836
rect 3310 3780 3314 3836
rect 3250 3776 3314 3780
rect 3330 3836 3394 3840
rect 3330 3780 3334 3836
rect 3334 3780 3390 3836
rect 3390 3780 3394 3836
rect 3330 3776 3394 3780
rect 3410 3836 3474 3840
rect 3410 3780 3414 3836
rect 3414 3780 3470 3836
rect 3470 3780 3474 3836
rect 3410 3776 3474 3780
rect 3490 3836 3554 3840
rect 3490 3780 3494 3836
rect 3494 3780 3550 3836
rect 3550 3780 3554 3836
rect 3490 3776 3554 3780
rect 7848 3836 7912 3840
rect 7848 3780 7852 3836
rect 7852 3780 7908 3836
rect 7908 3780 7912 3836
rect 7848 3776 7912 3780
rect 7928 3836 7992 3840
rect 7928 3780 7932 3836
rect 7932 3780 7988 3836
rect 7988 3780 7992 3836
rect 7928 3776 7992 3780
rect 8008 3836 8072 3840
rect 8008 3780 8012 3836
rect 8012 3780 8068 3836
rect 8068 3780 8072 3836
rect 8008 3776 8072 3780
rect 8088 3836 8152 3840
rect 8088 3780 8092 3836
rect 8092 3780 8148 3836
rect 8148 3780 8152 3836
rect 8088 3776 8152 3780
rect 12445 3836 12509 3840
rect 12445 3780 12449 3836
rect 12449 3780 12505 3836
rect 12505 3780 12509 3836
rect 12445 3776 12509 3780
rect 12525 3836 12589 3840
rect 12525 3780 12529 3836
rect 12529 3780 12585 3836
rect 12585 3780 12589 3836
rect 12525 3776 12589 3780
rect 12605 3836 12669 3840
rect 12605 3780 12609 3836
rect 12609 3780 12665 3836
rect 12665 3780 12669 3836
rect 12605 3776 12669 3780
rect 12685 3836 12749 3840
rect 12685 3780 12689 3836
rect 12689 3780 12745 3836
rect 12745 3780 12749 3836
rect 12685 3776 12749 3780
rect 5549 3292 5613 3296
rect 5549 3236 5553 3292
rect 5553 3236 5609 3292
rect 5609 3236 5613 3292
rect 5549 3232 5613 3236
rect 5629 3292 5693 3296
rect 5629 3236 5633 3292
rect 5633 3236 5689 3292
rect 5689 3236 5693 3292
rect 5629 3232 5693 3236
rect 5709 3292 5773 3296
rect 5709 3236 5713 3292
rect 5713 3236 5769 3292
rect 5769 3236 5773 3292
rect 5709 3232 5773 3236
rect 5789 3292 5853 3296
rect 5789 3236 5793 3292
rect 5793 3236 5849 3292
rect 5849 3236 5853 3292
rect 5789 3232 5853 3236
rect 10146 3292 10210 3296
rect 10146 3236 10150 3292
rect 10150 3236 10206 3292
rect 10206 3236 10210 3292
rect 10146 3232 10210 3236
rect 10226 3292 10290 3296
rect 10226 3236 10230 3292
rect 10230 3236 10286 3292
rect 10286 3236 10290 3292
rect 10226 3232 10290 3236
rect 10306 3292 10370 3296
rect 10306 3236 10310 3292
rect 10310 3236 10366 3292
rect 10366 3236 10370 3292
rect 10306 3232 10370 3236
rect 10386 3292 10450 3296
rect 10386 3236 10390 3292
rect 10390 3236 10446 3292
rect 10446 3236 10450 3292
rect 10386 3232 10450 3236
rect 3250 2748 3314 2752
rect 3250 2692 3254 2748
rect 3254 2692 3310 2748
rect 3310 2692 3314 2748
rect 3250 2688 3314 2692
rect 3330 2748 3394 2752
rect 3330 2692 3334 2748
rect 3334 2692 3390 2748
rect 3390 2692 3394 2748
rect 3330 2688 3394 2692
rect 3410 2748 3474 2752
rect 3410 2692 3414 2748
rect 3414 2692 3470 2748
rect 3470 2692 3474 2748
rect 3410 2688 3474 2692
rect 3490 2748 3554 2752
rect 3490 2692 3494 2748
rect 3494 2692 3550 2748
rect 3550 2692 3554 2748
rect 3490 2688 3554 2692
rect 7848 2748 7912 2752
rect 7848 2692 7852 2748
rect 7852 2692 7908 2748
rect 7908 2692 7912 2748
rect 7848 2688 7912 2692
rect 7928 2748 7992 2752
rect 7928 2692 7932 2748
rect 7932 2692 7988 2748
rect 7988 2692 7992 2748
rect 7928 2688 7992 2692
rect 8008 2748 8072 2752
rect 8008 2692 8012 2748
rect 8012 2692 8068 2748
rect 8068 2692 8072 2748
rect 8008 2688 8072 2692
rect 8088 2748 8152 2752
rect 8088 2692 8092 2748
rect 8092 2692 8148 2748
rect 8148 2692 8152 2748
rect 8088 2688 8152 2692
rect 12445 2748 12509 2752
rect 12445 2692 12449 2748
rect 12449 2692 12505 2748
rect 12505 2692 12509 2748
rect 12445 2688 12509 2692
rect 12525 2748 12589 2752
rect 12525 2692 12529 2748
rect 12529 2692 12585 2748
rect 12585 2692 12589 2748
rect 12525 2688 12589 2692
rect 12605 2748 12669 2752
rect 12605 2692 12609 2748
rect 12609 2692 12665 2748
rect 12665 2692 12669 2748
rect 12605 2688 12669 2692
rect 12685 2748 12749 2752
rect 12685 2692 12689 2748
rect 12689 2692 12745 2748
rect 12745 2692 12749 2748
rect 12685 2688 12749 2692
rect 5549 2204 5613 2208
rect 5549 2148 5553 2204
rect 5553 2148 5609 2204
rect 5609 2148 5613 2204
rect 5549 2144 5613 2148
rect 5629 2204 5693 2208
rect 5629 2148 5633 2204
rect 5633 2148 5689 2204
rect 5689 2148 5693 2204
rect 5629 2144 5693 2148
rect 5709 2204 5773 2208
rect 5709 2148 5713 2204
rect 5713 2148 5769 2204
rect 5769 2148 5773 2204
rect 5709 2144 5773 2148
rect 5789 2204 5853 2208
rect 5789 2148 5793 2204
rect 5793 2148 5849 2204
rect 5849 2148 5853 2204
rect 5789 2144 5853 2148
rect 10146 2204 10210 2208
rect 10146 2148 10150 2204
rect 10150 2148 10206 2204
rect 10206 2148 10210 2204
rect 10146 2144 10210 2148
rect 10226 2204 10290 2208
rect 10226 2148 10230 2204
rect 10230 2148 10286 2204
rect 10286 2148 10290 2204
rect 10226 2144 10290 2148
rect 10306 2204 10370 2208
rect 10306 2148 10310 2204
rect 10310 2148 10366 2204
rect 10366 2148 10370 2204
rect 10306 2144 10370 2148
rect 10386 2204 10450 2208
rect 10386 2148 10390 2204
rect 10390 2148 10446 2204
rect 10446 2148 10450 2204
rect 10386 2144 10450 2148
<< metal4 >>
rect 3242 13632 3563 13648
rect 3242 13568 3250 13632
rect 3314 13568 3330 13632
rect 3394 13568 3410 13632
rect 3474 13568 3490 13632
rect 3554 13568 3563 13632
rect 3242 12544 3563 13568
rect 3242 12480 3250 12544
rect 3314 12480 3330 12544
rect 3394 12480 3410 12544
rect 3474 12480 3490 12544
rect 3554 12480 3563 12544
rect 3242 11456 3563 12480
rect 3242 11392 3250 11456
rect 3314 11392 3330 11456
rect 3394 11392 3410 11456
rect 3474 11392 3490 11456
rect 3554 11392 3563 11456
rect 3242 10368 3563 11392
rect 3242 10304 3250 10368
rect 3314 10304 3330 10368
rect 3394 10304 3410 10368
rect 3474 10304 3490 10368
rect 3554 10304 3563 10368
rect 3242 9280 3563 10304
rect 3242 9216 3250 9280
rect 3314 9216 3330 9280
rect 3394 9216 3410 9280
rect 3474 9216 3490 9280
rect 3554 9216 3563 9280
rect 3242 8192 3563 9216
rect 3242 8128 3250 8192
rect 3314 8128 3330 8192
rect 3394 8128 3410 8192
rect 3474 8128 3490 8192
rect 3554 8128 3563 8192
rect 3242 7104 3563 8128
rect 3242 7040 3250 7104
rect 3314 7040 3330 7104
rect 3394 7040 3410 7104
rect 3474 7040 3490 7104
rect 3554 7040 3563 7104
rect 3242 6016 3563 7040
rect 3242 5952 3250 6016
rect 3314 5952 3330 6016
rect 3394 5952 3410 6016
rect 3474 5952 3490 6016
rect 3554 5952 3563 6016
rect 3242 4928 3563 5952
rect 3242 4864 3250 4928
rect 3314 4864 3330 4928
rect 3394 4864 3410 4928
rect 3474 4864 3490 4928
rect 3554 4864 3563 4928
rect 3242 3840 3563 4864
rect 3242 3776 3250 3840
rect 3314 3776 3330 3840
rect 3394 3776 3410 3840
rect 3474 3776 3490 3840
rect 3554 3776 3563 3840
rect 3242 2752 3563 3776
rect 3242 2688 3250 2752
rect 3314 2688 3330 2752
rect 3394 2688 3410 2752
rect 3474 2688 3490 2752
rect 3554 2688 3563 2752
rect 3242 2128 3563 2688
rect 5541 13088 5861 13648
rect 5541 13024 5549 13088
rect 5613 13024 5629 13088
rect 5693 13024 5709 13088
rect 5773 13024 5789 13088
rect 5853 13024 5861 13088
rect 5541 12000 5861 13024
rect 5541 11936 5549 12000
rect 5613 11936 5629 12000
rect 5693 11936 5709 12000
rect 5773 11936 5789 12000
rect 5853 11936 5861 12000
rect 5541 10912 5861 11936
rect 5541 10848 5549 10912
rect 5613 10848 5629 10912
rect 5693 10848 5709 10912
rect 5773 10848 5789 10912
rect 5853 10848 5861 10912
rect 5541 9824 5861 10848
rect 5541 9760 5549 9824
rect 5613 9760 5629 9824
rect 5693 9760 5709 9824
rect 5773 9760 5789 9824
rect 5853 9760 5861 9824
rect 5541 8736 5861 9760
rect 5541 8672 5549 8736
rect 5613 8672 5629 8736
rect 5693 8672 5709 8736
rect 5773 8672 5789 8736
rect 5853 8672 5861 8736
rect 5541 7648 5861 8672
rect 5541 7584 5549 7648
rect 5613 7584 5629 7648
rect 5693 7584 5709 7648
rect 5773 7584 5789 7648
rect 5853 7584 5861 7648
rect 5541 6560 5861 7584
rect 5541 6496 5549 6560
rect 5613 6496 5629 6560
rect 5693 6496 5709 6560
rect 5773 6496 5789 6560
rect 5853 6496 5861 6560
rect 5541 5472 5861 6496
rect 5541 5408 5549 5472
rect 5613 5408 5629 5472
rect 5693 5408 5709 5472
rect 5773 5408 5789 5472
rect 5853 5408 5861 5472
rect 5541 4384 5861 5408
rect 5541 4320 5549 4384
rect 5613 4320 5629 4384
rect 5693 4320 5709 4384
rect 5773 4320 5789 4384
rect 5853 4320 5861 4384
rect 5541 3296 5861 4320
rect 5541 3232 5549 3296
rect 5613 3232 5629 3296
rect 5693 3232 5709 3296
rect 5773 3232 5789 3296
rect 5853 3232 5861 3296
rect 5541 2208 5861 3232
rect 5541 2144 5549 2208
rect 5613 2144 5629 2208
rect 5693 2144 5709 2208
rect 5773 2144 5789 2208
rect 5853 2144 5861 2208
rect 5541 2128 5861 2144
rect 7840 13632 8160 13648
rect 7840 13568 7848 13632
rect 7912 13568 7928 13632
rect 7992 13568 8008 13632
rect 8072 13568 8088 13632
rect 8152 13568 8160 13632
rect 7840 12544 8160 13568
rect 7840 12480 7848 12544
rect 7912 12480 7928 12544
rect 7992 12480 8008 12544
rect 8072 12480 8088 12544
rect 8152 12480 8160 12544
rect 7840 11456 8160 12480
rect 7840 11392 7848 11456
rect 7912 11392 7928 11456
rect 7992 11392 8008 11456
rect 8072 11392 8088 11456
rect 8152 11392 8160 11456
rect 7840 10368 8160 11392
rect 7840 10304 7848 10368
rect 7912 10304 7928 10368
rect 7992 10304 8008 10368
rect 8072 10304 8088 10368
rect 8152 10304 8160 10368
rect 7840 9280 8160 10304
rect 7840 9216 7848 9280
rect 7912 9216 7928 9280
rect 7992 9216 8008 9280
rect 8072 9216 8088 9280
rect 8152 9216 8160 9280
rect 7840 8192 8160 9216
rect 7840 8128 7848 8192
rect 7912 8128 7928 8192
rect 7992 8128 8008 8192
rect 8072 8128 8088 8192
rect 8152 8128 8160 8192
rect 7840 7104 8160 8128
rect 7840 7040 7848 7104
rect 7912 7040 7928 7104
rect 7992 7040 8008 7104
rect 8072 7040 8088 7104
rect 8152 7040 8160 7104
rect 7840 6016 8160 7040
rect 7840 5952 7848 6016
rect 7912 5952 7928 6016
rect 7992 5952 8008 6016
rect 8072 5952 8088 6016
rect 8152 5952 8160 6016
rect 7840 4928 8160 5952
rect 7840 4864 7848 4928
rect 7912 4864 7928 4928
rect 7992 4864 8008 4928
rect 8072 4864 8088 4928
rect 8152 4864 8160 4928
rect 7840 3840 8160 4864
rect 7840 3776 7848 3840
rect 7912 3776 7928 3840
rect 7992 3776 8008 3840
rect 8072 3776 8088 3840
rect 8152 3776 8160 3840
rect 7840 2752 8160 3776
rect 7840 2688 7848 2752
rect 7912 2688 7928 2752
rect 7992 2688 8008 2752
rect 8072 2688 8088 2752
rect 8152 2688 8160 2752
rect 7840 2128 8160 2688
rect 10138 13088 10458 13648
rect 10138 13024 10146 13088
rect 10210 13024 10226 13088
rect 10290 13024 10306 13088
rect 10370 13024 10386 13088
rect 10450 13024 10458 13088
rect 10138 12000 10458 13024
rect 10138 11936 10146 12000
rect 10210 11936 10226 12000
rect 10290 11936 10306 12000
rect 10370 11936 10386 12000
rect 10450 11936 10458 12000
rect 10138 10912 10458 11936
rect 10138 10848 10146 10912
rect 10210 10848 10226 10912
rect 10290 10848 10306 10912
rect 10370 10848 10386 10912
rect 10450 10848 10458 10912
rect 10138 9824 10458 10848
rect 10138 9760 10146 9824
rect 10210 9760 10226 9824
rect 10290 9760 10306 9824
rect 10370 9760 10386 9824
rect 10450 9760 10458 9824
rect 10138 8736 10458 9760
rect 10138 8672 10146 8736
rect 10210 8672 10226 8736
rect 10290 8672 10306 8736
rect 10370 8672 10386 8736
rect 10450 8672 10458 8736
rect 10138 7648 10458 8672
rect 10138 7584 10146 7648
rect 10210 7584 10226 7648
rect 10290 7584 10306 7648
rect 10370 7584 10386 7648
rect 10450 7584 10458 7648
rect 10138 6560 10458 7584
rect 10138 6496 10146 6560
rect 10210 6496 10226 6560
rect 10290 6496 10306 6560
rect 10370 6496 10386 6560
rect 10450 6496 10458 6560
rect 10138 5472 10458 6496
rect 10138 5408 10146 5472
rect 10210 5408 10226 5472
rect 10290 5408 10306 5472
rect 10370 5408 10386 5472
rect 10450 5408 10458 5472
rect 10138 4384 10458 5408
rect 10138 4320 10146 4384
rect 10210 4320 10226 4384
rect 10290 4320 10306 4384
rect 10370 4320 10386 4384
rect 10450 4320 10458 4384
rect 10138 3296 10458 4320
rect 10138 3232 10146 3296
rect 10210 3232 10226 3296
rect 10290 3232 10306 3296
rect 10370 3232 10386 3296
rect 10450 3232 10458 3296
rect 10138 2208 10458 3232
rect 10138 2144 10146 2208
rect 10210 2144 10226 2208
rect 10290 2144 10306 2208
rect 10370 2144 10386 2208
rect 10450 2144 10458 2208
rect 10138 2128 10458 2144
rect 12437 13632 12757 13648
rect 12437 13568 12445 13632
rect 12509 13568 12525 13632
rect 12589 13568 12605 13632
rect 12669 13568 12685 13632
rect 12749 13568 12757 13632
rect 12437 12544 12757 13568
rect 12437 12480 12445 12544
rect 12509 12480 12525 12544
rect 12589 12480 12605 12544
rect 12669 12480 12685 12544
rect 12749 12480 12757 12544
rect 12437 11456 12757 12480
rect 12437 11392 12445 11456
rect 12509 11392 12525 11456
rect 12589 11392 12605 11456
rect 12669 11392 12685 11456
rect 12749 11392 12757 11456
rect 12437 10368 12757 11392
rect 12437 10304 12445 10368
rect 12509 10304 12525 10368
rect 12589 10304 12605 10368
rect 12669 10304 12685 10368
rect 12749 10304 12757 10368
rect 12437 9280 12757 10304
rect 12437 9216 12445 9280
rect 12509 9216 12525 9280
rect 12589 9216 12605 9280
rect 12669 9216 12685 9280
rect 12749 9216 12757 9280
rect 12437 8192 12757 9216
rect 12437 8128 12445 8192
rect 12509 8128 12525 8192
rect 12589 8128 12605 8192
rect 12669 8128 12685 8192
rect 12749 8128 12757 8192
rect 12437 7104 12757 8128
rect 12437 7040 12445 7104
rect 12509 7040 12525 7104
rect 12589 7040 12605 7104
rect 12669 7040 12685 7104
rect 12749 7040 12757 7104
rect 12437 6016 12757 7040
rect 12437 5952 12445 6016
rect 12509 5952 12525 6016
rect 12589 5952 12605 6016
rect 12669 5952 12685 6016
rect 12749 5952 12757 6016
rect 12437 4928 12757 5952
rect 12437 4864 12445 4928
rect 12509 4864 12525 4928
rect 12589 4864 12605 4928
rect 12669 4864 12685 4928
rect 12749 4864 12757 4928
rect 12437 3840 12757 4864
rect 12437 3776 12445 3840
rect 12509 3776 12525 3840
rect 12589 3776 12605 3840
rect 12669 3776 12685 3840
rect 12749 3776 12757 3840
rect 12437 2752 12757 3776
rect 12437 2688 12445 2752
rect 12509 2688 12525 2752
rect 12589 2688 12605 2752
rect 12669 2688 12685 2752
rect 12749 2688 12757 2752
rect 12437 2128 12757 2688
use sky130_fd_sc_hd__decap_8  FILLER_0_15 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 2484 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 3220 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 1380 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_15 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 2484 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_3
timestamp 1636915332
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1636915332
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1636915332
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtn_1  _448_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 2576 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__diode_2  ANTENNA__448__RESET_B $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 3864 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input3_A
timestamp 1636915332
transform -1 0 3680 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29
timestamp 1636915332
transform 1 0 3772 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_48
timestamp 1636915332
transform 1 0 5520 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_42 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__dfrtp_1  _453_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 4416 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__buf_12  input3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 4048 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__a21bo_1  _288_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform -1 0 7084 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_47
timestamp 1636915332
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_43
timestamp 1636915332
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_59
timestamp 1636915332
transform 1 0 6532 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__453__RESET_B
timestamp 1636915332
transform 1 0 6348 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__nor2_1  _360_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform -1 0 8004 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _274_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 7176 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_1_65
timestamp 1636915332
transform 1 0 7084 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_69
timestamp 1636915332
transform 1 0 7452 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__451__RESET_B
timestamp 1636915332
transform 1 0 7268 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__dfrtp_2  _451_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 7452 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__xor2_1  _361_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 8004 0 1 2176
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _340_
timestamp 1636915332
transform -1 0 9292 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_44
timestamp 1636915332
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_85
timestamp 1636915332
transform 1 0 8924 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_82 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 8648 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__nand3b_1  _341_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 9568 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _320_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform -1 0 9568 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _319_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 10120 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__445__RESET_B
timestamp 1636915332
transform 1 0 9384 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__dfrtp_1  _445_
timestamp 1636915332
transform 1 0 9568 0 1 2176
box -38 -48 1878 592
use sky130_fd_sc_hd__fill_1  FILLER_1_107
timestamp 1636915332
transform 1 0 10948 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_45
timestamp 1636915332
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_48
timestamp 1636915332
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _275_
timestamp 1636915332
transform 1 0 11500 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_1  _317_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform -1 0 11408 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__xor2_1  _318_
timestamp 1636915332
transform 1 0 11500 0 1 2176
box -38 -48 682 592
use sky130_fd_sc_hd__dfrtp_1  _446_
timestamp 1636915332
transform 1 0 12144 0 1 2176
box -38 -48 1878 592
use sky130_fd_sc_hd__buf_6  input1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform -1 0 12604 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__446__RESET_B
timestamp 1636915332
transform -1 0 14536 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_1_145
timestamp 1636915332
transform 1 0 14444 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1636915332
transform -1 0 14812 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1636915332
transform -1 0 14812 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_46
timestamp 1636915332
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _374_
timestamp 1636915332
transform 1 0 14076 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  _427_
timestamp 1636915332
transform -1 0 14444 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__diode_2  ANTENNA__449__SET_B
timestamp 1636915332
transform 1 0 2484 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_2_21
timestamp 1636915332
transform 1 0 3036 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_3
timestamp 1636915332
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1636915332
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__o21bai_1  _295_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 3128 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _303_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform -1 0 3036 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_49
timestamp 1636915332
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _280_
timestamp 1636915332
transform 1 0 5060 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _293_
timestamp 1636915332
transform 1 0 5336 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__nand3b_1  _296_
timestamp 1636915332
transform -1 0 5060 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__a21bo_1  _304_
timestamp 1636915332
transform -1 0 4508 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dfstp_1  _452_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 5612 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  _399_
timestamp 1636915332
transform 1 0 7544 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_2_83
timestamp 1636915332
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_94
timestamp 1636915332
transform 1 0 9752 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_50
timestamp 1636915332
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__nand3_1  _276_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform -1 0 8740 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _362_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 9844 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _363_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 10212 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _398_
timestamp 1636915332
transform 1 0 8924 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__427__RESET_B
timestamp 1636915332
transform 1 0 11684 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  _403_
timestamp 1636915332
transform 1 0 10856 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__dfrtp_4  _430_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform -1 0 13984 0 1 3264
box -38 -48 2154 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input1_A
timestamp 1636915332
transform -1 0 14260 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input7_A
timestamp 1636915332
transform -1 0 14536 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_2_143
timestamp 1636915332
transform 1 0 14260 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1636915332
transform -1 0 14812 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_51
timestamp 1636915332
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1636915332
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__o2bb2ai_1  _300_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 3312 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__dfstp_1  _449_
timestamp 1636915332
transform 1 0 1380 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__o21ai_1  _282_
timestamp 1636915332
transform -1 0 5980 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _294_
timestamp 1636915332
transform -1 0 4784 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _302_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform -1 0 4508 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _397_
timestamp 1636915332
transform 1 0 4784 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__452__SET_B
timestamp 1636915332
transform 1 0 5980 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_3_55
timestamp 1636915332
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_3_69
timestamp 1636915332
transform 1 0 7452 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_52
timestamp 1636915332
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__nand3_1  _287_
timestamp 1636915332
transform -1 0 7452 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__a21bo_1  _290_
timestamp 1636915332
transform 1 0 6348 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__a21bo_1  _292_
timestamp 1636915332
transform 1 0 7544 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__clkinv_2  _358_
timestamp 1636915332
transform 1 0 9936 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _404_
timestamp 1636915332
transform 1 0 9108 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _405_
timestamp 1636915332
transform 1 0 8280 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__428__SET_B
timestamp 1636915332
transform 1 0 12328 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__430__RESET_B
timestamp 1636915332
transform 1 0 11224 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_3_100
timestamp 1636915332
transform 1 0 10304 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_53
timestamp 1636915332
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _321_
timestamp 1636915332
transform 1 0 10396 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _400_
timestamp 1636915332
transform 1 0 11500 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__dfstp_1  _428_
timestamp 1636915332
transform -1 0 14444 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__fill_1  FILLER_3_145
timestamp 1636915332
transform 1 0 14444 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1636915332
transform -1 0 14812 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1636915332
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _297_
timestamp 1636915332
transform 1 0 3220 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtn_1  _450_
timestamp 1636915332
transform 1 0 1380 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__diode_2  ANTENNA__440__RESET_B
timestamp 1636915332
transform 1 0 3496 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_4_32
timestamp 1636915332
transform 1 0 4048 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_43
timestamp 1636915332
transform 1 0 5060 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_54
timestamp 1636915332
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _281_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 5612 0 1 4352
box -38 -48 958 592
use sky130_fd_sc_hd__nand2_2  _286_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 5152 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _298_
timestamp 1636915332
transform -1 0 4048 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__o211ai_1  _314_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform -1 0 5060 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_1_0_0_pll_clk $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform -1 0 4508 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__444__SET_B
timestamp 1636915332
transform 1 0 6900 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  _283_
timestamp 1636915332
transform 1 0 6532 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _359_
timestamp 1636915332
transform 1 0 7912 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _402_
timestamp 1636915332
transform 1 0 7084 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_4_94
timestamp 1636915332
transform 1 0 9752 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_55
timestamp 1636915332
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _345_
timestamp 1636915332
transform 1 0 8556 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _401_
timestamp 1636915332
transform 1 0 8924 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__dfstp_1  _444_
timestamp 1636915332
transform 1 0 9844 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__dfstp_4  _431_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform -1 0 13984 0 1 4352
box -38 -48 2246 592
use sky130_fd_sc_hd__diode_2  ANTENNA__431__SET_B
timestamp 1636915332
transform 1 0 14076 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1636915332
transform -1 0 14812 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_56
timestamp 1636915332
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp 1636915332
transform 1 0 14260 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__450__RESET_B
timestamp 1636915332
transform -1 0 2300 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_5_3
timestamp 1636915332
transform 1 0 1380 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_7 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 1748 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1636915332
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _299_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 3128 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _301__4
timestamp 1636915332
transform -1 0 1748 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _313_
timestamp 1636915332
transform -1 0 3128 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _337_
timestamp 1636915332
transform -1 0 2852 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _338_
timestamp 1636915332
transform 1 0 2300 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_5_25
timestamp 1636915332
transform 1 0 3404 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_5_38
timestamp 1636915332
transform 1 0 4600 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_1  _306_
timestamp 1636915332
transform 1 0 3496 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__o21bai_1  _315_
timestamp 1636915332
transform -1 0 5612 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _316_
timestamp 1636915332
transform 1 0 4692 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _330_
timestamp 1636915332
transform -1 0 5888 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _385_
timestamp 1636915332
transform 1 0 3772 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_57
timestamp 1636915332
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__nand3_1  _289_
timestamp 1636915332
transform 1 0 5888 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _307_
timestamp 1636915332
transform -1 0 6624 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _327_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 6624 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_pll_clk $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 7084 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__o21bai_1  _284_
timestamp 1636915332
transform -1 0 9476 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _322_
timestamp 1636915332
transform -1 0 9752 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _349_
timestamp 1636915332
transform 1 0 9752 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_58
timestamp 1636915332
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__nand3_1  _285_
timestamp 1636915332
transform -1 0 10764 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _342_
timestamp 1636915332
transform 1 0 10764 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _364_
timestamp 1636915332
transform -1 0 12604 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _411_
timestamp 1636915332
transform 1 0 11500 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1636915332
transform -1 0 14812 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__dfstp_1  _439_
timestamp 1636915332
transform 1 0 12604 0 -1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1636915332
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1636915332
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__nand3_1  _312_
timestamp 1636915332
transform -1 0 3588 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _339_
timestamp 1636915332
transform -1 0 3588 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__dfrtn_1  _440_
timestamp 1636915332
transform 1 0 1380 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtn_1  _442_
timestamp 1636915332
transform 1 0 1380 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__mux2_1  _386_
timestamp 1636915332
transform 1 0 3588 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _331_
timestamp 1636915332
transform -1 0 4692 0 1 5440
box -38 -48 958 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_59
timestamp 1636915332
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp 1636915332
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _407_
timestamp 1636915332
transform 1 0 4784 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _382_
timestamp 1636915332
transform 1 0 4692 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _332_
timestamp 1636915332
transform -1 0 4692 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_6_39
timestamp 1636915332
transform 1 0 4692 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__nand3_1  _309_
timestamp 1636915332
transform -1 0 5888 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__447__SET_B
timestamp 1636915332
transform 1 0 5612 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_7_55
timestamp 1636915332
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_62
timestamp 1636915332
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__nand3b_1  _279_
timestamp 1636915332
transform 1 0 7728 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _291_
timestamp 1636915332
transform 1 0 7176 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _305__5
timestamp 1636915332
transform 1 0 5888 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _406_
timestamp 1636915332
transform 1 0 6348 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__dfrtp_4  _443_
timestamp 1636915332
transform 1 0 7544 0 -1 6528
box -38 -48 2154 592
use sky130_fd_sc_hd__dfstp_1  _447_
timestamp 1636915332
transform 1 0 5796 0 1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_60
timestamp 1636915332
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _277_
timestamp 1636915332
transform -1 0 9936 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _278_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 8280 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _414_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 9936 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfstp_1  _454_
timestamp 1636915332
transform -1 0 10856 0 1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__diode_2  ANTENNA__424__RESET_B
timestamp 1636915332
transform 1 0 11500 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_6_119
timestamp 1636915332
transform 1 0 12052 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_63
timestamp 1636915332
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_1  _348_
timestamp 1636915332
transform -1 0 11960 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__o21bai_2  _351_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform -1 0 11684 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__dfrtp_1  _424_
timestamp 1636915332
transform -1 0 13800 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _429_
timestamp 1636915332
transform -1 0 13984 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_1_1_0_pll_clk
timestamp 1636915332
transform 1 0 11684 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__429__RESET_B
timestamp 1636915332
transform 1 0 14076 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__439__SET_B
timestamp 1636915332
transform 1 0 13800 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input4_A
timestamp 1636915332
transform -1 0 14536 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input5_A
timestamp 1636915332
transform -1 0 14352 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input8_A
timestamp 1636915332
transform -1 0 14168 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1636915332
transform -1 0 14812 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1636915332
transform -1 0 14812 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_61
timestamp 1636915332
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input8
timestamp 1636915332
transform 1 0 14260 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_8_17
timestamp 1636915332
transform 1 0 2668 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_8_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 1380 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_9
timestamp 1636915332
transform 1 0 1932 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1636915332
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _310_
timestamp 1636915332
transform -1 0 3036 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _333_
timestamp 1636915332
transform -1 0 2668 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _335_
timestamp 1636915332
transform 1 0 2024 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _357_
timestamp 1636915332
transform 1 0 3036 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__fill_1  FILLER_8_42
timestamp 1636915332
transform 1 0 4968 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_64
timestamp 1636915332
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__nor3b_2  _308_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 3772 0 1 6528
box -38 -48 958 592
use sky130_fd_sc_hd__inv_2  _311_
timestamp 1636915332
transform 1 0 4692 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _381_
timestamp 1636915332
transform 1 0 5060 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_8_52
timestamp 1636915332
transform 1 0 5888 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_1  _326_
timestamp 1636915332
transform 1 0 7452 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _329_
timestamp 1636915332
transform 1 0 7728 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _416_
timestamp 1636915332
transform 1 0 5980 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA__443__RESET_B
timestamp 1636915332
transform 1 0 8280 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__454__SET_B
timestamp 1636915332
transform 1 0 8924 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_0_pll_clk_A
timestamp 1636915332
transform -1 0 8648 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input9_A
timestamp 1636915332
transform -1 0 8832 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_8_87
timestamp 1636915332
transform 1 0 9108 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_65
timestamp 1636915332
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _415_
timestamp 1636915332
transform 1 0 9200 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_8_104
timestamp 1636915332
transform 1 0 10672 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_8_116
timestamp 1636915332
transform 1 0 11776 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__nand3_1  _325_
timestamp 1636915332
transform -1 0 11776 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__and2b_2  _350_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform -1 0 11408 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__dfrtp_4  _432_
timestamp 1636915332
transform -1 0 13984 0 1 6528
box -38 -48 2154 592
use sky130_fd_sc_hd__diode_2  ANTENNA__432__RESET_B
timestamp 1636915332
transform 1 0 14076 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1636915332
transform -1 0 14812 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_66
timestamp 1636915332
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input9
timestamp 1636915332
transform 1 0 14260 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_9_3
timestamp 1636915332
transform 1 0 1380 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1636915332
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__dfstp_1  _441_
timestamp 1636915332
transform 1 0 1932 0 -1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__fill_1  FILLER_9_30
timestamp 1636915332
transform 1 0 3864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_41
timestamp 1636915332
transform 1 0 4876 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__xnor2_1  _355_
timestamp 1636915332
transform 1 0 3956 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _356_
timestamp 1636915332
transform 1 0 4600 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__470__RESET_B
timestamp 1636915332
transform 1 0 6624 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_9_53
timestamp 1636915332
transform 1 0 5980 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_57
timestamp 1636915332
transform 1 0 6348 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_9_70
timestamp 1636915332
transform 1 0 7544 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_67
timestamp 1636915332
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__o21ai_1  _328_
timestamp 1636915332
transform 1 0 7176 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__nor3_1  _376_
timestamp 1636915332
transform -1 0 7176 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__dfrtp_1  _470_
timestamp 1636915332
transform -1 0 9476 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__fill_1  FILLER_9_91
timestamp 1636915332
transform 1 0 9476 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__or2b_1  _323_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 10120 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _324_
timestamp 1636915332
transform 1 0 9568 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_68
timestamp 1636915332
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__dfrtp_1  _426_
timestamp 1636915332
transform -1 0 13340 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform -1 0 11408 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_142
timestamp 1636915332
transform 1 0 14168 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1636915332
transform -1 0 14812 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _394_
timestamp 1636915332
transform 1 0 13340 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp 1636915332
transform 1 0 14260 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__442__RESET_B
timestamp 1636915332
transform 1 0 3220 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_13
timestamp 1636915332
transform 1 0 2300 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_19
timestamp 1636915332
transform 1 0 2852 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_10_3
timestamp 1636915332
transform 1 0 1380 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_9
timestamp 1636915332
transform 1 0 1932 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1636915332
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _334__6
timestamp 1636915332
transform -1 0 2300 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _336_
timestamp 1636915332
transform -1 0 2852 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__441__SET_B
timestamp 1636915332
transform 1 0 3864 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__468__SET_B
timestamp 1636915332
transform 1 0 5244 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_10_25
timestamp 1636915332
transform 1 0 3404 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_10_29
timestamp 1636915332
transform 1 0 3772 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_32
timestamp 1636915332
transform 1 0 4048 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_44
timestamp 1636915332
transform 1 0 5152 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_69
timestamp 1636915332
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__dfstp_1  _468_
timestamp 1636915332
transform 1 0 5428 0 1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__nor3b_2  _268_
timestamp 1636915332
transform 1 0 7360 0 1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__diode_2  ANTENNA__426__RESET_B
timestamp 1636915332
transform 1 0 10120 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__455__SET_B
timestamp 1636915332
transform 1 0 8648 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_78
timestamp 1636915332
transform 1 0 8280 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_97
timestamp 1636915332
transform 1 0 10028 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_70
timestamp 1636915332
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _270_
timestamp 1636915332
transform -1 0 10028 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _271_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform -1 0 9476 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _273_
timestamp 1636915332
transform -1 0 9752 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__343__S
timestamp 1636915332
transform 1 0 11776 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__425__RESET_B
timestamp 1636915332
transform 1 0 11960 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  _420_
timestamp 1636915332
transform 1 0 10304 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfrtp_1  _425_
timestamp 1636915332
transform 1 0 12144 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__diode_2  ANTENNA__433__RESET_B
timestamp 1636915332
transform 1 0 14076 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1636915332
transform -1 0 14812 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_71
timestamp 1636915332
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 1636915332
transform 1 0 14260 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_11_15
timestamp 1636915332
transform 1 0 2484 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_11_3
timestamp 1636915332
transform 1 0 1380 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1636915332
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtn_1  _460_
timestamp 1636915332
transform -1 0 4692 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__diode_2  ANTENNA__460__RESET_B
timestamp 1636915332
transform 1 0 5336 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_11_42
timestamp 1636915332
transform 1 0 4968 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_48
timestamp 1636915332
transform 1 0 5520 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  _205_
timestamp 1636915332
transform 1 0 5060 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _235_
timestamp 1636915332
transform -1 0 4968 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__469__RESET_B
timestamp 1636915332
transform 1 0 5704 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_11_55
timestamp 1636915332
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_72
timestamp 1636915332
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _206_
timestamp 1636915332
transform 1 0 6348 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _207_
timestamp 1636915332
transform 1 0 5888 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _373_
timestamp 1636915332
transform 1 0 7176 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _377_
timestamp 1636915332
transform 1 0 7820 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__nand3_1  _272_
timestamp 1636915332
transform -1 0 8832 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__dfstp_1  _455_
timestamp 1636915332
transform 1 0 8832 0 -1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_73
timestamp 1636915332
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_2  _343_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 11500 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _344_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform -1 0 11040 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _368_
timestamp 1636915332
transform -1 0 12696 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_1_0_0_ext_clk
timestamp 1636915332
transform 1 0 11040 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1636915332
transform -1 0 14812 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  _433_
timestamp 1636915332
transform -1 0 14536 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__fill_2  FILLER_12_15
timestamp 1636915332
transform 1 0 2484 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_12_21
timestamp 1636915332
transform 1 0 3036 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_3
timestamp 1636915332
transform 1 0 1380 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1636915332
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _239_
timestamp 1636915332
transform -1 0 3404 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _244_
timestamp 1636915332
transform -1 0 3036 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__461__SET_B
timestamp 1636915332
transform 1 0 3404 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_12_27
timestamp 1636915332
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_37
timestamp 1636915332
transform 1 0 4508 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_74
timestamp 1636915332
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__a21bo_1  _245_
timestamp 1636915332
transform -1 0 4508 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dfrtp_1  _469_
timestamp 1636915332
transform 1 0 4600 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__mux2_1  _204_
timestamp 1636915332
transform 1 0 6440 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _410_
timestamp 1636915332
transform 1 0 7268 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__463__RESET_B
timestamp 1636915332
transform 1 0 8924 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_12_80
timestamp 1636915332
transform 1 0 8464 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_75
timestamp 1636915332
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _269_
timestamp 1636915332
transform 1 0 8556 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _372_
timestamp 1636915332
transform 1 0 8096 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _413_
timestamp 1636915332
transform 1 0 9108 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__dfrtp_2  _463_
timestamp 1636915332
transform 1 0 9936 0 1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _436_
timestamp 1636915332
transform -1 0 13984 0 1 8704
box -38 -48 2154 592
use sky130_fd_sc_hd__diode_2  ANTENNA__436__RESET_B
timestamp 1636915332
transform -1 0 14536 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1636915332
transform -1 0 14812 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_76
timestamp 1636915332
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _347_
timestamp 1636915332
transform 1 0 14076 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_13_24
timestamp 1636915332
transform 1 0 3312 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1636915332
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1636915332
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _238_
timestamp 1636915332
transform 1 0 3220 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__dfstp_1  _461_
timestamp 1636915332
transform 1 0 1380 0 -1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtn_1  _462_
timestamp 1636915332
transform 1 0 1380 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__and2b_1  _243_
timestamp 1636915332
transform -1 0 3956 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__o2bb2ai_1  _241_
timestamp 1636915332
transform 1 0 3772 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__o21bai_1  _236_
timestamp 1636915332
transform 1 0 3956 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_79
timestamp 1636915332
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__462__RESET_B
timestamp 1636915332
transform 1 0 3496 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__o211ai_1  _255_
timestamp 1636915332
transform -1 0 5428 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__nand3b_1  _237_
timestamp 1636915332
transform 1 0 4508 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _234_
timestamp 1636915332
transform -1 0 4692 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_13_43
timestamp 1636915332
transform 1 0 5060 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_0_pll_clk90_A
timestamp 1636915332
transform 1 0 4692 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  _390_
timestamp 1636915332
transform 1 0 5336 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _216_
timestamp 1636915332
transform 1 0 5428 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_13_55
timestamp 1636915332
transform 1 0 6164 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_77
timestamp 1636915332
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__nand2_2  _217_
timestamp 1636915332
transform 1 0 6348 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _224_
timestamp 1636915332
transform 1 0 6808 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _247_
timestamp 1636915332
transform 1 0 7544 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _346_
timestamp 1636915332
transform -1 0 8096 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _387_
timestamp 1636915332
transform 1 0 7176 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_pll_clk90
timestamp 1636915332
transform 1 0 5704 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__nor2_1  _370_
timestamp 1636915332
transform -1 0 9108 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _353_
timestamp 1636915332
transform 1 0 8924 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _248_
timestamp 1636915332
transform -1 0 8740 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_2  _215_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform -1 0 8740 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_80
timestamp 1636915332
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_83
timestamp 1636915332
transform 1 0 8740 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_76
timestamp 1636915332
transform 1 0 8096 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_83
timestamp 1636915332
transform 1 0 8740 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_75
timestamp 1636915332
transform 1 0 8004 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__a21bo_1  _233_
timestamp 1636915332
transform 1 0 9568 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _225_
timestamp 1636915332
transform 1 0 10212 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__o2bb2ai_2  _354_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 9108 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_78
timestamp 1636915332
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__a21bo_1  _231_
timestamp 1636915332
transform 1 0 10304 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__nand3_1  _232_
timestamp 1636915332
transform -1 0 11868 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _352_
timestamp 1636915332
transform 1 0 11040 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _379_
timestamp 1636915332
transform 1 0 11868 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _380_
timestamp 1636915332
transform 1 0 11316 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _391_
timestamp 1636915332
transform 1 0 12144 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _412_
timestamp 1636915332
transform -1 0 11408 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__437__SET_B
timestamp 1636915332
transform 1 0 13800 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_14_141
timestamp 1636915332
transform 1 0 14076 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1636915332
transform -1 0 14812 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1636915332
transform -1 0 14812 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_81
timestamp 1636915332
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _393_
timestamp 1636915332
transform 1 0 12972 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_ext_clk
timestamp 1636915332
transform 1 0 12696 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_1_1_0_ext_clk
timestamp 1636915332
transform -1 0 14536 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_15_19
timestamp 1636915332
transform 1 0 2852 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_15_3
timestamp 1636915332
transform 1 0 1380 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_7
timestamp 1636915332
transform 1 0 1748 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1636915332
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _242__1
timestamp 1636915332
transform -1 0 1748 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_1_0_0_pll_clk90
timestamp 1636915332
transform -1 0 3496 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_44
timestamp 1636915332
transform 1 0 5152 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__nand2_1  _240_
timestamp 1636915332
transform 1 0 3496 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__nand3_1  _250_
timestamp 1636915332
transform 1 0 5336 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _254_
timestamp 1636915332
transform -1 0 4048 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _258_
timestamp 1636915332
transform 1 0 4048 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _384_
timestamp 1636915332
transform 1 0 4324 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__459__SET_B
timestamp 1636915332
transform 1 0 6348 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_82
timestamp 1636915332
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__o21bai_1  _256_
timestamp 1636915332
transform -1 0 6256 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__dfstp_1  _459_
timestamp 1636915332
transform 1 0 6532 0 -1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__diode_2  ANTENNA__464__SET_B
timestamp 1636915332
transform 1 0 9292 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_15_84
timestamp 1636915332
transform 1 0 8832 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__nand3_1  _227_
timestamp 1636915332
transform -1 0 9292 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__dfstp_1  _464_
timestamp 1636915332
transform 1 0 9476 0 -1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_1_1_0_pll_clk90
timestamp 1636915332
transform 1 0 8464 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_83
timestamp 1636915332
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _392_
timestamp 1636915332
transform 1 0 11500 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__dfstp_4  _437_
timestamp 1636915332
transform -1 0 14536 0 -1 10880
box -38 -48 2246 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1636915332
transform -1 0 14812 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_16_3
timestamp 1636915332
transform 1 0 1380 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_7
timestamp 1636915332
transform 1 0 1748 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1636915332
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtn_1  _456_
timestamp 1636915332
transform 1 0 1840 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_84
timestamp 1636915332
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _259_
timestamp 1636915332
transform 1 0 4140 0 1 10880
box -38 -48 958 592
use sky130_fd_sc_hd__o21ai_1  _267_
timestamp 1636915332
transform -1 0 4140 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _383_
timestamp 1636915332
transform 1 0 5060 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__466__SET_B
timestamp 1636915332
transform 1 0 5980 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_16_52
timestamp 1636915332
transform 1 0 5888 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_59
timestamp 1636915332
transform 1 0 6532 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _246__2
timestamp 1636915332
transform -1 0 6900 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__nand3_1  _257_
timestamp 1636915332
transform -1 0 6532 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__dfstp_1  _466_
timestamp 1636915332
transform 1 0 6900 0 1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__fill_1  FILLER_16_97
timestamp 1636915332
transform 1 0 10028 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_85
timestamp 1636915332
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__nand3b_1  _223_
timestamp 1636915332
transform -1 0 9476 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__o21bai_1  _226_
timestamp 1636915332
transform 1 0 9476 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _230_
timestamp 1636915332
transform 1 0 10120 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_118
timestamp 1636915332
transform 1 0 11960 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__xor2_1  _371_
timestamp 1636915332
transform 1 0 10488 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _389_
timestamp 1636915332
transform 1 0 11132 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__dfstp_1  _434_
timestamp 1636915332
transform 1 0 12052 0 1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_0_ext_clk_A
timestamp 1636915332
transform -1 0 14536 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1636915332
transform -1 0 14812 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_86
timestamp 1636915332
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _220_
timestamp 1636915332
transform 1 0 14076 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_17_15
timestamp 1636915332
transform 1 0 2484 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_17_3
timestamp 1636915332
transform 1 0 1380 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1636915332
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _261_
timestamp 1636915332
transform -1 0 3588 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__456__RESET_B
timestamp 1636915332
transform 1 0 4048 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__458__RESET_B
timestamp 1636915332
transform 1 0 3588 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_17_34
timestamp 1636915332
transform 1 0 4232 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_17_44
timestamp 1636915332
transform 1 0 5152 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _260_
timestamp 1636915332
transform -1 0 4048 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _265_
timestamp 1636915332
transform -1 0 4600 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _266_
timestamp 1636915332
transform -1 0 4876 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _366_
timestamp 1636915332
transform 1 0 4876 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _395_
timestamp 1636915332
transform 1 0 5428 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_87
timestamp 1636915332
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__and2_1  _212_
timestamp 1636915332
transform 1 0 7820 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__dfxtp_1  _419_
timestamp 1636915332
transform 1 0 6348 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_17_82
timestamp 1636915332
transform 1 0 8648 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_17_95
timestamp 1636915332
transform 1 0 9844 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_1  _211_
timestamp 1636915332
transform -1 0 9568 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _213_
timestamp 1636915332
transform -1 0 9292 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _214_
timestamp 1636915332
transform -1 0 8648 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _222_
timestamp 1636915332
transform 1 0 9568 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__nand3_1  _228_
timestamp 1636915332
transform -1 0 10304 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__434__SET_B
timestamp 1636915332
transform 1 0 11500 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_88
timestamp 1636915332
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__nand3_1  _221_
timestamp 1636915332
transform 1 0 11040 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__a21bo_1  _229_
timestamp 1636915332
transform 1 0 10304 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _388_
timestamp 1636915332
transform 1 0 11684 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__dfrtp_1  _435_
timestamp 1636915332
transform 1 0 12512 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__fill_2  FILLER_17_144
timestamp 1636915332
transform 1 0 14352 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1636915332
transform -1 0 14812 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_18_3
timestamp 1636915332
transform 1 0 1380 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1636915332
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtn_1  _458_
timestamp 1636915332
transform 1 0 1748 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__fill_1  FILLER_18_27
timestamp 1636915332
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_18_36
timestamp 1636915332
transform 1 0 4416 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_89
timestamp 1636915332
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _251_
timestamp 1636915332
transform -1 0 4416 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__nand3_1  _253_
timestamp 1636915332
transform 1 0 3772 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__xor2_1  _367_
timestamp 1636915332
transform 1 0 4508 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _396_
timestamp 1636915332
transform 1 0 5152 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_18_53
timestamp 1636915332
transform 1 0 5980 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_18_71
timestamp 1636915332
transform 1 0 7636 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__or2b_1  _209_
timestamp 1636915332
transform 1 0 7728 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _418_
timestamp 1636915332
transform 1 0 6164 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA__423__SET_B
timestamp 1636915332
transform 1 0 9292 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__465__RESET_B
timestamp 1636915332
transform 1 0 9660 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__467__RESET_B
timestamp 1636915332
transform 1 0 8648 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_85
timestamp 1636915332
transform 1 0 8924 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_91
timestamp 1636915332
transform 1 0 9476 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_90
timestamp 1636915332
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__nand3_1  _210_
timestamp 1636915332
transform -1 0 8648 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__dfrtp_1  _465_
timestamp 1636915332
transform 1 0 9844 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__diode_2  ANTENNA__435__RESET_B
timestamp 1636915332
transform 1 0 11684 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__dfrtp_4  _438_
timestamp 1636915332
transform -1 0 13984 0 1 11968
box -38 -48 2154 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input2_A
timestamp 1636915332
transform -1 0 14260 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1636915332
transform -1 0 14812 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_91
timestamp 1636915332
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 1636915332
transform 1 0 14260 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_19_3
timestamp 1636915332
transform 1 0 1380 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_15
timestamp 1636915332
transform 1 0 2484 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_20_22
timestamp 1636915332
transform 1 0 3128 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_20_3
timestamp 1636915332
transform 1 0 1380 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1636915332
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1636915332
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _262__3
timestamp 1636915332
transform -1 0 2852 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__dfstp_1  _457_
timestamp 1636915332
transform 1 0 2484 0 -1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__clkbuf_1  output10
timestamp 1636915332
transform 1 0 2852 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _264_
timestamp 1636915332
transform -1 0 4140 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _252_
timestamp 1636915332
transform -1 0 4416 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_94
timestamp 1636915332
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _409_
timestamp 1636915332
transform 1 0 5152 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _263_
timestamp 1636915332
transform -1 0 4692 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__nor3b_2  _249_
timestamp 1636915332
transform 1 0 4508 0 -1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__decap_3  FILLER_20_41
timestamp 1636915332
transform 1 0 4876 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_19_36
timestamp 1636915332
transform 1 0 4416 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__457__SET_B
timestamp 1636915332
transform -1 0 4876 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  _408_
timestamp 1636915332
transform 1 0 5428 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_20_53
timestamp 1636915332
transform 1 0 5980 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_20_57
timestamp 1636915332
transform 1 0 6348 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_92
timestamp 1636915332
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_95
timestamp 1636915332
transform 1 0 6256 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__or2b_1  _208_
timestamp 1636915332
transform 1 0 7452 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _365_
timestamp 1636915332
transform -1 0 6992 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__dfxtp_1  _417_
timestamp 1636915332
transform 1 0 6992 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_20_75
timestamp 1636915332
transform 1 0 8004 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_20_83
timestamp 1636915332
transform 1 0 8740 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_96
timestamp 1636915332
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__o21a_1  _218_
timestamp 1636915332
transform -1 0 8740 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  _378__13 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 9200 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__dfstp_1  _423_
timestamp 1636915332
transform 1 0 9476 0 1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _467_
timestamp 1636915332
transform 1 0 8464 0 -1 13056
box -38 -48 2154 592
use sky130_fd_sc_hd__clkbuf_1  output12
timestamp 1636915332
transform 1 0 8924 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _219_
timestamp 1636915332
transform 1 0 11132 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input6_A
timestamp 1636915332
transform -1 0 10764 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__438__RESET_B
timestamp 1636915332
transform 1 0 10764 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__422__SET_B
timestamp 1636915332
transform 1 0 10948 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 1636915332
transform -1 0 12052 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_97
timestamp 1636915332
transform 1 0 11408 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_93
timestamp 1636915332
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_20_113
timestamp 1636915332
transform 1 0 11500 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__421__SET_B
timestamp 1636915332
transform -1 0 11776 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__dfstp_1  _422_
timestamp 1636915332
transform 1 0 11500 0 -1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__dfstp_1  _421_
timestamp 1636915332
transform 1 0 12052 0 1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__fill_2  FILLER_19_144
timestamp 1636915332
transform 1 0 14352 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_20_145
timestamp 1636915332
transform 1 0 14444 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1636915332
transform -1 0 14812 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1636915332
transform -1 0 14812 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_98
timestamp 1636915332
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__xnor2_1  _369_
timestamp 1636915332
transform -1 0 14076 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _375_
timestamp 1636915332
transform 1 0 14076 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output11 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 14076 0 1 13056
box -38 -48 406 592
<< labels >>
rlabel metal4 s 5541 2128 5861 13648 6 VGND
port 0 nsew ground input
rlabel metal4 s 10138 2128 10458 13648 6 VGND
port 0 nsew ground input
rlabel metal4 s 3243 2128 3563 13648 6 VPWR
port 1 nsew power input
rlabel metal4 s 7840 2128 8160 13648 6 VPWR
port 1 nsew power input
rlabel metal4 s 12437 2128 12757 13648 6 VPWR
port 1 nsew power input
rlabel metal2 s 2686 15200 2742 16000 6 core_clk
port 2 nsew signal tristate
rlabel metal2 s 11978 0 12034 800 6 ext_clk
port 3 nsew signal input
rlabel metal3 s 15200 960 16000 1080 6 ext_clk_sel
port 4 nsew signal input
rlabel metal3 s 15200 14968 16000 15088 6 ext_reset
port 5 nsew signal input
rlabel metal3 s 0 3952 800 4072 6 pll_clk
port 6 nsew signal input
rlabel metal3 s 0 11976 800 12096 6 pll_clk90
port 7 nsew signal input
rlabel metal2 s 3974 0 4030 800 6 resetb
port 8 nsew signal input
rlabel metal2 s 13358 15200 13414 16000 6 resetb_sync
port 9 nsew signal tristate
rlabel metal3 s 15200 8984 16000 9104 6 sel2[0]
port 10 nsew signal input
rlabel metal3 s 15200 10888 16000 11008 6 sel2[1]
port 11 nsew signal input
rlabel metal3 s 15200 12928 16000 13048 6 sel2[2]
port 12 nsew signal input
rlabel metal3 s 15200 2864 16000 2984 6 sel[0]
port 13 nsew signal input
rlabel metal3 s 15200 4904 16000 5024 6 sel[1]
port 14 nsew signal input
rlabel metal3 s 15200 6944 16000 7064 6 sel[2]
port 15 nsew signal input
rlabel metal2 s 8022 15200 8078 16000 6 user_clk
port 16 nsew signal tristate
<< properties >>
string FIXED_BBOX 0 0 16000 16000
<< end >>
