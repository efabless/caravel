VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO gpio_control_block
  CLASS BLOCK ;
  FOREIGN gpio_control_block ;
  ORIGIN 0.000 0.000 ;
  SIZE 170.000 BY 65.000 ;
  PIN gpio_defaults[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 4.690 61.000 4.970 65.000 ;
    END
  END gpio_defaults[0]
  PIN gpio_defaults[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 27.690 61.000 27.970 65.000 ;
    END
  END gpio_defaults[10]
  PIN gpio_defaults[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.990 61.000 30.270 65.000 ;
    END
  END gpio_defaults[11]
  PIN gpio_defaults[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.290 61.000 32.570 65.000 ;
    END
  END gpio_defaults[12]
  PIN gpio_defaults[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.990 61.000 7.270 65.000 ;
    END
  END gpio_defaults[1]
  PIN gpio_defaults[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 9.290 61.000 9.570 65.000 ;
    END
  END gpio_defaults[2]
  PIN gpio_defaults[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 11.590 61.000 11.870 65.000 ;
    END
  END gpio_defaults[3]
  PIN gpio_defaults[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 13.890 61.000 14.170 65.000 ;
    END
  END gpio_defaults[4]
  PIN gpio_defaults[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.190 61.000 16.470 65.000 ;
    END
  END gpio_defaults[5]
  PIN gpio_defaults[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 18.490 61.000 18.770 65.000 ;
    END
  END gpio_defaults[6]
  PIN gpio_defaults[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 20.790 61.000 21.070 65.000 ;
    END
  END gpio_defaults[7]
  PIN gpio_defaults[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 23.090 61.000 23.370 65.000 ;
    END
  END gpio_defaults[8]
  PIN gpio_defaults[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 25.390 61.000 25.670 65.000 ;
    END
  END gpio_defaults[9]
  PIN mgmt_gpio_in
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 70.000 4.120 170.000 4.720 ;
    END
  END mgmt_gpio_in
  PIN mgmt_gpio_oeb
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 70.000 8.200 170.000 8.800 ;
    END
  END mgmt_gpio_oeb
  PIN mgmt_gpio_out
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 70.000 10.240 170.000 10.840 ;
    END
  END mgmt_gpio_out
  PIN one
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 70.000 6.160 170.000 6.760 ;
    END
  END one
  PIN pad_gpio_ana_en
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 70.000 12.280 170.000 12.880 ;
    END
  END pad_gpio_ana_en
  PIN pad_gpio_ana_pol
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 70.000 14.320 170.000 14.920 ;
    END
  END pad_gpio_ana_pol
  PIN pad_gpio_ana_sel
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 70.000 16.360 170.000 16.960 ;
    END
  END pad_gpio_ana_sel
  PIN pad_gpio_dm[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 70.000 18.400 170.000 19.000 ;
    END
  END pad_gpio_dm[0]
  PIN pad_gpio_dm[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 70.000 20.440 170.000 21.040 ;
    END
  END pad_gpio_dm[1]
  PIN pad_gpio_dm[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 70.000 22.480 170.000 23.080 ;
    END
  END pad_gpio_dm[2]
  PIN pad_gpio_holdover
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 70.000 24.520 170.000 25.120 ;
    END
  END pad_gpio_holdover
  PIN pad_gpio_ib_mode_sel
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 70.000 26.560 170.000 27.160 ;
    END
  END pad_gpio_ib_mode_sel
  PIN pad_gpio_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 70.000 28.600 170.000 29.200 ;
    END
  END pad_gpio_in
  PIN pad_gpio_inenb
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 70.000 30.640 170.000 31.240 ;
    END
  END pad_gpio_inenb
  PIN pad_gpio_out
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 70.000 32.680 170.000 33.280 ;
    END
  END pad_gpio_out
  PIN pad_gpio_outenb
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 70.000 34.720 170.000 35.320 ;
    END
  END pad_gpio_outenb
  PIN pad_gpio_slow_sel
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 70.000 36.760 170.000 37.360 ;
    END
  END pad_gpio_slow_sel
  PIN pad_gpio_vtrip_sel
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 70.000 38.800 170.000 39.400 ;
    END
  END pad_gpio_vtrip_sel
  PIN resetn
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 70.000 40.840 170.000 41.440 ;
    END
  END resetn
  PIN resetn_out
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 70.000 42.880 170.000 43.480 ;
    END
  END resetn_out
  PIN serial_clock
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 70.000 44.920 170.000 45.520 ;
    END
  END serial_clock
  PIN serial_clock_out
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 70.000 46.960 170.000 47.560 ;
    END
  END serial_clock_out
  PIN serial_data_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 70.000 49.000 170.000 49.600 ;
    END
  END serial_data_in
  PIN serial_data_out
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 70.000 51.040 170.000 51.640 ;
    END
  END serial_data_out
  PIN serial_load
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 70.000 53.080 170.000 53.680 ;
    END
  END serial_load
  PIN serial_load_out
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 70.000 55.120 170.000 55.720 ;
    END
  END serial_load_out
  PIN user_gpio_in
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 70.000 57.160 170.000 57.760 ;
    END
  END user_gpio_in
  PIN user_gpio_oeb
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 70.000 59.200 170.000 59.800 ;
    END
  END user_gpio_oeb
  PIN user_gpio_out
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 70.000 61.240 170.000 61.840 ;
    END
  END user_gpio_out
  PIN vccd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 12.800 2.480 14.400 60.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 37.800 2.480 39.400 60.080 ;
    END
    PORT
      LAYER met5 ;
        RECT 4.360 5.900 50.000 7.500 ;
    END
    PORT
      LAYER met5 ;
        RECT 4.360 22.800 50.000 24.400 ;
    END
    PORT
      LAYER met5 ;
        RECT 4.360 39.700 50.000 41.300 ;
    END
    PORT
      LAYER met5 ;
        RECT 4.360 56.600 50.000 58.200 ;
    END
  END vccd
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 17.800 2.480 19.400 60.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 42.800 2.480 44.400 60.080 ;
    END
    PORT
      LAYER met5 ;
        RECT 4.360 11.140 50.000 12.740 ;
    END
    PORT
      LAYER met5 ;
        RECT 4.360 28.040 50.000 29.640 ;
    END
    PORT
      LAYER met5 ;
        RECT 4.360 44.940 50.000 46.540 ;
    END
  END vccd1
  PIN vssd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 25.300 2.480 26.900 60.080 ;
    END
    PORT
      LAYER met5 ;
        RECT 4.360 14.350 50.000 15.950 ;
    END
    PORT
      LAYER met5 ;
        RECT 4.360 31.250 50.000 32.850 ;
    END
    PORT
      LAYER met5 ;
        RECT 4.360 48.150 50.000 49.750 ;
    END
  END vssd
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 30.300 2.480 31.900 60.080 ;
    END
    PORT
      LAYER met5 ;
        RECT 4.360 19.590 50.000 21.190 ;
    END
    PORT
      LAYER met5 ;
        RECT 4.360 36.490 50.000 38.090 ;
    END
    PORT
      LAYER met5 ;
        RECT 4.360 53.390 50.000 54.990 ;
    END
  END vssd1
  PIN zero
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 70.000 2.080 170.000 2.680 ;
    END
  END zero
  OBS
      LAYER li1 ;
        RECT 4.600 2.635 51.980 59.925 ;
      LAYER met1 ;
        RECT 4.600 2.480 103.890 60.480 ;
      LAYER met2 ;
        RECT 5.250 60.720 6.710 61.725 ;
        RECT 7.550 60.720 9.010 61.725 ;
        RECT 9.850 60.720 11.310 61.725 ;
        RECT 12.150 60.720 13.610 61.725 ;
        RECT 14.450 60.720 15.910 61.725 ;
        RECT 16.750 60.720 18.210 61.725 ;
        RECT 19.050 60.720 20.510 61.725 ;
        RECT 21.350 60.720 22.810 61.725 ;
        RECT 23.650 60.720 25.110 61.725 ;
        RECT 25.950 60.720 27.410 61.725 ;
        RECT 28.250 60.720 29.710 61.725 ;
        RECT 30.550 60.720 32.010 61.725 ;
        RECT 32.850 60.720 103.870 61.725 ;
        RECT 4.970 2.195 103.870 60.720 ;
      LAYER met3 ;
        RECT 6.045 60.840 69.600 61.705 ;
        RECT 6.045 60.200 70.000 60.840 ;
        RECT 6.045 58.800 69.600 60.200 ;
        RECT 6.045 58.160 70.000 58.800 ;
        RECT 6.045 56.760 69.600 58.160 ;
        RECT 6.045 56.120 70.000 56.760 ;
        RECT 6.045 54.720 69.600 56.120 ;
        RECT 6.045 54.080 70.000 54.720 ;
        RECT 6.045 52.680 69.600 54.080 ;
        RECT 6.045 52.040 70.000 52.680 ;
        RECT 6.045 50.640 69.600 52.040 ;
        RECT 6.045 50.000 70.000 50.640 ;
        RECT 6.045 48.600 69.600 50.000 ;
        RECT 6.045 47.960 70.000 48.600 ;
        RECT 6.045 46.560 69.600 47.960 ;
        RECT 6.045 45.920 70.000 46.560 ;
        RECT 6.045 44.520 69.600 45.920 ;
        RECT 6.045 43.880 70.000 44.520 ;
        RECT 6.045 42.480 69.600 43.880 ;
        RECT 6.045 41.840 70.000 42.480 ;
        RECT 6.045 40.440 69.600 41.840 ;
        RECT 6.045 39.800 70.000 40.440 ;
        RECT 6.045 38.400 69.600 39.800 ;
        RECT 6.045 37.760 70.000 38.400 ;
        RECT 6.045 36.360 69.600 37.760 ;
        RECT 6.045 35.720 70.000 36.360 ;
        RECT 6.045 34.320 69.600 35.720 ;
        RECT 6.045 33.680 70.000 34.320 ;
        RECT 6.045 32.280 69.600 33.680 ;
        RECT 6.045 31.640 70.000 32.280 ;
        RECT 6.045 30.240 69.600 31.640 ;
        RECT 6.045 29.600 70.000 30.240 ;
        RECT 6.045 28.200 69.600 29.600 ;
        RECT 6.045 27.560 70.000 28.200 ;
        RECT 6.045 26.160 69.600 27.560 ;
        RECT 6.045 25.520 70.000 26.160 ;
        RECT 6.045 24.120 69.600 25.520 ;
        RECT 6.045 23.480 70.000 24.120 ;
        RECT 6.045 22.080 69.600 23.480 ;
        RECT 6.045 21.440 70.000 22.080 ;
        RECT 6.045 20.040 69.600 21.440 ;
        RECT 6.045 19.400 70.000 20.040 ;
        RECT 6.045 18.000 69.600 19.400 ;
        RECT 6.045 17.360 70.000 18.000 ;
        RECT 6.045 15.960 69.600 17.360 ;
        RECT 6.045 15.320 70.000 15.960 ;
        RECT 6.045 13.920 69.600 15.320 ;
        RECT 6.045 13.280 70.000 13.920 ;
        RECT 6.045 11.880 69.600 13.280 ;
        RECT 6.045 11.240 70.000 11.880 ;
        RECT 6.045 9.840 69.600 11.240 ;
        RECT 6.045 9.200 70.000 9.840 ;
        RECT 6.045 7.800 69.600 9.200 ;
        RECT 6.045 7.160 70.000 7.800 ;
        RECT 6.045 5.760 69.600 7.160 ;
        RECT 6.045 5.120 70.000 5.760 ;
        RECT 6.045 3.720 69.600 5.120 ;
        RECT 6.045 3.080 70.000 3.720 ;
        RECT 6.045 2.215 69.600 3.080 ;
      LAYER met4 ;
        RECT 6.280 8.160 12.400 52.185 ;
        RECT 14.800 8.160 17.400 52.185 ;
        RECT 19.800 8.160 24.900 52.185 ;
        RECT 27.300 8.160 29.900 52.185 ;
        RECT 32.300 8.160 37.400 52.185 ;
        RECT 39.800 8.160 42.400 52.185 ;
        RECT 44.800 8.160 45.705 52.185 ;
  END
END gpio_control_block
END LIBRARY

