magic
tech sky130A
magscale 1 2
timestamp 1637524495
<< error_p >>
rect 45056 221322 46138 221346
rect 45056 220272 45080 221322
rect 46114 220272 46138 221322
rect 45056 220248 46138 220272
rect 41362 219704 42444 219728
rect 41362 218654 41386 219704
rect 42420 218654 42444 219704
rect 41362 218630 42444 218654
rect 31080 218031 31834 218032
rect 31080 216955 31081 218031
rect 31833 216955 31834 218031
rect 31080 216954 31834 216955
rect 37618 216463 38380 216464
rect 37618 215381 37619 216463
rect 38379 215381 38380 216463
rect 37618 215380 38380 215381
<< metal3 >>
rect 6032 221346 46270 221382
rect 6032 221338 45056 221346
rect 6032 220224 6162 221338
rect 6862 220248 45056 221338
rect 46138 220248 46270 221346
rect 6862 220224 46270 220248
rect 6032 220182 46270 220224
rect 7246 219742 42526 219782
rect 7246 218628 7360 219742
rect 8060 219728 42526 219742
rect 8060 218630 41362 219728
rect 42444 218630 42526 219728
rect 8060 218628 42526 218630
rect 7246 218582 42526 218628
rect 17838 218068 31922 218100
rect 17838 216936 17896 218068
rect 18646 218032 31922 218068
rect 18646 216954 31080 218032
rect 31834 216954 31922 218032
rect 18646 216936 31922 216954
rect 17838 216900 31922 216936
rect 19032 216470 38512 216500
rect 19032 215338 19100 216470
rect 19850 216464 38512 216470
rect 19850 215380 37618 216464
rect 38380 215380 38512 216464
rect 19850 215338 38512 215380
rect 19032 215300 38512 215338
<< via3 >>
rect 6162 220224 6862 221338
rect 45056 220248 46138 221346
rect 7360 218628 8060 219742
rect 41362 218630 42444 219728
rect 17896 216936 18646 218068
rect 31080 216954 31834 218032
rect 19100 215338 19850 216470
rect 37618 215380 38380 216464
<< metal4 >>
rect 6116 221338 6916 221470
rect 6116 220224 6162 221338
rect 6862 220224 6916 221338
rect 6116 211874 6916 220224
rect 44994 221346 46200 221388
rect 44994 220248 45056 221346
rect 46138 220248 46200 221346
rect 44994 220174 46200 220248
rect 6116 211604 6132 211874
rect 6898 211604 6916 211874
rect 6116 208514 6916 211604
rect 6116 208244 6138 208514
rect 6904 208244 6916 208514
rect 6116 205138 6916 208244
rect 7316 219742 8116 219842
rect 7316 218628 7360 219742
rect 8060 218628 8116 219742
rect 7316 213570 8116 218628
rect 41290 219728 42496 219788
rect 41290 218630 41362 219728
rect 42444 218630 42496 219728
rect 41290 218574 42496 218630
rect 7316 213300 7334 213570
rect 8100 213300 8116 213570
rect 7316 210186 8116 213300
rect 7316 209916 7332 210186
rect 8098 209916 8116 210186
rect 7316 206826 8116 209916
rect 7316 206528 7326 206826
rect 8100 206528 8116 206826
rect 7316 206476 8116 206528
rect 17880 218068 18680 218110
rect 17880 216936 17896 218068
rect 18646 217338 18680 218068
rect 18656 217056 18680 217338
rect 18646 216936 18680 217056
rect 17880 212534 18680 216936
rect 17880 212246 17896 212534
rect 18668 212246 18680 212534
rect 17880 209152 18680 212246
rect 17880 208864 17890 209152
rect 18662 208864 18680 209152
rect 17880 205770 18680 208864
rect 17880 205482 17892 205770
rect 18664 205482 18680 205770
rect 17880 205422 18680 205482
rect 19080 216634 19880 216732
rect 19080 215338 19100 216634
rect 19856 216352 19880 216634
rect 19850 215338 19880 216352
rect 19080 210844 19880 215338
rect 19080 210556 19092 210844
rect 19864 210556 19880 210844
rect 19080 207464 19880 210556
rect 19080 207176 19096 207464
rect 19868 207176 19880 207464
rect 6116 204840 6132 205138
rect 6906 204840 6916 205138
rect 6116 204746 6916 204840
rect 19080 204084 19880 207176
rect 19080 203796 19096 204084
rect 19868 203796 19880 204084
rect 19080 203748 19880 203796
<< via4 >>
rect 45056 220248 46138 221346
rect 6132 211604 6898 211874
rect 6138 208244 6904 208514
rect 41362 218630 42444 219728
rect 7334 213300 8100 213570
rect 7332 209916 8098 210186
rect 7326 206528 8100 206826
rect 17900 217056 18646 217338
rect 18646 217056 18656 217338
rect 17896 212246 18668 212534
rect 17890 208864 18662 209152
rect 17892 205482 18664 205770
rect 19100 216470 19856 216634
rect 19100 216352 19850 216470
rect 19850 216352 19856 216470
rect 19092 210556 19864 210844
rect 19096 207176 19868 207464
rect 6132 204840 6906 205138
rect 19096 203796 19868 204084
<< metal5 >>
rect 17862 217356 18688 217368
rect 14320 217338 18688 217356
rect 14320 217056 17900 217338
rect 18656 217056 18688 217338
rect 14320 217036 18688 217056
rect 17862 217025 18688 217036
rect 19073 216656 19899 216671
rect 14320 216634 19932 216656
rect 14320 216352 19100 216634
rect 19856 216352 19932 216634
rect 14320 216336 19932 216352
rect 19073 216328 19899 216336
rect 7293 213598 8130 213615
rect 7270 213570 8592 213598
rect 7270 213300 7334 213570
rect 8100 213300 8592 213570
rect 7270 213278 8592 213300
rect 7293 213260 8130 213278
rect 17855 212550 18720 212570
rect 17434 212534 18720 212550
rect 17434 212246 17896 212534
rect 18668 212246 18720 212534
rect 17434 212230 18720 212246
rect 17855 212216 18720 212230
rect 6092 211908 6929 211924
rect 6058 211874 8592 211908
rect 6058 211604 6132 211874
rect 6898 211604 8592 211874
rect 6058 211588 8592 211604
rect 6092 211569 6929 211588
rect 19052 210860 19917 210872
rect 17434 210844 19917 210860
rect 17434 210556 19092 210844
rect 19864 210556 19917 210844
rect 17434 210540 19917 210556
rect 19052 210518 19917 210540
rect 7298 210218 8135 210241
rect 7276 210186 8592 210218
rect 7276 209916 7332 210186
rect 8098 209916 8592 210186
rect 7276 209898 8592 209916
rect 7298 209886 8135 209898
rect 17832 209170 18697 209187
rect 17434 209152 18697 209170
rect 17434 208864 17890 209152
rect 18662 208864 18697 209152
rect 17434 208850 18697 208864
rect 17832 208833 18697 208850
rect 6058 208528 6940 208550
rect 6058 208514 8592 208528
rect 6058 208244 6138 208514
rect 6904 208244 8592 208514
rect 6058 208228 8592 208244
rect 6059 208212 8592 208228
rect 6060 208208 8592 208212
rect 19051 207480 19916 207492
rect 17434 207464 19916 207480
rect 17434 207176 19096 207464
rect 19868 207176 19916 207464
rect 17434 207160 19916 207176
rect 19051 207138 19916 207160
rect 7298 206838 8134 206856
rect 7298 206826 8624 206838
rect 7298 206528 7326 206826
rect 8100 206528 8624 206826
rect 7298 206518 8624 206528
rect 7298 206496 8134 206518
rect 17851 205790 18716 205811
rect 17434 205770 18716 205790
rect 17434 205482 17892 205770
rect 18664 205482 18716 205770
rect 17434 205470 18716 205482
rect 17851 205457 18716 205470
rect 6104 205148 6941 205164
rect 6104 205138 8624 205148
rect 6104 204840 6132 205138
rect 6906 204840 8624 205138
rect 6104 204828 8624 204840
rect 6104 204809 6941 204828
rect 19045 204100 19910 204120
rect 17434 204084 19910 204100
rect 17434 203796 19096 204084
rect 19868 203796 19910 204084
rect 17434 203780 19910 203796
rect 19045 203766 19910 203780
<< end >>
