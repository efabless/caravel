* NGSPICE file created from caravel_clocking.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_1 abstract view
.subckt sky130_fd_sc_hd__dfrtp_1 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_2 abstract view
.subckt sky130_fd_sc_hd__nor3b_2 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_2 abstract view
.subckt sky130_fd_sc_hd__dfstp_2 CLK D SET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_1 abstract view
.subckt sky130_fd_sc_hd__nand2b_1 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4bb_1 abstract view
.subckt sky130_fd_sc_hd__nand4bb_1 A_N B_N C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_1 abstract view
.subckt sky130_fd_sc_hd__dfstp_1 CLK D SET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_2 abstract view
.subckt sky130_fd_sc_hd__dfrtp_2 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2ai_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2ai_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_12 abstract view
.subckt sky130_fd_sc_hd__buf_12 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111ai_2 abstract view
.subckt sky130_fd_sc_hd__o2111ai_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_2 abstract view
.subckt sky130_fd_sc_hd__o31ai_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41oi_1 abstract view
.subckt sky130_fd_sc_hd__a41oi_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_4 abstract view
.subckt sky130_fd_sc_hd__clkinv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_2 abstract view
.subckt sky130_fd_sc_hd__nand2b_2 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_2 abstract view
.subckt sky130_fd_sc_hd__clkinv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtn_1 abstract view
.subckt sky130_fd_sc_hd__dfrtn_1 CLK_N D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_4 abstract view
.subckt sky130_fd_sc_hd__inv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111ai_1 abstract view
.subckt sky130_fd_sc_hd__o2111ai_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_2 abstract view
.subckt sky130_fd_sc_hd__nor3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_1 abstract view
.subckt sky130_fd_sc_hd__o21bai_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_4 abstract view
.subckt sky130_fd_sc_hd__dfrtp_4 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_1 abstract view
.subckt sky130_fd_sc_hd__nand3b_1 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_1 abstract view
.subckt sky130_fd_sc_hd__o31ai_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_4 abstract view
.subckt sky130_fd_sc_hd__o211ai_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_2 abstract view
.subckt sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_2 abstract view
.subckt sky130_fd_sc_hd__o21a_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_1 abstract view
.subckt sky130_fd_sc_hd__nor4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

.subckt caravel_clocking VGND VPWR core_clk ext_clk ext_clk_sel ext_reset pll_clk
+ pll_clk90 resetb resetb_sync sel2[0] sel2[1] sel2[2] sel[0] sel[1] sel[2] user_clk
XFILLER_22_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_432_ _204_/A1 _432_/D _372_/S VGND VGND VPWR VPWR _432_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_13_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_294_ _429_/Q _430_/Q VGND VGND VPWR VPWR _294_/Y sky130_fd_sc_hd__nor2_1
X_363_ _365_/A _429_/Q VGND VGND VPWR VPWR _363_/Y sky130_fd_sc_hd__nand2_1
XFILLER_8_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_415_ _204_/A1 _440_/Q _372_/S VGND VGND VPWR VPWR _415_/Q sky130_fd_sc_hd__dfrtp_1
X_346_ _416_/D _292_/Y _419_/Q VGND VGND VPWR VPWR _347_/B sky130_fd_sc_hd__o21ai_1
XFILLER_12_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_277_ _422_/Q _423_/Q _421_/Q VGND VGND VPWR VPWR _277_/Y sky130_fd_sc_hd__nor3b_2
XFILLER_5_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_79 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_329_ _329_/A _329_/B VGND VGND VPWR VPWR _329_/Y sky130_fd_sc_hd__nor2_1
XFILLER_18_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_1_1__f__037_ clkbuf_0__037_/X VGND VGND VPWR VPWR _208_/A0 sky130_fd_sc_hd__clkbuf_16
XFILLER_16_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_431_ _204_/A1 _431_/D _372_/S VGND VGND VPWR VPWR _431_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_13_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_293_ _223_/S _365_/A VGND VGND VPWR VPWR _293_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_9_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_362_ _295_/C _293_/Y _361_/Y VGND VGND VPWR VPWR _428_/D sky130_fd_sc_hd__o21ai_1
XANTENNA__265__A1 _327_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_104 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_345_ _311_/C _419_/Q _345_/C _431_/Q VGND VGND VPWR VPWR _347_/A sky130_fd_sc_hd__nand4bb_1
X_414_ _207_/A1 _414_/D fanout27/X VGND VGND VPWR VPWR _414_/Q sky130_fd_sc_hd__dfstp_1
X_276_ _426_/Q _210_/X _360_/S VGND VGND VPWR VPWR _426_/D sky130_fd_sc_hd__mux2_1
XFILLER_9_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_328_ _442_/D _441_/D _327_/A VGND VGND VPWR VPWR _329_/B sky130_fd_sc_hd__o21a_1
XFILLER_0_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__395__B1 _311_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_292_ _431_/Q _345_/C VGND VGND VPWR VPWR _292_/Y sky130_fd_sc_hd__nand2_1
XFILLER_13_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_430_ _456_/CLK _430_/D fanout26/X VGND VGND VPWR VPWR _430_/Q sky130_fd_sc_hd__dfrtp_2
X_361_ _223_/S _280_/X _219_/X VGND VGND VPWR VPWR _361_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_8_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_413_ _204_/A1 _413_/D _372_/S VGND VGND VPWR VPWR _413_/Q sky130_fd_sc_hd__dfrtp_1
X_344_ _414_/Q _342_/Y _343_/Y VGND VGND VPWR VPWR _414_/D sky130_fd_sc_hd__o21ai_1
X_275_ _232_/X _273_/Y _274_/Y _234_/S VGND VGND VPWR VPWR _447_/D sky130_fd_sc_hd__o2bb2ai_1
XFILLER_5_131 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_258_ _258_/A VGND VGND VPWR VPWR _258_/Y sky130_fd_sc_hd__inv_2
XFILLER_9_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_327_ _327_/A _442_/D _441_/D VGND VGND VPWR VPWR _329_/A sky130_fd_sc_hd__nor3_1
XFILLER_18_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__452__RESET_B fanout28/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_14 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput11 _341_/Y VGND VGND VPWR VPWR resetb_sync sky130_fd_sc_hd__buf_12
XFILLER_16_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_291_ _432_/Q _433_/Q VGND VGND VPWR VPWR _345_/C sky130_fd_sc_hd__nor2_1
XFILLER_26_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_360_ _427_/Q _211_/X _360_/S VGND VGND VPWR VPWR _427_/D sky130_fd_sc_hd__mux2_1
XFILLER_12_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_412_ _456_/CLK _412_/D fanout26/X VGND VGND VPWR VPWR _413_/D sky130_fd_sc_hd__dfrtp_1
X_343_ _342_/Y _414_/Q _234_/S VGND VGND VPWR VPWR _343_/Y sky130_fd_sc_hd__a21oi_1
X_274_ _385_/B _447_/Q VGND VGND VPWR VPWR _274_/Y sky130_fd_sc_hd__nand2_1
XFILLER_5_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_326_ _451_/Q _450_/Q VGND VGND VPWR VPWR _326_/Y sky130_fd_sc_hd__xnor2_1
X_257_ _257_/A VGND VGND VPWR VPWR _257_/Y sky130_fd_sc_hd__inv_2
XFILLER_18_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__395__A2 _311_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_309_ _311_/B _311_/C VGND VGND VPWR VPWR _309_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_29_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_0_divider.out _304_/Y VGND VGND VPWR VPWR clkbuf_0_divider.out/X sky130_fd_sc_hd__clkbuf_16
XFILLER_20_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_26 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_131 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_79 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input8_A sel[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_91 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_290_ _215_/X _288_/Y _289_/Y _219_/S VGND VGND VPWR VPWR _422_/D sky130_fd_sc_hd__o2bb2ai_1
Xclkbuf_0_pll_clk pll_clk VGND VGND VPWR VPWR clkbuf_0_pll_clk/X sky130_fd_sc_hd__clkbuf_16
XFILLER_12_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_411_ _411_/CLK _411_/D _372_/S VGND VGND VPWR VPWR _411_/Q sky130_fd_sc_hd__dfstp_1
X_273_ _234_/S _385_/B VGND VGND VPWR VPWR _273_/Y sky130_fd_sc_hd__nand2b_1
X_342_ _327_/A _442_/D _441_/D _453_/Q _299_/Y VGND VGND VPWR VPWR _342_/Y sky130_fd_sc_hd__o2111ai_2
XANTENNA__446__RESET_B fanout28/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_325_ _442_/D _441_/D VGND VGND VPWR VPWR _325_/Y sky130_fd_sc_hd__xnor2_1
X_308_ _307_/Y _298_/B _306_/X _305_/Y VGND VGND VPWR VPWR _308_/Y sky130_fd_sc_hd__o31ai_2
XFILLER_1_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_239_ _339_/Y _327_/A _300_/Y VGND VGND VPWR VPWR _239_/X sky130_fd_sc_hd__mux2_1
XFILLER_28_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__451__SET_B fanout28/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_1_0__f_pll_clk90 clkbuf_0_pll_clk90/X VGND VGND VPWR VPWR _455_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_12_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_341_ _341_/A _409_/Q VGND VGND VPWR VPWR _341_/Y sky130_fd_sc_hd__nor2_1
X_410_ _410_/CLK _411_/Q _372_/S VGND VGND VPWR VPWR _410_/Q sky130_fd_sc_hd__dfstp_1
X_272_ _263_/Y _265_/X _234_/S VGND VGND VPWR VPWR _272_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_4_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_324_ _432_/Q _431_/Q VGND VGND VPWR VPWR _324_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_9_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_255_ _255_/A VGND VGND VPWR VPWR _255_/Y sky130_fd_sc_hd__inv_2
XFILLER_1_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_307_ _449_/Q _414_/Q VGND VGND VPWR VPWR _307_/Y sky130_fd_sc_hd__nor2_1
X_238_ _237_/X _442_/D _240_/S VGND VGND VPWR VPWR _238_/X sky130_fd_sc_hd__mux2_1
XFILLER_29_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_92 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_340_ _458_/Q _457_/Q VGND VGND VPWR VPWR _340_/Y sky130_fd_sc_hd__xnor2_1
X_271_ _271_/A _271_/B VGND VGND VPWR VPWR _449_/D sky130_fd_sc_hd__nand2_1
XFILLER_5_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__455__RESET_B fanout28/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_323_ _321_/Y _323_/B VGND VGND VPWR VPWR _323_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_2_105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__240__A1 _327_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_306_ _449_/Q _414_/Q VGND VGND VPWR VPWR _306_/X sky130_fd_sc_hd__and2_1
X_237_ _336_/Y _442_/D _300_/Y VGND VGND VPWR VPWR _237_/X sky130_fd_sc_hd__mux2_1
XFILLER_20_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__213__A1 _311_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_118 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input6_A sel2[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_270_ _262_/Y _263_/Y _265_/X _243_/Y _234_/S VGND VGND VPWR VPWR _271_/B sky130_fd_sc_hd__a41oi_1
X_399_ _242_/X _458_/Q _400_/A VGND VGND VPWR VPWR _458_/D sky130_fd_sc_hd__mux2_1
XFILLER_4_40 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_322_ _428_/Q _429_/Q _430_/Q VGND VGND VPWR VPWR _323_/B sky130_fd_sc_hd__o21ai_1
XFILLER_2_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_1_0__f_net10 clkbuf_0_net10/X VGND VGND VPWR VPWR core_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_1_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_253_ _253_/A VGND VGND VPWR VPWR _412_/D sky130_fd_sc_hd__clkinv_4
XFILLER_24_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_305_ _441_/D _305_/B VGND VGND VPWR VPWR _305_/Y sky130_fd_sc_hd__nand2b_2
X_236_ _235_/X _441_/D _240_/S VGND VGND VPWR VPWR _236_/X sky130_fd_sc_hd__mux2_1
XFILLER_1_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_fanout27_A fanout28/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_219_ _218_/X _311_/C _219_/S VGND VGND VPWR VPWR _219_/X sky130_fd_sc_hd__mux2_1
XFILLER_31_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_0_pll_clk_A pll_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_398_ _241_/X _457_/Q _400_/A VGND VGND VPWR VPWR _457_/D sky130_fd_sc_hd__mux2_1
XFILLER_4_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_252_ _453_/Q VGND VGND VPWR VPWR _300_/C sky130_fd_sc_hd__clkinv_4
XFILLER_1_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_321_ _428_/Q _429_/Q _430_/Q VGND VGND VPWR VPWR _321_/Y sky130_fd_sc_hd__nor3_1
XFILLER_24_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_304_ _303_/Y _365_/A _302_/X _301_/Y VGND VGND VPWR VPWR _304_/Y sky130_fd_sc_hd__o31ai_2
X_235_ _300_/C _441_/D _300_/Y VGND VGND VPWR VPWR _235_/X sky130_fd_sc_hd__mux2_1
XFILLER_1_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_218_ _295_/C _311_/C _295_/Y VGND VGND VPWR VPWR _218_/X sky130_fd_sc_hd__mux2_1
XFILLER_24_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xuser_clk_out_buffer _208_/X VGND VGND VPWR VPWR user_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_21_186 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_397_ _456_/Q _395_/Y _396_/Y VGND VGND VPWR VPWR _456_/D sky130_fd_sc_hd__o21ai_1
XFILLER_4_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_251_ _446_/Q VGND VGND VPWR VPWR _251_/Y sky130_fd_sc_hd__clkinv_2
X_320_ _428_/Q _429_/Q VGND VGND VPWR VPWR _320_/Y sky130_fd_sc_hd__xnor2_1
X_449_ _449_/CLK _449_/D fanout27/X VGND VGND VPWR VPWR _449_/Q sky130_fd_sc_hd__dfstp_1
XANTENNA__234__A1 _327_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_1_1__f_divider.out clkbuf_0_divider.out/X VGND VGND VPWR VPWR _206_/A1 sky130_fd_sc_hd__clkbuf_16
X_303_ _424_/Q _456_/Q VGND VGND VPWR VPWR _303_/Y sky130_fd_sc_hd__nor2_1
X_234_ _233_/X _327_/A _234_/S VGND VGND VPWR VPWR _260_/A sky130_fd_sc_hd__mux2_1
XFILLER_1_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_217_ _216_/X _351_/A _223_/S VGND VGND VPWR VPWR _257_/A sky130_fd_sc_hd__mux2_1
XFILLER_25_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__328__B1 _327_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_465_ _208_/A1 _465_/D fanout27/X VGND VGND VPWR VPWR _465_/Q sky130_fd_sc_hd__dfrtp_1
X_396_ _395_/Y _456_/Q _223_/S VGND VGND VPWR VPWR _396_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_5_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout20 _437_/Q VGND VGND VPWR VPWR _416_/D sky130_fd_sc_hd__clkbuf_2
XANTENNA_input4_A sel2[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_63 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_250_ _450_/Q VGND VGND VPWR VPWR _250_/Y sky130_fd_sc_hd__inv_2
X_379_ _465_/Q _443_/Q VGND VGND VPWR VPWR _379_/Y sky130_fd_sc_hd__nor2_1
X_448_ _455_/CLK _448_/D fanout28/X VGND VGND VPWR VPWR _448_/Q sky130_fd_sc_hd__dfrtn_1
XFILLER_24_40 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_302_ _424_/Q _456_/Q VGND VGND VPWR VPWR _302_/X sky130_fd_sc_hd__and2_1
X_233_ _335_/Y _327_/A _262_/Y VGND VGND VPWR VPWR _233_/X sky130_fd_sc_hd__mux2_1
XFILLER_1_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_216_ _319_/Y _351_/A _277_/Y VGND VGND VPWR VPWR _216_/X sky130_fd_sc_hd__mux2_1
XFILLER_24_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__282__B1 _311_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_259__1 _455_/CLK VGND VGND VPWR VPWR _447_/CLK sky130_fd_sc_hd__inv_4
XFILLER_7_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_464_ _464_/CLK _464_/D fanout27/X VGND VGND VPWR VPWR _464_/Q sky130_fd_sc_hd__dfstp_1
X_395_ _351_/A _311_/B _311_/C _428_/Q _294_/Y VGND VGND VPWR VPWR _395_/Y sky130_fd_sc_hd__o2111ai_1
XFILLER_4_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout21 _234_/S VGND VGND VPWR VPWR _240_/S sky130_fd_sc_hd__clkbuf_4
X_447_ _447_/CLK _447_/D fanout28/X VGND VGND VPWR VPWR _447_/Q sky130_fd_sc_hd__dfstp_1
X_378_ _378_/A _378_/B _441_/Q VGND VGND VPWR VPWR _378_/Y sky130_fd_sc_hd__nand3_1
XFILLER_1_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_301_ _416_/D _301_/B VGND VGND VPWR VPWR _301_/Y sky130_fd_sc_hd__nand2b_2
XFILLER_24_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_232_ _231_/X _442_/D _234_/S VGND VGND VPWR VPWR _232_/X sky130_fd_sc_hd__mux2_1
Xclkbuf_1_0__f__037_ clkbuf_0__037_/X VGND VGND VPWR VPWR _206_/A0 sky130_fd_sc_hd__clkbuf_16
XFILLER_28_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_215_ _214_/X _311_/B _219_/S VGND VGND VPWR VPWR _215_/X sky130_fd_sc_hd__mux2_1
XFILLER_16_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_463_ _464_/CLK _463_/D fanout27/X VGND VGND VPWR VPWR _463_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_4_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_394_ _240_/S _455_/Q _265_/X _393_/Y VGND VGND VPWR VPWR _455_/D sky130_fd_sc_hd__o31a_1
XTAP_295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout22 _445_/Q VGND VGND VPWR VPWR _234_/S sky130_fd_sc_hd__clkbuf_4
Xclkbuf_1_1__f_pll_clk90 clkbuf_0_pll_clk90/X VGND VGND VPWR VPWR _207_/A1 sky130_fd_sc_hd__clkbuf_16
X_377_ _442_/Q _464_/Q VGND VGND VPWR VPWR _378_/B sky130_fd_sc_hd__nand2b_1
X_446_ _455_/CLK _446_/D fanout28/X VGND VGND VPWR VPWR _446_/Q sky130_fd_sc_hd__dfrtn_1
XFILLER_8_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__219__A1 _311_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_406__6 _204_/A1 VGND VGND VPWR VPWR _426_/CLK sky130_fd_sc_hd__inv_4
Xclkbuf_0_ext_clk ext_clk VGND VGND VPWR VPWR clkbuf_0_ext_clk/X sky130_fd_sc_hd__clkbuf_16
XFILLER_24_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_231_ _332_/Y _442_/D _262_/Y VGND VGND VPWR VPWR _231_/X sky130_fd_sc_hd__mux2_1
X_300_ _454_/Q _455_/Q _300_/C VGND VGND VPWR VPWR _300_/Y sky130_fd_sc_hd__nor3_2
X_429_ _456_/CLK _429_/D fanout26/X VGND VGND VPWR VPWR _429_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_1_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_90 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput1 ext_clk_sel VGND VGND VPWR VPWR _253_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_18_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_214_ _316_/Y _311_/B _277_/Y VGND VGND VPWR VPWR _214_/X sky130_fd_sc_hd__mux2_1
XFILLER_24_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__282__A2 _311_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_183 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_462_ _208_/A1 _462_/D fanout27/X VGND VGND VPWR VPWR _465_/D sky130_fd_sc_hd__dfrtp_1
XFILLER_27_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_393_ _240_/S _265_/X _240_/X VGND VGND VPWR VPWR _393_/Y sky130_fd_sc_hd__o21bai_1
XTAP_296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout23 _223_/S VGND VGND VPWR VPWR _219_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_1_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_445_ _207_/A1 _445_/D fanout28/X VGND VGND VPWR VPWR _445_/Q sky130_fd_sc_hd__dfrtp_1
X_376_ _464_/Q _442_/Q VGND VGND VPWR VPWR _378_/A sky130_fd_sc_hd__nand2b_1
X_256__4 _456_/CLK VGND VGND VPWR VPWR _422_/CLK sky130_fd_sc_hd__inv_4
XANTENNA_input2_A ext_reset VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_230_ _229_/X _441_/D _234_/S VGND VGND VPWR VPWR _258_/A sky130_fd_sc_hd__mux2_1
X_359_ _425_/Q _209_/X _360_/S VGND VGND VPWR VPWR _425_/D sky130_fd_sc_hd__mux2_1
X_428_ _456_/CLK _428_/D fanout26/X VGND VGND VPWR VPWR _428_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_1_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput2 ext_reset VGND VGND VPWR VPWR _341_/A sky130_fd_sc_hd__clkbuf_1
XTAP_80 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_91 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_213_ _212_/X _311_/C _219_/S VGND VGND VPWR VPWR _255_/A sky130_fd_sc_hd__mux2_1
X_403__8 _403__8/A VGND VGND VPWR VPWR _410_/CLK sky130_fd_sc_hd__inv_4
XFILLER_18_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_79 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_0_net10 _206_/X VGND VGND VPWR VPWR clkbuf_0_net10/X sky130_fd_sc_hd__clkbuf_16
XFILLER_21_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_66 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_461_ _464_/CLK _461_/D fanout27/X VGND VGND VPWR VPWR _464_/D sky130_fd_sc_hd__dfstp_1
X_392_ _240_/S _454_/Q _265_/X _391_/Y VGND VGND VPWR VPWR _454_/D sky130_fd_sc_hd__o31a_1
XFILLER_4_14 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout13 _465_/Q VGND VGND VPWR VPWR _327_/A sky130_fd_sc_hd__buf_4
Xfanout24 _420_/Q VGND VGND VPWR VPWR _223_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_1_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_444_ _207_/A1 _444_/D fanout27/X VGND VGND VPWR VPWR _444_/Q sky130_fd_sc_hd__dfstp_1
X_375_ _375_/A _375_/B VGND VGND VPWR VPWR _444_/D sky130_fd_sc_hd__nand2_1
XFILLER_24_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_427_ _456_/CLK _427_/D fanout26/X VGND VGND VPWR VPWR _427_/Q sky130_fd_sc_hd__dfrtn_1
XFILLER_1_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_358_ _257_/Y _287_/Y _357_/Y VGND VGND VPWR VPWR _423_/D sky130_fd_sc_hd__o21ai_1
Xinput3 resetb VGND VGND VPWR VPWR input3/X sky130_fd_sc_hd__clkbuf_1
XTAP_70 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_81 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_92 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__327__A _327_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_289_ _357_/B _422_/Q VGND VGND VPWR VPWR _289_/Y sky130_fd_sc_hd__nand2_1
XFILLER_27_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_212_ _247_/Y _311_/C _277_/Y VGND VGND VPWR VPWR _212_/X sky130_fd_sc_hd__mux2_1
XFILLER_32_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__267__A1 _327_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_411__30 VGND VGND VPWR VPWR _411__30/HI _411_/D sky130_fd_sc_hd__conb_1
XANTENNA__445__RESET_B fanout28/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_460_ _464_/CLK _460_/D fanout27/X VGND VGND VPWR VPWR _463_/D sky130_fd_sc_hd__dfrtp_1
XFILLER_27_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_391_ _240_/S _265_/X _238_/X VGND VGND VPWR VPWR _391_/Y sky130_fd_sc_hd__o21bai_1
XFILLER_4_26 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_144 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout25 fanout29/X VGND VGND VPWR VPWR _372_/S sky130_fd_sc_hd__buf_4
XTAP_298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout14 _464_/Q VGND VGND VPWR VPWR _442_/D sky130_fd_sc_hd__buf_4
XTAP_276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_374_ _400_/A _297_/Y _444_/Q VGND VGND VPWR VPWR _375_/B sky130_fd_sc_hd__o21ai_1
X_443_ _207_/A1 _465_/Q VGND VGND VPWR VPWR _443_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput4 sel2[0] VGND VGND VPWR VPWR _460_/D sky130_fd_sc_hd__clkbuf_1
X_426_ _426_/CLK _426_/D fanout26/X VGND VGND VPWR VPWR _426_/Q sky130_fd_sc_hd__dfstp_1
XTAP_71 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_82 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_93 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_288_ _219_/S _357_/B VGND VGND VPWR VPWR _288_/Y sky130_fd_sc_hd__nand2b_1
X_357_ _219_/S _357_/B _423_/Q VGND VGND VPWR VPWR _357_/Y sky130_fd_sc_hd__nand3b_1
XFILLER_27_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_211_ _315_/X _313_/B _223_/S VGND VGND VPWR VPWR _211_/X sky130_fd_sc_hd__mux2_1
XFILLER_10_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_409_ _409_/CLK _410_/Q fanout27/X VGND VGND VPWR VPWR _409_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_24_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_390_ _300_/C _298_/Y _389_/Y VGND VGND VPWR VPWR _453_/D sky130_fd_sc_hd__o21ai_1
XFILLER_4_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout15 _463_/Q VGND VGND VPWR VPWR _441_/D sky130_fd_sc_hd__buf_4
XTAP_255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_1__f_pll_clk clkbuf_0_pll_clk/X VGND VGND VPWR VPWR _204_/A1 sky130_fd_sc_hd__clkbuf_16
XTAP_200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout26 fanout29/X VGND VGND VPWR VPWR fanout26/X sky130_fd_sc_hd__buf_4
X_373_ _400_/A _444_/Q _373_/C _457_/Q VGND VGND VPWR VPWR _375_/A sky130_fd_sc_hd__nand4bb_1
XANTENNA__312__A1 _311_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_442_ _455_/CLK _442_/D VGND VGND VPWR VPWR _442_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_170 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_92 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__345__A_N _311_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__447__SET_B fanout28/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput5 sel2[1] VGND VGND VPWR VPWR _461_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_14_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_425_ _456_/CLK _425_/D fanout26/X VGND VGND VPWR VPWR _425_/Q sky130_fd_sc_hd__dfrtn_1
X_287_ _278_/Y _280_/X _219_/S VGND VGND VPWR VPWR _287_/Y sky130_fd_sc_hd__a21oi_1
X_356_ _255_/Y _287_/Y _355_/Y VGND VGND VPWR VPWR _421_/D sky130_fd_sc_hd__o21ai_1
XFILLER_27_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_35 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_72 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_83 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_94 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_210_ _310_/Y _313_/Y _223_/S VGND VGND VPWR VPWR _210_/X sky130_fd_sc_hd__mux2_1
Xclkbuf_1_0__f_divider2.out clkbuf_0_divider2.out/X VGND VGND VPWR VPWR _464_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_339_ _337_/Y _339_/B VGND VGND VPWR VPWR _339_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_2_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__264__A _327_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_92 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout16 _463_/Q VGND VGND VPWR VPWR _400_/A sky130_fd_sc_hd__clkbuf_2
XTAP_289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout27 fanout28/X VGND VGND VPWR VPWR fanout27/X sky130_fd_sc_hd__buf_4
XTAP_256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_372_ _440_/Q _372_/A1 _372_/S VGND VGND VPWR VPWR _440_/D sky130_fd_sc_hd__mux2_1
X_441_ _455_/CLK _441_/D VGND VGND VPWR VPWR _441_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_13_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__312__A2 _311_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_424_ _424_/CLK _424_/D fanout26/X VGND VGND VPWR VPWR _424_/Q sky130_fd_sc_hd__dfstp_1
X_286_ _286_/A _286_/B VGND VGND VPWR VPWR _424_/D sky130_fd_sc_hd__nand2_1
X_355_ _219_/S _357_/B _421_/Q VGND VGND VPWR VPWR _355_/Y sky130_fd_sc_hd__nand3b_1
Xinput6 sel2[2] VGND VGND VPWR VPWR _462_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_10_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_73 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_84 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_95 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__221__A1 _311_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__212__A1 _311_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_269_ _262_/Y _263_/Y _265_/X _243_/Y VGND VGND VPWR VPWR _271_/A sky130_fd_sc_hd__a31o_1
X_338_ _454_/Q _453_/Q _455_/Q VGND VGND VPWR VPWR _339_/B sky130_fd_sc_hd__o21ai_1
XFILLER_32_170 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_0__037_ _205_/X VGND VGND VPWR VPWR clkbuf_0__037_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_4_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout28 fanout29/X VGND VGND VPWR VPWR fanout28/X sky130_fd_sc_hd__buf_4
X_371_ _369_/Y _371_/B VGND VGND VPWR VPWR _433_/D sky130_fd_sc_hd__nand2b_1
X_440_ _204_/A1 _440_/D VGND VGND VPWR VPWR _440_/Q sky130_fd_sc_hd__dfxtp_1
Xfanout17 _439_/Q VGND VGND VPWR VPWR _351_/A sky130_fd_sc_hd__buf_4
XFILLER_13_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_354_ _223_/S _280_/X _352_/Y _353_/Y VGND VGND VPWR VPWR _420_/D sky130_fd_sc_hd__o22a_1
XFILLER_14_92 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_285_ _277_/Y _278_/Y _280_/X _244_/Y _223_/S VGND VGND VPWR VPWR _286_/B sky130_fd_sc_hd__a41oi_1
X_423_ _456_/CLK _423_/D fanout26/X VGND VGND VPWR VPWR _423_/Q sky130_fd_sc_hd__dfrtn_1
XANTENNA__448__RESET_B fanout28/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_85 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_74 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_96 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput7 sel[0] VGND VGND VPWR VPWR _434_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_27_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_268_ _385_/B VGND VGND VPWR VPWR _268_/Y sky130_fd_sc_hd__inv_2
X_337_ _454_/Q _453_/Q _455_/Q VGND VGND VPWR VPWR _337_/Y sky130_fd_sc_hd__nor3_1
XFILLER_2_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_0_pll_clk90_A pll_clk90 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_138 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_1_0__f_divider.out clkbuf_0_divider.out/X VGND VGND VPWR VPWR _439_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_11_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__342__A1 _327_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout29 input3/X VGND VGND VPWR VPWR fanout29/X sky130_fd_sc_hd__buf_2
Xfanout18 _438_/Q VGND VGND VPWR VPWR _311_/B sky130_fd_sc_hd__buf_4
X_370_ _416_/D _432_/Q _431_/Q _433_/Q VGND VGND VPWR VPWR _371_/B sky130_fd_sc_hd__o31ai_1
XANTENNA__242__A0 _327_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_353_ _353_/A _353_/B _416_/Q VGND VGND VPWR VPWR _353_/Y sky130_fd_sc_hd__nand3_1
X_284_ _277_/Y _278_/Y _280_/X _244_/Y VGND VGND VPWR VPWR _286_/A sky130_fd_sc_hd__a31o_1
X_422_ _422_/CLK _422_/D fanout26/X VGND VGND VPWR VPWR _422_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_30_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_1_0__f_pll_clk clkbuf_0_pll_clk/X VGND VGND VPWR VPWR _456_/CLK sky130_fd_sc_hd__clkbuf_16
Xinput8 sel[1] VGND VGND VPWR VPWR _435_/D sky130_fd_sc_hd__clkbuf_1
XTAP_86 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_75 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_97 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_267_ _327_/A _442_/D _441_/D _263_/Y VGND VGND VPWR VPWR _385_/B sky130_fd_sc_hd__o211ai_4
X_336_ _454_/Q _453_/Q VGND VGND VPWR VPWR _336_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_32_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_183 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_319_ _317_/Y _319_/B VGND VGND VPWR VPWR _319_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_32_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout19 _437_/Q VGND VGND VPWR VPWR _311_/C sky130_fd_sc_hd__buf_4
XTAP_259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_input9_A sel[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__233__A1 _327_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__215__A1 _311_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_421_ _456_/CLK _421_/D fanout26/X VGND VGND VPWR VPWR _421_/Q sky130_fd_sc_hd__dfrtn_1
X_352_ _350_/Y _351_/X _280_/X VGND VGND VPWR VPWR _352_/Y sky130_fd_sc_hd__o21ai_1
Xinput9 sel[2] VGND VGND VPWR VPWR _436_/D sky130_fd_sc_hd__clkbuf_1
X_283_ _357_/B VGND VGND VPWR VPWR _283_/Y sky130_fd_sc_hd__inv_2
XTAP_87 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_76 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_98 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_407__2 _207_/A1 VGND VGND VPWR VPWR _449_/CLK sky130_fd_sc_hd__inv_4
XPHY_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_266_ _327_/A _464_/Q _400_/A VGND VGND VPWR VPWR _298_/B sky130_fd_sc_hd__o21ai_2
XFILLER_18_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_335_ _333_/Y _335_/B VGND VGND VPWR VPWR _335_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_24_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_249_ _457_/Q VGND VGND VPWR VPWR _249_/Y sky130_fd_sc_hd__clkinv_2
X_318_ _422_/Q _421_/Q _423_/Q VGND VGND VPWR VPWR _319_/B sky130_fd_sc_hd__o21ai_1
XFILLER_22_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_0_divider2.out _308_/Y VGND VGND VPWR VPWR clkbuf_0_divider2.out/X sky130_fd_sc_hd__clkbuf_16
XFILLER_0_131 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_351_ _351_/A _418_/Q VGND VGND VPWR VPWR _351_/X sky130_fd_sc_hd__and2_1
X_420_ _204_/A1 _420_/D _372_/S VGND VGND VPWR VPWR _420_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_14_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_282_ _351_/A _311_/B _311_/C _278_/Y VGND VGND VPWR VPWR _357_/B sky130_fd_sc_hd__o211ai_4
XFILLER_27_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_77 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_66 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_88 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_99 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_334_ _447_/Q _446_/Q _448_/Q VGND VGND VPWR VPWR _335_/B sky130_fd_sc_hd__o21ai_1
XFILLER_32_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_265_ _327_/A _442_/D _441_/D VGND VGND VPWR VPWR _265_/X sky130_fd_sc_hd__o21a_2
XFILLER_23_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_248_ _428_/Q VGND VGND VPWR VPWR _295_/C sky130_fd_sc_hd__clkinv_4
X_317_ _422_/Q _421_/Q _423_/Q VGND VGND VPWR VPWR _317_/Y sky130_fd_sc_hd__nor3_1
XFILLER_2_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__281__B1 _311_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_281_ _351_/A _311_/B _311_/C VGND VGND VPWR VPWR _365_/A sky130_fd_sc_hd__o21ai_2
X_350_ _351_/A _418_/Q VGND VGND VPWR VPWR _350_/Y sky130_fd_sc_hd__nor2_1
XFILLER_14_74 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_78 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_67 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_89 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_402_ _400_/Y _402_/B VGND VGND VPWR VPWR _459_/D sky130_fd_sc_hd__nand2b_1
X_264_ _327_/A _464_/Q VGND VGND VPWR VPWR _264_/Y sky130_fd_sc_hd__nor2_1
XPHY_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_333_ _447_/Q _446_/Q _448_/Q VGND VGND VPWR VPWR _333_/Y sky130_fd_sc_hd__nor3_1
XFILLER_2_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_316_ _422_/Q _421_/Q VGND VGND VPWR VPWR _316_/Y sky130_fd_sc_hd__xnor2_1
X_247_ _421_/Q VGND VGND VPWR VPWR _247_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_28_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_167 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_144 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__218__A1 _311_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_280_ _351_/A _311_/B _311_/C VGND VGND VPWR VPWR _280_/X sky130_fd_sc_hd__o21a_1
XFILLER_14_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input7_A sel[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_1_1__f_divider2.out clkbuf_0_divider2.out/X VGND VGND VPWR VPWR _208_/A1 sky130_fd_sc_hd__clkbuf_16
XTAP_79 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_68 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_401_ _400_/A _458_/Q _457_/Q _459_/Q VGND VGND VPWR VPWR _402_/B sky130_fd_sc_hd__o31ai_1
XPHY_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_332_ _447_/Q _446_/Q VGND VGND VPWR VPWR _332_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_18_118 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_263_ _451_/Q _452_/Q VGND VGND VPWR VPWR _263_/Y sky130_fd_sc_hd__nor2_2
XFILLER_23_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__281__A2 _311_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_315_ _246_/Y _278_/Y _314_/X VGND VGND VPWR VPWR _315_/X sky130_fd_sc_hd__a21o_1
X_246_ _425_/Q VGND VGND VPWR VPWR _246_/Y sky130_fd_sc_hd__inv_2
XFILLER_22_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__454__SET_B fanout28/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_229_ _251_/Y _441_/D _262_/Y VGND VGND VPWR VPWR _229_/X sky130_fd_sc_hd__mux2_1
XANTENNA__450__RESET_B fanout28/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_69 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_1_1__f_ext_clk clkbuf_0_ext_clk/X VGND VGND VPWR VPWR _205_/A0 sky130_fd_sc_hd__clkbuf_16
XPHY_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_400_ _400_/A _458_/Q _457_/Q _459_/Q VGND VGND VPWR VPWR _400_/Y sky130_fd_sc_hd__nor4_1
XFILLER_25_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_262_ _447_/Q _448_/Q _446_/Q VGND VGND VPWR VPWR _262_/Y sky130_fd_sc_hd__nor3b_2
XPHY_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_331_ _250_/Y _263_/Y _330_/X VGND VGND VPWR VPWR _331_/X sky130_fd_sc_hd__a21o_1
XFILLER_32_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_144 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_245_ _431_/Q VGND VGND VPWR VPWR _245_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_14_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_314_ _426_/Q _425_/Q _427_/Q VGND VGND VPWR VPWR _314_/X sky130_fd_sc_hd__o21a_1
XFILLER_11_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__309__A _311_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_228_ _331_/X _329_/B _240_/S VGND VGND VPWR VPWR _228_/X sky130_fd_sc_hd__mux2_1
XFILLER_6_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__311__B _311_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_330_ _451_/Q _450_/Q _452_/Q VGND VGND VPWR VPWR _330_/X sky130_fd_sc_hd__o21a_1
XPHY_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_261_ _451_/Q _227_/X _388_/S VGND VGND VPWR VPWR _451_/D sky130_fd_sc_hd__mux2_1
X_459_ _207_/A1 _459_/D fanout28/X VGND VGND VPWR VPWR _459_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_17_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__266__A1 _327_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_313_ _313_/A _313_/B VGND VGND VPWR VPWR _313_/Y sky130_fd_sc_hd__nor2_1
XFILLER_14_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_244_ _424_/Q VGND VGND VPWR VPWR _244_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_20_126 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__309__B _311_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_227_ _326_/Y _329_/Y _240_/S VGND VGND VPWR VPWR _227_/X sky130_fd_sc_hd__mux2_1
XANTENNA__239__A1 _327_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__311__C _311_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input5_A sel2[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_260_ _260_/A VGND VGND VPWR VPWR _260_/Y sky130_fd_sc_hd__inv_2
XPHY_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_458_ _207_/A1 _458_/D fanout27/X VGND VGND VPWR VPWR _458_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_17_143 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_389_ _234_/S _265_/X _236_/X VGND VGND VPWR VPWR _389_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_23_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_243_ _449_/Q VGND VGND VPWR VPWR _243_/Y sky130_fd_sc_hd__clkinv_4
XTAP_190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_312_ _311_/B _311_/C _351_/A VGND VGND VPWR VPWR _313_/B sky130_fd_sc_hd__o21a_1
XFILLER_11_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_404__9 core_clk VGND VGND VPWR VPWR _411_/CLK sky130_fd_sc_hd__inv_4
XFILLER_20_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_226_ _250_/Y _325_/Y _240_/S VGND VGND VPWR VPWR _226_/X sky130_fd_sc_hd__mux2_1
XFILLER_3_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_209_ _246_/Y _309_/Y _219_/S VGND VGND VPWR VPWR _209_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__453__RESET_B fanout28/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_457_ _207_/A1 _457_/D fanout27/X VGND VGND VPWR VPWR _457_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_23_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_388_ _452_/Q _228_/X _388_/S VGND VGND VPWR VPWR _452_/D sky130_fd_sc_hd__mux2_1
X_242_ _327_/A _340_/Y _297_/Y VGND VGND VPWR VPWR _242_/X sky130_fd_sc_hd__mux2_1
X_311_ _351_/A _311_/B _311_/C VGND VGND VPWR VPWR _313_/A sky130_fd_sc_hd__nor3_1
XTAP_191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_254__7 _403__8/A VGND VGND VPWR VPWR _409_/CLK sky130_fd_sc_hd__inv_4
XFILLER_9_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_1_0__f_ext_clk clkbuf_0_ext_clk/X VGND VGND VPWR VPWR _372_/A1 sky130_fd_sc_hd__clkbuf_16
XFILLER_22_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_225_ _439_/Q _324_/Y _292_/Y VGND VGND VPWR VPWR _225_/X sky130_fd_sc_hd__mux2_1
XFILLER_12_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_208_ _208_/A0 _208_/A1 _413_/Q VGND VGND VPWR VPWR _208_/X sky130_fd_sc_hd__mux2_1
XFILLER_31_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_14 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__220__A1 _311_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_17 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_456_ _456_/CLK _456_/D fanout26/X VGND VGND VPWR VPWR _456_/Q sky130_fd_sc_hd__dfstp_1
X_387_ _450_/Q _226_/X _388_/S VGND VGND VPWR VPWR _450_/D sky130_fd_sc_hd__mux2_1
X_310_ _426_/Q _425_/Q VGND VGND VPWR VPWR _310_/Y sky130_fd_sc_hd__xnor2_1
XTAP_192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_104 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_241_ _442_/D _249_/Y _297_/Y VGND VGND VPWR VPWR _241_/X sky130_fd_sc_hd__mux2_1
XFILLER_22_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_439_ _439_/CLK _439_/D fanout29/X VGND VGND VPWR VPWR _439_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_20_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_14 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_224_ _438_/Q _245_/Y _292_/Y VGND VGND VPWR VPWR _224_/X sky130_fd_sc_hd__mux2_1
XFILLER_10_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_207_ _444_/Q _207_/A1 _264_/Y VGND VGND VPWR VPWR _305_/B sky130_fd_sc_hd__mux2_1
XFILLER_24_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_91 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_386_ _260_/Y _272_/Y _385_/Y VGND VGND VPWR VPWR _448_/D sky130_fd_sc_hd__o21ai_1
X_455_ _455_/CLK _455_/D fanout28/X VGND VGND VPWR VPWR _455_/Q sky130_fd_sc_hd__dfrtp_2
XANTENNA_input3_A resetb VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_240_ _239_/X _327_/A _240_/S VGND VGND VPWR VPWR _240_/X sky130_fd_sc_hd__mux2_1
X_369_ _416_/D _432_/Q _431_/Q _433_/Q VGND VGND VPWR VPWR _369_/Y sky130_fd_sc_hd__nor4_1
X_438_ _206_/A1 _438_/D fanout29/X VGND VGND VPWR VPWR _438_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_13_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_26 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_223_ _222_/X _351_/A _223_/S VGND VGND VPWR VPWR _223_/X sky130_fd_sc_hd__mux2_1
XFILLER_12_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_206_ _206_/A0 _206_/A1 _413_/Q VGND VGND VPWR VPWR _206_/X sky130_fd_sc_hd__mux2_1
XFILLER_2_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_118 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_40 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__434__D _434_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_385_ _234_/S _385_/B _448_/Q VGND VGND VPWR VPWR _385_/Y sky130_fd_sc_hd__nand3b_1
X_454_ _455_/CLK _454_/D fanout28/X VGND VGND VPWR VPWR _454_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_31_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_368_ _225_/X _432_/Q _416_/D VGND VGND VPWR VPWR _432_/D sky130_fd_sc_hd__mux2_1
X_437_ _206_/A1 _437_/D fanout29/X VGND VGND VPWR VPWR _437_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_13_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_299_ _454_/Q _455_/Q VGND VGND VPWR VPWR _299_/Y sky130_fd_sc_hd__nor2_1
XFILLER_22_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_222_ _323_/Y _351_/A _295_/Y VGND VGND VPWR VPWR _222_/X sky130_fd_sc_hd__mux2_1
XFILLER_6_102 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_205_ _205_/A0 _415_/Q _413_/D VGND VGND VPWR VPWR _205_/X sky130_fd_sc_hd__mux2_1
XFILLER_3_105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_0_pll_clk90 pll_clk90 VGND VGND VPWR VPWR clkbuf_0_pll_clk90/X sky130_fd_sc_hd__clkbuf_16
XFILLER_18_92 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__214__A1 _311_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_51 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_384_ _258_/Y _272_/Y _383_/Y VGND VGND VPWR VPWR _446_/D sky130_fd_sc_hd__o21ai_1
X_453_ _455_/CLK _453_/D fanout28/X VGND VGND VPWR VPWR _453_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_23_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_170 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_0_ext_clk_A ext_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_367_ _224_/X _431_/Q _416_/D VGND VGND VPWR VPWR _431_/D sky130_fd_sc_hd__mux2_1
XANTENNA__279__B _311_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_436_ _439_/CLK _436_/D fanout29/X VGND VGND VPWR VPWR _439_/D sky130_fd_sc_hd__dfrtp_1
XFILLER_9_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_298_ _240_/S _298_/B VGND VGND VPWR VPWR _298_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_3_30 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_221_ _220_/X _311_/B _223_/S VGND VGND VPWR VPWR _221_/X sky130_fd_sc_hd__mux2_1
XFILLER_6_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_419_ _204_/A1 _419_/D _372_/S VGND VGND VPWR VPWR _419_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_5_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_204_ _419_/Q _204_/A1 _279_/Y VGND VGND VPWR VPWR _301_/B sky130_fd_sc_hd__mux2_1
XFILLER_3_117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_1_1__f_net10 clkbuf_0_net10/X VGND VGND VPWR VPWR _403__8/A sky130_fd_sc_hd__clkbuf_16
XTAP_322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_383_ _234_/S _385_/B _446_/Q VGND VGND VPWR VPWR _383_/Y sky130_fd_sc_hd__nand3b_1
X_452_ _455_/CLK _452_/D fanout28/X VGND VGND VPWR VPWR _452_/Q sky130_fd_sc_hd__dfrtn_1
XFILLER_31_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_182 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_297_ _457_/Q _373_/C VGND VGND VPWR VPWR _297_/Y sky130_fd_sc_hd__nand2_1
X_435_ _439_/CLK _435_/D _372_/S VGND VGND VPWR VPWR _438_/D sky130_fd_sc_hd__dfstp_1
X_366_ _219_/S _365_/Y _293_/Y _223_/X VGND VGND VPWR VPWR _430_/D sky130_fd_sc_hd__a2bb2o_1
XFILLER_9_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__280__B1 _311_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_input1_A ext_clk_sel VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_220_ _320_/Y _311_/B _295_/Y VGND VGND VPWR VPWR _220_/X sky130_fd_sc_hd__mux2_1
XFILLER_6_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_418_ _204_/A1 _439_/Q VGND VGND VPWR VPWR _418_/Q sky130_fd_sc_hd__dfxtp_1
X_349_ _417_/Q _438_/Q VGND VGND VPWR VPWR _353_/B sky130_fd_sc_hd__nand2b_1
XFILLER_3_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_203_ _298_/Y _240_/S _268_/Y VGND VGND VPWR VPWR _388_/S sky130_fd_sc_hd__mux2_1
XFILLER_0_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_382_ _445_/Q _265_/X _378_/Y _381_/Y VGND VGND VPWR VPWR _445_/D sky130_fd_sc_hd__o22a_1
X_451_ _451_/CLK _451_/D fanout28/X VGND VGND VPWR VPWR _451_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_31_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_408__3 _455_/CLK VGND VGND VPWR VPWR _451_/CLK sky130_fd_sc_hd__inv_4
XTAP_120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_296_ _458_/Q _459_/Q VGND VGND VPWR VPWR _373_/C sky130_fd_sc_hd__nor2_1
X_434_ _206_/A1 _434_/D _372_/S VGND VGND VPWR VPWR _437_/D sky130_fd_sc_hd__dfrtp_1
XFILLER_13_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_365_ _365_/A _430_/Q VGND VGND VPWR VPWR _365_/Y sky130_fd_sc_hd__nand2_1
XFILLER_9_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_279_ _439_/Q _311_/B VGND VGND VPWR VPWR _279_/Y sky130_fd_sc_hd__nor2_1
X_417_ _204_/A1 _438_/Q VGND VGND VPWR VPWR _417_/Q sky130_fd_sc_hd__dfxtp_1
X_348_ _438_/Q _417_/Q VGND VGND VPWR VPWR _353_/A sky130_fd_sc_hd__nand2b_1
XFILLER_5_160 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_202_ _293_/Y _219_/S _283_/Y VGND VGND VPWR VPWR _360_/S sky130_fd_sc_hd__mux2_1
XFILLER_0_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_381_ _379_/Y _380_/X _265_/X VGND VGND VPWR VPWR _381_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_17_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_450_ _455_/CLK _450_/D fanout28/X VGND VGND VPWR VPWR _450_/Q sky130_fd_sc_hd__dfrtn_1
XTAP_198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_433_ _204_/A1 _433_/D _372_/S VGND VGND VPWR VPWR _433_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_26_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__280__A2 _311_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_364_ _219_/S _363_/Y _293_/Y _221_/X VGND VGND VPWR VPWR _429_/D sky130_fd_sc_hd__a2bb2o_1
XFILLER_9_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_295_ _429_/Q _430_/Q _295_/C VGND VGND VPWR VPWR _295_/Y sky130_fd_sc_hd__nor3_2
XFILLER_3_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_347_ _347_/A _347_/B VGND VGND VPWR VPWR _419_/D sky130_fd_sc_hd__nand2_1
XANTENNA__459__RESET_B fanout28/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_416_ _204_/A1 _416_/D VGND VGND VPWR VPWR _416_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_12_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_278_ _426_/Q _427_/Q VGND VGND VPWR VPWR _278_/Y sky130_fd_sc_hd__nor2_2
XFILLER_5_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_405__5 _456_/CLK VGND VGND VPWR VPWR _424_/CLK sky130_fd_sc_hd__inv_4
XFILLER_5_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_66 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_380_ _465_/Q _443_/Q VGND VGND VPWR VPWR _380_/X sky130_fd_sc_hd__and2_1
XFILLER_15_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
.ends

