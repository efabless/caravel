magic
tech sky130A
magscale 1 2
timestamp 1681219932
<< obsli1 >>
rect 2024 2159 630936 950929
<< obsm1 >>
rect 934 2048 631842 952536
<< metal2 >>
rect 34749 952600 34805 953787
rect 35393 952600 35449 953787
rect 36037 952600 36093 953787
rect 37877 952600 37933 953787
rect 38429 952600 38485 953787
rect 39073 952600 39129 953787
rect 39717 952600 39773 953787
rect 42201 952600 42257 953787
rect 42753 952600 42809 953787
rect 43397 952600 43453 953787
rect 44041 952600 44097 953787
rect 45237 952600 45293 953787
rect 46433 952600 46489 953787
rect 47077 952600 47133 953787
rect 47721 952600 47777 953787
rect 48917 952600 48973 953787
rect 86149 952600 86205 953787
rect 86793 952600 86849 953787
rect 87437 952600 87493 953787
rect 89277 952600 89333 953787
rect 89829 952600 89885 953787
rect 90473 952600 90529 953787
rect 91117 952600 91173 953787
rect 93601 952600 93657 953787
rect 94153 952600 94209 953787
rect 94797 952600 94853 953787
rect 95441 952600 95497 953787
rect 96637 952600 96693 953787
rect 97833 952600 97889 953787
rect 98477 952600 98533 953787
rect 99121 952600 99177 953787
rect 100317 952600 100373 953787
rect 137549 952600 137605 953787
rect 138193 952600 138249 953787
rect 138837 952600 138893 953787
rect 140677 952600 140733 953787
rect 141229 952600 141285 953787
rect 141873 952600 141929 953787
rect 142517 952600 142573 953787
rect 145001 952600 145057 953787
rect 145553 952600 145609 953787
rect 146197 952600 146253 953787
rect 146841 952600 146897 953787
rect 148037 952600 148093 953787
rect 149233 952600 149289 953787
rect 149877 952600 149933 953787
rect 150521 952600 150577 953787
rect 151717 952600 151773 953787
rect 188949 952600 189005 953787
rect 189593 952600 189649 953787
rect 190237 952600 190293 953787
rect 192077 952600 192133 953787
rect 192629 952600 192685 953787
rect 193273 952600 193329 953787
rect 193917 952600 193973 953787
rect 196401 952600 196457 953787
rect 196953 952600 197009 953787
rect 197597 952600 197653 953787
rect 198241 952600 198297 953787
rect 199437 952600 199493 953787
rect 200633 952600 200689 953787
rect 201277 952600 201333 953787
rect 201921 952600 201977 953787
rect 203117 952600 203173 953787
rect 240549 952600 240605 953787
rect 241193 952600 241249 953787
rect 241837 952600 241893 953787
rect 243677 952600 243733 953787
rect 244229 952600 244285 953787
rect 244873 952600 244929 953787
rect 245517 952600 245573 953787
rect 248001 952600 248057 953787
rect 248553 952600 248609 953787
rect 249197 952600 249253 953787
rect 249841 952600 249897 953787
rect 251037 952600 251093 953787
rect 252233 952600 252289 953787
rect 252877 952600 252933 953787
rect 253521 952600 253577 953787
rect 254717 952600 254773 953787
rect 342349 952600 342405 953787
rect 342993 952600 343049 953787
rect 343637 952600 343693 953787
rect 345477 952600 345533 953787
rect 346029 952600 346085 953787
rect 346673 952600 346729 953787
rect 347317 952600 347373 953787
rect 349801 952600 349857 953787
rect 350353 952600 350409 953787
rect 350997 952600 351053 953787
rect 351641 952600 351697 953787
rect 352837 952600 352893 953787
rect 354033 952600 354089 953787
rect 354677 952600 354733 953787
rect 355321 952600 355377 953787
rect 356517 952600 356573 953787
rect 431349 952600 431405 953787
rect 431993 952600 432049 953787
rect 432637 952600 432693 953787
rect 434477 952600 434533 953787
rect 435029 952600 435085 953787
rect 435673 952600 435729 953787
rect 436317 952600 436373 953787
rect 438801 952600 438857 953787
rect 439353 952600 439409 953787
rect 439997 952600 440053 953787
rect 440641 952600 440697 953787
rect 441837 952600 441893 953787
rect 443033 952600 443089 953787
rect 443677 952600 443733 953787
rect 444321 952600 444377 953787
rect 445517 952600 445573 953787
rect 482749 952600 482805 953787
rect 483393 952600 483449 953787
rect 484037 952600 484093 953787
rect 485877 952600 485933 953787
rect 486429 952600 486485 953787
rect 487073 952600 487129 953787
rect 487717 952600 487773 953787
rect 490201 952600 490257 953787
rect 490753 952600 490809 953787
rect 491397 952600 491453 953787
rect 492041 952600 492097 953787
rect 493237 952600 493293 953787
rect 494433 952600 494489 953787
rect 495077 952600 495133 953787
rect 495721 952600 495777 953787
rect 496917 952600 496973 953787
rect 584549 952600 584605 953787
rect 585193 952600 585249 953787
rect 585837 952600 585893 953787
rect 587677 952600 587733 953787
rect 588229 952600 588285 953787
rect 588873 952600 588929 953787
rect 589517 952600 589573 953787
rect 592001 952600 592057 953787
rect 592553 952600 592609 953787
rect 593197 952600 593253 953787
rect 593841 952600 593897 953787
rect 595037 952600 595093 953787
rect 596233 952600 596289 953787
rect 596877 952600 596933 953787
rect 597521 952600 597577 953787
rect 598717 952600 598773 953787
rect 99367 -2105 99423 800
rect 145027 -400 145083 800
rect 151743 -400 151799 800
rect 264667 -400 264723 800
rect 265955 -400 266011 800
rect 267795 -400 267851 800
rect 319467 -400 319523 800
rect 322595 -400 322651 800
rect 363227 -400 363283 800
rect 369943 -400 369999 800
rect 374267 -400 374323 800
rect 377395 -400 377451 800
rect 418027 -400 418083 800
rect 424743 -400 424799 800
rect 429067 -400 429123 800
rect 432195 -400 432251 800
rect 472827 -400 472883 800
rect 478347 -400 478403 800
rect 479543 -400 479599 800
rect 482671 -400 482727 800
rect 483867 -400 483923 800
rect 486995 -400 487051 800
<< obsm2 >>
rect 938 952544 34693 952762
rect 34861 952544 35337 952762
rect 35505 952544 35981 952762
rect 36149 952544 37821 952762
rect 37989 952544 38373 952762
rect 38541 952544 39017 952762
rect 39185 952544 39661 952762
rect 39829 952544 42145 952762
rect 42313 952544 42697 952762
rect 42865 952544 43341 952762
rect 43509 952544 43985 952762
rect 44153 952544 45181 952762
rect 45349 952544 46377 952762
rect 46545 952544 47021 952762
rect 47189 952544 47665 952762
rect 47833 952544 48861 952762
rect 49029 952544 86093 952762
rect 86261 952544 86737 952762
rect 86905 952544 87381 952762
rect 87549 952544 89221 952762
rect 89389 952544 89773 952762
rect 89941 952544 90417 952762
rect 90585 952544 91061 952762
rect 91229 952544 93545 952762
rect 93713 952544 94097 952762
rect 94265 952544 94741 952762
rect 94909 952544 95385 952762
rect 95553 952544 96581 952762
rect 96749 952544 97777 952762
rect 97945 952544 98421 952762
rect 98589 952544 99065 952762
rect 99233 952544 100261 952762
rect 100429 952544 137493 952762
rect 137661 952544 138137 952762
rect 138305 952544 138781 952762
rect 138949 952544 140621 952762
rect 140789 952544 141173 952762
rect 141341 952544 141817 952762
rect 141985 952544 142461 952762
rect 142629 952544 144945 952762
rect 145113 952544 145497 952762
rect 145665 952544 146141 952762
rect 146309 952544 146785 952762
rect 146953 952544 147981 952762
rect 148149 952544 149177 952762
rect 149345 952544 149821 952762
rect 149989 952544 150465 952762
rect 150633 952544 151661 952762
rect 151829 952544 188893 952762
rect 189061 952544 189537 952762
rect 189705 952544 190181 952762
rect 190349 952544 192021 952762
rect 192189 952544 192573 952762
rect 192741 952544 193217 952762
rect 193385 952544 193861 952762
rect 194029 952544 196345 952762
rect 196513 952544 196897 952762
rect 197065 952544 197541 952762
rect 197709 952544 198185 952762
rect 198353 952544 199381 952762
rect 199549 952544 200577 952762
rect 200745 952544 201221 952762
rect 201389 952544 201865 952762
rect 202033 952544 203061 952762
rect 203229 952544 240493 952762
rect 240661 952544 241137 952762
rect 241305 952544 241781 952762
rect 241949 952544 243621 952762
rect 243789 952544 244173 952762
rect 244341 952544 244817 952762
rect 244985 952544 245461 952762
rect 245629 952544 247945 952762
rect 248113 952544 248497 952762
rect 248665 952544 249141 952762
rect 249309 952544 249785 952762
rect 249953 952544 250981 952762
rect 251149 952544 252177 952762
rect 252345 952544 252821 952762
rect 252989 952544 253465 952762
rect 253633 952544 254661 952762
rect 254829 952544 342293 952762
rect 342461 952544 342937 952762
rect 343105 952544 343581 952762
rect 343749 952544 345421 952762
rect 345589 952544 345973 952762
rect 346141 952544 346617 952762
rect 346785 952544 347261 952762
rect 347429 952544 349745 952762
rect 349913 952544 350297 952762
rect 350465 952544 350941 952762
rect 351109 952544 351585 952762
rect 351753 952544 352781 952762
rect 352949 952544 353977 952762
rect 354145 952544 354621 952762
rect 354789 952544 355265 952762
rect 355433 952544 356461 952762
rect 356629 952544 431293 952762
rect 431461 952544 431937 952762
rect 432105 952544 432581 952762
rect 432749 952544 434421 952762
rect 434589 952544 434973 952762
rect 435141 952544 435617 952762
rect 435785 952544 436261 952762
rect 436429 952544 438745 952762
rect 438913 952544 439297 952762
rect 439465 952544 439941 952762
rect 440109 952544 440585 952762
rect 440753 952544 441781 952762
rect 441949 952544 442977 952762
rect 443145 952544 443621 952762
rect 443789 952544 444265 952762
rect 444433 952544 445461 952762
rect 445629 952544 482693 952762
rect 482861 952544 483337 952762
rect 483505 952544 483981 952762
rect 484149 952544 485821 952762
rect 485989 952544 486373 952762
rect 486541 952544 487017 952762
rect 487185 952544 487661 952762
rect 487829 952544 490145 952762
rect 490313 952544 490697 952762
rect 490865 952544 491341 952762
rect 491509 952544 491985 952762
rect 492153 952544 493181 952762
rect 493349 952544 494377 952762
rect 494545 952544 495021 952762
rect 495189 952544 495665 952762
rect 495833 952544 496861 952762
rect 497029 952544 584493 952762
rect 584661 952544 585137 952762
rect 585305 952544 585781 952762
rect 585949 952544 587621 952762
rect 587789 952544 588173 952762
rect 588341 952544 588817 952762
rect 588985 952544 589461 952762
rect 589629 952544 591945 952762
rect 592113 952544 592497 952762
rect 592665 952544 593141 952762
rect 593309 952544 593785 952762
rect 593953 952544 594981 952762
rect 595149 952544 596177 952762
rect 596345 952544 596821 952762
rect 596989 952544 597465 952762
rect 597633 952544 598661 952762
rect 598829 952544 631838 952762
rect 938 856 631838 952544
rect 938 734 99311 856
rect 99479 734 144971 856
rect 145139 734 151687 856
rect 151855 734 264611 856
rect 264779 734 265899 856
rect 266067 734 267739 856
rect 267907 734 319411 856
rect 319579 734 322539 856
rect 322707 734 363171 856
rect 363339 734 369887 856
rect 370055 734 374211 856
rect 374379 734 377339 856
rect 377507 734 417971 856
rect 418139 734 424687 856
rect 424855 734 429011 856
rect 429179 734 432139 856
rect 432307 734 472771 856
rect 472939 734 478291 856
rect 478459 734 479487 856
rect 479655 734 482615 856
rect 482783 734 483811 856
rect 483979 734 486939 856
rect 487107 734 631838 856
<< metal3 >>
rect -437 927085 800 927205
rect -437 925889 800 926009
rect -437 925245 800 925365
rect -437 924601 800 924721
rect 632200 924563 633437 924683
rect 632200 923919 633437 924039
rect -437 923405 800 923525
rect 632200 923275 633437 923395
rect -437 922209 800 922329
rect -437 921565 800 921685
rect 632200 921435 633437 921555
rect -437 920921 800 921041
rect 632200 920883 633437 921003
rect -437 920369 800 920489
rect 632200 920239 633437 920359
rect 632200 919595 633437 919715
rect -437 917885 800 918005
rect -437 917241 800 917361
rect 632200 917111 633437 917231
rect -437 916597 800 916717
rect 632200 916559 633437 916679
rect -437 916045 800 916165
rect 632200 915915 633437 916035
rect 632200 915271 633437 915391
rect -437 914205 800 914325
rect 632200 914075 633437 914195
rect -437 913561 800 913681
rect -437 912917 800 913037
rect 632200 912879 633437 912999
rect 632200 912235 633437 912355
rect 632200 911591 633437 911711
rect 632200 910395 633437 910515
rect 632200 835363 633437 835483
rect 632200 834719 633437 834839
rect 632200 834075 633437 834195
rect 632200 832235 633437 832355
rect 632200 831683 633437 831803
rect 632200 831039 633437 831159
rect 632200 830395 633437 830515
rect 632200 827911 633437 828031
rect 632200 827359 633437 827479
rect 632200 826715 633437 826835
rect 632200 826071 633437 826191
rect 632200 824875 633437 824995
rect 632200 823679 633437 823799
rect 632200 823035 633437 823155
rect 632200 822391 633437 822511
rect 632200 821195 633437 821315
rect -437 757285 800 757405
rect -437 756089 800 756209
rect -437 755445 800 755565
rect -437 754801 800 754921
rect -437 753605 800 753725
rect -437 752409 800 752529
rect -437 751765 800 751885
rect -437 751121 800 751241
rect -437 750569 800 750689
rect -437 748085 800 748205
rect -437 747441 800 747561
rect -437 746797 800 746917
rect -437 746245 800 746365
rect 632200 746163 633437 746283
rect 632200 745519 633437 745639
rect 632200 744875 633437 744995
rect -437 744405 800 744525
rect -437 743761 800 743881
rect -437 743117 800 743237
rect 632200 743035 633437 743155
rect 632200 742483 633437 742603
rect 632200 741839 633437 741959
rect 632200 741195 633437 741315
rect 632200 738711 633437 738831
rect 632200 738159 633437 738279
rect 632200 737515 633437 737635
rect 632200 736871 633437 736991
rect 632200 735675 633437 735795
rect 632200 734479 633437 734599
rect 632200 733835 633437 733955
rect 632200 733191 633437 733311
rect 632200 731995 633437 732115
rect -437 714085 800 714205
rect -437 712889 800 713009
rect -437 712245 800 712365
rect -437 711601 800 711721
rect -437 710405 800 710525
rect -437 709209 800 709329
rect -437 708565 800 708685
rect -437 707921 800 708041
rect -437 707369 800 707489
rect -437 704885 800 705005
rect -437 704241 800 704361
rect -437 703597 800 703717
rect -437 703045 800 703165
rect -437 701205 800 701325
rect 632200 701163 633437 701283
rect -437 700561 800 700681
rect 632200 700519 633437 700639
rect -437 699917 800 700037
rect 632200 699875 633437 699995
rect 632200 698035 633437 698155
rect 632200 697483 633437 697603
rect 632200 696839 633437 696959
rect 632200 696195 633437 696315
rect 632200 693711 633437 693831
rect 632200 693159 633437 693279
rect 632200 692515 633437 692635
rect 632200 691871 633437 691991
rect 632200 690675 633437 690795
rect 632200 689479 633437 689599
rect 632200 688835 633437 688955
rect 632200 688191 633437 688311
rect 632200 686995 633437 687115
rect -437 670885 800 671005
rect -437 669689 800 669809
rect -437 669045 800 669165
rect -437 668401 800 668521
rect -437 667205 800 667325
rect -437 666009 800 666129
rect -437 665365 800 665485
rect -437 664721 800 664841
rect -437 664169 800 664289
rect -437 661685 800 661805
rect -437 661041 800 661161
rect -437 660397 800 660517
rect -437 659845 800 659965
rect -437 658005 800 658125
rect -437 657361 800 657481
rect -437 656717 800 656837
rect 632200 656163 633437 656283
rect 632200 655519 633437 655639
rect 632200 654875 633437 654995
rect 632200 653035 633437 653155
rect 632200 652483 633437 652603
rect 632200 651839 633437 651959
rect 632200 651195 633437 651315
rect 632200 648711 633437 648831
rect 632200 648159 633437 648279
rect 632200 647515 633437 647635
rect 632200 646871 633437 646991
rect 632200 645675 633437 645795
rect 632200 644479 633437 644599
rect 632200 643835 633437 643955
rect 632200 643191 633437 643311
rect 632200 641995 633437 642115
rect -437 627685 800 627805
rect -437 626489 800 626609
rect -437 625845 800 625965
rect -437 625201 800 625321
rect -437 624005 800 624125
rect -437 622809 858 622929
rect -437 622165 800 622285
rect -437 621521 800 621641
rect -437 620969 800 621089
rect -437 618485 800 618605
rect -437 617841 800 617961
rect -437 617197 800 617317
rect -437 616645 800 616765
rect -437 614805 800 614925
rect -437 614161 800 614281
rect -437 613517 800 613637
rect 632200 610963 633437 611083
rect 632200 610319 633437 610439
rect 632200 609675 633437 609795
rect 632200 607835 633437 607955
rect 632200 607283 633437 607403
rect 632200 606639 633437 606759
rect 632200 605995 633437 606115
rect 632200 603511 633437 603631
rect 632200 602959 633437 603079
rect 632200 602315 633437 602435
rect 632200 601671 633437 601791
rect 632200 600475 633437 600595
rect 632200 599279 633437 599399
rect 632200 598635 633437 598755
rect 632200 597991 633437 598111
rect 632200 596795 633437 596915
rect -437 584485 800 584605
rect -437 583289 800 583409
rect -437 582645 800 582765
rect -437 582001 800 582121
rect -437 580805 800 580925
rect -437 579609 800 579729
rect -437 578965 800 579085
rect -437 578321 800 578441
rect -437 577769 800 577889
rect -437 575285 800 575405
rect -437 574641 800 574761
rect -437 573997 800 574117
rect -437 573445 800 573565
rect -437 571605 800 571725
rect -437 570961 800 571081
rect -437 570317 800 570437
rect 632200 565963 633437 566083
rect 632200 565319 633437 565439
rect 632200 564675 633437 564795
rect 632200 562835 633437 562955
rect 632200 562283 633437 562403
rect 632200 561639 633437 561759
rect 632200 560995 633437 561115
rect 632200 558511 633437 558631
rect 632200 557959 633437 558079
rect 632200 557315 633437 557435
rect 632200 556671 633437 556791
rect 632200 555475 633437 555595
rect 632200 554279 633437 554399
rect 632200 553635 633437 553755
rect 632200 552991 633437 553111
rect 632200 551795 633437 551915
rect -437 541285 800 541405
rect -437 540089 800 540209
rect -437 539445 800 539565
rect -437 538801 800 538921
rect -437 537605 800 537725
rect -437 536409 800 536529
rect -437 535765 800 535885
rect -437 535121 800 535241
rect -437 534569 800 534689
rect -437 532085 800 532205
rect -437 531441 800 531561
rect -437 530797 800 530917
rect -437 530245 800 530365
rect -437 528405 800 528525
rect -437 527761 800 527881
rect -437 527117 800 527237
rect 632200 520763 633437 520883
rect 632200 520119 633437 520239
rect 632200 519475 633437 519595
rect 632200 517635 633437 517755
rect 632200 517083 633437 517203
rect 632200 516439 633437 516559
rect 632200 515795 633437 515915
rect 632200 513311 633437 513431
rect 632200 512759 633437 512879
rect 632200 512115 633437 512235
rect 632200 511471 633437 511591
rect 632200 510275 633437 510395
rect 632200 509079 633437 509199
rect 632200 508435 633437 508555
rect 632200 507791 633437 507911
rect 632200 506595 633437 506715
rect -437 498085 800 498205
rect -437 496889 800 497009
rect -437 496245 800 496365
rect -437 495601 800 495721
rect -437 494405 800 494525
rect -437 493209 800 493329
rect -437 492565 800 492685
rect -437 491921 800 492041
rect -437 491369 800 491489
rect -437 488885 800 489005
rect -437 488241 800 488361
rect -437 487597 800 487717
rect -437 487045 800 487165
rect -437 485205 800 485325
rect -437 484561 800 484681
rect -437 483917 800 484037
rect -437 370485 800 370605
rect -437 369289 800 369409
rect -437 368645 800 368765
rect -437 368001 800 368121
rect -437 366805 800 366925
rect -437 365609 800 365729
rect -437 364965 800 365085
rect -437 364321 800 364441
rect -437 363769 800 363889
rect -437 361285 800 361405
rect -437 360641 800 360761
rect -437 359997 800 360117
rect -437 359445 800 359565
rect -437 357605 800 357725
rect -437 356961 800 357081
rect -437 356317 800 356437
rect 632200 343563 633437 343683
rect 632200 342919 633437 343039
rect 632200 342275 633437 342395
rect 632200 340435 633437 340555
rect 632200 339883 633437 340003
rect 632200 339239 633437 339359
rect 632200 338595 633437 338715
rect 632200 336111 633437 336231
rect 632200 335559 633437 335679
rect 632200 334915 633437 335035
rect 632200 334271 633437 334391
rect 632200 333075 633437 333195
rect 632200 331235 633437 331355
rect 632200 330591 633437 330711
rect 632200 329395 633437 329515
rect -437 327285 800 327405
rect -437 326089 800 326209
rect -437 325445 800 325565
rect -437 324801 800 324921
rect -437 323605 800 323725
rect -437 322409 800 322529
rect -437 321765 800 321885
rect -437 321121 800 321241
rect -437 320569 800 320689
rect -437 318085 800 318205
rect -437 317441 800 317561
rect -437 316797 800 316917
rect -437 316245 800 316365
rect -437 314405 800 314525
rect -437 313761 800 313881
rect -437 313117 800 313237
rect 632200 298363 633437 298483
rect 632200 297719 633437 297839
rect 632200 297075 633437 297195
rect 632200 295235 633437 295355
rect 632200 294683 633437 294803
rect 632200 294039 633437 294159
rect 632200 293395 633437 293515
rect 632200 290911 633437 291031
rect 632200 290359 633437 290479
rect 632200 289715 633437 289835
rect 632200 289071 633437 289191
rect 632200 287875 633437 287995
rect 632200 286035 633437 286155
rect 632200 285391 633437 285511
rect -437 284085 800 284205
rect 632200 284195 633437 284315
rect -437 282889 800 283009
rect -437 282245 800 282365
rect -437 281601 800 281721
rect -437 280405 800 280525
rect -437 279209 800 279329
rect -437 278565 800 278685
rect -437 277921 800 278041
rect -437 277369 800 277489
rect -437 274885 800 275005
rect -437 274241 800 274361
rect -437 273597 800 273717
rect -437 273045 800 273165
rect -437 271205 800 271325
rect -437 270561 800 270681
rect -437 269917 800 270037
rect 632200 253363 633437 253483
rect 632200 252719 633437 252839
rect 632200 252075 633437 252195
rect 632200 250235 633437 250355
rect 632200 249683 633437 249803
rect 632200 249039 633437 249159
rect 632200 248395 633437 248515
rect 632200 245911 633437 246031
rect 632200 245359 633437 245479
rect 632200 244715 633437 244835
rect 632200 244071 633437 244191
rect 632200 242875 633437 242995
rect -437 240885 800 241005
rect 632200 241035 633437 241155
rect 632200 240391 633437 240511
rect -437 239689 858 239809
rect -437 239045 800 239165
rect 632200 239195 633437 239315
rect -437 238401 800 238521
rect -437 237205 800 237325
rect -437 236009 800 236129
rect -437 235365 858 235485
rect -437 234721 800 234841
rect -437 234169 800 234289
rect -437 231685 800 231805
rect -437 231041 800 231161
rect -437 230397 800 230517
rect -437 229845 800 229965
rect -437 228005 800 228125
rect -437 227361 800 227481
rect -437 226717 800 226837
rect 632200 208363 633437 208483
rect 632200 207719 633437 207839
rect 632200 207075 633437 207195
rect 632200 205235 633437 205355
rect 632200 204683 633437 204803
rect 632200 204039 633437 204159
rect 632200 203395 633437 203515
rect 632200 200911 633437 201031
rect 632200 200359 633437 200479
rect 632200 199715 633437 199835
rect 632200 199071 633437 199191
rect -437 197685 800 197805
rect 632200 197875 633437 197995
rect -437 196489 800 196609
rect -437 195845 800 195965
rect 632200 196035 633437 196155
rect 632200 195391 633437 195511
rect -437 194005 800 194125
rect 632200 194195 633437 194315
rect -437 192809 800 192929
rect -437 192165 800 192285
rect -437 191521 800 191641
rect -437 190969 800 191089
rect -437 188485 800 188605
rect -437 187841 800 187961
rect -437 187197 800 187317
rect -437 186645 800 186765
rect -437 184805 800 184925
rect -437 184161 800 184281
rect -437 183517 800 183637
rect 632200 163163 633437 163283
rect 632200 162519 633437 162639
rect 632200 161875 633437 161995
rect 632200 160035 633437 160155
rect 632200 159483 633437 159603
rect 632200 158839 633437 158959
rect 632200 158195 633437 158315
rect 632200 155711 633437 155831
rect 632200 155159 633437 155279
rect -437 154485 800 154605
rect 632200 154515 633437 154635
rect 632200 153871 633437 153991
rect -437 153289 800 153409
rect -437 152645 800 152765
rect 632200 152675 633437 152795
rect -437 150805 800 150925
rect 632200 150835 633437 150955
rect 632200 150191 633437 150311
rect -437 149609 800 149729
rect -437 148965 800 149085
rect 632200 148995 633437 149115
rect -437 148321 800 148441
rect -437 147769 800 147889
rect -437 145285 800 145405
rect -437 144641 800 144761
rect -437 143997 800 144117
rect -437 143445 800 143565
rect -437 141605 800 141725
rect -437 140961 800 141081
rect -437 140317 800 140437
rect 632200 118163 633437 118283
rect 632200 117519 633437 117639
rect 632200 116875 633437 116995
rect 632200 115035 633437 115155
rect 632200 114483 633437 114603
rect 632200 113839 633437 113959
rect 632200 113195 633437 113315
rect 632200 110711 633437 110831
rect 632200 110159 633437 110279
rect 632200 109515 633437 109635
rect 632200 108871 633437 108991
rect 632200 107675 633437 107795
rect 632200 105835 633437 105955
rect 632200 105191 633437 105311
rect 632200 103995 633437 104115
rect 632200 72963 633437 73083
rect 632200 72319 633437 72439
rect 632200 71675 633437 71795
rect 632200 69835 633437 69955
rect 632200 69283 633437 69403
rect 632200 68639 633437 68759
rect 632200 67995 633437 68115
rect 632200 65511 633437 65631
rect 632200 64959 633437 65079
rect 632200 64315 633437 64435
rect 632200 63671 633437 63791
rect 632200 62475 633437 62595
rect 632200 60635 633437 60755
rect 632200 59991 633437 60111
rect 632200 58795 633437 58915
<< obsm3 >>
rect 533387 953400 538193 955596
rect 543368 953400 548174 955596
rect 0 927285 633000 953400
rect 880 927005 633000 927285
rect 0 926089 633000 927005
rect 880 925809 633000 926089
rect 0 925445 633000 925809
rect 880 925165 633000 925445
rect 0 924801 633000 925165
rect 880 924763 633000 924801
rect 880 924521 632120 924763
rect 0 924483 632120 924521
rect 0 924119 633000 924483
rect 0 923839 632120 924119
rect 0 923605 633000 923839
rect 880 923475 633000 923605
rect 880 923325 632120 923475
rect 0 923195 632120 923325
rect 0 922409 633000 923195
rect 880 922129 633000 922409
rect 0 921765 633000 922129
rect 880 921635 633000 921765
rect 880 921485 632120 921635
rect 0 921355 632120 921485
rect 0 921121 633000 921355
rect 880 921083 633000 921121
rect 880 920841 632120 921083
rect 0 920803 632120 920841
rect 0 920569 633000 920803
rect 880 920439 633000 920569
rect 880 920289 632120 920439
rect 0 920159 632120 920289
rect 0 919795 633000 920159
rect 0 919515 632120 919795
rect 0 918085 633000 919515
rect 880 917805 633000 918085
rect 0 917441 633000 917805
rect 880 917311 633000 917441
rect 880 917161 632120 917311
rect 0 917031 632120 917161
rect 0 916797 633000 917031
rect 880 916759 633000 916797
rect 880 916517 632120 916759
rect 0 916479 632120 916517
rect 0 916245 633000 916479
rect 880 916115 633000 916245
rect 880 915965 632120 916115
rect 0 915835 632120 915965
rect 0 915471 633000 915835
rect 0 915191 632120 915471
rect 0 914405 633000 915191
rect 880 914275 633000 914405
rect 880 914125 632120 914275
rect 0 913995 632120 914125
rect 0 913761 633000 913995
rect 880 913481 633000 913761
rect 0 913117 633000 913481
rect 880 913079 633000 913117
rect 880 912837 632120 913079
rect 0 912799 632120 912837
rect 0 912435 633000 912799
rect 0 912155 632120 912435
rect 0 911791 633000 912155
rect 0 911511 632120 911791
rect 0 910595 633000 911511
rect 0 910315 632120 910595
rect 0 884840 633000 910315
rect -3216 880400 633000 884840
rect -3216 880051 635604 880400
rect 0 879730 635604 880051
rect -2200 875611 635604 879730
rect -2200 875290 633000 875611
rect -2200 875120 635204 875290
rect 0 874800 635204 875120
rect -3216 870669 635204 874800
rect -3216 870349 633000 870669
rect -3216 870011 635604 870349
rect 0 865560 635604 870011
rect 0 835563 633000 865560
rect 0 835283 632120 835563
rect 0 834919 633000 835283
rect 0 834639 632120 834919
rect 0 834275 633000 834639
rect 0 833995 632120 834275
rect 0 832435 633000 833995
rect 0 832155 632120 832435
rect 0 831883 633000 832155
rect 0 831603 632120 831883
rect 0 831239 633000 831603
rect 0 830959 632120 831239
rect 0 830595 633000 830959
rect 0 830315 632120 830595
rect 0 828111 633000 830315
rect 0 827831 632120 828111
rect 0 827559 633000 827831
rect 0 827279 632120 827559
rect 0 826915 633000 827279
rect 0 826635 632120 826915
rect 0 826271 633000 826635
rect 0 825991 632120 826271
rect 0 825075 633000 825991
rect 0 824795 632120 825075
rect 0 823879 633000 824795
rect 0 823599 632120 823879
rect 0 823235 633000 823599
rect 0 822955 632120 823235
rect 0 822591 633000 822955
rect 0 822311 632120 822591
rect 0 821395 633000 822311
rect 0 821115 632120 821395
rect 0 800358 633000 821115
rect -3216 795569 633000 800358
rect 0 791201 633000 795569
rect 0 790379 635604 791201
rect -3216 786412 635604 790379
rect -3216 785590 633000 786412
rect 0 781218 633000 785590
rect 0 776429 635604 781218
rect 0 757485 633000 776429
rect 880 757205 633000 757485
rect 0 756289 633000 757205
rect 880 756009 633000 756289
rect 0 755645 633000 756009
rect 880 755365 633000 755645
rect 0 755001 633000 755365
rect 880 754721 633000 755001
rect 0 753805 633000 754721
rect 880 753525 633000 753805
rect 0 752609 633000 753525
rect 880 752329 633000 752609
rect 0 751965 633000 752329
rect 880 751685 633000 751965
rect 0 751321 633000 751685
rect 880 751041 633000 751321
rect 0 750769 633000 751041
rect 880 750489 633000 750769
rect 0 748285 633000 750489
rect 880 748005 633000 748285
rect 0 747641 633000 748005
rect 880 747361 633000 747641
rect 0 746997 633000 747361
rect 880 746717 633000 746997
rect 0 746445 633000 746717
rect 880 746363 633000 746445
rect 880 746165 632120 746363
rect 0 746083 632120 746165
rect 0 745719 633000 746083
rect 0 745439 632120 745719
rect 0 745075 633000 745439
rect 0 744795 632120 745075
rect 0 744605 633000 744795
rect 880 744325 633000 744605
rect 0 743961 633000 744325
rect 880 743681 633000 743961
rect 0 743317 633000 743681
rect 880 743235 633000 743317
rect 880 743037 632120 743235
rect 0 742955 632120 743037
rect 0 742683 633000 742955
rect 0 742403 632120 742683
rect 0 742039 633000 742403
rect 0 741759 632120 742039
rect 0 741395 633000 741759
rect 0 741115 632120 741395
rect 0 738911 633000 741115
rect 0 738631 632120 738911
rect 0 738359 633000 738631
rect 0 738079 632120 738359
rect 0 737715 633000 738079
rect 0 737435 632120 737715
rect 0 737071 633000 737435
rect 0 736791 632120 737071
rect 0 735875 633000 736791
rect 0 735595 632120 735875
rect 0 734679 633000 735595
rect 0 734399 632120 734679
rect 0 734035 633000 734399
rect 0 733755 632120 734035
rect 0 733391 633000 733755
rect 0 733111 632120 733391
rect 0 732195 633000 733111
rect 0 731915 632120 732195
rect 0 714285 633000 731915
rect 880 714005 633000 714285
rect 0 713089 633000 714005
rect 880 712809 633000 713089
rect 0 712445 633000 712809
rect 880 712165 633000 712445
rect 0 711801 633000 712165
rect 880 711521 633000 711801
rect 0 710605 633000 711521
rect 880 710325 633000 710605
rect 0 709409 633000 710325
rect 880 709129 633000 709409
rect 0 708765 633000 709129
rect 880 708485 633000 708765
rect 0 708121 633000 708485
rect 880 707841 633000 708121
rect 0 707569 633000 707841
rect 880 707289 633000 707569
rect 0 705085 633000 707289
rect 880 704805 633000 705085
rect 0 704441 633000 704805
rect 880 704161 633000 704441
rect 0 703797 633000 704161
rect 880 703517 633000 703797
rect 0 703245 633000 703517
rect 880 702965 633000 703245
rect 0 701405 633000 702965
rect 880 701363 633000 701405
rect 880 701125 632120 701363
rect 0 701083 632120 701125
rect 0 700761 633000 701083
rect 880 700719 633000 700761
rect 880 700481 632120 700719
rect 0 700439 632120 700481
rect 0 700117 633000 700439
rect 880 700075 633000 700117
rect 880 699837 632120 700075
rect 0 699795 632120 699837
rect 0 698235 633000 699795
rect 0 697955 632120 698235
rect 0 697683 633000 697955
rect 0 697403 632120 697683
rect 0 697039 633000 697403
rect 0 696759 632120 697039
rect 0 696395 633000 696759
rect 0 696115 632120 696395
rect 0 693911 633000 696115
rect 0 693631 632120 693911
rect 0 693359 633000 693631
rect 0 693079 632120 693359
rect 0 692715 633000 693079
rect 0 692435 632120 692715
rect 0 692071 633000 692435
rect 0 691791 632120 692071
rect 0 690875 633000 691791
rect 0 690595 632120 690875
rect 0 689679 633000 690595
rect 0 689399 632120 689679
rect 0 689035 633000 689399
rect 0 688755 632120 689035
rect 0 688391 633000 688755
rect 0 688111 632120 688391
rect 0 687195 633000 688111
rect 0 686915 632120 687195
rect 0 671085 633000 686915
rect 880 670805 633000 671085
rect 0 669889 633000 670805
rect 880 669609 633000 669889
rect 0 669245 633000 669609
rect 880 668965 633000 669245
rect 0 668601 633000 668965
rect 880 668321 633000 668601
rect 0 667405 633000 668321
rect 880 667125 633000 667405
rect 0 666209 633000 667125
rect 880 665929 633000 666209
rect 0 665565 633000 665929
rect 880 665285 633000 665565
rect 0 664921 633000 665285
rect 880 664641 633000 664921
rect 0 664369 633000 664641
rect 880 664089 633000 664369
rect 0 661885 633000 664089
rect 880 661605 633000 661885
rect 0 661241 633000 661605
rect 880 660961 633000 661241
rect 0 660597 633000 660961
rect 880 660317 633000 660597
rect 0 660045 633000 660317
rect 880 659765 633000 660045
rect 0 658205 633000 659765
rect 880 657925 633000 658205
rect 0 657561 633000 657925
rect 880 657281 633000 657561
rect 0 656917 633000 657281
rect 880 656637 633000 656917
rect 0 656363 633000 656637
rect 0 656083 632120 656363
rect 0 655719 633000 656083
rect 0 655439 632120 655719
rect 0 655075 633000 655439
rect 0 654795 632120 655075
rect 0 653235 633000 654795
rect 0 652955 632120 653235
rect 0 652683 633000 652955
rect 0 652403 632120 652683
rect 0 652039 633000 652403
rect 0 651759 632120 652039
rect 0 651395 633000 651759
rect 0 651115 632120 651395
rect 0 648911 633000 651115
rect 0 648631 632120 648911
rect 0 648359 633000 648631
rect 0 648079 632120 648359
rect 0 647715 633000 648079
rect 0 647435 632120 647715
rect 0 647071 633000 647435
rect 0 646791 632120 647071
rect 0 645875 633000 646791
rect 0 645595 632120 645875
rect 0 644679 633000 645595
rect 0 644399 632120 644679
rect 0 644035 633000 644399
rect 0 643755 632120 644035
rect 0 643391 633000 643755
rect 0 643111 632120 643391
rect 0 642195 633000 643111
rect 0 641915 632120 642195
rect 0 627885 633000 641915
rect 880 627605 633000 627885
rect 0 626689 633000 627605
rect 880 626409 633000 626689
rect 0 626045 633000 626409
rect 880 625765 633000 626045
rect 0 625401 633000 625765
rect 880 625121 633000 625401
rect 0 624205 633000 625121
rect 880 623925 633000 624205
rect 0 623009 633000 623925
rect 938 622729 633000 623009
rect 0 622365 633000 622729
rect 880 622085 633000 622365
rect 0 621721 633000 622085
rect 880 621441 633000 621721
rect 0 621169 633000 621441
rect 880 620889 633000 621169
rect 0 618685 633000 620889
rect 880 618405 633000 618685
rect 0 618041 633000 618405
rect 880 617761 633000 618041
rect 0 617397 633000 617761
rect 880 617117 633000 617397
rect 0 616845 633000 617117
rect 880 616565 633000 616845
rect 0 615005 633000 616565
rect 880 614725 633000 615005
rect 0 614361 633000 614725
rect 880 614081 633000 614361
rect 0 613717 633000 614081
rect 880 613437 633000 613717
rect 0 611163 633000 613437
rect 0 610883 632120 611163
rect 0 610519 633000 610883
rect 0 610239 632120 610519
rect 0 609875 633000 610239
rect 0 609595 632120 609875
rect 0 608035 633000 609595
rect 0 607755 632120 608035
rect 0 607483 633000 607755
rect 0 607203 632120 607483
rect 0 606839 633000 607203
rect 0 606559 632120 606839
rect 0 606195 633000 606559
rect 0 605915 632120 606195
rect 0 603711 633000 605915
rect 0 603431 632120 603711
rect 0 603159 633000 603431
rect 0 602879 632120 603159
rect 0 602515 633000 602879
rect 0 602235 632120 602515
rect 0 601871 633000 602235
rect 0 601591 632120 601871
rect 0 600675 633000 601591
rect 0 600395 632120 600675
rect 0 599479 633000 600395
rect 0 599199 632120 599479
rect 0 598835 633000 599199
rect 0 598555 632120 598835
rect 0 598191 633000 598555
rect 0 597911 632120 598191
rect 0 596995 633000 597911
rect 0 596715 632120 596995
rect 0 584685 633000 596715
rect 880 584405 633000 584685
rect 0 583489 633000 584405
rect 880 583209 633000 583489
rect 0 582845 633000 583209
rect 880 582565 633000 582845
rect 0 582201 633000 582565
rect 880 581921 633000 582201
rect 0 581005 633000 581921
rect 880 580725 633000 581005
rect 0 579809 633000 580725
rect 880 579529 633000 579809
rect 0 579165 633000 579529
rect 880 578885 633000 579165
rect 0 578521 633000 578885
rect 880 578241 633000 578521
rect 0 577969 633000 578241
rect 880 577689 633000 577969
rect 0 575485 633000 577689
rect 880 575205 633000 575485
rect 0 574841 633000 575205
rect 880 574561 633000 574841
rect 0 574197 633000 574561
rect 880 573917 633000 574197
rect 0 573645 633000 573917
rect 880 573365 633000 573645
rect 0 571805 633000 573365
rect 880 571525 633000 571805
rect 0 571161 633000 571525
rect 880 570881 633000 571161
rect 0 570517 633000 570881
rect 880 570237 633000 570517
rect 0 566163 633000 570237
rect 0 565883 632120 566163
rect 0 565519 633000 565883
rect 0 565239 632120 565519
rect 0 564875 633000 565239
rect 0 564595 632120 564875
rect 0 563035 633000 564595
rect 0 562755 632120 563035
rect 0 562483 633000 562755
rect 0 562203 632120 562483
rect 0 561839 633000 562203
rect 0 561559 632120 561839
rect 0 561195 633000 561559
rect 0 560915 632120 561195
rect 0 558711 633000 560915
rect 0 558431 632120 558711
rect 0 558159 633000 558431
rect 0 557879 632120 558159
rect 0 557515 633000 557879
rect 0 557235 632120 557515
rect 0 556871 633000 557235
rect 0 556591 632120 556871
rect 0 555675 633000 556591
rect 0 555395 632120 555675
rect 0 554479 633000 555395
rect 0 554199 632120 554479
rect 0 553835 633000 554199
rect 0 553555 632120 553835
rect 0 553191 633000 553555
rect 0 552911 632120 553191
rect 0 551995 633000 552911
rect 0 551715 632120 551995
rect 0 541485 633000 551715
rect 880 541205 633000 541485
rect 0 540289 633000 541205
rect 880 540009 633000 540289
rect 0 539645 633000 540009
rect 880 539365 633000 539645
rect 0 539001 633000 539365
rect 880 538721 633000 539001
rect 0 537805 633000 538721
rect 880 537525 633000 537805
rect 0 536609 633000 537525
rect 880 536329 633000 536609
rect 0 535965 633000 536329
rect 880 535685 633000 535965
rect 0 535321 633000 535685
rect 880 535041 633000 535321
rect 0 534769 633000 535041
rect 880 534489 633000 534769
rect 0 532285 633000 534489
rect 880 532005 633000 532285
rect 0 531641 633000 532005
rect 880 531361 633000 531641
rect 0 530997 633000 531361
rect 880 530717 633000 530997
rect 0 530445 633000 530717
rect 880 530165 633000 530445
rect 0 528605 633000 530165
rect 880 528325 633000 528605
rect 0 527961 633000 528325
rect 880 527681 633000 527961
rect 0 527317 633000 527681
rect 880 527037 633000 527317
rect 0 520963 633000 527037
rect 0 520683 632120 520963
rect 0 520319 633000 520683
rect 0 520039 632120 520319
rect 0 519675 633000 520039
rect 0 519395 632120 519675
rect 0 517835 633000 519395
rect 0 517555 632120 517835
rect 0 517283 633000 517555
rect 0 517003 632120 517283
rect 0 516639 633000 517003
rect 0 516359 632120 516639
rect 0 515995 633000 516359
rect 0 515715 632120 515995
rect 0 513511 633000 515715
rect 0 513231 632120 513511
rect 0 512959 633000 513231
rect 0 512679 632120 512959
rect 0 512315 633000 512679
rect 0 512035 632120 512315
rect 0 511671 633000 512035
rect 0 511391 632120 511671
rect 0 510475 633000 511391
rect 0 510195 632120 510475
rect 0 509279 633000 510195
rect 0 508999 632120 509279
rect 0 508635 633000 508999
rect 0 508355 632120 508635
rect 0 507991 633000 508355
rect 0 507711 632120 507991
rect 0 506795 633000 507711
rect 0 506515 632120 506795
rect 0 498285 633000 506515
rect 880 498005 633000 498285
rect 0 497089 633000 498005
rect 880 496809 633000 497089
rect 0 496445 633000 496809
rect 880 496165 633000 496445
rect 0 495801 633000 496165
rect 880 495521 633000 495801
rect 0 494605 633000 495521
rect 880 494325 633000 494605
rect 0 493409 633000 494325
rect 880 493129 633000 493409
rect 0 492765 633000 493129
rect 880 492485 633000 492765
rect 0 492121 633000 492485
rect 880 491841 633000 492121
rect 0 491569 633000 491841
rect 880 491289 633000 491569
rect 0 489085 633000 491289
rect 880 488805 633000 489085
rect 0 488441 633000 488805
rect 880 488161 633000 488441
rect 0 487797 633000 488161
rect 880 487517 633000 487797
rect 0 487245 633000 487517
rect 880 486965 633000 487245
rect 0 485405 633000 486965
rect 880 485125 633000 485405
rect 0 484761 633000 485125
rect 880 484481 633000 484761
rect 0 484117 633000 484481
rect 880 483837 633000 484117
rect 0 476601 633000 483837
rect 0 471812 635604 476601
rect 0 466618 633000 471812
rect 0 461829 635604 466618
rect 0 455758 633000 461829
rect -3216 450969 633000 455758
rect 0 445779 633000 450969
rect -3216 440990 633000 445779
rect 0 432600 633000 440990
rect 0 427811 635604 432600
rect 0 427490 633000 427811
rect 0 422869 635204 427490
rect 0 422549 633000 422869
rect 0 417760 635604 422549
rect 0 413640 633000 417760
rect -3216 408851 633000 413640
rect 0 408530 633000 408851
rect -2216 403920 633000 408530
rect 0 403600 633000 403920
rect -3216 398811 633000 403600
rect 0 388409 633000 398811
rect 0 383620 635604 388409
rect 0 378426 633000 383620
rect 0 373637 635604 378426
rect 0 370685 633000 373637
rect 880 370405 633000 370685
rect 0 369489 633000 370405
rect 880 369209 633000 369489
rect 0 368845 633000 369209
rect 880 368565 633000 368845
rect 0 368201 633000 368565
rect 880 367921 633000 368201
rect 0 367005 633000 367921
rect 880 366725 633000 367005
rect 0 365809 633000 366725
rect 880 365529 633000 365809
rect 0 365165 633000 365529
rect 880 364885 633000 365165
rect 0 364521 633000 364885
rect 880 364241 633000 364521
rect 0 363969 633000 364241
rect 880 363689 633000 363969
rect 0 361485 633000 363689
rect 880 361205 633000 361485
rect 0 360841 633000 361205
rect 880 360561 633000 360841
rect 0 360197 633000 360561
rect 880 359917 633000 360197
rect 0 359645 633000 359917
rect 880 359365 633000 359645
rect 0 357805 633000 359365
rect 880 357525 633000 357805
rect 0 357161 633000 357525
rect 880 356881 633000 357161
rect 0 356517 633000 356881
rect 880 356237 633000 356517
rect 0 343763 633000 356237
rect 0 343483 632120 343763
rect 0 343119 633000 343483
rect 0 342839 632120 343119
rect 0 342475 633000 342839
rect 0 342195 632120 342475
rect 0 340635 633000 342195
rect 0 340355 632120 340635
rect 0 340083 633000 340355
rect 0 339803 632120 340083
rect 0 339439 633000 339803
rect 0 339159 632120 339439
rect 0 338795 633000 339159
rect 0 338515 632120 338795
rect 0 336311 633000 338515
rect 0 336031 632120 336311
rect 0 335759 633000 336031
rect 0 335479 632120 335759
rect 0 335115 633000 335479
rect 0 334835 632120 335115
rect 0 334471 633000 334835
rect 0 334191 632120 334471
rect 0 333275 633000 334191
rect 0 332995 632120 333275
rect 0 331435 633000 332995
rect 0 331155 632120 331435
rect 0 330791 633000 331155
rect 0 330511 632120 330791
rect 0 329595 633000 330511
rect 0 329315 632120 329595
rect 0 327485 633000 329315
rect 880 327205 633000 327485
rect 0 326289 633000 327205
rect 880 326009 633000 326289
rect 0 325645 633000 326009
rect 880 325365 633000 325645
rect 0 325001 633000 325365
rect 880 324721 633000 325001
rect 0 323805 633000 324721
rect 880 323525 633000 323805
rect 0 322609 633000 323525
rect 880 322329 633000 322609
rect 0 321965 633000 322329
rect 880 321685 633000 321965
rect 0 321321 633000 321685
rect 880 321041 633000 321321
rect 0 320769 633000 321041
rect 880 320489 633000 320769
rect 0 318285 633000 320489
rect 880 318005 633000 318285
rect 0 317641 633000 318005
rect 880 317361 633000 317641
rect 0 316997 633000 317361
rect 880 316717 633000 316997
rect 0 316445 633000 316717
rect 880 316165 633000 316445
rect 0 314605 633000 316165
rect 880 314325 633000 314605
rect 0 313961 633000 314325
rect 880 313681 633000 313961
rect 0 313317 633000 313681
rect 880 313037 633000 313317
rect 0 298563 633000 313037
rect 0 298283 632120 298563
rect 0 297919 633000 298283
rect 0 297639 632120 297919
rect 0 297275 633000 297639
rect 0 296995 632120 297275
rect 0 295435 633000 296995
rect 0 295155 632120 295435
rect 0 294883 633000 295155
rect 0 294603 632120 294883
rect 0 294239 633000 294603
rect 0 293959 632120 294239
rect 0 293595 633000 293959
rect 0 293315 632120 293595
rect 0 291111 633000 293315
rect 0 290831 632120 291111
rect 0 290559 633000 290831
rect 0 290279 632120 290559
rect 0 289915 633000 290279
rect 0 289635 632120 289915
rect 0 289271 633000 289635
rect 0 288991 632120 289271
rect 0 288075 633000 288991
rect 0 287795 632120 288075
rect 0 286235 633000 287795
rect 0 285955 632120 286235
rect 0 285591 633000 285955
rect 0 285311 632120 285591
rect 0 284395 633000 285311
rect 0 284285 632120 284395
rect 880 284115 632120 284285
rect 880 284005 633000 284115
rect 0 283089 633000 284005
rect 880 282809 633000 283089
rect 0 282445 633000 282809
rect 880 282165 633000 282445
rect 0 281801 633000 282165
rect 880 281521 633000 281801
rect 0 280605 633000 281521
rect 880 280325 633000 280605
rect 0 279409 633000 280325
rect 880 279129 633000 279409
rect 0 278765 633000 279129
rect 880 278485 633000 278765
rect 0 278121 633000 278485
rect 880 277841 633000 278121
rect 0 277569 633000 277841
rect 880 277289 633000 277569
rect 0 275085 633000 277289
rect 880 274805 633000 275085
rect 0 274441 633000 274805
rect 880 274161 633000 274441
rect 0 273797 633000 274161
rect 880 273517 633000 273797
rect 0 273245 633000 273517
rect 880 272965 633000 273245
rect 0 271405 633000 272965
rect 880 271125 633000 271405
rect 0 270761 633000 271125
rect 880 270481 633000 270761
rect 0 270117 633000 270481
rect 880 269837 633000 270117
rect 0 253563 633000 269837
rect 0 253283 632120 253563
rect 0 252919 633000 253283
rect 0 252639 632120 252919
rect 0 252275 633000 252639
rect 0 251995 632120 252275
rect 0 250435 633000 251995
rect 0 250155 632120 250435
rect 0 249883 633000 250155
rect 0 249603 632120 249883
rect 0 249239 633000 249603
rect 0 248959 632120 249239
rect 0 248595 633000 248959
rect 0 248315 632120 248595
rect 0 246111 633000 248315
rect 0 245831 632120 246111
rect 0 245559 633000 245831
rect 0 245279 632120 245559
rect 0 244915 633000 245279
rect 0 244635 632120 244915
rect 0 244271 633000 244635
rect 0 243991 632120 244271
rect 0 243075 633000 243991
rect 0 242795 632120 243075
rect 0 241235 633000 242795
rect 0 241085 632120 241235
rect 880 240955 632120 241085
rect 880 240805 633000 240955
rect 0 240591 633000 240805
rect 0 240311 632120 240591
rect 0 239889 633000 240311
rect 938 239609 633000 239889
rect 0 239395 633000 239609
rect 0 239245 632120 239395
rect 880 239115 632120 239245
rect 880 238965 633000 239115
rect 0 238601 633000 238965
rect 880 238321 633000 238601
rect 0 237405 633000 238321
rect 880 237125 633000 237405
rect 0 236209 633000 237125
rect 880 235929 633000 236209
rect 0 235565 633000 235929
rect 938 235285 633000 235565
rect 0 234921 633000 235285
rect 880 234641 633000 234921
rect 0 234369 633000 234641
rect 880 234089 633000 234369
rect 0 231885 633000 234089
rect 880 231605 633000 231885
rect 0 231241 633000 231605
rect 880 230961 633000 231241
rect 0 230597 633000 230961
rect 880 230317 633000 230597
rect 0 230045 633000 230317
rect 880 229765 633000 230045
rect 0 228205 633000 229765
rect 880 227925 633000 228205
rect 0 227561 633000 227925
rect 880 227281 633000 227561
rect 0 226917 633000 227281
rect 880 226637 633000 226917
rect 0 208563 633000 226637
rect 0 208283 632120 208563
rect 0 207919 633000 208283
rect 0 207639 632120 207919
rect 0 207275 633000 207639
rect 0 206995 632120 207275
rect 0 205435 633000 206995
rect 0 205155 632120 205435
rect 0 204883 633000 205155
rect 0 204603 632120 204883
rect 0 204239 633000 204603
rect 0 203959 632120 204239
rect 0 203595 633000 203959
rect 0 203315 632120 203595
rect 0 201111 633000 203315
rect 0 200831 632120 201111
rect 0 200559 633000 200831
rect 0 200279 632120 200559
rect 0 199915 633000 200279
rect 0 199635 632120 199915
rect 0 199271 633000 199635
rect 0 198991 632120 199271
rect 0 198075 633000 198991
rect 0 197885 632120 198075
rect 880 197795 632120 197885
rect 880 197605 633000 197795
rect 0 196689 633000 197605
rect 880 196409 633000 196689
rect 0 196235 633000 196409
rect 0 196045 632120 196235
rect 880 195955 632120 196045
rect 880 195765 633000 195955
rect 0 195591 633000 195765
rect 0 195311 632120 195591
rect 0 194395 633000 195311
rect 0 194205 632120 194395
rect 880 194115 632120 194205
rect 880 193925 633000 194115
rect 0 193009 633000 193925
rect 880 192729 633000 193009
rect 0 192365 633000 192729
rect 880 192085 633000 192365
rect 0 191721 633000 192085
rect 880 191441 633000 191721
rect 0 191169 633000 191441
rect 880 190889 633000 191169
rect 0 188685 633000 190889
rect 880 188405 633000 188685
rect 0 188041 633000 188405
rect 880 187761 633000 188041
rect 0 187397 633000 187761
rect 880 187117 633000 187397
rect 0 186845 633000 187117
rect 880 186565 633000 186845
rect 0 185005 633000 186565
rect 880 184725 633000 185005
rect 0 184361 633000 184725
rect 880 184081 633000 184361
rect 0 183717 633000 184081
rect 880 183437 633000 183717
rect 0 163363 633000 183437
rect 0 163083 632120 163363
rect 0 162719 633000 163083
rect 0 162439 632120 162719
rect 0 162075 633000 162439
rect 0 161795 632120 162075
rect 0 160235 633000 161795
rect 0 159955 632120 160235
rect 0 159683 633000 159955
rect 0 159403 632120 159683
rect 0 159039 633000 159403
rect 0 158759 632120 159039
rect 0 158395 633000 158759
rect 0 158115 632120 158395
rect 0 155911 633000 158115
rect 0 155631 632120 155911
rect 0 155359 633000 155631
rect 0 155079 632120 155359
rect 0 154715 633000 155079
rect 0 154685 632120 154715
rect 880 154435 632120 154685
rect 880 154405 633000 154435
rect 0 154071 633000 154405
rect 0 153791 632120 154071
rect 0 153489 633000 153791
rect 880 153209 633000 153489
rect 0 152875 633000 153209
rect 0 152845 632120 152875
rect 880 152595 632120 152845
rect 880 152565 633000 152595
rect 0 151035 633000 152565
rect 0 151005 632120 151035
rect 880 150755 632120 151005
rect 880 150725 633000 150755
rect 0 150391 633000 150725
rect 0 150111 632120 150391
rect 0 149809 633000 150111
rect 880 149529 633000 149809
rect 0 149195 633000 149529
rect 0 149165 632120 149195
rect 880 148915 632120 149165
rect 880 148885 633000 148915
rect 0 148521 633000 148885
rect 880 148241 633000 148521
rect 0 147969 633000 148241
rect 880 147689 633000 147969
rect 0 145485 633000 147689
rect 880 145205 633000 145485
rect 0 144841 633000 145205
rect 880 144561 633000 144841
rect 0 144197 633000 144561
rect 880 143917 633000 144197
rect 0 143645 633000 143917
rect 880 143365 633000 143645
rect 0 141805 633000 143365
rect 880 141525 633000 141805
rect 0 141161 633000 141525
rect 880 140881 633000 141161
rect 0 140517 633000 140881
rect 880 140237 633000 140517
rect 0 118363 633000 140237
rect 0 118083 632120 118363
rect 0 117719 633000 118083
rect 0 117439 632120 117719
rect 0 117075 633000 117439
rect 0 116795 632120 117075
rect 0 115235 633000 116795
rect 0 114955 632120 115235
rect 0 114683 633000 114955
rect 0 114403 632120 114683
rect 0 114039 633000 114403
rect 0 113759 632120 114039
rect 0 113395 633000 113759
rect 0 113115 632120 113395
rect 0 110911 633000 113115
rect 0 110631 632120 110911
rect 0 110359 633000 110631
rect 0 110079 632120 110359
rect 0 109715 633000 110079
rect 0 109435 632120 109715
rect 0 109071 633000 109435
rect 0 108791 632120 109071
rect 0 107875 633000 108791
rect 0 107595 632120 107875
rect 0 106035 633000 107595
rect 0 105755 632120 106035
rect 0 105391 633000 105755
rect 0 105111 632120 105391
rect 0 104195 633000 105111
rect 0 103915 632120 104195
rect 0 73163 633000 103915
rect 0 72883 632120 73163
rect 0 72519 633000 72883
rect 0 72239 632120 72519
rect 0 71875 633000 72239
rect 0 71595 632120 71875
rect 0 70035 633000 71595
rect 0 69755 632120 70035
rect 0 69483 633000 69755
rect 0 69203 632120 69483
rect 0 68839 633000 69203
rect 0 68559 632120 68839
rect 0 68195 633000 68559
rect 0 67915 632120 68195
rect 0 65711 633000 67915
rect 0 65431 632120 65711
rect 0 65159 633000 65431
rect 0 64879 632120 65159
rect 0 64515 633000 64879
rect 0 64235 632120 64515
rect 0 63871 633000 64235
rect 0 63591 632120 63871
rect 0 62675 633000 63591
rect 0 62395 632120 62675
rect 0 60835 633000 62395
rect 0 60555 632120 60835
rect 0 60191 633000 60555
rect 0 59911 632120 60191
rect 0 58995 633000 59911
rect 0 58715 632120 58995
rect 0 40840 633000 58715
rect -3216 36051 633000 40840
rect 0 30800 633000 36051
rect -3216 26011 633000 30800
rect 0 0 633000 26011
rect 171700 -6251 175302 -135
rect 193205 -8197 195949 -135
rect 198943 -2938 203749 -22
rect 208994 -2938 213800 -22
<< metal4 >>
rect 2184 2128 3184 950960
rect 3384 2128 4384 950960
rect 4584 2128 5584 950960
rect 5784 2128 6784 950960
rect 6984 2128 7984 950960
rect 8184 2128 9184 950960
rect 9384 2128 10384 950960
rect 10584 2128 11584 950960
rect 11784 2128 12784 950960
rect 12984 2128 13984 950960
rect 14184 2128 14584 950960
rect 14784 2128 15184 950960
rect 24784 919260 26064 950960
rect 26304 919260 27584 950960
rect 44784 919260 46064 950960
rect 46304 919260 47584 950960
rect 51208 919260 52488 950960
rect 52728 919260 54008 950960
rect 64784 919260 66064 950960
rect 66304 919260 67584 950960
rect 84784 919260 86064 950960
rect 86304 919260 87584 950960
rect 104784 919260 106064 950960
rect 106304 919260 107584 950960
rect 111208 919260 112488 950960
rect 112728 919260 114008 950960
rect 124784 919260 126064 950960
rect 126304 919260 127584 950960
rect 144784 919260 146064 950960
rect 146304 919260 147584 950960
rect 164784 919260 166064 950960
rect 166304 919260 167584 950960
rect 184784 919260 186064 950960
rect 186304 919260 187584 950960
rect 191208 919260 192488 950960
rect 192728 919260 194008 950960
rect 204784 919260 206064 950960
rect 206304 919260 207584 950960
rect 224784 919260 226064 950960
rect 226304 919260 227584 950960
rect 231208 919260 232488 950960
rect 232728 919260 234008 950960
rect 244784 919260 246064 950960
rect 246304 919260 247584 950960
rect 264784 919260 266064 950960
rect 266304 919260 267584 950960
rect 284784 919260 286064 950960
rect 286304 919260 287584 950960
rect 291208 919260 292488 950960
rect 292728 919260 294008 950960
rect 295144 919260 296104 950960
rect 304784 919260 306064 950960
rect 306304 919260 307584 950960
rect 324784 919260 326064 950960
rect 326304 919260 327584 950960
rect 344784 919260 346064 950960
rect 346304 919260 347584 950960
rect 351208 919260 352488 950960
rect 352728 919260 354008 950960
rect 364784 919260 366064 950960
rect 366304 919260 367584 950960
rect 384784 919260 386064 950960
rect 386304 919260 387584 950960
rect 404784 919260 406064 950960
rect 406304 919260 407584 950960
rect 411208 919260 412488 950960
rect 412728 919260 414008 950960
rect 424784 919260 426064 950960
rect 426304 919260 427584 950960
rect 444784 919260 446064 950960
rect 446304 919260 447584 950960
rect 464784 919260 466064 950960
rect 466304 919260 467584 950960
rect 471208 919260 472488 950960
rect 472728 919260 474008 950960
rect 484784 919260 486064 950960
rect 486304 919260 487584 950960
rect 504784 919260 506064 950960
rect 506304 919260 507584 950960
rect 524784 919260 526064 950960
rect 526304 919260 527584 950960
rect 530064 928016 531064 938448
rect 531352 928016 532352 938448
rect 544784 919260 546064 920600
rect 546304 919260 547584 920600
rect 551208 919260 552488 950960
rect 552728 919260 554008 950960
rect 564784 919260 566064 950960
rect 566304 919260 567584 950960
rect 584784 919260 586064 950960
rect 586304 919260 587584 950960
rect 604784 919260 606064 950960
rect 606304 919260 607584 950960
rect 24784 2128 26064 197800
rect 26304 2128 27584 197800
rect 44784 124073 46064 197800
rect 46304 124073 47584 197800
rect 64784 124073 66064 197800
rect 66304 124073 67584 197800
rect 84784 124073 86064 197800
rect 86304 124073 87584 197800
rect 44784 2128 46064 34735
rect 46304 2128 47584 34735
rect 64784 2128 66064 34735
rect 66304 2128 67584 34735
rect 84784 2128 86064 34735
rect 86304 2128 87584 34735
rect 104784 2128 106064 197800
rect 106304 2128 107584 197800
rect 111208 2128 112488 197800
rect 112728 2128 114008 197800
rect 124784 124073 126064 197800
rect 126304 124073 127584 197800
rect 144784 124073 146064 197800
rect 146304 124073 147584 197800
rect 164784 124073 166064 197800
rect 166304 124073 167584 197800
rect 170144 124073 171104 197800
rect 171744 124073 172704 197800
rect 124784 2128 126064 34735
rect 126304 2128 127584 34735
rect 130944 2128 131904 34735
rect 132304 2128 133264 33836
rect 144784 2128 146064 34735
rect 146304 2128 147584 33836
rect 164784 2128 166064 34735
rect 166304 2128 167584 34735
rect 180144 2128 181104 197800
rect 181744 2128 182704 197800
rect 184784 2128 186064 197800
rect 186304 2128 187584 197800
rect 191208 2128 192488 197800
rect 204784 6816 206064 197800
rect 206304 6816 207584 197800
rect 208144 6816 209104 37800
rect 209504 6816 210464 37800
rect 224784 2128 226064 197800
rect 226304 2128 227584 197800
rect 231208 2128 232488 197800
rect 232728 2128 234008 197800
rect 244784 2128 246064 197800
rect 246304 2128 247584 197800
rect 255144 2128 256104 197800
rect 256744 2128 257704 197800
rect 264784 2128 266064 197800
rect 266304 2128 267584 197800
rect 275144 2128 276104 197800
rect 276744 2128 277704 197800
rect 284784 2128 286064 197800
rect 286304 2128 287584 197800
rect 291208 2128 292488 197800
rect 292728 2128 294008 197800
rect 295144 2128 296104 197800
rect 296744 2128 297704 197800
rect 304784 2128 306064 197800
rect 306304 2128 307584 197800
rect 324784 56804 326064 197800
rect 326304 56804 327584 197800
rect 324784 2128 326064 35436
rect 326304 2128 327584 35436
rect 344784 2128 346064 197800
rect 346304 2128 347584 197800
rect 351208 2128 352488 197800
rect 352728 2128 354008 197800
rect 364784 114073 366064 197800
rect 366304 114073 367584 197800
rect 368744 114073 369704 197800
rect 370344 114073 371304 197800
rect 371944 114073 372904 197800
rect 373544 114073 374504 197800
rect 376744 114073 377704 197800
rect 378344 114073 379304 197800
rect 379944 114073 380904 197800
rect 381544 114073 382504 197800
rect 384784 114073 386064 197800
rect 386304 114073 387584 197800
rect 404784 114073 406064 197800
rect 406304 114073 407584 197800
rect 364784 2128 366064 24735
rect 366304 2128 367584 24735
rect 384784 2128 386064 24735
rect 386304 2128 387584 24735
rect 404784 2128 406064 24735
rect 406304 2128 407584 23836
rect 424784 2128 426064 197800
rect 426304 2128 427584 197800
rect 444784 2128 446064 197800
rect 446304 2128 447584 197800
rect 464784 2128 466064 197800
rect 466304 2128 467584 197800
rect 471208 2128 472488 197800
rect 472728 2128 474008 197800
rect 484784 2128 486064 197800
rect 486304 2128 487584 197800
rect 504784 2128 506064 197800
rect 506304 2128 507584 197800
rect 524784 2128 526064 197800
rect 526304 2128 527584 197800
rect 544784 146657 546064 197800
rect 546304 146657 547584 197800
rect 564784 147420 566064 197800
rect 566304 146657 567584 197800
rect 584784 146657 586064 197800
rect 586304 146657 587584 197800
rect 604784 146657 606064 197800
rect 606304 146657 607584 197800
rect 544784 2128 546064 38687
rect 546304 2128 547584 38687
rect 564784 2128 566064 38468
rect 566304 2128 567584 38687
rect 584784 2128 586064 38687
rect 586304 2128 587584 38687
rect 604784 2128 606064 38687
rect 606304 2128 607584 38687
rect 617436 2128 617836 950960
rect 618036 2128 618436 950960
rect 618636 2128 619636 950960
rect 619836 2128 620836 950960
rect 621036 2128 622036 950960
rect 622236 2128 623236 950960
rect 623436 2128 624436 950960
rect 624636 2128 625636 950960
rect 625836 2128 626836 950960
rect 627036 2128 628036 950960
rect 628236 2128 629236 950960
rect 629436 2128 630436 950960
<< obsm4 >>
rect 533387 953400 538193 954482
rect 543368 953400 548174 954482
rect 0 951040 633000 953400
rect 0 884840 2104 951040
rect -1858 880051 2104 884840
rect 0 879730 2104 880051
rect -1858 875120 2104 879730
rect 0 874800 2104 875120
rect -1858 870011 2104 874800
rect 0 800358 2104 870011
rect -1858 795569 2104 800358
rect 0 790318 2104 795569
rect -1858 785589 2104 790318
rect 0 455758 2104 785589
rect -1858 450969 2104 455758
rect 0 445718 2104 450969
rect -1858 440989 2104 445718
rect 0 413640 2104 440989
rect -1858 408851 2104 413640
rect 0 408530 2104 408851
rect -1858 403920 2104 408530
rect 0 403600 2104 403920
rect -1858 398811 2104 403600
rect 0 40840 2104 398811
rect -1858 36051 2104 40840
rect 0 30800 2104 36051
rect -1858 26011 2104 30800
rect 0 2048 2104 26011
rect 3264 2048 3304 951040
rect 4464 2048 4504 951040
rect 5664 2048 5704 951040
rect 6864 2048 6904 951040
rect 8064 2048 8104 951040
rect 9264 2048 9304 951040
rect 10464 2048 10504 951040
rect 11664 2048 11704 951040
rect 12864 2048 12904 951040
rect 14064 2048 14104 951040
rect 14664 2048 14704 951040
rect 15264 919180 24704 951040
rect 26144 919180 26224 951040
rect 27664 919180 44704 951040
rect 46144 919180 46224 951040
rect 47664 919180 51128 951040
rect 52568 919180 52648 951040
rect 54088 919180 64704 951040
rect 66144 919180 66224 951040
rect 67664 919180 84704 951040
rect 86144 919180 86224 951040
rect 87664 919180 104704 951040
rect 106144 919180 106224 951040
rect 107664 919180 111128 951040
rect 112568 919180 112648 951040
rect 114088 919180 124704 951040
rect 126144 919180 126224 951040
rect 127664 919180 144704 951040
rect 146144 919180 146224 951040
rect 147664 919180 164704 951040
rect 166144 919180 166224 951040
rect 167664 919180 184704 951040
rect 186144 919180 186224 951040
rect 187664 919180 191128 951040
rect 192568 919180 192648 951040
rect 194088 919180 204704 951040
rect 206144 919180 206224 951040
rect 207664 919180 224704 951040
rect 226144 919180 226224 951040
rect 227664 919180 231128 951040
rect 232568 919180 232648 951040
rect 234088 919180 244704 951040
rect 246144 919180 246224 951040
rect 247664 919180 264704 951040
rect 266144 919180 266224 951040
rect 267664 919180 284704 951040
rect 286144 919180 286224 951040
rect 287664 919180 291128 951040
rect 292568 919180 292648 951040
rect 294088 919180 295064 951040
rect 296184 919180 304704 951040
rect 306144 919180 306224 951040
rect 307664 919180 324704 951040
rect 326144 919180 326224 951040
rect 327664 919180 344704 951040
rect 346144 919180 346224 951040
rect 347664 919180 351128 951040
rect 352568 919180 352648 951040
rect 354088 919180 364704 951040
rect 366144 919180 366224 951040
rect 367664 919180 384704 951040
rect 386144 919180 386224 951040
rect 387664 919180 404704 951040
rect 406144 919180 406224 951040
rect 407664 919180 411128 951040
rect 412568 919180 412648 951040
rect 414088 919180 424704 951040
rect 426144 919180 426224 951040
rect 427664 919180 444704 951040
rect 446144 919180 446224 951040
rect 447664 919180 464704 951040
rect 466144 919180 466224 951040
rect 467664 919180 471128 951040
rect 472568 919180 472648 951040
rect 474088 919180 484704 951040
rect 486144 919180 486224 951040
rect 487664 919180 504704 951040
rect 506144 919180 506224 951040
rect 507664 919180 524704 951040
rect 526144 919180 526224 951040
rect 527664 938528 551128 951040
rect 527664 927936 529984 938528
rect 531144 927936 531272 938528
rect 532432 927936 551128 938528
rect 527664 920680 551128 927936
rect 527664 919180 544704 920680
rect 546144 919180 546224 920680
rect 547664 919180 551128 920680
rect 552568 919180 552648 951040
rect 554088 919180 564704 951040
rect 566144 919180 566224 951040
rect 567664 919180 584704 951040
rect 586144 919180 586224 951040
rect 587664 919180 604704 951040
rect 606144 919180 606224 951040
rect 607664 919180 617356 951040
rect 15264 197880 617356 919180
rect 15264 2048 24704 197880
rect 26144 2048 26224 197880
rect 27664 123993 44704 197880
rect 46144 123993 46224 197880
rect 47664 123993 64704 197880
rect 66144 123993 66224 197880
rect 67664 123993 84704 197880
rect 86144 123993 86224 197880
rect 87664 123993 104704 197880
rect 27664 34815 104704 123993
rect 27664 2048 44704 34815
rect 46144 2048 46224 34815
rect 47664 2048 64704 34815
rect 66144 2048 66224 34815
rect 67664 2048 84704 34815
rect 86144 2048 86224 34815
rect 87664 2048 104704 34815
rect 106144 2048 106224 197880
rect 107664 2048 111128 197880
rect 112568 2048 112648 197880
rect 114088 123993 124704 197880
rect 126144 123993 126224 197880
rect 127664 123993 144704 197880
rect 146144 123993 146224 197880
rect 147664 123993 164704 197880
rect 166144 123993 166224 197880
rect 167664 123993 170064 197880
rect 171184 123993 171664 197880
rect 172784 123993 180064 197880
rect 114088 34815 180064 123993
rect 114088 2048 124704 34815
rect 126144 2048 126224 34815
rect 127664 2048 130864 34815
rect 131984 33916 144704 34815
rect 131984 2048 132224 33916
rect 133344 2048 144704 33916
rect 146144 33916 164704 34815
rect 146144 2048 146224 33916
rect 147664 2048 164704 33916
rect 166144 2048 166224 34815
rect 167664 2048 180064 34815
rect 181184 2048 181664 197880
rect 182784 2048 184704 197880
rect 186144 2048 186224 197880
rect 187664 2048 191128 197880
rect 192568 6736 204704 197880
rect 206144 6736 206224 197880
rect 207664 37880 224704 197880
rect 207664 6736 208064 37880
rect 209184 6736 209424 37880
rect 210544 6736 224704 37880
rect 192568 2048 224704 6736
rect 226144 2048 226224 197880
rect 227664 2048 231128 197880
rect 232568 2048 232648 197880
rect 234088 2048 244704 197880
rect 246144 2048 246224 197880
rect 247664 2048 255064 197880
rect 256184 2048 256664 197880
rect 257784 2048 264704 197880
rect 266144 2048 266224 197880
rect 267664 2048 275064 197880
rect 276184 2048 276664 197880
rect 277784 2048 284704 197880
rect 286144 2048 286224 197880
rect 287664 2048 291128 197880
rect 292568 2048 292648 197880
rect 294088 2048 295064 197880
rect 296184 2048 296664 197880
rect 297784 2048 304704 197880
rect 306144 2048 306224 197880
rect 307664 56724 324704 197880
rect 326144 56724 326224 197880
rect 327664 56724 344704 197880
rect 307664 35516 344704 56724
rect 307664 2048 324704 35516
rect 326144 2048 326224 35516
rect 327664 2048 344704 35516
rect 346144 2048 346224 197880
rect 347664 2048 351128 197880
rect 352568 2048 352648 197880
rect 354088 113993 364704 197880
rect 366144 113993 366224 197880
rect 367664 113993 368664 197880
rect 369784 113993 370264 197880
rect 371384 113993 371864 197880
rect 372984 113993 373464 197880
rect 374584 113993 376664 197880
rect 377784 113993 378264 197880
rect 379384 113993 379864 197880
rect 380984 113993 381464 197880
rect 382584 113993 384704 197880
rect 386144 113993 386224 197880
rect 387664 113993 404704 197880
rect 406144 113993 406224 197880
rect 407664 113993 424704 197880
rect 354088 24815 424704 113993
rect 354088 2048 364704 24815
rect 366144 2048 366224 24815
rect 367664 2048 384704 24815
rect 386144 2048 386224 24815
rect 387664 2048 404704 24815
rect 406144 23916 424704 24815
rect 406144 2048 406224 23916
rect 407664 2048 424704 23916
rect 426144 2048 426224 197880
rect 427664 2048 444704 197880
rect 446144 2048 446224 197880
rect 447664 2048 464704 197880
rect 466144 2048 466224 197880
rect 467664 2048 471128 197880
rect 472568 2048 472648 197880
rect 474088 2048 484704 197880
rect 486144 2048 486224 197880
rect 487664 2048 504704 197880
rect 506144 2048 506224 197880
rect 507664 2048 524704 197880
rect 526144 2048 526224 197880
rect 527664 146577 544704 197880
rect 546144 146577 546224 197880
rect 547664 147340 564704 197880
rect 566144 147340 566224 197880
rect 547664 146577 566224 147340
rect 567664 146577 584704 197880
rect 586144 146577 586224 197880
rect 587664 146577 604704 197880
rect 606144 146577 606224 197880
rect 607664 146577 617356 197880
rect 527664 38767 617356 146577
rect 527664 2048 544704 38767
rect 546144 2048 546224 38767
rect 547664 38548 566224 38767
rect 547664 2048 564704 38548
rect 566144 2048 566224 38548
rect 567664 2048 584704 38767
rect 586144 2048 586224 38767
rect 587664 2048 604704 38767
rect 606144 2048 606224 38767
rect 607664 2048 617356 38767
rect 617916 2048 617956 951040
rect 618516 2048 618556 951040
rect 619716 2048 619756 951040
rect 620916 2048 620956 951040
rect 622116 2048 622156 951040
rect 623316 2048 623356 951040
rect 624516 2048 624556 951040
rect 625716 2048 625756 951040
rect 626916 2048 626956 951040
rect 628116 2048 628156 951040
rect 629316 2048 629356 951040
rect 630516 880400 633000 951040
rect 630516 875611 634246 880400
rect 630516 875290 633000 875611
rect 630516 870669 634246 875290
rect 630516 870349 633000 870669
rect 630516 865560 634246 870349
rect 630516 791201 633000 865560
rect 630516 786412 634246 791201
rect 630516 781218 633000 786412
rect 630516 776429 634246 781218
rect 630516 476601 633000 776429
rect 630516 471812 634246 476601
rect 630516 466618 633000 471812
rect 630516 461829 634246 466618
rect 630516 432600 633000 461829
rect 630516 427811 634246 432600
rect 630516 427490 633000 427811
rect 630516 422869 634246 427490
rect 630516 422549 633000 422869
rect 630516 417760 634246 422549
rect 630516 388409 633000 417760
rect 630516 383620 634246 388409
rect 630516 378426 633000 383620
rect 630516 373637 634246 378426
rect 630516 2048 633000 373637
rect 0 0 633000 2048
rect 171700 -1937 175302 0
rect 193205 -1937 195949 0
rect 198943 -1824 203749 0
rect 208994 -1824 213800 0
rect 193308 -8126 195772 -7342
<< metal5 >>
rect 1976 947012 630984 949612
rect 1976 944092 630984 946692
rect 1976 941172 630984 943772
rect 1976 938252 630984 940852
rect 1976 935332 630984 937932
rect 1976 932412 630984 935012
rect 1976 929492 630984 932092
rect 1976 926572 630984 929172
rect 1976 923652 630984 926252
rect 1976 920732 630984 923332
rect 524784 919540 567584 919860
rect 1976 903496 15184 904776
rect 1976 901736 15184 903016
rect 617436 903496 630984 904776
rect 617436 901736 630984 903016
rect 1976 855496 15184 856776
rect 1976 853736 15184 855016
rect 617436 855496 630984 856776
rect 617436 853736 630984 855016
rect 1976 831496 15184 832776
rect 1976 829736 15184 831016
rect 617436 831496 630984 832776
rect 617436 829736 630984 831016
rect 1976 807496 15184 808776
rect 1976 805736 15184 807016
rect 617436 807496 630984 808776
rect 617436 805736 630984 807016
rect 1976 783496 15184 784776
rect 1976 781736 15184 783016
rect 1976 759496 15184 760776
rect 1976 757736 15184 759016
rect 617436 759496 630984 760776
rect 617436 757736 630984 759016
rect 1976 735496 15184 736776
rect 1976 733736 15184 735016
rect 617436 735496 630984 736776
rect 617436 733736 630984 735016
rect 1976 711496 15184 712776
rect 1976 709736 15184 711016
rect 617436 711496 630984 712776
rect 617436 709736 630984 711016
rect 1976 687496 15184 688776
rect 1976 685736 15184 687016
rect 617436 687496 630984 688776
rect 617436 685736 630984 687016
rect 1976 663496 15184 664776
rect 1976 661736 15184 663016
rect 617436 663496 630984 664776
rect 617436 661736 630984 663016
rect 1976 639496 15184 640776
rect 1976 637736 15184 639016
rect 617436 639496 630984 640776
rect 617436 637736 630984 639016
rect 1976 615496 15184 616776
rect 1976 613736 15184 615016
rect 617436 615496 630984 616776
rect 617436 613736 630984 615016
rect 1976 591496 15184 592776
rect 1976 589736 15184 591016
rect 617436 591496 630984 592776
rect 617436 589736 630984 591016
rect 1976 567496 15184 568776
rect 1976 565736 15184 567016
rect 617436 567496 630984 568776
rect 617436 565736 630984 567016
rect 1976 543496 15184 544776
rect 1976 541736 15184 543016
rect 617436 543496 630984 544776
rect 617436 541736 630984 543016
rect 1976 519496 15184 520776
rect 1976 517736 15184 519016
rect 617436 519496 630984 520776
rect 617436 517736 630984 519016
rect 1976 495496 15184 496776
rect 1976 493736 15184 495016
rect 617436 495496 630984 496776
rect 617436 493736 630984 495016
rect 1976 471496 15184 472776
rect 1976 469736 15184 471016
rect 617436 447496 630984 448776
rect 617436 445736 630984 447016
rect 1976 423496 15184 424776
rect 1976 421736 15184 423016
rect 617436 399496 630984 400776
rect 617436 397736 630984 399016
rect 1976 375496 15184 376776
rect 1976 373736 15184 375016
rect 1976 351496 15184 352776
rect 1976 349736 15184 351016
rect 617436 351496 630984 352776
rect 617436 349736 630984 351016
rect 1976 327496 15184 328776
rect 1976 325736 15184 327016
rect 617436 327496 630984 328776
rect 617436 325736 630984 327016
rect 1976 303496 15184 304776
rect 1976 301736 15184 303016
rect 617436 303496 630984 304776
rect 617436 301736 630984 303016
rect 1976 279496 15184 280776
rect 1976 277736 15184 279016
rect 617436 279496 630984 280776
rect 617436 277736 630984 279016
rect 1976 255496 15184 256776
rect 1976 253736 15184 255016
rect 617436 255496 630984 256776
rect 617436 253736 630984 255016
rect 1976 231496 15184 232776
rect 1976 229736 15184 231016
rect 617436 231496 630984 232776
rect 617436 229736 630984 231016
rect 1976 207496 15184 208776
rect 1976 205736 15184 207016
rect 617436 207496 630984 208776
rect 617436 205736 630984 207016
rect 1976 193960 630984 196840
rect 1976 190600 630984 193480
rect 1976 183496 630984 184776
rect 1976 181736 630984 183016
rect 1976 174296 630984 175256
rect 1976 172696 630984 173656
rect 1976 171096 630984 172056
rect 1976 169496 630984 170456
rect 1976 167896 630984 168856
rect 1976 166296 630984 167256
rect 1976 164696 630984 165656
rect 1976 163096 630984 164056
rect 1976 159496 630984 160776
rect 1976 157736 630984 159016
rect 1976 147896 630984 150776
rect 1976 144536 630984 147416
rect 1976 135496 630984 136776
rect 1976 133736 630984 135016
rect 1976 123896 630984 126776
rect 1976 120536 630984 123416
rect 1976 111496 630984 112776
rect 1976 109736 630984 111016
rect 1976 99896 630984 102776
rect 1976 96536 630984 99416
rect 1976 87496 630984 88776
rect 1976 85736 630984 87016
rect 1976 75896 630984 78776
rect 1976 72536 630984 75416
rect 1976 63496 630984 64776
rect 1976 61736 630984 63016
rect 1976 51896 630984 54776
rect 1976 48536 630984 51416
rect 5600 39496 630984 40776
rect 5600 37736 630984 39016
rect 130000 33276 216423 34276
rect 130000 31876 216423 32876
rect 130000 30476 216423 31476
rect 130000 29076 216423 30076
rect 1976 23056 630984 25056
rect 1976 20736 630984 22736
rect 1976 18416 630984 20416
rect 1976 16096 630984 18096
rect 1976 13776 630984 15776
rect 1976 11456 630984 13456
rect 1976 9136 630984 11136
rect 1976 6816 630984 8816
rect 1976 4496 630984 6496
rect 1976 2176 630984 4176
<< obsm5 >>
rect 0 905096 633000 918990
rect 0 901416 1656 905096
rect 15504 901416 617116 905096
rect 631304 901416 633000 905096
rect 0 884840 633000 901416
rect -1858 880400 633000 884840
rect -1858 880050 634246 880400
rect 0 879730 634246 880050
rect -1858 875610 634246 879730
rect -1858 875290 633000 875610
rect -1858 875120 634246 875290
rect 0 874800 634246 875120
rect -1858 870669 634246 874800
rect -1858 870349 633000 870669
rect -1858 870010 634246 870349
rect 0 865559 634246 870010
rect 0 857096 633000 865559
rect 0 853416 1656 857096
rect 15504 853416 617116 857096
rect 631304 853416 633000 857096
rect 0 833096 633000 853416
rect 0 829416 1656 833096
rect 15504 829416 617116 833096
rect 631304 829416 633000 833096
rect 0 809096 633000 829416
rect 0 805416 1656 809096
rect 15504 805416 617116 809096
rect 631304 805416 633000 809096
rect 0 800358 633000 805416
rect -1858 795568 633000 800358
rect 0 791201 633000 795568
rect 0 790379 634246 791201
rect -1858 786411 634246 790379
rect -1858 785589 633000 786411
rect 0 785096 633000 785589
rect 0 781416 1656 785096
rect 15504 781416 633000 785096
rect 0 781218 633000 781416
rect 0 776428 634246 781218
rect 0 761096 633000 776428
rect 0 757416 1656 761096
rect 15504 757416 617116 761096
rect 631304 757416 633000 761096
rect 0 737096 633000 757416
rect 0 733416 1656 737096
rect 15504 733416 617116 737096
rect 631304 733416 633000 737096
rect 0 713096 633000 733416
rect 0 709416 1656 713096
rect 15504 709416 617116 713096
rect 631304 709416 633000 713096
rect 0 689096 633000 709416
rect 0 685416 1656 689096
rect 15504 685416 617116 689096
rect 631304 685416 633000 689096
rect 0 665096 633000 685416
rect 0 661416 1656 665096
rect 15504 661416 617116 665096
rect 631304 661416 633000 665096
rect 0 641096 633000 661416
rect 0 637416 1656 641096
rect 15504 637416 617116 641096
rect 631304 637416 633000 641096
rect 0 617096 633000 637416
rect 0 613416 1656 617096
rect 15504 613416 617116 617096
rect 631304 613416 633000 617096
rect 0 593096 633000 613416
rect 0 589416 1656 593096
rect 15504 589416 617116 593096
rect 631304 589416 633000 593096
rect 0 569096 633000 589416
rect 0 565416 1656 569096
rect 15504 565416 617116 569096
rect 631304 565416 633000 569096
rect 0 545096 633000 565416
rect 0 541416 1656 545096
rect 15504 541416 617116 545096
rect 631304 541416 633000 545096
rect 0 521096 633000 541416
rect 0 517416 1656 521096
rect 15504 517416 617116 521096
rect 631304 517416 633000 521096
rect 0 497096 633000 517416
rect 0 493416 1656 497096
rect 15504 493416 617116 497096
rect 631304 493416 633000 497096
rect 0 476601 633000 493416
rect 0 473096 634246 476601
rect 0 469416 1656 473096
rect 15504 471811 634246 473096
rect 15504 469416 633000 471811
rect 0 466618 633000 469416
rect 0 461828 634246 466618
rect 0 455758 633000 461828
rect -1858 450968 633000 455758
rect 0 449096 633000 450968
rect 0 445779 617116 449096
rect -1858 445416 617116 445779
rect 631304 445416 633000 449096
rect -1858 440989 633000 445416
rect 0 432600 633000 440989
rect 0 427810 634246 432600
rect 0 427490 633000 427810
rect 0 425096 634246 427490
rect 0 421416 1656 425096
rect 15504 422869 634246 425096
rect 15504 422549 633000 422869
rect 15504 421416 634246 422549
rect 0 417759 634246 421416
rect 0 413640 633000 417759
rect -1858 408850 633000 413640
rect 0 408530 633000 408850
rect -1858 403920 633000 408530
rect 0 403600 633000 403920
rect -1858 401096 633000 403600
rect -1858 398810 617116 401096
rect 0 397416 617116 398810
rect 631304 397416 633000 401096
rect 0 388409 633000 397416
rect 0 383619 634246 388409
rect 0 378426 633000 383619
rect 0 377096 634246 378426
rect 0 373416 1656 377096
rect 15504 373636 634246 377096
rect 15504 373416 633000 373636
rect 0 353096 633000 373416
rect 0 349416 1656 353096
rect 15504 349416 617116 353096
rect 631304 349416 633000 353096
rect 0 329096 633000 349416
rect 0 325416 1656 329096
rect 15504 325416 617116 329096
rect 631304 325416 633000 329096
rect 0 305096 633000 325416
rect 0 301416 1656 305096
rect 15504 301416 617116 305096
rect 631304 301416 633000 305096
rect 0 281096 633000 301416
rect 0 277416 1656 281096
rect 15504 277416 617116 281096
rect 631304 277416 633000 281096
rect 0 257096 633000 277416
rect 0 253416 1656 257096
rect 15504 253416 617116 257096
rect 631304 253416 633000 257096
rect 0 233096 633000 253416
rect 0 229416 1656 233096
rect 15504 229416 617116 233096
rect 631304 229416 633000 233096
rect 0 209096 633000 229416
rect 0 205416 1656 209096
rect 15504 205416 617116 209096
rect 631304 205416 633000 209096
rect 0 197160 633000 205416
rect 0 190280 1656 197160
rect 631304 190280 633000 197160
rect 0 185096 633000 190280
rect 0 181416 1656 185096
rect 631304 181416 633000 185096
rect 0 175576 633000 181416
rect 0 162776 1656 175576
rect 631304 162776 633000 175576
rect 0 161096 633000 162776
rect 0 157416 1656 161096
rect 631304 157416 633000 161096
rect 0 151096 633000 157416
rect 0 144216 1656 151096
rect 631304 144216 633000 151096
rect 0 137096 633000 144216
rect 0 133416 1656 137096
rect 631304 133416 633000 137096
rect 0 127096 633000 133416
rect 0 120216 1656 127096
rect 631304 120216 633000 127096
rect 0 113096 633000 120216
rect 0 109416 1656 113096
rect 631304 109416 633000 113096
rect 0 103096 633000 109416
rect 0 96216 1656 103096
rect 631304 96216 633000 103096
rect 0 89096 633000 96216
rect 0 85416 1656 89096
rect 631304 85416 633000 89096
rect 0 79096 633000 85416
rect 0 72216 1656 79096
rect 631304 72216 633000 79096
rect 0 65096 633000 72216
rect 0 61416 1656 65096
rect 631304 61416 633000 65096
rect 0 55096 633000 61416
rect 0 48216 1656 55096
rect 631304 48216 633000 55096
rect 0 41096 633000 48216
rect 0 40840 5280 41096
rect -1858 37416 5280 40840
rect 631304 37416 633000 41096
rect -1858 36050 633000 37416
rect 0 34596 633000 36050
rect 0 30800 129680 34596
rect -1858 28756 129680 30800
rect 216743 28756 633000 34596
rect -1858 26010 633000 28756
<< labels >>
rlabel metal2 s 145027 -400 145083 800 6 clock_core
port 1 nsew signal input
rlabel metal2 s 319467 -400 319523 800 6 flash_clk_frame
port 2 nsew signal output
rlabel metal2 s 322595 -400 322651 800 6 flash_clk_oeb
port 3 nsew signal output
rlabel metal2 s 264667 -400 264723 800 6 flash_csb_frame
port 4 nsew signal output
rlabel metal2 s 267795 -400 267851 800 6 flash_csb_oeb
port 5 nsew signal output
rlabel metal2 s 363227 -400 363283 800 6 flash_io0_di
port 6 nsew signal input
rlabel metal2 s 374267 -400 374323 800 6 flash_io0_do
port 7 nsew signal output
rlabel metal2 s 369943 -400 369999 800 6 flash_io0_ieb
port 8 nsew signal output
rlabel metal2 s 377395 -400 377451 800 6 flash_io0_oeb
port 9 nsew signal output
rlabel metal2 s 418027 -400 418083 800 6 flash_io1_di
port 10 nsew signal input
rlabel metal2 s 429067 -400 429123 800 6 flash_io1_do
port 11 nsew signal output
rlabel metal2 s 424743 -400 424799 800 6 flash_io1_ieb
port 12 nsew signal output
rlabel metal2 s 432195 -400 432251 800 6 flash_io1_oeb
port 13 nsew signal output
rlabel metal2 s 472827 -400 472883 800 6 gpio_in_core
port 14 nsew signal input
rlabel metal2 s 479543 -400 479599 800 6 gpio_inenb_core
port 15 nsew signal output
rlabel metal2 s 478347 -400 478403 800 6 gpio_mode0_core
port 16 nsew signal output
rlabel metal2 s 482671 -400 482727 800 6 gpio_mode1_core
port 17 nsew signal output
rlabel metal2 s 483867 -400 483923 800 6 gpio_out_core
port 18 nsew signal output
rlabel metal2 s 486995 -400 487051 800 6 gpio_outenb_core
port 19 nsew signal output
rlabel metal3 s 632200 509079 633437 509199 6 mprj_analog_io[0]
port 20 nsew signal bidirectional
rlabel metal2 s 443033 952600 443089 953787 6 mprj_analog_io[10]
port 21 nsew signal bidirectional
rlabel metal2 s 354033 952600 354089 953787 6 mprj_analog_io[11]
port 22 nsew signal bidirectional
rlabel metal2 s 252233 952600 252289 953787 6 mprj_analog_io[12]
port 23 nsew signal bidirectional
rlabel metal2 s 200633 952600 200689 953787 6 mprj_analog_io[13]
port 24 nsew signal bidirectional
rlabel metal2 s 149233 952600 149289 953787 6 mprj_analog_io[14]
port 25 nsew signal bidirectional
rlabel metal2 s 97833 952600 97889 953787 6 mprj_analog_io[15]
port 26 nsew signal bidirectional
rlabel metal2 s 46433 952600 46489 953787 6 mprj_analog_io[16]
port 27 nsew signal bidirectional
rlabel metal3 s -437 924601 800 924721 6 mprj_analog_io[17]
port 28 nsew signal bidirectional
rlabel metal3 s -437 754801 800 754921 6 mprj_analog_io[18]
port 29 nsew signal bidirectional
rlabel metal3 s -437 711601 800 711721 6 mprj_analog_io[19]
port 30 nsew signal bidirectional
rlabel metal3 s 632200 554279 633437 554399 6 mprj_analog_io[1]
port 31 nsew signal bidirectional
rlabel metal3 s -437 668401 800 668521 6 mprj_analog_io[20]
port 32 nsew signal bidirectional
rlabel metal3 s -437 625201 800 625321 6 mprj_analog_io[21]
port 33 nsew signal bidirectional
rlabel metal3 s -437 582001 800 582121 6 mprj_analog_io[22]
port 34 nsew signal bidirectional
rlabel metal3 s -437 538801 800 538921 6 mprj_analog_io[23]
port 35 nsew signal bidirectional
rlabel metal3 s -437 495601 800 495721 6 mprj_analog_io[24]
port 36 nsew signal bidirectional
rlabel metal3 s -437 368001 800 368121 6 mprj_analog_io[25]
port 37 nsew signal bidirectional
rlabel metal3 s -437 324801 800 324921 6 mprj_analog_io[26]
port 38 nsew signal bidirectional
rlabel metal3 s -437 281601 800 281721 6 mprj_analog_io[27]
port 39 nsew signal bidirectional
rlabel metal3 s -437 238401 800 238521 6 mprj_analog_io[28]
port 40 nsew signal bidirectional
rlabel metal3 s 632200 599279 633437 599399 6 mprj_analog_io[2]
port 41 nsew signal bidirectional
rlabel metal3 s 632200 644479 633437 644599 6 mprj_analog_io[3]
port 42 nsew signal bidirectional
rlabel metal3 s 632200 689479 633437 689599 6 mprj_analog_io[4]
port 43 nsew signal bidirectional
rlabel metal3 s 632200 734479 633437 734599 6 mprj_analog_io[5]
port 44 nsew signal bidirectional
rlabel metal3 s 632200 823679 633437 823799 6 mprj_analog_io[6]
port 45 nsew signal bidirectional
rlabel metal3 s 632200 912879 633437 912999 6 mprj_analog_io[7]
port 46 nsew signal bidirectional
rlabel metal2 s 596233 952600 596289 953787 6 mprj_analog_io[8]
port 47 nsew signal bidirectional
rlabel metal2 s 494433 952600 494489 953787 6 mprj_analog_io[9]
port 48 nsew signal bidirectional
rlabel metal3 s 632200 63671 633437 63791 6 mprj_io_analog_en[0]
port 49 nsew signal output
rlabel metal3 s 632200 646871 633437 646991 6 mprj_io_analog_en[10]
port 50 nsew signal output
rlabel metal3 s 632200 691871 633437 691991 6 mprj_io_analog_en[11]
port 51 nsew signal output
rlabel metal3 s 632200 736871 633437 736991 6 mprj_io_analog_en[12]
port 52 nsew signal output
rlabel metal3 s 632200 826071 633437 826191 6 mprj_io_analog_en[13]
port 53 nsew signal output
rlabel metal3 s 632200 915271 633437 915391 6 mprj_io_analog_en[14]
port 54 nsew signal output
rlabel metal2 s 593841 952600 593897 953787 6 mprj_io_analog_en[15]
port 55 nsew signal output
rlabel metal2 s 492041 952600 492097 953787 6 mprj_io_analog_en[16]
port 56 nsew signal output
rlabel metal2 s 440641 952600 440697 953787 6 mprj_io_analog_en[17]
port 57 nsew signal output
rlabel metal2 s 351641 952600 351697 953787 6 mprj_io_analog_en[18]
port 58 nsew signal output
rlabel metal2 s 249841 952600 249897 953787 6 mprj_io_analog_en[19]
port 59 nsew signal output
rlabel metal3 s 632200 108871 633437 108991 6 mprj_io_analog_en[1]
port 60 nsew signal output
rlabel metal2 s 198241 952600 198297 953787 6 mprj_io_analog_en[20]
port 61 nsew signal output
rlabel metal2 s 146841 952600 146897 953787 6 mprj_io_analog_en[21]
port 62 nsew signal output
rlabel metal2 s 95441 952600 95497 953787 6 mprj_io_analog_en[22]
port 63 nsew signal output
rlabel metal2 s 44041 952600 44097 953787 6 mprj_io_analog_en[23]
port 64 nsew signal output
rlabel metal3 s -437 922209 800 922329 6 mprj_io_analog_en[24]
port 65 nsew signal output
rlabel metal3 s -437 752409 800 752529 6 mprj_io_analog_en[25]
port 66 nsew signal output
rlabel metal3 s -437 709209 800 709329 6 mprj_io_analog_en[26]
port 67 nsew signal output
rlabel metal3 s -437 666009 800 666129 6 mprj_io_analog_en[27]
port 68 nsew signal output
rlabel metal3 s -437 622809 858 622929 6 mprj_io_analog_en[28]
port 69 nsew signal output
rlabel metal3 s -437 579609 800 579729 6 mprj_io_analog_en[29]
port 70 nsew signal output
rlabel metal3 s 632200 153871 633437 153991 6 mprj_io_analog_en[2]
port 71 nsew signal output
rlabel metal3 s -437 536409 800 536529 6 mprj_io_analog_en[30]
port 72 nsew signal output
rlabel metal3 s -437 493209 800 493329 6 mprj_io_analog_en[31]
port 73 nsew signal output
rlabel metal3 s -437 365609 800 365729 6 mprj_io_analog_en[32]
port 74 nsew signal output
rlabel metal3 s -437 322409 800 322529 6 mprj_io_analog_en[33]
port 75 nsew signal output
rlabel metal3 s -437 279209 800 279329 6 mprj_io_analog_en[34]
port 76 nsew signal output
rlabel metal3 s -437 236009 800 236129 6 mprj_io_analog_en[35]
port 77 nsew signal output
rlabel metal3 s -437 192809 800 192929 6 mprj_io_analog_en[36]
port 78 nsew signal output
rlabel metal3 s -437 149609 800 149729 6 mprj_io_analog_en[37]
port 79 nsew signal output
rlabel metal3 s 632200 199071 633437 199191 6 mprj_io_analog_en[3]
port 80 nsew signal output
rlabel metal3 s 632200 244071 633437 244191 6 mprj_io_analog_en[4]
port 81 nsew signal output
rlabel metal3 s 632200 289071 633437 289191 6 mprj_io_analog_en[5]
port 82 nsew signal output
rlabel metal3 s 632200 334271 633437 334391 6 mprj_io_analog_en[6]
port 83 nsew signal output
rlabel metal3 s 632200 511471 633437 511591 6 mprj_io_analog_en[7]
port 84 nsew signal output
rlabel metal3 s 632200 556671 633437 556791 6 mprj_io_analog_en[8]
port 85 nsew signal output
rlabel metal3 s 632200 601671 633437 601791 6 mprj_io_analog_en[9]
port 86 nsew signal output
rlabel metal3 s 632200 64959 633437 65079 6 mprj_io_analog_pol[0]
port 87 nsew signal output
rlabel metal3 s 632200 648159 633437 648279 6 mprj_io_analog_pol[10]
port 88 nsew signal output
rlabel metal3 s 632200 693159 633437 693279 6 mprj_io_analog_pol[11]
port 89 nsew signal output
rlabel metal3 s 632200 738159 633437 738279 6 mprj_io_analog_pol[12]
port 90 nsew signal output
rlabel metal3 s 632200 827359 633437 827479 6 mprj_io_analog_pol[13]
port 91 nsew signal output
rlabel metal3 s 632200 916559 633437 916679 6 mprj_io_analog_pol[14]
port 92 nsew signal output
rlabel metal2 s 592553 952600 592609 953787 6 mprj_io_analog_pol[15]
port 93 nsew signal output
rlabel metal2 s 490753 952600 490809 953787 6 mprj_io_analog_pol[16]
port 94 nsew signal output
rlabel metal2 s 439353 952600 439409 953787 6 mprj_io_analog_pol[17]
port 95 nsew signal output
rlabel metal2 s 350353 952600 350409 953787 6 mprj_io_analog_pol[18]
port 96 nsew signal output
rlabel metal2 s 248553 952600 248609 953787 6 mprj_io_analog_pol[19]
port 97 nsew signal output
rlabel metal3 s 632200 110159 633437 110279 6 mprj_io_analog_pol[1]
port 98 nsew signal output
rlabel metal2 s 196953 952600 197009 953787 6 mprj_io_analog_pol[20]
port 99 nsew signal output
rlabel metal2 s 145553 952600 145609 953787 6 mprj_io_analog_pol[21]
port 100 nsew signal output
rlabel metal2 s 94153 952600 94209 953787 6 mprj_io_analog_pol[22]
port 101 nsew signal output
rlabel metal2 s 42753 952600 42809 953787 6 mprj_io_analog_pol[23]
port 102 nsew signal output
rlabel metal3 s -437 920921 800 921041 6 mprj_io_analog_pol[24]
port 103 nsew signal output
rlabel metal3 s -437 751121 800 751241 6 mprj_io_analog_pol[25]
port 104 nsew signal output
rlabel metal3 s -437 707921 800 708041 6 mprj_io_analog_pol[26]
port 105 nsew signal output
rlabel metal3 s -437 664721 800 664841 6 mprj_io_analog_pol[27]
port 106 nsew signal output
rlabel metal3 s -437 621521 800 621641 6 mprj_io_analog_pol[28]
port 107 nsew signal output
rlabel metal3 s -437 578321 800 578441 6 mprj_io_analog_pol[29]
port 108 nsew signal output
rlabel metal3 s 632200 155159 633437 155279 6 mprj_io_analog_pol[2]
port 109 nsew signal output
rlabel metal3 s -437 535121 800 535241 6 mprj_io_analog_pol[30]
port 110 nsew signal output
rlabel metal3 s -437 491921 800 492041 6 mprj_io_analog_pol[31]
port 111 nsew signal output
rlabel metal3 s -437 364321 800 364441 6 mprj_io_analog_pol[32]
port 112 nsew signal output
rlabel metal3 s -437 321121 800 321241 6 mprj_io_analog_pol[33]
port 113 nsew signal output
rlabel metal3 s -437 277921 800 278041 6 mprj_io_analog_pol[34]
port 114 nsew signal output
rlabel metal3 s -437 234721 800 234841 6 mprj_io_analog_pol[35]
port 115 nsew signal output
rlabel metal3 s -437 191521 800 191641 6 mprj_io_analog_pol[36]
port 116 nsew signal output
rlabel metal3 s -437 148321 800 148441 6 mprj_io_analog_pol[37]
port 117 nsew signal output
rlabel metal3 s 632200 200359 633437 200479 6 mprj_io_analog_pol[3]
port 118 nsew signal output
rlabel metal3 s 632200 245359 633437 245479 6 mprj_io_analog_pol[4]
port 119 nsew signal output
rlabel metal3 s 632200 290359 633437 290479 6 mprj_io_analog_pol[5]
port 120 nsew signal output
rlabel metal3 s 632200 335559 633437 335679 6 mprj_io_analog_pol[6]
port 121 nsew signal output
rlabel metal3 s 632200 512759 633437 512879 6 mprj_io_analog_pol[7]
port 122 nsew signal output
rlabel metal3 s 632200 557959 633437 558079 6 mprj_io_analog_pol[8]
port 123 nsew signal output
rlabel metal3 s 632200 602959 633437 603079 6 mprj_io_analog_pol[9]
port 124 nsew signal output
rlabel metal3 s 632200 67995 633437 68115 6 mprj_io_analog_sel[0]
port 125 nsew signal output
rlabel metal3 s 632200 651195 633437 651315 6 mprj_io_analog_sel[10]
port 126 nsew signal output
rlabel metal3 s 632200 696195 633437 696315 6 mprj_io_analog_sel[11]
port 127 nsew signal output
rlabel metal3 s 632200 741195 633437 741315 6 mprj_io_analog_sel[12]
port 128 nsew signal output
rlabel metal3 s 632200 830395 633437 830515 6 mprj_io_analog_sel[13]
port 129 nsew signal output
rlabel metal3 s 632200 919595 633437 919715 6 mprj_io_analog_sel[14]
port 130 nsew signal output
rlabel metal2 s 589517 952600 589573 953787 6 mprj_io_analog_sel[15]
port 131 nsew signal output
rlabel metal2 s 487717 952600 487773 953787 6 mprj_io_analog_sel[16]
port 132 nsew signal output
rlabel metal2 s 436317 952600 436373 953787 6 mprj_io_analog_sel[17]
port 133 nsew signal output
rlabel metal2 s 347317 952600 347373 953787 6 mprj_io_analog_sel[18]
port 134 nsew signal output
rlabel metal2 s 245517 952600 245573 953787 6 mprj_io_analog_sel[19]
port 135 nsew signal output
rlabel metal3 s 632200 113195 633437 113315 6 mprj_io_analog_sel[1]
port 136 nsew signal output
rlabel metal2 s 193917 952600 193973 953787 6 mprj_io_analog_sel[20]
port 137 nsew signal output
rlabel metal2 s 142517 952600 142573 953787 6 mprj_io_analog_sel[21]
port 138 nsew signal output
rlabel metal2 s 91117 952600 91173 953787 6 mprj_io_analog_sel[22]
port 139 nsew signal output
rlabel metal2 s 39717 952600 39773 953787 6 mprj_io_analog_sel[23]
port 140 nsew signal output
rlabel metal3 s -437 917885 800 918005 6 mprj_io_analog_sel[24]
port 141 nsew signal output
rlabel metal3 s -437 748085 800 748205 6 mprj_io_analog_sel[25]
port 142 nsew signal output
rlabel metal3 s -437 704885 800 705005 6 mprj_io_analog_sel[26]
port 143 nsew signal output
rlabel metal3 s -437 661685 800 661805 6 mprj_io_analog_sel[27]
port 144 nsew signal output
rlabel metal3 s -437 618485 800 618605 6 mprj_io_analog_sel[28]
port 145 nsew signal output
rlabel metal3 s -437 575285 800 575405 6 mprj_io_analog_sel[29]
port 146 nsew signal output
rlabel metal3 s 632200 158195 633437 158315 6 mprj_io_analog_sel[2]
port 147 nsew signal output
rlabel metal3 s -437 532085 800 532205 6 mprj_io_analog_sel[30]
port 148 nsew signal output
rlabel metal3 s -437 488885 800 489005 6 mprj_io_analog_sel[31]
port 149 nsew signal output
rlabel metal3 s -437 361285 800 361405 6 mprj_io_analog_sel[32]
port 150 nsew signal output
rlabel metal3 s -437 318085 800 318205 6 mprj_io_analog_sel[33]
port 151 nsew signal output
rlabel metal3 s -437 274885 800 275005 6 mprj_io_analog_sel[34]
port 152 nsew signal output
rlabel metal3 s -437 231685 800 231805 6 mprj_io_analog_sel[35]
port 153 nsew signal output
rlabel metal3 s -437 188485 800 188605 6 mprj_io_analog_sel[36]
port 154 nsew signal output
rlabel metal3 s -437 145285 800 145405 6 mprj_io_analog_sel[37]
port 155 nsew signal output
rlabel metal3 s 632200 203395 633437 203515 6 mprj_io_analog_sel[3]
port 156 nsew signal output
rlabel metal3 s 632200 248395 633437 248515 6 mprj_io_analog_sel[4]
port 157 nsew signal output
rlabel metal3 s 632200 293395 633437 293515 6 mprj_io_analog_sel[5]
port 158 nsew signal output
rlabel metal3 s 632200 338595 633437 338715 6 mprj_io_analog_sel[6]
port 159 nsew signal output
rlabel metal3 s 632200 515795 633437 515915 6 mprj_io_analog_sel[7]
port 160 nsew signal output
rlabel metal3 s 632200 560995 633437 561115 6 mprj_io_analog_sel[8]
port 161 nsew signal output
rlabel metal3 s 632200 605995 633437 606115 6 mprj_io_analog_sel[9]
port 162 nsew signal output
rlabel metal3 s 632200 64315 633437 64435 6 mprj_io_dm[0]
port 163 nsew signal output
rlabel metal3 s -437 323605 800 323725 6 mprj_io_dm[100]
port 164 nsew signal output
rlabel metal3 s -437 317441 800 317561 6 mprj_io_dm[101]
port 165 nsew signal output
rlabel metal3 s -437 278565 800 278685 6 mprj_io_dm[102]
port 166 nsew signal output
rlabel metal3 s -437 280405 800 280525 6 mprj_io_dm[103]
port 167 nsew signal output
rlabel metal3 s -437 274241 800 274361 6 mprj_io_dm[104]
port 168 nsew signal output
rlabel metal3 s -437 235365 858 235485 6 mprj_io_dm[105]
port 169 nsew signal output
rlabel metal3 s -437 237205 800 237325 6 mprj_io_dm[106]
port 170 nsew signal output
rlabel metal3 s -437 231041 800 231161 6 mprj_io_dm[107]
port 171 nsew signal output
rlabel metal3 s -437 192165 800 192285 6 mprj_io_dm[108]
port 172 nsew signal output
rlabel metal3 s -437 194005 800 194125 6 mprj_io_dm[109]
port 173 nsew signal output
rlabel metal3 s 632200 197875 633437 197995 6 mprj_io_dm[10]
port 174 nsew signal output
rlabel metal3 s -437 187841 800 187961 6 mprj_io_dm[110]
port 175 nsew signal output
rlabel metal3 s -437 148965 800 149085 6 mprj_io_dm[111]
port 176 nsew signal output
rlabel metal3 s -437 150805 800 150925 6 mprj_io_dm[112]
port 177 nsew signal output
rlabel metal3 s -437 144641 800 144761 6 mprj_io_dm[113]
port 178 nsew signal output
rlabel metal3 s 632200 204039 633437 204159 6 mprj_io_dm[11]
port 179 nsew signal output
rlabel metal3 s 632200 244715 633437 244835 6 mprj_io_dm[12]
port 180 nsew signal output
rlabel metal3 s 632200 242875 633437 242995 6 mprj_io_dm[13]
port 181 nsew signal output
rlabel metal3 s 632200 249039 633437 249159 6 mprj_io_dm[14]
port 182 nsew signal output
rlabel metal3 s 632200 289715 633437 289835 6 mprj_io_dm[15]
port 183 nsew signal output
rlabel metal3 s 632200 287875 633437 287995 6 mprj_io_dm[16]
port 184 nsew signal output
rlabel metal3 s 632200 294039 633437 294159 6 mprj_io_dm[17]
port 185 nsew signal output
rlabel metal3 s 632200 334915 633437 335035 6 mprj_io_dm[18]
port 186 nsew signal output
rlabel metal3 s 632200 333075 633437 333195 6 mprj_io_dm[19]
port 187 nsew signal output
rlabel metal3 s 632200 62475 633437 62595 6 mprj_io_dm[1]
port 188 nsew signal output
rlabel metal3 s 632200 339239 633437 339359 6 mprj_io_dm[20]
port 189 nsew signal output
rlabel metal3 s 632200 512115 633437 512235 6 mprj_io_dm[21]
port 190 nsew signal output
rlabel metal3 s 632200 510275 633437 510395 6 mprj_io_dm[22]
port 191 nsew signal output
rlabel metal3 s 632200 516439 633437 516559 6 mprj_io_dm[23]
port 192 nsew signal output
rlabel metal3 s 632200 557315 633437 557435 6 mprj_io_dm[24]
port 193 nsew signal output
rlabel metal3 s 632200 555475 633437 555595 6 mprj_io_dm[25]
port 194 nsew signal output
rlabel metal3 s 632200 561639 633437 561759 6 mprj_io_dm[26]
port 195 nsew signal output
rlabel metal3 s 632200 602315 633437 602435 6 mprj_io_dm[27]
port 196 nsew signal output
rlabel metal3 s 632200 600475 633437 600595 6 mprj_io_dm[28]
port 197 nsew signal output
rlabel metal3 s 632200 606639 633437 606759 6 mprj_io_dm[29]
port 198 nsew signal output
rlabel metal3 s 632200 68639 633437 68759 6 mprj_io_dm[2]
port 199 nsew signal output
rlabel metal3 s 632200 647515 633437 647635 6 mprj_io_dm[30]
port 200 nsew signal output
rlabel metal3 s 632200 645675 633437 645795 6 mprj_io_dm[31]
port 201 nsew signal output
rlabel metal3 s 632200 651839 633437 651959 6 mprj_io_dm[32]
port 202 nsew signal output
rlabel metal3 s 632200 692515 633437 692635 6 mprj_io_dm[33]
port 203 nsew signal output
rlabel metal3 s 632200 690675 633437 690795 6 mprj_io_dm[34]
port 204 nsew signal output
rlabel metal3 s 632200 696839 633437 696959 6 mprj_io_dm[35]
port 205 nsew signal output
rlabel metal3 s 632200 737515 633437 737635 6 mprj_io_dm[36]
port 206 nsew signal output
rlabel metal3 s 632200 735675 633437 735795 6 mprj_io_dm[37]
port 207 nsew signal output
rlabel metal3 s 632200 741839 633437 741959 6 mprj_io_dm[38]
port 208 nsew signal output
rlabel metal3 s 632200 826715 633437 826835 6 mprj_io_dm[39]
port 209 nsew signal output
rlabel metal3 s 632200 109515 633437 109635 6 mprj_io_dm[3]
port 210 nsew signal output
rlabel metal3 s 632200 824875 633437 824995 6 mprj_io_dm[40]
port 211 nsew signal output
rlabel metal3 s 632200 831039 633437 831159 6 mprj_io_dm[41]
port 212 nsew signal output
rlabel metal3 s 632200 915915 633437 916035 6 mprj_io_dm[42]
port 213 nsew signal output
rlabel metal3 s 632200 914075 633437 914195 6 mprj_io_dm[43]
port 214 nsew signal output
rlabel metal3 s 632200 920239 633437 920359 6 mprj_io_dm[44]
port 215 nsew signal output
rlabel metal2 s 593197 952600 593253 953787 6 mprj_io_dm[45]
port 216 nsew signal output
rlabel metal2 s 595037 952600 595093 953787 6 mprj_io_dm[46]
port 217 nsew signal output
rlabel metal2 s 588873 952600 588929 953787 6 mprj_io_dm[47]
port 218 nsew signal output
rlabel metal2 s 491397 952600 491453 953787 6 mprj_io_dm[48]
port 219 nsew signal output
rlabel metal2 s 493237 952600 493293 953787 6 mprj_io_dm[49]
port 220 nsew signal output
rlabel metal3 s 632200 107675 633437 107795 6 mprj_io_dm[4]
port 221 nsew signal output
rlabel metal2 s 487073 952600 487129 953787 6 mprj_io_dm[50]
port 222 nsew signal output
rlabel metal2 s 439997 952600 440053 953787 6 mprj_io_dm[51]
port 223 nsew signal output
rlabel metal2 s 441837 952600 441893 953787 6 mprj_io_dm[52]
port 224 nsew signal output
rlabel metal2 s 435673 952600 435729 953787 6 mprj_io_dm[53]
port 225 nsew signal output
rlabel metal2 s 350997 952600 351053 953787 6 mprj_io_dm[54]
port 226 nsew signal output
rlabel metal2 s 352837 952600 352893 953787 6 mprj_io_dm[55]
port 227 nsew signal output
rlabel metal2 s 346673 952600 346729 953787 6 mprj_io_dm[56]
port 228 nsew signal output
rlabel metal2 s 249197 952600 249253 953787 6 mprj_io_dm[57]
port 229 nsew signal output
rlabel metal2 s 251037 952600 251093 953787 6 mprj_io_dm[58]
port 230 nsew signal output
rlabel metal2 s 244873 952600 244929 953787 6 mprj_io_dm[59]
port 231 nsew signal output
rlabel metal3 s 632200 113839 633437 113959 6 mprj_io_dm[5]
port 232 nsew signal output
rlabel metal2 s 197597 952600 197653 953787 6 mprj_io_dm[60]
port 233 nsew signal output
rlabel metal2 s 199437 952600 199493 953787 6 mprj_io_dm[61]
port 234 nsew signal output
rlabel metal2 s 193273 952600 193329 953787 6 mprj_io_dm[62]
port 235 nsew signal output
rlabel metal2 s 146197 952600 146253 953787 6 mprj_io_dm[63]
port 236 nsew signal output
rlabel metal2 s 148037 952600 148093 953787 6 mprj_io_dm[64]
port 237 nsew signal output
rlabel metal2 s 141873 952600 141929 953787 6 mprj_io_dm[65]
port 238 nsew signal output
rlabel metal2 s 94797 952600 94853 953787 6 mprj_io_dm[66]
port 239 nsew signal output
rlabel metal2 s 96637 952600 96693 953787 6 mprj_io_dm[67]
port 240 nsew signal output
rlabel metal2 s 90473 952600 90529 953787 6 mprj_io_dm[68]
port 241 nsew signal output
rlabel metal2 s 43397 952600 43453 953787 6 mprj_io_dm[69]
port 242 nsew signal output
rlabel metal3 s 632200 154515 633437 154635 6 mprj_io_dm[6]
port 243 nsew signal output
rlabel metal2 s 45237 952600 45293 953787 6 mprj_io_dm[70]
port 244 nsew signal output
rlabel metal2 s 39073 952600 39129 953787 6 mprj_io_dm[71]
port 245 nsew signal output
rlabel metal3 s -437 921565 800 921685 6 mprj_io_dm[72]
port 246 nsew signal output
rlabel metal3 s -437 923405 800 923525 6 mprj_io_dm[73]
port 247 nsew signal output
rlabel metal3 s -437 917241 800 917361 6 mprj_io_dm[74]
port 248 nsew signal output
rlabel metal3 s -437 751765 800 751885 6 mprj_io_dm[75]
port 249 nsew signal output
rlabel metal3 s -437 753605 800 753725 6 mprj_io_dm[76]
port 250 nsew signal output
rlabel metal3 s -437 747441 800 747561 6 mprj_io_dm[77]
port 251 nsew signal output
rlabel metal3 s -437 708565 800 708685 6 mprj_io_dm[78]
port 252 nsew signal output
rlabel metal3 s -437 710405 800 710525 6 mprj_io_dm[79]
port 253 nsew signal output
rlabel metal3 s 632200 152675 633437 152795 6 mprj_io_dm[7]
port 254 nsew signal output
rlabel metal3 s -437 704241 800 704361 6 mprj_io_dm[80]
port 255 nsew signal output
rlabel metal3 s -437 665365 800 665485 6 mprj_io_dm[81]
port 256 nsew signal output
rlabel metal3 s -437 667205 800 667325 6 mprj_io_dm[82]
port 257 nsew signal output
rlabel metal3 s -437 661041 800 661161 6 mprj_io_dm[83]
port 258 nsew signal output
rlabel metal3 s -437 622165 800 622285 6 mprj_io_dm[84]
port 259 nsew signal output
rlabel metal3 s -437 624005 800 624125 6 mprj_io_dm[85]
port 260 nsew signal output
rlabel metal3 s -437 617841 800 617961 6 mprj_io_dm[86]
port 261 nsew signal output
rlabel metal3 s -437 578965 800 579085 6 mprj_io_dm[87]
port 262 nsew signal output
rlabel metal3 s -437 580805 800 580925 6 mprj_io_dm[88]
port 263 nsew signal output
rlabel metal3 s -437 574641 800 574761 6 mprj_io_dm[89]
port 264 nsew signal output
rlabel metal3 s 632200 158839 633437 158959 6 mprj_io_dm[8]
port 265 nsew signal output
rlabel metal3 s -437 535765 800 535885 6 mprj_io_dm[90]
port 266 nsew signal output
rlabel metal3 s -437 537605 800 537725 6 mprj_io_dm[91]
port 267 nsew signal output
rlabel metal3 s -437 531441 800 531561 6 mprj_io_dm[92]
port 268 nsew signal output
rlabel metal3 s -437 492565 800 492685 6 mprj_io_dm[93]
port 269 nsew signal output
rlabel metal3 s -437 494405 800 494525 6 mprj_io_dm[94]
port 270 nsew signal output
rlabel metal3 s -437 488241 800 488361 6 mprj_io_dm[95]
port 271 nsew signal output
rlabel metal3 s -437 364965 800 365085 6 mprj_io_dm[96]
port 272 nsew signal output
rlabel metal3 s -437 366805 800 366925 6 mprj_io_dm[97]
port 273 nsew signal output
rlabel metal3 s -437 360641 800 360761 6 mprj_io_dm[98]
port 274 nsew signal output
rlabel metal3 s -437 321765 800 321885 6 mprj_io_dm[99]
port 275 nsew signal output
rlabel metal3 s 632200 199715 633437 199835 6 mprj_io_dm[9]
port 276 nsew signal output
rlabel metal3 s 632200 69283 633437 69403 6 mprj_io_holdover[0]
port 277 nsew signal output
rlabel metal3 s 632200 652483 633437 652603 6 mprj_io_holdover[10]
port 278 nsew signal output
rlabel metal3 s 632200 697483 633437 697603 6 mprj_io_holdover[11]
port 279 nsew signal output
rlabel metal3 s 632200 742483 633437 742603 6 mprj_io_holdover[12]
port 280 nsew signal output
rlabel metal3 s 632200 831683 633437 831803 6 mprj_io_holdover[13]
port 281 nsew signal output
rlabel metal3 s 632200 920883 633437 921003 6 mprj_io_holdover[14]
port 282 nsew signal output
rlabel metal2 s 588229 952600 588285 953787 6 mprj_io_holdover[15]
port 283 nsew signal output
rlabel metal2 s 486429 952600 486485 953787 6 mprj_io_holdover[16]
port 284 nsew signal output
rlabel metal2 s 435029 952600 435085 953787 6 mprj_io_holdover[17]
port 285 nsew signal output
rlabel metal2 s 346029 952600 346085 953787 6 mprj_io_holdover[18]
port 286 nsew signal output
rlabel metal2 s 244229 952600 244285 953787 6 mprj_io_holdover[19]
port 287 nsew signal output
rlabel metal3 s 632200 114483 633437 114603 6 mprj_io_holdover[1]
port 288 nsew signal output
rlabel metal2 s 192629 952600 192685 953787 6 mprj_io_holdover[20]
port 289 nsew signal output
rlabel metal2 s 141229 952600 141285 953787 6 mprj_io_holdover[21]
port 290 nsew signal output
rlabel metal2 s 89829 952600 89885 953787 6 mprj_io_holdover[22]
port 291 nsew signal output
rlabel metal2 s 38429 952600 38485 953787 6 mprj_io_holdover[23]
port 292 nsew signal output
rlabel metal3 s -437 916597 800 916717 6 mprj_io_holdover[24]
port 293 nsew signal output
rlabel metal3 s -437 746797 800 746917 6 mprj_io_holdover[25]
port 294 nsew signal output
rlabel metal3 s -437 703597 800 703717 6 mprj_io_holdover[26]
port 295 nsew signal output
rlabel metal3 s -437 660397 800 660517 6 mprj_io_holdover[27]
port 296 nsew signal output
rlabel metal3 s -437 617197 800 617317 6 mprj_io_holdover[28]
port 297 nsew signal output
rlabel metal3 s -437 573997 800 574117 6 mprj_io_holdover[29]
port 298 nsew signal output
rlabel metal3 s 632200 159483 633437 159603 6 mprj_io_holdover[2]
port 299 nsew signal output
rlabel metal3 s -437 530797 800 530917 6 mprj_io_holdover[30]
port 300 nsew signal output
rlabel metal3 s -437 487597 800 487717 6 mprj_io_holdover[31]
port 301 nsew signal output
rlabel metal3 s -437 359997 800 360117 6 mprj_io_holdover[32]
port 302 nsew signal output
rlabel metal3 s -437 316797 800 316917 6 mprj_io_holdover[33]
port 303 nsew signal output
rlabel metal3 s -437 273597 800 273717 6 mprj_io_holdover[34]
port 304 nsew signal output
rlabel metal3 s -437 230397 800 230517 6 mprj_io_holdover[35]
port 305 nsew signal output
rlabel metal3 s -437 187197 800 187317 6 mprj_io_holdover[36]
port 306 nsew signal output
rlabel metal3 s -437 143997 800 144117 6 mprj_io_holdover[37]
port 307 nsew signal output
rlabel metal3 s 632200 204683 633437 204803 6 mprj_io_holdover[3]
port 308 nsew signal output
rlabel metal3 s 632200 249683 633437 249803 6 mprj_io_holdover[4]
port 309 nsew signal output
rlabel metal3 s 632200 294683 633437 294803 6 mprj_io_holdover[5]
port 310 nsew signal output
rlabel metal3 s 632200 339883 633437 340003 6 mprj_io_holdover[6]
port 311 nsew signal output
rlabel metal3 s 632200 517083 633437 517203 6 mprj_io_holdover[7]
port 312 nsew signal output
rlabel metal3 s 632200 562283 633437 562403 6 mprj_io_holdover[8]
port 313 nsew signal output
rlabel metal3 s 632200 607283 633437 607403 6 mprj_io_holdover[9]
port 314 nsew signal output
rlabel metal3 s 632200 72319 633437 72439 6 mprj_io_ib_mode_sel[0]
port 315 nsew signal output
rlabel metal3 s 632200 655519 633437 655639 6 mprj_io_ib_mode_sel[10]
port 316 nsew signal output
rlabel metal3 s 632200 700519 633437 700639 6 mprj_io_ib_mode_sel[11]
port 317 nsew signal output
rlabel metal3 s 632200 745519 633437 745639 6 mprj_io_ib_mode_sel[12]
port 318 nsew signal output
rlabel metal3 s 632200 834719 633437 834839 6 mprj_io_ib_mode_sel[13]
port 319 nsew signal output
rlabel metal3 s 632200 923919 633437 924039 6 mprj_io_ib_mode_sel[14]
port 320 nsew signal output
rlabel metal2 s 585193 952600 585249 953787 6 mprj_io_ib_mode_sel[15]
port 321 nsew signal output
rlabel metal2 s 483393 952600 483449 953787 6 mprj_io_ib_mode_sel[16]
port 322 nsew signal output
rlabel metal2 s 431993 952600 432049 953787 6 mprj_io_ib_mode_sel[17]
port 323 nsew signal output
rlabel metal2 s 342993 952600 343049 953787 6 mprj_io_ib_mode_sel[18]
port 324 nsew signal output
rlabel metal2 s 241193 952600 241249 953787 6 mprj_io_ib_mode_sel[19]
port 325 nsew signal output
rlabel metal3 s 632200 117519 633437 117639 6 mprj_io_ib_mode_sel[1]
port 326 nsew signal output
rlabel metal2 s 189593 952600 189649 953787 6 mprj_io_ib_mode_sel[20]
port 327 nsew signal output
rlabel metal2 s 138193 952600 138249 953787 6 mprj_io_ib_mode_sel[21]
port 328 nsew signal output
rlabel metal2 s 86793 952600 86849 953787 6 mprj_io_ib_mode_sel[22]
port 329 nsew signal output
rlabel metal2 s 35393 952600 35449 953787 6 mprj_io_ib_mode_sel[23]
port 330 nsew signal output
rlabel metal3 s -437 913561 800 913681 6 mprj_io_ib_mode_sel[24]
port 331 nsew signal output
rlabel metal3 s -437 743761 800 743881 6 mprj_io_ib_mode_sel[25]
port 332 nsew signal output
rlabel metal3 s -437 700561 800 700681 6 mprj_io_ib_mode_sel[26]
port 333 nsew signal output
rlabel metal3 s -437 657361 800 657481 6 mprj_io_ib_mode_sel[27]
port 334 nsew signal output
rlabel metal3 s -437 614161 800 614281 6 mprj_io_ib_mode_sel[28]
port 335 nsew signal output
rlabel metal3 s -437 570961 800 571081 6 mprj_io_ib_mode_sel[29]
port 336 nsew signal output
rlabel metal3 s 632200 162519 633437 162639 6 mprj_io_ib_mode_sel[2]
port 337 nsew signal output
rlabel metal3 s -437 527761 800 527881 6 mprj_io_ib_mode_sel[30]
port 338 nsew signal output
rlabel metal3 s -437 484561 800 484681 6 mprj_io_ib_mode_sel[31]
port 339 nsew signal output
rlabel metal3 s -437 356961 800 357081 6 mprj_io_ib_mode_sel[32]
port 340 nsew signal output
rlabel metal3 s -437 313761 800 313881 6 mprj_io_ib_mode_sel[33]
port 341 nsew signal output
rlabel metal3 s -437 270561 800 270681 6 mprj_io_ib_mode_sel[34]
port 342 nsew signal output
rlabel metal3 s -437 227361 800 227481 6 mprj_io_ib_mode_sel[35]
port 343 nsew signal output
rlabel metal3 s -437 184161 800 184281 6 mprj_io_ib_mode_sel[36]
port 344 nsew signal output
rlabel metal3 s -437 140961 800 141081 6 mprj_io_ib_mode_sel[37]
port 345 nsew signal output
rlabel metal3 s 632200 207719 633437 207839 6 mprj_io_ib_mode_sel[3]
port 346 nsew signal output
rlabel metal3 s 632200 252719 633437 252839 6 mprj_io_ib_mode_sel[4]
port 347 nsew signal output
rlabel metal3 s 632200 297719 633437 297839 6 mprj_io_ib_mode_sel[5]
port 348 nsew signal output
rlabel metal3 s 632200 342919 633437 343039 6 mprj_io_ib_mode_sel[6]
port 349 nsew signal output
rlabel metal3 s 632200 520119 633437 520239 6 mprj_io_ib_mode_sel[7]
port 350 nsew signal output
rlabel metal3 s 632200 565319 633437 565439 6 mprj_io_ib_mode_sel[8]
port 351 nsew signal output
rlabel metal3 s 632200 610319 633437 610439 6 mprj_io_ib_mode_sel[9]
port 352 nsew signal output
rlabel metal3 s 632200 58795 633437 58915 6 mprj_io_in[0]
port 353 nsew signal input
rlabel metal3 s 632200 641995 633437 642115 6 mprj_io_in[10]
port 354 nsew signal input
rlabel metal3 s 632200 686995 633437 687115 6 mprj_io_in[11]
port 355 nsew signal input
rlabel metal3 s 632200 731995 633437 732115 6 mprj_io_in[12]
port 356 nsew signal input
rlabel metal3 s 632200 821195 633437 821315 6 mprj_io_in[13]
port 357 nsew signal input
rlabel metal3 s 632200 910395 633437 910515 6 mprj_io_in[14]
port 358 nsew signal input
rlabel metal2 s 598717 952600 598773 953787 6 mprj_io_in[15]
port 359 nsew signal input
rlabel metal2 s 496917 952600 496973 953787 6 mprj_io_in[16]
port 360 nsew signal input
rlabel metal2 s 445517 952600 445573 953787 6 mprj_io_in[17]
port 361 nsew signal input
rlabel metal2 s 356517 952600 356573 953787 6 mprj_io_in[18]
port 362 nsew signal input
rlabel metal2 s 254717 952600 254773 953787 6 mprj_io_in[19]
port 363 nsew signal input
rlabel metal3 s 632200 103995 633437 104115 6 mprj_io_in[1]
port 364 nsew signal input
rlabel metal2 s 203117 952600 203173 953787 6 mprj_io_in[20]
port 365 nsew signal input
rlabel metal2 s 151717 952600 151773 953787 6 mprj_io_in[21]
port 366 nsew signal input
rlabel metal2 s 100317 952600 100373 953787 6 mprj_io_in[22]
port 367 nsew signal input
rlabel metal2 s 48917 952600 48973 953787 6 mprj_io_in[23]
port 368 nsew signal input
rlabel metal3 s -437 927085 800 927205 6 mprj_io_in[24]
port 369 nsew signal input
rlabel metal3 s -437 757285 800 757405 6 mprj_io_in[25]
port 370 nsew signal input
rlabel metal3 s -437 714085 800 714205 6 mprj_io_in[26]
port 371 nsew signal input
rlabel metal3 s -437 670885 800 671005 6 mprj_io_in[27]
port 372 nsew signal input
rlabel metal3 s -437 627685 800 627805 6 mprj_io_in[28]
port 373 nsew signal input
rlabel metal3 s -437 584485 800 584605 6 mprj_io_in[29]
port 374 nsew signal input
rlabel metal3 s 632200 148995 633437 149115 6 mprj_io_in[2]
port 375 nsew signal input
rlabel metal3 s -437 541285 800 541405 6 mprj_io_in[30]
port 376 nsew signal input
rlabel metal3 s -437 498085 800 498205 6 mprj_io_in[31]
port 377 nsew signal input
rlabel metal3 s -437 370485 800 370605 6 mprj_io_in[32]
port 378 nsew signal input
rlabel metal3 s -437 327285 800 327405 6 mprj_io_in[33]
port 379 nsew signal input
rlabel metal3 s -437 284085 800 284205 6 mprj_io_in[34]
port 380 nsew signal input
rlabel metal3 s -437 240885 800 241005 6 mprj_io_in[35]
port 381 nsew signal input
rlabel metal3 s -437 197685 800 197805 6 mprj_io_in[36]
port 382 nsew signal input
rlabel metal3 s -437 154485 800 154605 6 mprj_io_in[37]
port 383 nsew signal input
rlabel metal3 s 632200 194195 633437 194315 6 mprj_io_in[3]
port 384 nsew signal input
rlabel metal3 s 632200 239195 633437 239315 6 mprj_io_in[4]
port 385 nsew signal input
rlabel metal3 s 632200 284195 633437 284315 6 mprj_io_in[5]
port 386 nsew signal input
rlabel metal3 s 632200 329395 633437 329515 6 mprj_io_in[6]
port 387 nsew signal input
rlabel metal3 s 632200 506595 633437 506715 6 mprj_io_in[7]
port 388 nsew signal input
rlabel metal3 s 632200 551795 633437 551915 6 mprj_io_in[8]
port 389 nsew signal input
rlabel metal3 s 632200 596795 633437 596915 6 mprj_io_in[9]
port 390 nsew signal input
rlabel metal3 s 632200 65511 633437 65631 6 mprj_io_inp_dis[0]
port 391 nsew signal output
rlabel metal3 s 632200 648711 633437 648831 6 mprj_io_inp_dis[10]
port 392 nsew signal output
rlabel metal3 s 632200 693711 633437 693831 6 mprj_io_inp_dis[11]
port 393 nsew signal output
rlabel metal3 s 632200 738711 633437 738831 6 mprj_io_inp_dis[12]
port 394 nsew signal output
rlabel metal3 s 632200 827911 633437 828031 6 mprj_io_inp_dis[13]
port 395 nsew signal output
rlabel metal3 s 632200 917111 633437 917231 6 mprj_io_inp_dis[14]
port 396 nsew signal output
rlabel metal2 s 592001 952600 592057 953787 6 mprj_io_inp_dis[15]
port 397 nsew signal output
rlabel metal2 s 490201 952600 490257 953787 6 mprj_io_inp_dis[16]
port 398 nsew signal output
rlabel metal2 s 438801 952600 438857 953787 6 mprj_io_inp_dis[17]
port 399 nsew signal output
rlabel metal2 s 349801 952600 349857 953787 6 mprj_io_inp_dis[18]
port 400 nsew signal output
rlabel metal2 s 248001 952600 248057 953787 6 mprj_io_inp_dis[19]
port 401 nsew signal output
rlabel metal3 s 632200 110711 633437 110831 6 mprj_io_inp_dis[1]
port 402 nsew signal output
rlabel metal2 s 196401 952600 196457 953787 6 mprj_io_inp_dis[20]
port 403 nsew signal output
rlabel metal2 s 145001 952600 145057 953787 6 mprj_io_inp_dis[21]
port 404 nsew signal output
rlabel metal2 s 93601 952600 93657 953787 6 mprj_io_inp_dis[22]
port 405 nsew signal output
rlabel metal2 s 42201 952600 42257 953787 6 mprj_io_inp_dis[23]
port 406 nsew signal output
rlabel metal3 s -437 920369 800 920489 6 mprj_io_inp_dis[24]
port 407 nsew signal output
rlabel metal3 s -437 750569 800 750689 6 mprj_io_inp_dis[25]
port 408 nsew signal output
rlabel metal3 s -437 707369 800 707489 6 mprj_io_inp_dis[26]
port 409 nsew signal output
rlabel metal3 s -437 664169 800 664289 6 mprj_io_inp_dis[27]
port 410 nsew signal output
rlabel metal3 s -437 620969 800 621089 6 mprj_io_inp_dis[28]
port 411 nsew signal output
rlabel metal3 s -437 577769 800 577889 6 mprj_io_inp_dis[29]
port 412 nsew signal output
rlabel metal3 s 632200 155711 633437 155831 6 mprj_io_inp_dis[2]
port 413 nsew signal output
rlabel metal3 s -437 534569 800 534689 6 mprj_io_inp_dis[30]
port 414 nsew signal output
rlabel metal3 s -437 491369 800 491489 6 mprj_io_inp_dis[31]
port 415 nsew signal output
rlabel metal3 s -437 363769 800 363889 6 mprj_io_inp_dis[32]
port 416 nsew signal output
rlabel metal3 s -437 320569 800 320689 6 mprj_io_inp_dis[33]
port 417 nsew signal output
rlabel metal3 s -437 277369 800 277489 6 mprj_io_inp_dis[34]
port 418 nsew signal output
rlabel metal3 s -437 234169 800 234289 6 mprj_io_inp_dis[35]
port 419 nsew signal output
rlabel metal3 s -437 190969 800 191089 6 mprj_io_inp_dis[36]
port 420 nsew signal output
rlabel metal3 s -437 147769 800 147889 6 mprj_io_inp_dis[37]
port 421 nsew signal output
rlabel metal3 s 632200 200911 633437 201031 6 mprj_io_inp_dis[3]
port 422 nsew signal output
rlabel metal3 s 632200 245911 633437 246031 6 mprj_io_inp_dis[4]
port 423 nsew signal output
rlabel metal3 s 632200 290911 633437 291031 6 mprj_io_inp_dis[5]
port 424 nsew signal output
rlabel metal3 s 632200 336111 633437 336231 6 mprj_io_inp_dis[6]
port 425 nsew signal output
rlabel metal3 s 632200 513311 633437 513431 6 mprj_io_inp_dis[7]
port 426 nsew signal output
rlabel metal3 s 632200 558511 633437 558631 6 mprj_io_inp_dis[8]
port 427 nsew signal output
rlabel metal3 s 632200 603511 633437 603631 6 mprj_io_inp_dis[9]
port 428 nsew signal output
rlabel metal3 s 632200 72963 633437 73083 6 mprj_io_oeb[0]
port 429 nsew signal output
rlabel metal3 s 632200 656163 633437 656283 6 mprj_io_oeb[10]
port 430 nsew signal output
rlabel metal3 s 632200 701163 633437 701283 6 mprj_io_oeb[11]
port 431 nsew signal output
rlabel metal3 s 632200 746163 633437 746283 6 mprj_io_oeb[12]
port 432 nsew signal output
rlabel metal3 s 632200 835363 633437 835483 6 mprj_io_oeb[13]
port 433 nsew signal output
rlabel metal3 s 632200 924563 633437 924683 6 mprj_io_oeb[14]
port 434 nsew signal output
rlabel metal2 s 584549 952600 584605 953787 6 mprj_io_oeb[15]
port 435 nsew signal output
rlabel metal2 s 482749 952600 482805 953787 6 mprj_io_oeb[16]
port 436 nsew signal output
rlabel metal2 s 431349 952600 431405 953787 6 mprj_io_oeb[17]
port 437 nsew signal output
rlabel metal2 s 342349 952600 342405 953787 6 mprj_io_oeb[18]
port 438 nsew signal output
rlabel metal2 s 240549 952600 240605 953787 6 mprj_io_oeb[19]
port 439 nsew signal output
rlabel metal3 s 632200 118163 633437 118283 6 mprj_io_oeb[1]
port 440 nsew signal output
rlabel metal2 s 188949 952600 189005 953787 6 mprj_io_oeb[20]
port 441 nsew signal output
rlabel metal2 s 137549 952600 137605 953787 6 mprj_io_oeb[21]
port 442 nsew signal output
rlabel metal2 s 86149 952600 86205 953787 6 mprj_io_oeb[22]
port 443 nsew signal output
rlabel metal2 s 34749 952600 34805 953787 6 mprj_io_oeb[23]
port 444 nsew signal output
rlabel metal3 s -437 912917 800 913037 6 mprj_io_oeb[24]
port 445 nsew signal output
rlabel metal3 s -437 743117 800 743237 6 mprj_io_oeb[25]
port 446 nsew signal output
rlabel metal3 s -437 699917 800 700037 6 mprj_io_oeb[26]
port 447 nsew signal output
rlabel metal3 s -437 656717 800 656837 6 mprj_io_oeb[27]
port 448 nsew signal output
rlabel metal3 s -437 613517 800 613637 6 mprj_io_oeb[28]
port 449 nsew signal output
rlabel metal3 s -437 570317 800 570437 6 mprj_io_oeb[29]
port 450 nsew signal output
rlabel metal3 s 632200 163163 633437 163283 6 mprj_io_oeb[2]
port 451 nsew signal output
rlabel metal3 s -437 527117 800 527237 6 mprj_io_oeb[30]
port 452 nsew signal output
rlabel metal3 s -437 483917 800 484037 6 mprj_io_oeb[31]
port 453 nsew signal output
rlabel metal3 s -437 356317 800 356437 6 mprj_io_oeb[32]
port 454 nsew signal output
rlabel metal3 s -437 313117 800 313237 6 mprj_io_oeb[33]
port 455 nsew signal output
rlabel metal3 s -437 269917 800 270037 6 mprj_io_oeb[34]
port 456 nsew signal output
rlabel metal3 s -437 226717 800 226837 6 mprj_io_oeb[35]
port 457 nsew signal output
rlabel metal3 s -437 183517 800 183637 6 mprj_io_oeb[36]
port 458 nsew signal output
rlabel metal3 s -437 140317 800 140437 6 mprj_io_oeb[37]
port 459 nsew signal output
rlabel metal3 s 632200 208363 633437 208483 6 mprj_io_oeb[3]
port 460 nsew signal output
rlabel metal3 s 632200 253363 633437 253483 6 mprj_io_oeb[4]
port 461 nsew signal output
rlabel metal3 s 632200 298363 633437 298483 6 mprj_io_oeb[5]
port 462 nsew signal output
rlabel metal3 s 632200 343563 633437 343683 6 mprj_io_oeb[6]
port 463 nsew signal output
rlabel metal3 s 632200 520763 633437 520883 6 mprj_io_oeb[7]
port 464 nsew signal output
rlabel metal3 s 632200 565963 633437 566083 6 mprj_io_oeb[8]
port 465 nsew signal output
rlabel metal3 s 632200 610963 633437 611083 6 mprj_io_oeb[9]
port 466 nsew signal output
rlabel metal3 s 632200 59991 633437 60111 6 mprj_io_one[0]
port 467 nsew signal output
rlabel metal3 s 632200 643191 633437 643311 6 mprj_io_one[10]
port 468 nsew signal output
rlabel metal3 s 632200 688191 633437 688311 6 mprj_io_one[11]
port 469 nsew signal output
rlabel metal3 s 632200 733191 633437 733311 6 mprj_io_one[12]
port 470 nsew signal output
rlabel metal3 s 632200 822391 633437 822511 6 mprj_io_one[13]
port 471 nsew signal output
rlabel metal3 s 632200 911591 633437 911711 6 mprj_io_one[14]
port 472 nsew signal output
rlabel metal2 s 597521 952600 597577 953787 6 mprj_io_one[15]
port 473 nsew signal output
rlabel metal2 s 495721 952600 495777 953787 6 mprj_io_one[16]
port 474 nsew signal output
rlabel metal2 s 444321 952600 444377 953787 6 mprj_io_one[17]
port 475 nsew signal output
rlabel metal2 s 355321 952600 355377 953787 6 mprj_io_one[18]
port 476 nsew signal output
rlabel metal2 s 253521 952600 253577 953787 6 mprj_io_one[19]
port 477 nsew signal output
rlabel metal3 s 632200 105191 633437 105311 6 mprj_io_one[1]
port 478 nsew signal output
rlabel metal2 s 201921 952600 201977 953787 6 mprj_io_one[20]
port 479 nsew signal output
rlabel metal2 s 150521 952600 150577 953787 6 mprj_io_one[21]
port 480 nsew signal output
rlabel metal2 s 99121 952600 99177 953787 6 mprj_io_one[22]
port 481 nsew signal output
rlabel metal2 s 47721 952600 47777 953787 6 mprj_io_one[23]
port 482 nsew signal output
rlabel metal3 s -437 925889 800 926009 6 mprj_io_one[24]
port 483 nsew signal output
rlabel metal3 s -437 756089 800 756209 6 mprj_io_one[25]
port 484 nsew signal output
rlabel metal3 s -437 712889 800 713009 6 mprj_io_one[26]
port 485 nsew signal output
rlabel metal3 s -437 669689 800 669809 6 mprj_io_one[27]
port 486 nsew signal output
rlabel metal3 s -437 626489 800 626609 6 mprj_io_one[28]
port 487 nsew signal output
rlabel metal3 s -437 583289 800 583409 6 mprj_io_one[29]
port 488 nsew signal output
rlabel metal3 s 632200 150191 633437 150311 6 mprj_io_one[2]
port 489 nsew signal output
rlabel metal3 s -437 540089 800 540209 6 mprj_io_one[30]
port 490 nsew signal output
rlabel metal3 s -437 496889 800 497009 6 mprj_io_one[31]
port 491 nsew signal output
rlabel metal3 s -437 369289 800 369409 6 mprj_io_one[32]
port 492 nsew signal output
rlabel metal3 s -437 326089 800 326209 6 mprj_io_one[33]
port 493 nsew signal output
rlabel metal3 s -437 282889 800 283009 6 mprj_io_one[34]
port 494 nsew signal output
rlabel metal3 s -437 239689 858 239809 6 mprj_io_one[35]
port 495 nsew signal output
rlabel metal3 s -437 196489 800 196609 6 mprj_io_one[36]
port 496 nsew signal output
rlabel metal3 s -437 153289 800 153409 6 mprj_io_one[37]
port 497 nsew signal output
rlabel metal3 s 632200 195391 633437 195511 6 mprj_io_one[3]
port 498 nsew signal output
rlabel metal3 s 632200 240391 633437 240511 6 mprj_io_one[4]
port 499 nsew signal output
rlabel metal3 s 632200 285391 633437 285511 6 mprj_io_one[5]
port 500 nsew signal output
rlabel metal3 s 632200 330591 633437 330711 6 mprj_io_one[6]
port 501 nsew signal output
rlabel metal3 s 632200 507791 633437 507911 6 mprj_io_one[7]
port 502 nsew signal output
rlabel metal3 s 632200 552991 633437 553111 6 mprj_io_one[8]
port 503 nsew signal output
rlabel metal3 s 632200 597991 633437 598111 6 mprj_io_one[9]
port 504 nsew signal output
rlabel metal3 s 632200 69835 633437 69955 6 mprj_io_out[0]
port 505 nsew signal output
rlabel metal3 s 632200 653035 633437 653155 6 mprj_io_out[10]
port 506 nsew signal output
rlabel metal3 s 632200 698035 633437 698155 6 mprj_io_out[11]
port 507 nsew signal output
rlabel metal3 s 632200 743035 633437 743155 6 mprj_io_out[12]
port 508 nsew signal output
rlabel metal3 s 632200 832235 633437 832355 6 mprj_io_out[13]
port 509 nsew signal output
rlabel metal3 s 632200 921435 633437 921555 6 mprj_io_out[14]
port 510 nsew signal output
rlabel metal2 s 587677 952600 587733 953787 6 mprj_io_out[15]
port 511 nsew signal output
rlabel metal2 s 485877 952600 485933 953787 6 mprj_io_out[16]
port 512 nsew signal output
rlabel metal2 s 434477 952600 434533 953787 6 mprj_io_out[17]
port 513 nsew signal output
rlabel metal2 s 345477 952600 345533 953787 6 mprj_io_out[18]
port 514 nsew signal output
rlabel metal2 s 243677 952600 243733 953787 6 mprj_io_out[19]
port 515 nsew signal output
rlabel metal3 s 632200 115035 633437 115155 6 mprj_io_out[1]
port 516 nsew signal output
rlabel metal2 s 192077 952600 192133 953787 6 mprj_io_out[20]
port 517 nsew signal output
rlabel metal2 s 140677 952600 140733 953787 6 mprj_io_out[21]
port 518 nsew signal output
rlabel metal2 s 89277 952600 89333 953787 6 mprj_io_out[22]
port 519 nsew signal output
rlabel metal2 s 37877 952600 37933 953787 6 mprj_io_out[23]
port 520 nsew signal output
rlabel metal3 s -437 916045 800 916165 6 mprj_io_out[24]
port 521 nsew signal output
rlabel metal3 s -437 746245 800 746365 6 mprj_io_out[25]
port 522 nsew signal output
rlabel metal3 s -437 703045 800 703165 6 mprj_io_out[26]
port 523 nsew signal output
rlabel metal3 s -437 659845 800 659965 6 mprj_io_out[27]
port 524 nsew signal output
rlabel metal3 s -437 616645 800 616765 6 mprj_io_out[28]
port 525 nsew signal output
rlabel metal3 s -437 573445 800 573565 6 mprj_io_out[29]
port 526 nsew signal output
rlabel metal3 s 632200 160035 633437 160155 6 mprj_io_out[2]
port 527 nsew signal output
rlabel metal3 s -437 530245 800 530365 6 mprj_io_out[30]
port 528 nsew signal output
rlabel metal3 s -437 487045 800 487165 6 mprj_io_out[31]
port 529 nsew signal output
rlabel metal3 s -437 359445 800 359565 6 mprj_io_out[32]
port 530 nsew signal output
rlabel metal3 s -437 316245 800 316365 6 mprj_io_out[33]
port 531 nsew signal output
rlabel metal3 s -437 273045 800 273165 6 mprj_io_out[34]
port 532 nsew signal output
rlabel metal3 s -437 229845 800 229965 6 mprj_io_out[35]
port 533 nsew signal output
rlabel metal3 s -437 186645 800 186765 6 mprj_io_out[36]
port 534 nsew signal output
rlabel metal3 s -437 143445 800 143565 6 mprj_io_out[37]
port 535 nsew signal output
rlabel metal3 s 632200 205235 633437 205355 6 mprj_io_out[3]
port 536 nsew signal output
rlabel metal3 s 632200 250235 633437 250355 6 mprj_io_out[4]
port 537 nsew signal output
rlabel metal3 s 632200 295235 633437 295355 6 mprj_io_out[5]
port 538 nsew signal output
rlabel metal3 s 632200 340435 633437 340555 6 mprj_io_out[6]
port 539 nsew signal output
rlabel metal3 s 632200 517635 633437 517755 6 mprj_io_out[7]
port 540 nsew signal output
rlabel metal3 s 632200 562835 633437 562955 6 mprj_io_out[8]
port 541 nsew signal output
rlabel metal3 s 632200 607835 633437 607955 6 mprj_io_out[9]
port 542 nsew signal output
rlabel metal3 s 632200 60635 633437 60755 6 mprj_io_slow_sel[0]
port 543 nsew signal output
rlabel metal3 s 632200 643835 633437 643955 6 mprj_io_slow_sel[10]
port 544 nsew signal output
rlabel metal3 s 632200 688835 633437 688955 6 mprj_io_slow_sel[11]
port 545 nsew signal output
rlabel metal3 s 632200 733835 633437 733955 6 mprj_io_slow_sel[12]
port 546 nsew signal output
rlabel metal3 s 632200 823035 633437 823155 6 mprj_io_slow_sel[13]
port 547 nsew signal output
rlabel metal3 s 632200 912235 633437 912355 6 mprj_io_slow_sel[14]
port 548 nsew signal output
rlabel metal2 s 596877 952600 596933 953787 6 mprj_io_slow_sel[15]
port 549 nsew signal output
rlabel metal2 s 495077 952600 495133 953787 6 mprj_io_slow_sel[16]
port 550 nsew signal output
rlabel metal2 s 443677 952600 443733 953787 6 mprj_io_slow_sel[17]
port 551 nsew signal output
rlabel metal2 s 354677 952600 354733 953787 6 mprj_io_slow_sel[18]
port 552 nsew signal output
rlabel metal2 s 252877 952600 252933 953787 6 mprj_io_slow_sel[19]
port 553 nsew signal output
rlabel metal3 s 632200 105835 633437 105955 6 mprj_io_slow_sel[1]
port 554 nsew signal output
rlabel metal2 s 201277 952600 201333 953787 6 mprj_io_slow_sel[20]
port 555 nsew signal output
rlabel metal2 s 149877 952600 149933 953787 6 mprj_io_slow_sel[21]
port 556 nsew signal output
rlabel metal2 s 98477 952600 98533 953787 6 mprj_io_slow_sel[22]
port 557 nsew signal output
rlabel metal2 s 47077 952600 47133 953787 6 mprj_io_slow_sel[23]
port 558 nsew signal output
rlabel metal3 s -437 925245 800 925365 6 mprj_io_slow_sel[24]
port 559 nsew signal output
rlabel metal3 s -437 755445 800 755565 6 mprj_io_slow_sel[25]
port 560 nsew signal output
rlabel metal3 s -437 712245 800 712365 6 mprj_io_slow_sel[26]
port 561 nsew signal output
rlabel metal3 s -437 669045 800 669165 6 mprj_io_slow_sel[27]
port 562 nsew signal output
rlabel metal3 s -437 625845 800 625965 6 mprj_io_slow_sel[28]
port 563 nsew signal output
rlabel metal3 s -437 582645 800 582765 6 mprj_io_slow_sel[29]
port 564 nsew signal output
rlabel metal3 s 632200 150835 633437 150955 6 mprj_io_slow_sel[2]
port 565 nsew signal output
rlabel metal3 s -437 539445 800 539565 6 mprj_io_slow_sel[30]
port 566 nsew signal output
rlabel metal3 s -437 496245 800 496365 6 mprj_io_slow_sel[31]
port 567 nsew signal output
rlabel metal3 s -437 368645 800 368765 6 mprj_io_slow_sel[32]
port 568 nsew signal output
rlabel metal3 s -437 325445 800 325565 6 mprj_io_slow_sel[33]
port 569 nsew signal output
rlabel metal3 s -437 282245 800 282365 6 mprj_io_slow_sel[34]
port 570 nsew signal output
rlabel metal3 s -437 239045 800 239165 6 mprj_io_slow_sel[35]
port 571 nsew signal output
rlabel metal3 s -437 195845 800 195965 6 mprj_io_slow_sel[36]
port 572 nsew signal output
rlabel metal3 s -437 152645 800 152765 6 mprj_io_slow_sel[37]
port 573 nsew signal output
rlabel metal3 s 632200 196035 633437 196155 6 mprj_io_slow_sel[3]
port 574 nsew signal output
rlabel metal3 s 632200 241035 633437 241155 6 mprj_io_slow_sel[4]
port 575 nsew signal output
rlabel metal3 s 632200 286035 633437 286155 6 mprj_io_slow_sel[5]
port 576 nsew signal output
rlabel metal3 s 632200 331235 633437 331355 6 mprj_io_slow_sel[6]
port 577 nsew signal output
rlabel metal3 s 632200 508435 633437 508555 6 mprj_io_slow_sel[7]
port 578 nsew signal output
rlabel metal3 s 632200 553635 633437 553755 6 mprj_io_slow_sel[8]
port 579 nsew signal output
rlabel metal3 s 632200 598635 633437 598755 6 mprj_io_slow_sel[9]
port 580 nsew signal output
rlabel metal3 s 632200 71675 633437 71795 6 mprj_io_vtrip_sel[0]
port 581 nsew signal output
rlabel metal3 s 632200 654875 633437 654995 6 mprj_io_vtrip_sel[10]
port 582 nsew signal output
rlabel metal3 s 632200 699875 633437 699995 6 mprj_io_vtrip_sel[11]
port 583 nsew signal output
rlabel metal3 s 632200 744875 633437 744995 6 mprj_io_vtrip_sel[12]
port 584 nsew signal output
rlabel metal3 s 632200 834075 633437 834195 6 mprj_io_vtrip_sel[13]
port 585 nsew signal output
rlabel metal3 s 632200 923275 633437 923395 6 mprj_io_vtrip_sel[14]
port 586 nsew signal output
rlabel metal2 s 585837 952600 585893 953787 6 mprj_io_vtrip_sel[15]
port 587 nsew signal output
rlabel metal2 s 484037 952600 484093 953787 6 mprj_io_vtrip_sel[16]
port 588 nsew signal output
rlabel metal2 s 432637 952600 432693 953787 6 mprj_io_vtrip_sel[17]
port 589 nsew signal output
rlabel metal2 s 343637 952600 343693 953787 6 mprj_io_vtrip_sel[18]
port 590 nsew signal output
rlabel metal2 s 241837 952600 241893 953787 6 mprj_io_vtrip_sel[19]
port 591 nsew signal output
rlabel metal3 s 632200 116875 633437 116995 6 mprj_io_vtrip_sel[1]
port 592 nsew signal output
rlabel metal2 s 190237 952600 190293 953787 6 mprj_io_vtrip_sel[20]
port 593 nsew signal output
rlabel metal2 s 138837 952600 138893 953787 6 mprj_io_vtrip_sel[21]
port 594 nsew signal output
rlabel metal2 s 87437 952600 87493 953787 6 mprj_io_vtrip_sel[22]
port 595 nsew signal output
rlabel metal2 s 36037 952600 36093 953787 6 mprj_io_vtrip_sel[23]
port 596 nsew signal output
rlabel metal3 s -437 914205 800 914325 6 mprj_io_vtrip_sel[24]
port 597 nsew signal output
rlabel metal3 s -437 744405 800 744525 6 mprj_io_vtrip_sel[25]
port 598 nsew signal output
rlabel metal3 s -437 701205 800 701325 6 mprj_io_vtrip_sel[26]
port 599 nsew signal output
rlabel metal3 s -437 658005 800 658125 6 mprj_io_vtrip_sel[27]
port 600 nsew signal output
rlabel metal3 s -437 614805 800 614925 6 mprj_io_vtrip_sel[28]
port 601 nsew signal output
rlabel metal3 s -437 571605 800 571725 6 mprj_io_vtrip_sel[29]
port 602 nsew signal output
rlabel metal3 s 632200 161875 633437 161995 6 mprj_io_vtrip_sel[2]
port 603 nsew signal output
rlabel metal3 s -437 528405 800 528525 6 mprj_io_vtrip_sel[30]
port 604 nsew signal output
rlabel metal3 s -437 485205 800 485325 6 mprj_io_vtrip_sel[31]
port 605 nsew signal output
rlabel metal3 s -437 357605 800 357725 6 mprj_io_vtrip_sel[32]
port 606 nsew signal output
rlabel metal3 s -437 314405 800 314525 6 mprj_io_vtrip_sel[33]
port 607 nsew signal output
rlabel metal3 s -437 271205 800 271325 6 mprj_io_vtrip_sel[34]
port 608 nsew signal output
rlabel metal3 s -437 228005 800 228125 6 mprj_io_vtrip_sel[35]
port 609 nsew signal output
rlabel metal3 s -437 184805 800 184925 6 mprj_io_vtrip_sel[36]
port 610 nsew signal output
rlabel metal3 s -437 141605 800 141725 6 mprj_io_vtrip_sel[37]
port 611 nsew signal output
rlabel metal3 s 632200 207075 633437 207195 6 mprj_io_vtrip_sel[3]
port 612 nsew signal output
rlabel metal3 s 632200 252075 633437 252195 6 mprj_io_vtrip_sel[4]
port 613 nsew signal output
rlabel metal3 s 632200 297075 633437 297195 6 mprj_io_vtrip_sel[5]
port 614 nsew signal output
rlabel metal3 s 632200 342275 633437 342395 6 mprj_io_vtrip_sel[6]
port 615 nsew signal output
rlabel metal3 s 632200 519475 633437 519595 6 mprj_io_vtrip_sel[7]
port 616 nsew signal output
rlabel metal3 s 632200 564675 633437 564795 6 mprj_io_vtrip_sel[8]
port 617 nsew signal output
rlabel metal3 s 632200 609675 633437 609795 6 mprj_io_vtrip_sel[9]
port 618 nsew signal output
rlabel metal2 s 151743 -400 151799 800 6 por_l
port 619 nsew signal output
rlabel metal2 s 265955 -400 266011 800 6 porb_h
port 620 nsew signal output
rlabel metal2 s 99367 -2105 99423 800 8 rstb_h
port 621 nsew signal input
rlabel metal4 s 2184 2128 3184 950960 6 vccd
port 622 nsew power bidirectional
rlabel metal4 s 629436 2128 630436 950960 6 vccd
port 622 nsew power bidirectional
rlabel metal5 s 1976 2176 630984 4176 6 vccd
port 622 nsew power bidirectional
rlabel metal5 s 1976 947012 630984 949612 6 vccd
port 622 nsew power bidirectional
rlabel metal4 s 14184 2128 14584 950960 6 vccd
port 622 nsew power bidirectional
rlabel metal4 s 617436 2128 617836 950960 6 vccd
port 622 nsew power bidirectional
rlabel metal4 s 24784 2128 26064 197800 6 vccd
port 622 nsew power bidirectional
rlabel metal4 s 24784 919260 26064 950960 6 vccd
port 622 nsew power bidirectional
rlabel metal4 s 44784 2128 46064 34735 6 vccd
port 622 nsew power bidirectional
rlabel metal4 s 44784 124073 46064 197800 6 vccd
port 622 nsew power bidirectional
rlabel metal4 s 44784 919260 46064 950960 6 vccd
port 622 nsew power bidirectional
rlabel metal4 s 64784 2128 66064 34735 6 vccd
port 622 nsew power bidirectional
rlabel metal4 s 64784 124073 66064 197800 6 vccd
port 622 nsew power bidirectional
rlabel metal4 s 64784 919260 66064 950960 6 vccd
port 622 nsew power bidirectional
rlabel metal4 s 84784 2128 86064 34735 6 vccd
port 622 nsew power bidirectional
rlabel metal4 s 84784 124073 86064 197800 6 vccd
port 622 nsew power bidirectional
rlabel metal4 s 84784 919260 86064 950960 6 vccd
port 622 nsew power bidirectional
rlabel metal4 s 104784 2128 106064 197800 6 vccd
port 622 nsew power bidirectional
rlabel metal4 s 104784 919260 106064 950960 6 vccd
port 622 nsew power bidirectional
rlabel metal4 s 124784 2128 126064 34735 6 vccd
port 622 nsew power bidirectional
rlabel metal4 s 124784 124073 126064 197800 6 vccd
port 622 nsew power bidirectional
rlabel metal4 s 124784 919260 126064 950960 6 vccd
port 622 nsew power bidirectional
rlabel metal4 s 144784 2128 146064 34735 6 vccd
port 622 nsew power bidirectional
rlabel metal4 s 144784 124073 146064 197800 6 vccd
port 622 nsew power bidirectional
rlabel metal4 s 144784 919260 146064 950960 6 vccd
port 622 nsew power bidirectional
rlabel metal4 s 164784 2128 166064 34735 6 vccd
port 622 nsew power bidirectional
rlabel metal4 s 164784 124073 166064 197800 6 vccd
port 622 nsew power bidirectional
rlabel metal4 s 164784 919260 166064 950960 6 vccd
port 622 nsew power bidirectional
rlabel metal4 s 184784 2128 186064 197800 6 vccd
port 622 nsew power bidirectional
rlabel metal4 s 184784 919260 186064 950960 6 vccd
port 622 nsew power bidirectional
rlabel metal4 s 204784 6816 206064 197800 6 vccd
port 622 nsew power bidirectional
rlabel metal4 s 204784 919260 206064 950960 6 vccd
port 622 nsew power bidirectional
rlabel metal4 s 224784 2128 226064 197800 6 vccd
port 622 nsew power bidirectional
rlabel metal4 s 224784 919260 226064 950960 6 vccd
port 622 nsew power bidirectional
rlabel metal4 s 244784 2128 246064 197800 6 vccd
port 622 nsew power bidirectional
rlabel metal4 s 244784 919260 246064 950960 6 vccd
port 622 nsew power bidirectional
rlabel metal4 s 264784 2128 266064 197800 6 vccd
port 622 nsew power bidirectional
rlabel metal4 s 264784 919260 266064 950960 6 vccd
port 622 nsew power bidirectional
rlabel metal4 s 284784 2128 286064 197800 6 vccd
port 622 nsew power bidirectional
rlabel metal4 s 284784 919260 286064 950960 6 vccd
port 622 nsew power bidirectional
rlabel metal4 s 304784 2128 306064 197800 6 vccd
port 622 nsew power bidirectional
rlabel metal4 s 304784 919260 306064 950960 6 vccd
port 622 nsew power bidirectional
rlabel metal4 s 324784 2128 326064 35436 6 vccd
port 622 nsew power bidirectional
rlabel metal4 s 324784 56804 326064 197800 6 vccd
port 622 nsew power bidirectional
rlabel metal4 s 324784 919260 326064 950960 6 vccd
port 622 nsew power bidirectional
rlabel metal4 s 344784 2128 346064 197800 6 vccd
port 622 nsew power bidirectional
rlabel metal4 s 344784 919260 346064 950960 6 vccd
port 622 nsew power bidirectional
rlabel metal4 s 364784 2128 366064 24735 6 vccd
port 622 nsew power bidirectional
rlabel metal4 s 364784 114073 366064 197800 6 vccd
port 622 nsew power bidirectional
rlabel metal4 s 364784 919260 366064 950960 6 vccd
port 622 nsew power bidirectional
rlabel metal4 s 384784 2128 386064 24735 6 vccd
port 622 nsew power bidirectional
rlabel metal4 s 384784 114073 386064 197800 6 vccd
port 622 nsew power bidirectional
rlabel metal4 s 384784 919260 386064 950960 6 vccd
port 622 nsew power bidirectional
rlabel metal4 s 404784 2128 406064 24735 6 vccd
port 622 nsew power bidirectional
rlabel metal4 s 404784 114073 406064 197800 6 vccd
port 622 nsew power bidirectional
rlabel metal4 s 404784 919260 406064 950960 6 vccd
port 622 nsew power bidirectional
rlabel metal4 s 424784 2128 426064 197800 6 vccd
port 622 nsew power bidirectional
rlabel metal4 s 424784 919260 426064 950960 6 vccd
port 622 nsew power bidirectional
rlabel metal4 s 444784 2128 446064 197800 6 vccd
port 622 nsew power bidirectional
rlabel metal4 s 444784 919260 446064 950960 6 vccd
port 622 nsew power bidirectional
rlabel metal4 s 464784 2128 466064 197800 6 vccd
port 622 nsew power bidirectional
rlabel metal4 s 464784 919260 466064 950960 6 vccd
port 622 nsew power bidirectional
rlabel metal4 s 484784 2128 486064 197800 6 vccd
port 622 nsew power bidirectional
rlabel metal4 s 484784 919260 486064 950960 6 vccd
port 622 nsew power bidirectional
rlabel metal4 s 504784 2128 506064 197800 6 vccd
port 622 nsew power bidirectional
rlabel metal4 s 504784 919260 506064 950960 6 vccd
port 622 nsew power bidirectional
rlabel metal4 s 524784 2128 526064 197800 6 vccd
port 622 nsew power bidirectional
rlabel metal4 s 524784 919260 526064 950960 6 vccd
port 622 nsew power bidirectional
rlabel metal4 s 544784 2128 546064 38687 6 vccd
port 622 nsew power bidirectional
rlabel metal4 s 544784 146657 546064 197800 6 vccd
port 622 nsew power bidirectional
rlabel metal4 s 544784 919260 546064 920600 6 vccd
port 622 nsew power bidirectional
rlabel metal4 s 564784 2128 566064 38468 6 vccd
port 622 nsew power bidirectional
rlabel metal4 s 564784 147420 566064 197800 6 vccd
port 622 nsew power bidirectional
rlabel metal4 s 564784 919260 566064 950960 6 vccd
port 622 nsew power bidirectional
rlabel metal4 s 584784 2128 586064 38687 6 vccd
port 622 nsew power bidirectional
rlabel metal4 s 584784 146657 586064 197800 6 vccd
port 622 nsew power bidirectional
rlabel metal4 s 584784 919260 586064 950960 6 vccd
port 622 nsew power bidirectional
rlabel metal4 s 604784 2128 606064 38687 6 vccd
port 622 nsew power bidirectional
rlabel metal4 s 604784 146657 606064 197800 6 vccd
port 622 nsew power bidirectional
rlabel metal4 s 604784 919260 606064 950960 6 vccd
port 622 nsew power bidirectional
rlabel metal5 s 1976 61736 630984 63016 6 vccd
port 622 nsew power bidirectional
rlabel metal5 s 1976 85736 630984 87016 6 vccd
port 622 nsew power bidirectional
rlabel metal5 s 1976 109736 630984 111016 6 vccd
port 622 nsew power bidirectional
rlabel metal5 s 1976 133736 630984 135016 6 vccd
port 622 nsew power bidirectional
rlabel metal5 s 1976 157736 630984 159016 6 vccd
port 622 nsew power bidirectional
rlabel metal5 s 1976 181736 630984 183016 6 vccd
port 622 nsew power bidirectional
rlabel metal5 s 1976 205736 15184 207016 6 vccd
port 622 nsew power bidirectional
rlabel metal5 s 1976 229736 15184 231016 6 vccd
port 622 nsew power bidirectional
rlabel metal5 s 1976 253736 15184 255016 6 vccd
port 622 nsew power bidirectional
rlabel metal5 s 1976 277736 15184 279016 6 vccd
port 622 nsew power bidirectional
rlabel metal5 s 1976 301736 15184 303016 6 vccd
port 622 nsew power bidirectional
rlabel metal5 s 1976 325736 15184 327016 6 vccd
port 622 nsew power bidirectional
rlabel metal5 s 1976 349736 15184 351016 6 vccd
port 622 nsew power bidirectional
rlabel metal5 s 1976 373736 15184 375016 6 vccd
port 622 nsew power bidirectional
rlabel metal5 s 1976 421736 15184 423016 6 vccd
port 622 nsew power bidirectional
rlabel metal5 s 1976 469736 15184 471016 6 vccd
port 622 nsew power bidirectional
rlabel metal5 s 1976 493736 15184 495016 6 vccd
port 622 nsew power bidirectional
rlabel metal5 s 1976 517736 15184 519016 6 vccd
port 622 nsew power bidirectional
rlabel metal5 s 1976 541736 15184 543016 6 vccd
port 622 nsew power bidirectional
rlabel metal5 s 1976 565736 15184 567016 6 vccd
port 622 nsew power bidirectional
rlabel metal5 s 1976 589736 15184 591016 6 vccd
port 622 nsew power bidirectional
rlabel metal5 s 1976 613736 15184 615016 6 vccd
port 622 nsew power bidirectional
rlabel metal5 s 1976 637736 15184 639016 6 vccd
port 622 nsew power bidirectional
rlabel metal5 s 1976 661736 15184 663016 6 vccd
port 622 nsew power bidirectional
rlabel metal5 s 1976 685736 15184 687016 6 vccd
port 622 nsew power bidirectional
rlabel metal5 s 1976 709736 15184 711016 6 vccd
port 622 nsew power bidirectional
rlabel metal5 s 1976 733736 15184 735016 6 vccd
port 622 nsew power bidirectional
rlabel metal5 s 1976 757736 15184 759016 6 vccd
port 622 nsew power bidirectional
rlabel metal5 s 1976 781736 15184 783016 6 vccd
port 622 nsew power bidirectional
rlabel metal5 s 1976 805736 15184 807016 6 vccd
port 622 nsew power bidirectional
rlabel metal5 s 1976 829736 15184 831016 6 vccd
port 622 nsew power bidirectional
rlabel metal5 s 1976 853736 15184 855016 6 vccd
port 622 nsew power bidirectional
rlabel metal5 s 1976 901736 15184 903016 6 vccd
port 622 nsew power bidirectional
rlabel metal5 s 5600 37736 630984 39016 6 vccd
port 622 nsew power bidirectional
rlabel metal5 s 617436 205736 630984 207016 6 vccd
port 622 nsew power bidirectional
rlabel metal5 s 617436 229736 630984 231016 6 vccd
port 622 nsew power bidirectional
rlabel metal5 s 617436 253736 630984 255016 6 vccd
port 622 nsew power bidirectional
rlabel metal5 s 617436 277736 630984 279016 6 vccd
port 622 nsew power bidirectional
rlabel metal5 s 617436 301736 630984 303016 6 vccd
port 622 nsew power bidirectional
rlabel metal5 s 617436 325736 630984 327016 6 vccd
port 622 nsew power bidirectional
rlabel metal5 s 617436 349736 630984 351016 6 vccd
port 622 nsew power bidirectional
rlabel metal5 s 617436 397736 630984 399016 6 vccd
port 622 nsew power bidirectional
rlabel metal5 s 617436 445736 630984 447016 6 vccd
port 622 nsew power bidirectional
rlabel metal5 s 617436 493736 630984 495016 6 vccd
port 622 nsew power bidirectional
rlabel metal5 s 617436 517736 630984 519016 6 vccd
port 622 nsew power bidirectional
rlabel metal5 s 617436 541736 630984 543016 6 vccd
port 622 nsew power bidirectional
rlabel metal5 s 617436 565736 630984 567016 6 vccd
port 622 nsew power bidirectional
rlabel metal5 s 617436 589736 630984 591016 6 vccd
port 622 nsew power bidirectional
rlabel metal5 s 617436 613736 630984 615016 6 vccd
port 622 nsew power bidirectional
rlabel metal5 s 617436 637736 630984 639016 6 vccd
port 622 nsew power bidirectional
rlabel metal5 s 617436 661736 630984 663016 6 vccd
port 622 nsew power bidirectional
rlabel metal5 s 617436 685736 630984 687016 6 vccd
port 622 nsew power bidirectional
rlabel metal5 s 617436 709736 630984 711016 6 vccd
port 622 nsew power bidirectional
rlabel metal5 s 617436 733736 630984 735016 6 vccd
port 622 nsew power bidirectional
rlabel metal5 s 617436 757736 630984 759016 6 vccd
port 622 nsew power bidirectional
rlabel metal5 s 617436 805736 630984 807016 6 vccd
port 622 nsew power bidirectional
rlabel metal5 s 617436 829736 630984 831016 6 vccd
port 622 nsew power bidirectional
rlabel metal5 s 617436 853736 630984 855016 6 vccd
port 622 nsew power bidirectional
rlabel metal5 s 617436 901736 630984 903016 6 vccd
port 622 nsew power bidirectional
rlabel metal5 s 1976 48536 630984 51416 6 vccd
port 622 nsew power bidirectional
rlabel metal5 s 1976 72536 630984 75416 6 vccd
port 622 nsew power bidirectional
rlabel metal5 s 1976 96536 630984 99416 6 vccd
port 622 nsew power bidirectional
rlabel metal5 s 1976 120536 630984 123416 6 vccd
port 622 nsew power bidirectional
rlabel metal5 s 1976 144536 630984 147416 6 vccd
port 622 nsew power bidirectional
rlabel metal5 s 1976 190600 630984 193480 6 vccd
port 622 nsew power bidirectional
rlabel metal4 s 530064 928016 531064 938448 6 vccd
port 622 nsew power bidirectional
rlabel metal5 s 524784 919540 567584 919860 6 vccd
port 622 nsew power bidirectional
rlabel metal4 s 4584 2128 5584 950960 6 vccd1
port 623 nsew power bidirectional
rlabel metal4 s 627036 2128 628036 950960 6 vccd1
port 623 nsew power bidirectional
rlabel metal5 s 1976 6816 630984 8816 6 vccd1
port 623 nsew power bidirectional
rlabel metal5 s 1976 941172 630984 943772 6 vccd1
port 623 nsew power bidirectional
rlabel metal5 s 1976 163096 630984 164056 6 vccd1
port 623 nsew power bidirectional
rlabel metal4 s 255144 2128 256104 197800 6 vccd1
port 623 nsew power bidirectional
rlabel metal4 s 275144 2128 276104 197800 6 vccd1
port 623 nsew power bidirectional
rlabel metal4 s 295144 2128 296104 197800 6 vccd1
port 623 nsew power bidirectional
rlabel metal4 s 295144 919260 296104 950960 6 vccd1
port 623 nsew power bidirectional
rlabel metal4 s 52728 919260 54008 950960 6 vccd1
port 623 nsew power bidirectional
rlabel metal4 s 112728 2128 114008 197800 6 vccd1
port 623 nsew power bidirectional
rlabel metal4 s 112728 919260 114008 950960 6 vccd1
port 623 nsew power bidirectional
rlabel metal4 s 232728 2128 234008 197800 6 vccd1
port 623 nsew power bidirectional
rlabel metal4 s 232728 919260 234008 950960 6 vccd1
port 623 nsew power bidirectional
rlabel metal4 s 292728 2128 294008 197800 6 vccd1
port 623 nsew power bidirectional
rlabel metal4 s 292728 919260 294008 950960 6 vccd1
port 623 nsew power bidirectional
rlabel metal4 s 352728 2128 354008 197800 6 vccd1
port 623 nsew power bidirectional
rlabel metal4 s 352728 919260 354008 950960 6 vccd1
port 623 nsew power bidirectional
rlabel metal4 s 412728 919260 414008 950960 6 vccd1
port 623 nsew power bidirectional
rlabel metal4 s 472728 2128 474008 197800 6 vccd1
port 623 nsew power bidirectional
rlabel metal4 s 472728 919260 474008 950960 6 vccd1
port 623 nsew power bidirectional
rlabel metal4 s 552728 919260 554008 950960 6 vccd1
port 623 nsew power bidirectional
rlabel metal4 s 192728 919260 194008 950960 6 vccd1
port 623 nsew power bidirectional
rlabel metal4 s 12984 2128 13984 950960 6 vccd2
port 624 nsew power bidirectional
rlabel metal4 s 618636 2128 619636 950960 6 vccd2
port 624 nsew power bidirectional
rlabel metal5 s 1976 23056 630984 25056 6 vccd2
port 624 nsew power bidirectional
rlabel metal5 s 1976 920732 630984 923332 6 vccd2
port 624 nsew power bidirectional
rlabel metal5 s 1976 166296 630984 167256 6 vccd2
port 624 nsew power bidirectional
rlabel metal4 s 170144 124073 171104 197800 6 vccd2
port 624 nsew power bidirectional
rlabel metal4 s 180144 2128 181104 197800 6 vccd2
port 624 nsew power bidirectional
rlabel metal4 s 10584 2128 11584 950960 6 vdda1
port 625 nsew power bidirectional
rlabel metal4 s 621036 2128 622036 950960 6 vdda1
port 625 nsew power bidirectional
rlabel metal5 s 1976 18416 630984 20416 6 vdda1
port 625 nsew power bidirectional
rlabel metal5 s 1976 926572 630984 929172 6 vdda1
port 625 nsew power bidirectional
rlabel metal5 s 1976 169496 630984 170456 6 vdda1
port 625 nsew power bidirectional
rlabel metal4 s 368744 114073 369704 197800 6 vdda1
port 625 nsew power bidirectional
rlabel metal4 s 376744 114073 377704 197800 6 vdda1
port 625 nsew power bidirectional
rlabel metal4 s 8184 2128 9184 950960 6 vdda2
port 626 nsew power bidirectional
rlabel metal4 s 623436 2128 624436 950960 6 vdda2
port 626 nsew power bidirectional
rlabel metal5 s 1976 13776 630984 15776 6 vdda2
port 626 nsew power bidirectional
rlabel metal5 s 1976 932412 630984 935012 6 vdda2
port 626 nsew power bidirectional
rlabel metal5 s 1976 172696 630984 173656 6 vdda2
port 626 nsew power bidirectional
rlabel metal4 s 371944 114073 372904 197800 6 vdda2
port 626 nsew power bidirectional
rlabel metal4 s 379944 114073 380904 197800 6 vdda2
port 626 nsew power bidirectional
rlabel metal5 s 130000 29076 216423 30076 6 vddio
port 627 nsew power bidirectional
rlabel metal5 s 130000 31876 216423 32876 6 vddio
port 627 nsew power bidirectional
rlabel metal4 s 130944 2128 131904 34735 6 vddio
port 627 nsew power bidirectional
rlabel metal4 s 208144 6816 209104 37800 6 vddio
port 627 nsew power bidirectional
rlabel metal4 s 9384 2128 10384 950960 6 vssa1
port 628 nsew ground bidirectional
rlabel metal4 s 622236 2128 623236 950960 6 vssa1
port 628 nsew ground bidirectional
rlabel metal5 s 1976 16096 630984 18096 6 vssa1
port 628 nsew ground bidirectional
rlabel metal5 s 1976 929492 630984 932092 6 vssa1
port 628 nsew ground bidirectional
rlabel metal5 s 1976 171096 630984 172056 6 vssa1
port 628 nsew ground bidirectional
rlabel metal4 s 370344 114073 371304 197800 6 vssa1
port 628 nsew ground bidirectional
rlabel metal4 s 378344 114073 379304 197800 6 vssa1
port 628 nsew ground bidirectional
rlabel metal4 s 6984 2128 7984 950960 6 vssa2
port 629 nsew ground bidirectional
rlabel metal4 s 624636 2128 625636 950960 6 vssa2
port 629 nsew ground bidirectional
rlabel metal5 s 1976 11456 630984 13456 6 vssa2
port 629 nsew ground bidirectional
rlabel metal5 s 1976 935332 630984 937932 6 vssa2
port 629 nsew ground bidirectional
rlabel metal5 s 1976 174296 630984 175256 6 vssa2
port 629 nsew ground bidirectional
rlabel metal4 s 373544 114073 374504 197800 6 vssa2
port 629 nsew ground bidirectional
rlabel metal4 s 381544 114073 382504 197800 6 vssa2
port 629 nsew ground bidirectional
rlabel metal4 s 3384 2128 4384 950960 6 vssd
port 630 nsew ground bidirectional
rlabel metal4 s 628236 2128 629236 950960 6 vssd
port 630 nsew ground bidirectional
rlabel metal5 s 1976 4496 630984 6496 6 vssd
port 630 nsew ground bidirectional
rlabel metal5 s 1976 944092 630984 946692 6 vssd
port 630 nsew ground bidirectional
rlabel metal4 s 14784 2128 15184 950960 6 vssd
port 630 nsew ground bidirectional
rlabel metal4 s 618036 2128 618436 950960 6 vssd
port 630 nsew ground bidirectional
rlabel metal4 s 26304 2128 27584 197800 6 vssd
port 630 nsew ground bidirectional
rlabel metal4 s 26304 919260 27584 950960 6 vssd
port 630 nsew ground bidirectional
rlabel metal4 s 46304 2128 47584 34735 6 vssd
port 630 nsew ground bidirectional
rlabel metal4 s 46304 124073 47584 197800 6 vssd
port 630 nsew ground bidirectional
rlabel metal4 s 46304 919260 47584 950960 6 vssd
port 630 nsew ground bidirectional
rlabel metal4 s 66304 2128 67584 34735 6 vssd
port 630 nsew ground bidirectional
rlabel metal4 s 66304 124073 67584 197800 6 vssd
port 630 nsew ground bidirectional
rlabel metal4 s 66304 919260 67584 950960 6 vssd
port 630 nsew ground bidirectional
rlabel metal4 s 86304 2128 87584 34735 6 vssd
port 630 nsew ground bidirectional
rlabel metal4 s 86304 124073 87584 197800 6 vssd
port 630 nsew ground bidirectional
rlabel metal4 s 86304 919260 87584 950960 6 vssd
port 630 nsew ground bidirectional
rlabel metal4 s 106304 2128 107584 197800 6 vssd
port 630 nsew ground bidirectional
rlabel metal4 s 106304 919260 107584 950960 6 vssd
port 630 nsew ground bidirectional
rlabel metal4 s 126304 2128 127584 34735 6 vssd
port 630 nsew ground bidirectional
rlabel metal4 s 126304 124073 127584 197800 6 vssd
port 630 nsew ground bidirectional
rlabel metal4 s 126304 919260 127584 950960 6 vssd
port 630 nsew ground bidirectional
rlabel metal4 s 146304 2128 147584 33836 6 vssd
port 630 nsew ground bidirectional
rlabel metal4 s 146304 124073 147584 197800 6 vssd
port 630 nsew ground bidirectional
rlabel metal4 s 146304 919260 147584 950960 6 vssd
port 630 nsew ground bidirectional
rlabel metal4 s 166304 2128 167584 34735 6 vssd
port 630 nsew ground bidirectional
rlabel metal4 s 166304 124073 167584 197800 6 vssd
port 630 nsew ground bidirectional
rlabel metal4 s 166304 919260 167584 950960 6 vssd
port 630 nsew ground bidirectional
rlabel metal4 s 186304 2128 187584 197800 6 vssd
port 630 nsew ground bidirectional
rlabel metal4 s 186304 919260 187584 950960 6 vssd
port 630 nsew ground bidirectional
rlabel metal4 s 206304 6816 207584 197800 6 vssd
port 630 nsew ground bidirectional
rlabel metal4 s 206304 919260 207584 950960 6 vssd
port 630 nsew ground bidirectional
rlabel metal4 s 226304 2128 227584 197800 6 vssd
port 630 nsew ground bidirectional
rlabel metal4 s 226304 919260 227584 950960 6 vssd
port 630 nsew ground bidirectional
rlabel metal4 s 246304 2128 247584 197800 6 vssd
port 630 nsew ground bidirectional
rlabel metal4 s 246304 919260 247584 950960 6 vssd
port 630 nsew ground bidirectional
rlabel metal4 s 266304 2128 267584 197800 6 vssd
port 630 nsew ground bidirectional
rlabel metal4 s 266304 919260 267584 950960 6 vssd
port 630 nsew ground bidirectional
rlabel metal4 s 286304 2128 287584 197800 6 vssd
port 630 nsew ground bidirectional
rlabel metal4 s 286304 919260 287584 950960 6 vssd
port 630 nsew ground bidirectional
rlabel metal4 s 306304 2128 307584 197800 6 vssd
port 630 nsew ground bidirectional
rlabel metal4 s 306304 919260 307584 950960 6 vssd
port 630 nsew ground bidirectional
rlabel metal4 s 326304 2128 327584 35436 6 vssd
port 630 nsew ground bidirectional
rlabel metal4 s 326304 56804 327584 197800 6 vssd
port 630 nsew ground bidirectional
rlabel metal4 s 326304 919260 327584 950960 6 vssd
port 630 nsew ground bidirectional
rlabel metal4 s 346304 2128 347584 197800 6 vssd
port 630 nsew ground bidirectional
rlabel metal4 s 346304 919260 347584 950960 6 vssd
port 630 nsew ground bidirectional
rlabel metal4 s 366304 2128 367584 24735 6 vssd
port 630 nsew ground bidirectional
rlabel metal4 s 366304 114073 367584 197800 6 vssd
port 630 nsew ground bidirectional
rlabel metal4 s 366304 919260 367584 950960 6 vssd
port 630 nsew ground bidirectional
rlabel metal4 s 386304 2128 387584 24735 6 vssd
port 630 nsew ground bidirectional
rlabel metal4 s 386304 114073 387584 197800 6 vssd
port 630 nsew ground bidirectional
rlabel metal4 s 386304 919260 387584 950960 6 vssd
port 630 nsew ground bidirectional
rlabel metal4 s 406304 2128 407584 23836 6 vssd
port 630 nsew ground bidirectional
rlabel metal4 s 406304 114073 407584 197800 6 vssd
port 630 nsew ground bidirectional
rlabel metal4 s 406304 919260 407584 950960 6 vssd
port 630 nsew ground bidirectional
rlabel metal4 s 426304 2128 427584 197800 6 vssd
port 630 nsew ground bidirectional
rlabel metal4 s 426304 919260 427584 950960 6 vssd
port 630 nsew ground bidirectional
rlabel metal4 s 446304 2128 447584 197800 6 vssd
port 630 nsew ground bidirectional
rlabel metal4 s 446304 919260 447584 950960 6 vssd
port 630 nsew ground bidirectional
rlabel metal4 s 466304 2128 467584 197800 6 vssd
port 630 nsew ground bidirectional
rlabel metal4 s 466304 919260 467584 950960 6 vssd
port 630 nsew ground bidirectional
rlabel metal4 s 486304 2128 487584 197800 6 vssd
port 630 nsew ground bidirectional
rlabel metal4 s 486304 919260 487584 950960 6 vssd
port 630 nsew ground bidirectional
rlabel metal4 s 506304 2128 507584 197800 6 vssd
port 630 nsew ground bidirectional
rlabel metal4 s 506304 919260 507584 950960 6 vssd
port 630 nsew ground bidirectional
rlabel metal4 s 526304 2128 527584 197800 6 vssd
port 630 nsew ground bidirectional
rlabel metal4 s 526304 919260 527584 950960 6 vssd
port 630 nsew ground bidirectional
rlabel metal4 s 546304 2128 547584 38687 6 vssd
port 630 nsew ground bidirectional
rlabel metal4 s 546304 146657 547584 197800 6 vssd
port 630 nsew ground bidirectional
rlabel metal4 s 546304 919260 547584 920600 6 vssd
port 630 nsew ground bidirectional
rlabel metal4 s 566304 2128 567584 38687 6 vssd
port 630 nsew ground bidirectional
rlabel metal4 s 566304 146657 567584 197800 6 vssd
port 630 nsew ground bidirectional
rlabel metal4 s 566304 919260 567584 950960 6 vssd
port 630 nsew ground bidirectional
rlabel metal4 s 586304 2128 587584 38687 6 vssd
port 630 nsew ground bidirectional
rlabel metal4 s 586304 146657 587584 197800 6 vssd
port 630 nsew ground bidirectional
rlabel metal4 s 586304 919260 587584 950960 6 vssd
port 630 nsew ground bidirectional
rlabel metal4 s 606304 2128 607584 38687 6 vssd
port 630 nsew ground bidirectional
rlabel metal4 s 606304 146657 607584 197800 6 vssd
port 630 nsew ground bidirectional
rlabel metal4 s 606304 919260 607584 950960 6 vssd
port 630 nsew ground bidirectional
rlabel metal5 s 1976 63496 630984 64776 6 vssd
port 630 nsew ground bidirectional
rlabel metal5 s 1976 87496 630984 88776 6 vssd
port 630 nsew ground bidirectional
rlabel metal5 s 1976 111496 630984 112776 6 vssd
port 630 nsew ground bidirectional
rlabel metal5 s 1976 135496 630984 136776 6 vssd
port 630 nsew ground bidirectional
rlabel metal5 s 1976 159496 630984 160776 6 vssd
port 630 nsew ground bidirectional
rlabel metal5 s 1976 183496 630984 184776 6 vssd
port 630 nsew ground bidirectional
rlabel metal5 s 1976 207496 15184 208776 6 vssd
port 630 nsew ground bidirectional
rlabel metal5 s 1976 231496 15184 232776 6 vssd
port 630 nsew ground bidirectional
rlabel metal5 s 1976 255496 15184 256776 6 vssd
port 630 nsew ground bidirectional
rlabel metal5 s 1976 279496 15184 280776 6 vssd
port 630 nsew ground bidirectional
rlabel metal5 s 1976 303496 15184 304776 6 vssd
port 630 nsew ground bidirectional
rlabel metal5 s 1976 327496 15184 328776 6 vssd
port 630 nsew ground bidirectional
rlabel metal5 s 1976 351496 15184 352776 6 vssd
port 630 nsew ground bidirectional
rlabel metal5 s 1976 375496 15184 376776 6 vssd
port 630 nsew ground bidirectional
rlabel metal5 s 1976 423496 15184 424776 6 vssd
port 630 nsew ground bidirectional
rlabel metal5 s 1976 471496 15184 472776 6 vssd
port 630 nsew ground bidirectional
rlabel metal5 s 1976 495496 15184 496776 6 vssd
port 630 nsew ground bidirectional
rlabel metal5 s 1976 519496 15184 520776 6 vssd
port 630 nsew ground bidirectional
rlabel metal5 s 1976 543496 15184 544776 6 vssd
port 630 nsew ground bidirectional
rlabel metal5 s 1976 567496 15184 568776 6 vssd
port 630 nsew ground bidirectional
rlabel metal5 s 1976 591496 15184 592776 6 vssd
port 630 nsew ground bidirectional
rlabel metal5 s 1976 615496 15184 616776 6 vssd
port 630 nsew ground bidirectional
rlabel metal5 s 1976 639496 15184 640776 6 vssd
port 630 nsew ground bidirectional
rlabel metal5 s 1976 663496 15184 664776 6 vssd
port 630 nsew ground bidirectional
rlabel metal5 s 1976 687496 15184 688776 6 vssd
port 630 nsew ground bidirectional
rlabel metal5 s 1976 711496 15184 712776 6 vssd
port 630 nsew ground bidirectional
rlabel metal5 s 1976 735496 15184 736776 6 vssd
port 630 nsew ground bidirectional
rlabel metal5 s 1976 759496 15184 760776 6 vssd
port 630 nsew ground bidirectional
rlabel metal5 s 1976 783496 15184 784776 6 vssd
port 630 nsew ground bidirectional
rlabel metal5 s 1976 807496 15184 808776 6 vssd
port 630 nsew ground bidirectional
rlabel metal5 s 1976 831496 15184 832776 6 vssd
port 630 nsew ground bidirectional
rlabel metal5 s 1976 855496 15184 856776 6 vssd
port 630 nsew ground bidirectional
rlabel metal5 s 1976 903496 15184 904776 6 vssd
port 630 nsew ground bidirectional
rlabel metal5 s 5600 39496 630984 40776 6 vssd
port 630 nsew ground bidirectional
rlabel metal5 s 617436 207496 630984 208776 6 vssd
port 630 nsew ground bidirectional
rlabel metal5 s 617436 231496 630984 232776 6 vssd
port 630 nsew ground bidirectional
rlabel metal5 s 617436 255496 630984 256776 6 vssd
port 630 nsew ground bidirectional
rlabel metal5 s 617436 279496 630984 280776 6 vssd
port 630 nsew ground bidirectional
rlabel metal5 s 617436 303496 630984 304776 6 vssd
port 630 nsew ground bidirectional
rlabel metal5 s 617436 327496 630984 328776 6 vssd
port 630 nsew ground bidirectional
rlabel metal5 s 617436 351496 630984 352776 6 vssd
port 630 nsew ground bidirectional
rlabel metal5 s 617436 399496 630984 400776 6 vssd
port 630 nsew ground bidirectional
rlabel metal5 s 617436 447496 630984 448776 6 vssd
port 630 nsew ground bidirectional
rlabel metal5 s 617436 495496 630984 496776 6 vssd
port 630 nsew ground bidirectional
rlabel metal5 s 617436 519496 630984 520776 6 vssd
port 630 nsew ground bidirectional
rlabel metal5 s 617436 543496 630984 544776 6 vssd
port 630 nsew ground bidirectional
rlabel metal5 s 617436 567496 630984 568776 6 vssd
port 630 nsew ground bidirectional
rlabel metal5 s 617436 591496 630984 592776 6 vssd
port 630 nsew ground bidirectional
rlabel metal5 s 617436 615496 630984 616776 6 vssd
port 630 nsew ground bidirectional
rlabel metal5 s 617436 639496 630984 640776 6 vssd
port 630 nsew ground bidirectional
rlabel metal5 s 617436 663496 630984 664776 6 vssd
port 630 nsew ground bidirectional
rlabel metal5 s 617436 687496 630984 688776 6 vssd
port 630 nsew ground bidirectional
rlabel metal5 s 617436 711496 630984 712776 6 vssd
port 630 nsew ground bidirectional
rlabel metal5 s 617436 735496 630984 736776 6 vssd
port 630 nsew ground bidirectional
rlabel metal5 s 617436 759496 630984 760776 6 vssd
port 630 nsew ground bidirectional
rlabel metal5 s 617436 807496 630984 808776 6 vssd
port 630 nsew ground bidirectional
rlabel metal5 s 617436 831496 630984 832776 6 vssd
port 630 nsew ground bidirectional
rlabel metal5 s 617436 855496 630984 856776 6 vssd
port 630 nsew ground bidirectional
rlabel metal5 s 617436 903496 630984 904776 6 vssd
port 630 nsew ground bidirectional
rlabel metal5 s 1976 51896 630984 54776 6 vssd
port 630 nsew ground bidirectional
rlabel metal5 s 1976 75896 630984 78776 6 vssd
port 630 nsew ground bidirectional
rlabel metal5 s 1976 99896 630984 102776 6 vssd
port 630 nsew ground bidirectional
rlabel metal5 s 1976 123896 630984 126776 6 vssd
port 630 nsew ground bidirectional
rlabel metal5 s 1976 147896 630984 150776 6 vssd
port 630 nsew ground bidirectional
rlabel metal5 s 1976 193960 630984 196840 6 vssd
port 630 nsew ground bidirectional
rlabel metal4 s 531352 928016 532352 938448 6 vssd
port 630 nsew ground bidirectional
rlabel metal4 s 5784 2128 6784 950960 6 vssd1
port 631 nsew ground bidirectional
rlabel metal4 s 625836 2128 626836 950960 6 vssd1
port 631 nsew ground bidirectional
rlabel metal5 s 1976 9136 630984 11136 6 vssd1
port 631 nsew ground bidirectional
rlabel metal5 s 1976 938252 630984 940852 6 vssd1
port 631 nsew ground bidirectional
rlabel metal5 s 1976 164696 630984 165656 6 vssd1
port 631 nsew ground bidirectional
rlabel metal4 s 256744 2128 257704 197800 6 vssd1
port 631 nsew ground bidirectional
rlabel metal4 s 276744 2128 277704 197800 6 vssd1
port 631 nsew ground bidirectional
rlabel metal4 s 296744 2128 297704 197800 6 vssd1
port 631 nsew ground bidirectional
rlabel metal4 s 51208 919260 52488 950960 6 vssd1
port 631 nsew ground bidirectional
rlabel metal4 s 111208 2128 112488 197800 6 vssd1
port 631 nsew ground bidirectional
rlabel metal4 s 111208 919260 112488 950960 6 vssd1
port 631 nsew ground bidirectional
rlabel metal4 s 231208 2128 232488 197800 6 vssd1
port 631 nsew ground bidirectional
rlabel metal4 s 231208 919260 232488 950960 6 vssd1
port 631 nsew ground bidirectional
rlabel metal4 s 291208 2128 292488 197800 6 vssd1
port 631 nsew ground bidirectional
rlabel metal4 s 291208 919260 292488 950960 6 vssd1
port 631 nsew ground bidirectional
rlabel metal4 s 351208 2128 352488 197800 6 vssd1
port 631 nsew ground bidirectional
rlabel metal4 s 351208 919260 352488 950960 6 vssd1
port 631 nsew ground bidirectional
rlabel metal4 s 411208 919260 412488 950960 6 vssd1
port 631 nsew ground bidirectional
rlabel metal4 s 471208 2128 472488 197800 6 vssd1
port 631 nsew ground bidirectional
rlabel metal4 s 471208 919260 472488 950960 6 vssd1
port 631 nsew ground bidirectional
rlabel metal4 s 551208 919260 552488 950960 6 vssd1
port 631 nsew ground bidirectional
rlabel metal4 s 191208 2128 192488 197800 6 vssd1
port 631 nsew ground bidirectional
rlabel metal4 s 191208 919260 192488 950960 6 vssd1
port 631 nsew ground bidirectional
rlabel metal4 s 11784 2128 12784 950960 6 vssd2
port 632 nsew ground bidirectional
rlabel metal4 s 619836 2128 620836 950960 6 vssd2
port 632 nsew ground bidirectional
rlabel metal5 s 1976 20736 630984 22736 6 vssd2
port 632 nsew ground bidirectional
rlabel metal5 s 1976 923652 630984 926252 6 vssd2
port 632 nsew ground bidirectional
rlabel metal5 s 1976 167896 630984 168856 6 vssd2
port 632 nsew ground bidirectional
rlabel metal4 s 171744 124073 172704 197800 6 vssd2
port 632 nsew ground bidirectional
rlabel metal4 s 181744 2128 182704 197800 6 vssd2
port 632 nsew ground bidirectional
rlabel metal5 s 130000 30476 216423 31476 6 vssio
port 633 nsew ground bidirectional
rlabel metal5 s 130000 33276 216423 34276 6 vssio
port 633 nsew ground bidirectional
rlabel metal4 s 132304 2128 133264 33836 6 vssio
port 633 nsew ground bidirectional
rlabel metal4 s 209504 6816 210464 37800 6 vssio
port 633 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 633000 953400
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 256243992
string GDS_FILE /home/hosni/caravel-redesign-2/caravel/openlane/caravel_core/runs/23_04_11_05_23/results/signoff/caravel_core.magic.gds
string GDS_START 63666460
<< end >>

