VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO digital_locked_loop
  CLASS BLOCK ;
  FOREIGN digital_locked_loop ;
  ORIGIN 0.000 0.000 ;
  SIZE 100.000 BY 75.000 ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met2 ;
        RECT 41.040 5.200 42.640 68.240 ;
    END
    PORT
      LAYER met2 ;
        RECT 81.040 5.200 82.640 68.240 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.280 41.050 94.540 42.650 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met2 ;
        RECT 21.040 5.200 22.640 68.240 ;
    END
    PORT
      LAYER met2 ;
        RECT 61.040 5.200 62.640 68.240 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.280 21.050 94.540 22.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.280 61.050 94.540 62.650 ;
    END
  END VPWR
  PIN clockp[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 5.480 4.000 6.080 ;
    END
  END clockp[0]
  PIN clockp[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 9.560 4.000 10.160 ;
    END
  END clockp[1]
  PIN dco
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 38.120 4.000 38.720 ;
    END
  END dco
  PIN div[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 13.640 4.000 14.240 ;
    END
  END div[0]
  PIN div[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 17.720 4.000 18.320 ;
    END
  END div[1]
  PIN div[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 21.800 4.000 22.400 ;
    END
  END div[2]
  PIN div[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 25.880 4.000 26.480 ;
    END
  END div[3]
  PIN div[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 29.960 4.000 30.560 ;
    END
  END div[4]
  PIN enable
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 34.040 4.000 34.640 ;
    END
  END enable
  PIN ext_trim[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 42.200 4.000 42.800 ;
    END
  END ext_trim[0]
  PIN ext_trim[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 27.690 71.000 27.970 75.000 ;
    END
  END ext_trim[10]
  PIN ext_trim[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.050 71.000 35.330 75.000 ;
    END
  END ext_trim[11]
  PIN ext_trim[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 42.410 71.000 42.690 75.000 ;
    END
  END ext_trim[12]
  PIN ext_trim[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 49.770 71.000 50.050 75.000 ;
    END
  END ext_trim[13]
  PIN ext_trim[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 57.130 71.000 57.410 75.000 ;
    END
  END ext_trim[14]
  PIN ext_trim[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.490 71.000 64.770 75.000 ;
    END
  END ext_trim[15]
  PIN ext_trim[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 71.850 71.000 72.130 75.000 ;
    END
  END ext_trim[16]
  PIN ext_trim[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 79.210 71.000 79.490 75.000 ;
    END
  END ext_trim[17]
  PIN ext_trim[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 86.570 71.000 86.850 75.000 ;
    END
  END ext_trim[18]
  PIN ext_trim[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.930 71.000 94.210 75.000 ;
    END
  END ext_trim[19]
  PIN ext_trim[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 46.280 4.000 46.880 ;
    END
  END ext_trim[1]
  PIN ext_trim[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 66.680 100.000 67.280 ;
    END
  END ext_trim[20]
  PIN ext_trim[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 54.440 100.000 55.040 ;
    END
  END ext_trim[21]
  PIN ext_trim[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 42.200 100.000 42.800 ;
    END
  END ext_trim[22]
  PIN ext_trim[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 29.960 100.000 30.560 ;
    END
  END ext_trim[23]
  PIN ext_trim[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 17.720 100.000 18.320 ;
    END
  END ext_trim[24]
  PIN ext_trim[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 5.480 100.000 6.080 ;
    END
  END ext_trim[25]
  PIN ext_trim[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 50.360 4.000 50.960 ;
    END
  END ext_trim[2]
  PIN ext_trim[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 54.440 4.000 55.040 ;
    END
  END ext_trim[3]
  PIN ext_trim[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 58.520 4.000 59.120 ;
    END
  END ext_trim[4]
  PIN ext_trim[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 62.600 4.000 63.200 ;
    END
  END ext_trim[5]
  PIN ext_trim[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 66.680 4.000 67.280 ;
    END
  END ext_trim[6]
  PIN ext_trim[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 5.610 71.000 5.890 75.000 ;
    END
  END ext_trim[7]
  PIN ext_trim[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.970 71.000 13.250 75.000 ;
    END
  END ext_trim[8]
  PIN ext_trim[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 20.330 71.000 20.610 75.000 ;
    END
  END ext_trim[9]
  PIN osc
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 74.610 0.000 74.890 4.000 ;
    END
  END osc
  PIN resetb
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 24.930 0.000 25.210 4.000 ;
    END
  END resetb
  OBS
      LAYER li1 ;
        RECT 5.520 5.355 94.300 68.085 ;
      LAYER met1 ;
        RECT 4.670 4.800 94.600 69.660 ;
      LAYER met2 ;
        RECT 4.690 70.720 5.330 71.810 ;
        RECT 6.170 70.720 12.690 71.810 ;
        RECT 13.530 70.720 20.050 71.810 ;
        RECT 20.890 70.720 27.410 71.810 ;
        RECT 28.250 70.720 34.770 71.810 ;
        RECT 35.610 70.720 42.130 71.810 ;
        RECT 42.970 70.720 49.490 71.810 ;
        RECT 50.330 70.720 56.850 71.810 ;
        RECT 57.690 70.720 64.210 71.810 ;
        RECT 65.050 70.720 71.570 71.810 ;
        RECT 72.410 70.720 78.930 71.810 ;
        RECT 79.770 70.720 86.290 71.810 ;
        RECT 87.130 70.720 93.650 71.810 ;
        RECT 4.690 68.520 94.210 70.720 ;
        RECT 4.690 4.920 20.760 68.520 ;
        RECT 22.920 4.920 40.760 68.520 ;
        RECT 42.920 4.920 60.760 68.520 ;
        RECT 62.920 4.920 80.760 68.520 ;
        RECT 82.920 4.920 94.210 68.520 ;
        RECT 4.690 4.280 94.210 4.920 ;
        RECT 4.690 4.000 24.650 4.280 ;
        RECT 25.490 4.000 74.330 4.280 ;
        RECT 75.170 4.000 94.210 4.280 ;
      LAYER met3 ;
        RECT 4.400 66.280 95.600 67.145 ;
        RECT 3.990 63.600 96.000 66.280 ;
        RECT 4.400 63.050 96.000 63.600 ;
        RECT 4.400 62.200 4.880 63.050 ;
        RECT 3.990 60.650 4.880 62.200 ;
        RECT 94.940 60.650 96.000 63.050 ;
        RECT 3.990 59.520 96.000 60.650 ;
        RECT 4.400 58.120 96.000 59.520 ;
        RECT 3.990 55.440 96.000 58.120 ;
        RECT 4.400 54.040 95.600 55.440 ;
        RECT 3.990 51.360 96.000 54.040 ;
        RECT 4.400 49.960 96.000 51.360 ;
        RECT 3.990 47.280 96.000 49.960 ;
        RECT 4.400 45.880 96.000 47.280 ;
        RECT 3.990 43.200 96.000 45.880 ;
        RECT 4.400 43.050 95.600 43.200 ;
        RECT 4.400 41.800 4.880 43.050 ;
        RECT 3.990 40.650 4.880 41.800 ;
        RECT 94.940 41.800 95.600 43.050 ;
        RECT 94.940 40.650 96.000 41.800 ;
        RECT 3.990 39.120 96.000 40.650 ;
        RECT 4.400 37.720 96.000 39.120 ;
        RECT 3.990 35.040 96.000 37.720 ;
        RECT 4.400 33.640 96.000 35.040 ;
        RECT 3.990 30.960 96.000 33.640 ;
        RECT 4.400 29.560 95.600 30.960 ;
        RECT 3.990 26.880 96.000 29.560 ;
        RECT 4.400 25.480 96.000 26.880 ;
        RECT 3.990 23.050 96.000 25.480 ;
        RECT 3.990 22.800 4.880 23.050 ;
        RECT 4.400 21.400 4.880 22.800 ;
        RECT 3.990 20.650 4.880 21.400 ;
        RECT 94.940 20.650 96.000 23.050 ;
        RECT 3.990 18.720 96.000 20.650 ;
        RECT 4.400 17.320 95.600 18.720 ;
        RECT 3.990 14.640 96.000 17.320 ;
        RECT 4.400 13.240 96.000 14.640 ;
        RECT 3.990 10.560 96.000 13.240 ;
        RECT 4.400 9.160 96.000 10.560 ;
        RECT 3.990 6.480 96.000 9.160 ;
        RECT 4.400 5.615 95.600 6.480 ;
  END
END digital_locked_loop
END LIBRARY

